// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bxhwJ15ctlkvAv/cg4c3IYNDpCujFd7zKSTl3KkmYOKmRko+5DM1O6wHBLE8GSrx
TKKupGTdmfWhol3FBoxe3+s2O/2rOacIp0wj7dC9df34s/sswmPVGWJuXK0dbNsw
0+2FAum4jTO6RHNpw2oC8a3hpHb9RJ1Gp8KdWEUH0k0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6240)
ND+goM141MCiWT+gM6+zrnxAzCgZMkrvCilCpyYAxng9iTOXwGWrzMzixAIdGaQN
EJoQ6nguOUtbMXpeap+Xqj8qm4JCnUwdoQ1k2Tn6CZOUY0CpcLRPtQlaYROoyNqI
qXMPHBlSWu0Am0CHcPto+owsULf7tRpQ15I2cFXvM3istwge9UgZThiQFkigKXJP
QGJxKhgSlynNuXlBJyRmSbEvL/IrcM3mKciY4NMmGQeubxuX6pBQP9vct3uhT8tr
zf1bb8FDhTEub3881d3O+pVK8qOjnM8pFw4HzWP9geH1n5iRv2yIHgXD8DzQmUE+
jd6zFmfk8jyfm68Qv3fW5LXGkrnikAY2N6CiDmKSRVjR5s9ORy0gvoNKA2FHVHXu
F9YZsqBkiWTvQeBuDqyz+YIMG9MJBH9jRh0PCjfeEyd0/CsIP6bZhTdFITJl2egN
FVf7vtUWFE2+DrwOPiANePDSQBvAj4VKcAQSNAOYAiYBo6OCdixpPh4B5pAcsHyT
ZfGnaOlZ5WQYkXaoXujOSEEfZr+yNZ8GCQfa0oJ/BvXsP07+UOARdOrR4+IFhG7g
a9K5uFnpioPTS0C7IdmftcCqnjWHpcqkUT1VaHcMajw8BkSHmyLR9CRRVki3ZXTQ
dZOBF5ukF/erWXhsjiPn9sXGNUTfXoGgAKcVu32oIfBUgyT94az1YbNKMqTyMW5f
FMGLXe7PWBLAojuoKTv/6acr5M3s3lYKQmMsWr59+/6c5nGno7yXuO2kYsJGYxMe
HtB0CTyOrOJb9pL8tO6XgwouVsl7tbcbLYbUhE1VYHL2/TY4b/N1rjSTIYh2nwFn
Bn8SQ5F3Q+cU1ihNon5msuV4MWysbxSagFlMaF7CAPt3Ol1BWGIRwxQmaoJjQkxM
2y9+K8++5dk1q8C8XhRG2D+mKT7WH77xf7S8rmnsiUYmM61SaYwtmaw/KsRdI/Qt
4x+GiDz5hlHWAUfxHb01ctceIVvdKAgGSAQaF3fy6/uxAC8klN1Qj2yYH3OUH1Ca
B3NamNKK3UzHHscUKIbuncDFFFwIVAXQ4rXlIHMndwmE9DIXmNoYCZbVlKhMnaHY
0qLalpL/O1n0xo4ciVsmXoB0Rm88gEa5wm2cR2wM9t0JYFbSDBwz3uOj+0VyCgxK
O1B4H7eqdidSMd1X5m4J/Z1R9b9c/wyGMn7FE7UtJi+YyC+g5F0/leZ7rrgpP7bR
nE3T8N7pqrffQoj9ck0s3FaRtUaX13ZFU+8hbKYvUcyWre8lYO4wQTJ19Us8SAAi
PY6kkiNiXq3q8CsfOUA/++4H5pvKybsRx9ruyWdRPBBwrRStl9YYMayV/SqCR1KM
7dtXIB5UW2txhkltrQXezhkCip6sGvdmbyhcjYMn1qGs/xlTO5Og1KGGaZfLt3os
xGQsqT4sVJp8tHZ3ksHWehDwhiMVkLXScrXtNm/HqrLAtcQ8vRQghJisNRecZ3wz
oyzlreE5AFS3Wq/AYoceYcjvYqZ982T5yeihVCJFXBRmQTnpqHREk69rsZU3miDG
9AbLBY8u0UV4c3JDBgahvL2lcezUqBo2vXrWx+UGh4srNfnnHLyMAFvDLHh/wxFl
Ajjq9DwjhTByGC5DUPapGPjnriTUHM3EdAn356CrSH9Fbpmq83Ef3Az8Y0dWr5+e
A2QdrFNDwJPyFmWVSxj+vTN694INJkDQxj5P373579sGGP9GPv+trPzaQg0YYcbl
ybPXTE/RctznMH/ih7mXa7unEWe7RbyRkhFtL/03OkrlCsYYRFDALj1ZU8ZyDVpy
li65pdtjNA6uf08jWyVEVgquoEfYsiHj+YjRZRankYXoQ69r70Q0C8Wc2ci5seT5
L/kb+b5uczTLwkU7Ct24ACIoFuPtwUg1MssHSskfHlsbzVr6KaV4V5rjFWysgdlB
bIa4VE/RTIJijaxUKWJJi07O4XO0V9oXPTwKLgWx4GmyU+BgKKzqSdo/JJVwCo8J
8G1MBOWGHT7jWYWUShj4jSYUlepXlHBhye1HNuQ4gGryMBb3AfQsE2H5DaXY+H9z
VN1FkbOafTf+ac5wQCMvKJAx1/rKEpY0KrsTOpC2Jq9AEk5olc7xRpnj7qovsIfF
lZ5BW0uc9qWfEpsM8IEE9tKAhbr68mJNAcBvdg9tcLve/dd2w9iI6E2OL2tY9I5R
TSrhqaZeZ3uhRZPToX+mhCcgzt8X33fSUV71AWr9seTJHOc/cE6Czcg6F+YXJD9V
2Svz9vg4bBVIeFow+DTzNkBxj0+fRFVN/LvTEEdl4NWYmv5+Lz7uplp+zDve6g0s
xQwEiouhMSMUawAOPzsDzU6QVfgw5/RgLC44IAu/YSTXq8IhhqSvjp9tsZWR2hPd
OeGmElJAsvAdPbOPHprPJLxkFxsTEs6rOuT7ItsTdR71I3QpbfylnrKvR0gWZGto
WpQu22zApkEjDY6Z1PWkivPbykqn59e2ZurTRWtgzKSt1G6psCcfWJQsmBPapIpQ
EPtVxjKam4VLpaBsbQVzN/KpNHYv6sG0NjfNczR8lfs/GOpIIIDa5p++Ul1kJTBX
r41OtrewCWF6RnmL/B1Psmrr9E1xpUX2b6YJNodmNYaJyel4vKoBq0L7KVPh47TY
YlxbwtXINAevtmTA49bsRAgBOdFc2Z5GKs8Jhm1tuljDlbN67lVi6j6K38rwX04c
90e5SoTAQ4ENgXmjucVWOtYmV/U/vhuzpyeaabzcwFF3eyKAM60KlhbFjTDfFFkn
S2JArvOkz/D8qCiZr/iwYsHf5JMo3qJR1fTmW1wpp+eyDoidqGPPUf+Cy/l4B6rK
rW0jYi3ax45FSBluSe/0FVUfyA9yoM8eRA1eevD61tW59pqH429XQMXG5whcrh0P
5BqUe1ynYf/2TO3VcS1nwAcY7MsKyXE+ti+n/0TBkWuHCwHI0kQ52pt3EEaNje45
qLbpiclRxTavkLYNd6BvNqC6nGFNRLnKAmMJh8dwtFJldULxxEq0tndwKmfwfBGm
fstGXuuEKXzR/nWiv+GQNnR97ZIYCtnVqk/RsKOksg2kNLDvHKumG1J4aJzRC6/Y
cw1bZ5koxKQfBLJrLl8YncePScQlGyeKZb8XjVTeo9UvWrmbf3JDDxioyTenZJFq
AhgD2dHJ1X00b5WgwosF4xVHxqy6gsb1KqxAzmoObDOJrgPMfnjWrXExNsIAHy8B
iaXpVioDoLu6acOMlvVzRkEHFqDZqvRi9iyUdCnGWRpHGQQoGyDn1QwWFasZ6G/O
sgZ0RCl+e12G+7LPCh9zNSpnX4gTjo+cE4zRQnm2SFtF8zFuDxrHn6BRF2/JHhoK
cQOYi4Omx9BCmwpKiPnc1BaKjev/bOumGeb5N1HHyPm6anCOL+vWNUplmNklSjuh
y5Hcrq0/46UGu9oPRLj1MvCTriFr1aIrU3KfT3/M6bzmIOwQWMRm2ITAi06dRJIY
ZRcEQtdji6Q2qEORGfub3fa0YaJRMEovLZ2G3UZ+utmCrFMWLzvLetEeY1NbNLRX
l+DkA7ixDI+Xx+Is1H5+CBgk0aMcB8IpdWWmujQLVy43fH4qunX/lpVll3MSPJvt
m1XroWcaFLexS/KGjyiNymhxLctg8MQcWIa4GieWTvaeUDlXNSaNKbmj0dwCp1eC
Zdim2RO9Upn/XvbgShTeh3DgCKSKi4GgxUfbwgYf8oVjmarpndSA1QhHItuQuKH3
bS6dphLc6BC8eN/Dl49hqrcWs5mPLy/w792J67tNEmeTuzu8GxvSFF4dHRMBQklk
LCreKBakhFNwa7GgA9pXfHTs5GlQOju7rPCG55532Nyp7R5Lqjd1Z1z67KVHRtwY
q7Yt0G9narRBou2iifpA6GTVYTxjlgG2I0hpfRJR6tXxnegTInodC3x9xAMkNBo+
HgeD8QYX7HC+pduEHeUyBllrQG1QPI9udX596gm3Fpdn6WsKnN1GLQTutZbEp3bh
3ds1UXWY+XObHvCY0fBWYqG+9ThZ8dVXzr+zkOtUlWZfwzZ8YJSsyoAeR12ditS0
q20mGhrVmQHt5E104t/Fl+Oeb8VItP1pqckkPkAZKEWKBlD/Z/Qw0cxzlMN8FwmP
Wdfqvbvl4n3lUD1nTjKgNTr5Sge3veUgGzWbwEQYgkMfJ0TXEI9e+MixzbxOYFDe
/tzr44xoirAvvtBmF0m75zILflQ3e10VEyTGW3P5M57ivm6lcfnJ31OMVkur//eG
JHrwMdcWXcmox3V6jHV5Gfe3iyVP/tuMhmTBWHaDiN+QNL9vyqSJoFDt2w/HhbH3
ks/KCe7Eu6Qfg88DrfgnIzsVFFjBsLi2pHysV83QsSzfizdK9OIUVQnxsTYveRfY
2jNjHNVdZJ0O/dlpMQQwrENACmsYnjogosjE2hnuCx4H6cIMetV6ecB6pwBy4h33
N43xIpgQWWDHgnyMtbYbrb8Pqy16bWr5wvwU6+vwc1MyUC8i1H8peV/IQzcWeFNF
o81LGGT9jn1hIcnjALsFuKrHk6AZvEppN57lqEKtqV63KF/0vx4j9Adl27ZiXmjr
Bkc/EzNW+0IIfmA0kA6GFsLPnMc37QuPoCpBLMbw41QYa7XqS6cknUDCt/zHVh6R
U7z3ZRrYPs0XYEy8RvRk9RNEjiDlGRCILIsTLR6OwXORMxt4fyHGiemRv3F+2bL5
E1drv4mflORUD2+f6Q19rOk3CVfuEFCnoln5/lsc9ETvqps8262BHX7R3d/rUyEA
fUsiVphtiXjxdFw+SXyuK00kkymT6oBhE+SRWJ4bxa+rGLMxn8DmHH7c1UbsKti9
7Euai8hRObwnCLoTjCRVqyg4sYFOAvBjFVW5iILN5EN+jdIe/f8MRHkQYeWbWre9
c+VLV9LzVyTHWoiNxG/Z/KnBbGBoFomed1jRqjeS68JNroJHvi+X6M5GsE2i9Rdj
MG7JNzo4cSf+NPHYMa/6giOQ4GAB2502NB/hiPtf6trqy8+Odk+J+NFmnR3SUBbL
SAapW9zZR+KQXXe5+E1xB689X9VhoRkeXjxGKLi26AzgT43h5+q7LIVoaR9nstPZ
SCb3B7Hw6vdJ5JN6wL5JesbolqvmdTj6TWXQMuwmYQWDVEcjzz12p8/9bWPqU89A
x9npUGHYYvx1Jvxmh9i34D+dN9HprLN4EVvQWTkd/Jn5YGVcVO5VsrrfbmWdvsFF
XMblcZEN4iu3eGKZwQQV+2Mh+eR24PHuN3wd3WXgSB7uWWUuw+x1hH8fXH+o3Kox
kqccbTfnxZRwvt55UXT4AhzHgEk/6uNatfPh92bX5AQTKttFR/3cjAAIDXQvl7nY
S7JsfjF9PxqCPtkMVk+oXP+zszK/KLNvNc5cGRrURKyUzYF1Q0HUjAA2snf4201W
YxBLUzj9awefIiRQLg77a7toD/Z8lHYSTk0/3zK0zta8veR1RxCrFSjbvJ+2/Vvh
hojhBt0Rx8YfE0KEKb3XOuGEWe73+6TaWj/QXiDGYHgnGdCNuwFQfqqh85ClRKfz
aawlPEIawLm/kcL3+DbuLicFWBAETauHqej6gLo9rq5qmbJxoKP5xDgESJI4bmAs
ysX7UJeGr51s+5CEXbu+Ns7DeFExYTya7ODpENcSRPxs0+Z22DaGtxNIechA7hYP
rmlvKthV5MO9CjqMTggPzgQYeSq/xRA2giQoirRf/2zmlnN0OGjHNXk/yCe2sSYY
0jmrgz4vtbDQFqLnDYS5mfmQPiUly+NN2VQOdZUW3sI803+twyzr7Tp2d+ZT3+pZ
7Oc5HBZcqH9XNzXVBwwEU1kXr9TDkrEF1IF2k0/n5ijxtYLr1M6d1hE1VVYt9L+p
P+L6PwchdeI8+x/yULq0UMFAO9LMheujSLn73N/Utz8wDcxrS3FKXfj3c2PcGAQS
3lXCoKMAWQkpK0mAzIhd1QE/0dDVV/Qpr8vz0rNQwmF/PULg1llb3tTR6i/BNFqa
NINMxBkDlUJ06TgQeeQKwHfJzKX12CybYowSjDe3my1g3e2BjpzPcKEY0H/s1L4U
AiznL63+NtYuoKsf957RYUfT/W1i3QmGduMNECZFwMEj35s8i0Z0krAtBqwmuX22
yOYkmmLssLj/ccjqu7xZeDzWuQdcZuVrHADuQkHlKjKgs7W7vASQS7E+Nnt+z+qr
Nsz3IK9E4CakWa9TdtGxYO9CgH5C/BzEUYYqT/JKsFgYk0PIXKvZplQ6iaQr8nZi
EuqaFnNcG9CG5pLjNDUH7FaIFHOoQHvJD+WwZTVZZOyL9ENL4noMb3AzL6wrEvzz
fxufYKfAmLq16yuxk7vCZ8BgFd2h0sHOrpWBfGRPP1HUgjI4zMMpIyBDXuIl7qmQ
Yd5L/d0aD7RpWqOieh91N6JPDn3v8seJlG68Tc4gx2uFIBLxBLyhegR5yXnX2y0G
a53/3HEosH2kJcbY5RR5iswwEaG6mo0EeXB+iZCHShMrR9Ut4XrYcuE9PE2eu5HM
26UcsQJ/mXAoyLmJcxCQl02jA6/k9c5aW0EjzqPhxb4hCNM4hg3UqsxbAcz++/U6
p+Gee5V8SnpJgT1PNTyN3B8Dgf4T77h+l4bN/OCLHqPlaB8mzhjQpz6GUCph1jsg
FfPiLmAyGZORceVCjvFn+BvrmFV3pZ0zVXmSAtmhBr+ZRBbg514BcBPxYH0ORySk
XcLXuhEhiTbz0p81+Udu0Kr4oD5aQTRuR/iNH5yqdsj34WDHG5GQVEdGWxbeXZZQ
aEh8yoQkwt/k6TTj8jrZ5OBg0xnJb8O/CJisIBl7HkysIkKQcX1xN1HBsIqmi+g7
lA9OAGnjnffge2YRiFfolDLx8lYfY3uEjjF10mKkjQBAztF+jI2xlkG0BlljyHWO
gG6+hy9Ow91iXqK22+AsCSWnxVZCzBNOAIYBpFFncGqp97YFE+LYaKFRLwPfnLzD
PRjibimtc3PhfaIVS9vj4XFE1bl24yHt0F7X0zj04kCRv8u2hz3N8uICsLiLJ71y
yyDdaKhbzMNBpVFm4un3FZ/pK+1pfPJ0uK+n8aYQ5AIMT6wp00ceBlo0VV1zo7A7
0Pqz4Gb0YgirwM59FdGQPoN5rvB+yzMAG1p13BOImE5pl6OstsgzIKHIfkgCZRa0
Sr44Gg7R+qqRvDDAoh1G2ZO3qFOB11hhgJMovr+0oEAIFlosxnV6BHBpjuTN+lrJ
Z1h5ijHGy84tfkfWldPeNtGcfcPawNJy2GwCNxbwTytzMRyJaf2zidMdsjGzjYcj
FHDfrzmz4z1vnB1W3e90EBZ7zX5ItWxA5HoU2n445oei+BSpb/VfkyiuCvrnebI7
N3yF0wsGXug87TKUaOO411pzVbbA4EBNEFzgbUj897ag1LJvzeV0PdJk32A4BCtc
rgyO0WzJiVDUXWfuDK+SA2FHe5sXkf2QL+LfAnTdMJALRHPgn5SAJCzOCodD+/Tz
NntJ3AqDGTmc6H5LGPW0ZA2gLT52es3nGEV4laZvWYwFRf747w3ll+/TdrFgIQWi
hcZ9YEnWoqvmQv6vQDWpqKVpp4rdPg6HYtB5bEU2gp1T+Gq4uEYnwsLL4h/vJQc1
J1LUOHlgnZrMRM3qi/srIWLhEbvsrz8E0/ljn5EtbO/rpCqE4YOG0wu02aRmLMeI
f5plakvIP0TwPqAjFCaBD3RpRpbloujpFMILBacdb3lGXj+HOnWZxZinfdY/letz
Jpj4FHEfHxJP7PCEX/YY8X864PPkOh23YS2YnU4R/N/Q281Nrwsic8EDPPinZPCp
rVAIYvHxVoL2dnUhR182YEo9E3/jbMAvRUHc2rbeD4Jm2VZNNO8VDAjxQaQDX/w1
7VsH0oC/C93uytlCYeNRdmFOtwBRzIOav+70zk7buMzANK/8TAEEu0PqoZKnONDv
oy0WiPzj+j2ZD0xTfH8M+Vwcrh4FSe/f+R+fIEapG/wGnsiG0Di2Ucz5COHIXpc0
QaMBn6i4EZ5e4VS3ANKWTGcw3wl2bNyRD3XQNYwA7lz/hrUsYekbDkzCfXzuQ4BN
iVqroKt0akwyoWyibUpopO6M2cPacBaSxIimk3tNZUf/lrVQq+FactBfbOIeXZjQ
qRFn9ZV0fEBQoVu7Rx6wUspS42hGDS/8ZZNeOXVbr0OPE3uzXPLEuPQarvXfSFXA
d1XOLoCS9E9rYVEL2eYoBLkCMIINSXmkwM2Csz3Fz5NLoLEpI1E9om3aOLdYHG5j
wyaP5ZM0v6MH5LeQ1br/tVaNpzwmSjpwSVbliDs2Sba+wvH1IF89aRjZnrKjxOOm
lw02dX+hmh83CpJ9f2Qu2ReNHlmqYOcE4N4sT9rI9FuxW9N50bbeAPKtjOVyjAkm
`pragma protect end_protected

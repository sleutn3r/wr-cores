// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
PJSX6HkHWxFfxS5G8NpmArq1ET1NRWCeIQhxtS020cIK40KYIdmNiB+DufUV+FJq
MCUpptRfi/0W/VVYV/PPIiM75yT9BYYvtoJdG5cM1Vig+tKCb+hvBu326Snjor7U
XW+pqu3NjAjgHiDHgYfhp9RwSibaX4BaTraNnI/N17Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8272)
Y5gzeKI8YLlIC1n4zCi6LAEAGnPvxzRZv8kYwiEFoLl/UCGnX7z+wWCb73QP+me9
k8FCk2ZYHziLRLeBDbxlJlQzCsoTiy3T4kGG2GJrvzDarMx8c6UrQ/bsUM2pSNAf
v1NpITJ2W9bh+KZ4bDhDlPbhJpAna+rNSb2MnRE7440peUiEdO0ynaOfIm2eJ/ey
LWeTOmr8bhIYqZ+34wKuoRFqdgv6oD0ju1N/pxtJF7+ttd4qFs6/DJYv+5jqxHyv
n0zWJi5DGB8y2h4VTrqRhvrhf/3ExvY74PWcMf44MWrtYj0TZqb53w0UPm4cKhiF
zCP+Z9keRS/6RH75+VOiKKCt3aAABPge7UiKLtOp1o3+aysol1GgATylpO7hkX7X
bT15n8ODSMwNB6AY5llP62j+sX/KI24BsjGUYuVpyhP2azLJcJIstzHoYVWZTTvZ
wEgiR0T1EkJHWsSu0hCn1UiKAzMbHSvktQRrWMpPqypMHt9UNN0txaGzd+/zwFua
/68XojY8eXZ7JUh68yHJbJlobefbfIJy0Cz0NFcyO6IZ5vJ9NJ5CydmPMogViPYL
QmvEUGqbMyuIcPGVDX3sHItH4ua1vA3m70I00BaccElwEg8rQ/OZw72mSYl6d4Dj
JFj3evSns7sBhK1t2NAoP2pS5FC+BLktc3F3dNzzHwK0FmSeoM/KFfaMDKLV1uhE
fqoyRoKVuD8FOCRtm+5S0iviebCbsnjEcAr7QMJzgkRFwX5Sx5l2sfan22a2+i4U
Ix88VZoaI4RJATtxgXlrsUOsfVVsAo3RfKsUlitg0rcA9CWe9wykotJFC/Sbl6T3
hWMhq7zSLBeRMpf9Bgh9hoRqGz6A4WlCWVT4IQIi0Ae0KeCSlAA6xJh5Mb3aSUsl
Gu/iF0yvjLWBvxMV1JkCvZR1kry0alhYFfwyNPGjruNaHCUM1C9ukFJAak+NppD8
cFtwFD83KopQApo8AuxjiJ8ffsEvp56fQj7L0gqRZqh2HrcH3NnfBN3K49weV/EW
Xi1YCEsKejE1QUuYMNky4yMTF6gGoFQtZJ0KYqvruvNtosAVqIC5+x4cO/jEM78V
mL5GkTDoqi0T0BnzFpJt2Rv/UTNGNx5AEp2XlGTIG2/xXa/8a9gSMhjWfGKlDQg8
jz7CJKRxcNmZPWRnzFDJ7GpEgbogNEitooKtrBHBFZBGINFYDV01c7gFegMqjX1i
W212OM1KqnPACw0yvhvMpjUd6FMC7m5spHpIQv471iHOc1NzjSeDMoFtDVPDUuQT
HaL18HvzQlw6QKwBsKEZrnlMq5sWF4Ha1zbaI+GK2D69chElkEAn1E8IjP1oRKvm
JVMaHG6GpYia7mzRjzbNk5epZEffsvjBdqsuAfehb51Kk6T3gzkB1yiqFCpD7roe
q8W9fpH2XOrbbK319CKM2dvhqYnwpz+9mavA1xhlB6lPZyulC6CDP/dwToWOChqX
x9g+SxsF6EOcG57e6fNvqhcedukZkcowRGZ0TpRbi/eEeCVh8z437O3YGliM91SO
WsC95EjxMbLa6GKQocY8tAmVogYWXOJmw4D4lb1/cMH6NifkynxV4AowcBZTX26a
q9RAlfT65P5bHnc5X/4q6tUS18KDn1G6nMgLT9oN7yk1os3ZpA0uKcDD14T2URpw
sh7pFaO1i+VTysi6YQZtkj7M7IGGEBJ3p2hUB9AsLakMYXvAceCUEg9+wDbscw90
VSlTAncQy7QlukddOtUnLfiD3rJ24P/7ND0b8rSdhGBS+JYlc+M5wEU67UO/joCu
oyJJegKtjqkOEzwLFLjpO1tirCEbl2a17Bp7lmL7gMLXqzhQqhamib9TMNTiEplX
6eoHHsZoT16CLaHib3/mdFvq4+IlVJGR48VMRBfVWSyav+QjYas3u7v778BcqZe4
yqzVS6RrIw7JBiVF+sWulHJN9nnuzSI1/NPq1tr5IQZc2bWzDbG1820opJbn3yhs
r80nAV5pBpGa9/3EWZ+drtn2hohIXsYzFay//zHASjMcb4f2UrF4QMJubszlyGaS
oCOhFR536tIHQqFvjqqus0UKOr7lhzpl1LAMJcx7h+jZxYpebuRH17tgxsLvEVcJ
WCbA/quSI5nd215GzezM5XiMKVnvQUsyTAuSv63K8BnP0hECrhbIU5RZSn/ivMNN
7S1np+H0mueNvv7YiluKswDPawtZFOG8HxVvo/LrtkFvl7dzV3PRPYF1Rb9bwhak
IBK4GpXkIxFVj33Es/a9ckLF0VpS7+XRkd4lWGnYqMV0I5hTgyArc/zsVUCJ83AG
8BcjjOB2gnb963eg5o7a1zg6j8VzDbRPm0C5KJfgfedmTV3ADFxnLWUMDDX2ivHB
O7rQQ1sIx54q/ulk5TMGmDfvQ77o8hNqZ+kyely1mop53TtqX0q5leI0Ve6/3rto
jNStg3KK5gJhjgw04FylKRKxehklNBTRBJfgoU5PtuWgE3pI45NyCPZFRtDDkONQ
p8LKROxHlzSCBuVILyVa8+rJhzkX4UelZCHZsHVZqrzeD8C2bf+85nNcHmzCAUbu
TmN93eDKkKAIEID3Gh1Kat0ghdlQDdGc1x3rWR4kiL4u78eFHR6xe8wg70Jm5NnQ
kwk6DI6mfpRG4I2X/0agsOicE+8GI302i9IYeeJiaK49oausNVXEMX9sqm+dh/Yt
l1u9UIQttO0jh+1JWdrofF1bL3vXES3YUrYJisTChS7HMGLIBKLgksdu8oOfTmdL
dFW07NuP26Yci0gZoZ/4O4LOuuVDK8WzNh71tVnA160wNeqpOGCaORDFx0t6sJad
W9oNYZkoPCrRD6DTHVMRZly2VttrWn09L6WOjg8g/JEsvmGd0FqPmV0pDW7b88BX
rL23cvk287L5iFRMP8BXmZTDfBpbap9XfMQXsG7ZZq3f942GJToUI6Fcg7DctHNR
0EqLv+qX5wMKHBNCmETCBHKmoksQA+3t5VQekuK67pMIfcxqUS0IqUXriAM4K0z8
S0Qwq4RRidLoj+w9DwMNV91AMG26Tlz4cuo+LUse3t2AkVHc/rKC+c56ISTIhBJ7
UFuGwV7skKRGtJb1NK+zNuF9qrz65xhTEJhGLtdJO8SwVQTFhBYov0dhGiCqrvWm
l1aplOwBjxBbWpU5oNIWSvmbeloKL2GMJLtYPtNcEslGEzKNgq5axWWFCfhESJka
bpoAKy+alz3Oharh0iDCFs86uW035u60gbUgMkaq5B63Tp5YxhRZBqIar2EGda9p
QJln+3RPEKP3sePGjZK9C899Sd0tJMMYMOXXiefpmUk4IhuvkAuozaTxHGM5opOH
IXNwIVmFo0kelVizUxozzkgXx/Dt6ZnI/tNvkzzWhmYPWa0oJLVR5iqUFxzK8HCC
qedFznGENrm1F/jheS3nXoyP4lijRUzG7LyB7khkQxjVRFzh2E0G1d4g8xgzLF0f
mYAjWzdPkh5xp9KO4kurokEglJ4jNYAmTqaCyrkiTPxKZxFtUu9AmRyQcjrmVbVr
oh7Ip2a0g2MNOXsigYOgQJDB2YGomUeJDpycOxGg3Zqe4SPEEGZHsldIA+hm0W1u
ydbdluapqGhWD7NdnUZ5inzdwslnkpkqPm6YqtGg/XbhsBJfGvAXjQftbcP6jHje
rSbUZIC85FdJgNRvgT5lO978FQjXQniGrZAPGQXhliGD7GmQgZgqr/wjutvEUCvt
IlvvvjcPbeGTpyYACi56oRs3Cc9JEN9wMV98cNybhASPQHcTIT7rzrFMmtzLfiad
JtGCjlRwmbNTEmZEUeBExUdN4EPkm9YhDiYNJNhbpaFeU/WGRu2NWy1EoxjZlOA1
BVfkwWKT0f7VTlbgJEzzbxfQMymzqQUVZUeA5lExb+9lFWBAuRVjC5FUCgtCFKlE
J/WiVgf46xH3cjyNuvtcgy1/CrNk1Fe/TFF//Iqb8qpDZvNpIPTTFrkyl/2dxB6u
pG1+7PL5+CI9Y16ul9Vh+OegT7+OqFD6x3cSrZ2w+PE+Arc6Ium/j4WEdvxR0w4J
eNo7FburK0NoA93NAPrfmD/uXfxk3M636IBnpbyoIOdIFuj9RPa7GUYg2fCa7eun
zUmTgCt77OZQ9W1KOQxQbaqoJl382FZyU6tvznudwuRxyNJSRUInfmy8arBecC6K
X8H2foSatE4/3JIJLuJlYc+NW418WGcCRsfi8EojlwVhE+6uTP0B6/J4I06DMVS9
zbc6ykaKC+Yh6N/AHVul6sgo+V2DCA+pEWFCmd6ckaiyW6GVW2blzXTg6t1eOqF9
r+QWbfufXLvrOeJmk9nYclanHHMGKwpzf8aziHuvKeMq6BMnWfuh9NiSi9BirWJU
HskwvWY/gp1cuyCmBJklgTlqLKa26L8OvsEcWvjoKbtCFgQeHkmGoGC7ia1CSK65
mEHyFRy29HM+IuJIdty2AjdDA6FZPYIfK0NNosoZ0eEU1hqB7i/GuFVAoX0JBo3Q
khH03Vdm0PCwF8AYMirEpNtaXaI+Z2OuTjiMGRsqTrIR6YrFwiW2H/KPM6oSCnIz
lYSASrw9nV2wJQfHYQ0aO60cjNnVzPkg+6LEtGlMSn732J3+mODxmaLK6sbnuZb7
00HmTpTuSNiacAeL1uwQGzRcx9buW/3LhFXL3K7NEE14yLmROTu4IJC+npXMM9gR
uhEr1RHn+eADFsUP8GPzJdcNKpmK1L87rv11Um5OAjNRR099bZPzT6twKzoMA16H
55cEwXlz3DEejABFqPuCXesnyWLC7xPaHJ60M7MUf71nwpqxCONnkts3tgwZJNrQ
PPS2mWBQ4OhCYfR6oCLY45w107gB20o1q9pToHJLhh7dwMpiqzTUQY3fkMmf0Pwo
3lu2ZJ4agadmfRTRk397ZAq9TEa+zmxxdGSjGfNCwx07r3YPQxH/pZYze2JBYp4v
GCHdN/v3pVXIwKIbULhDev9MCbxB9c3pX9w5m+nphJcYv+SAnZVEimlhs9oQMuft
Yq9pCjd5C6GkyS3nOPj5cujVlnxYkEWsjUePiq9/63dSrjhsC7fkiCOQ4eSHhw3n
osK0llC859UORYnk1YZVO5Dx+/Ymq9Q2VfrvHFbApMEAq8TC/LhBp0yPYZ8Z8rmU
rPq6RXvACXHPzqcZKyAB5nPZTfmjcjXZRjNoJ35yqB06dlFEZe5yE9uEKNdcvhRp
N50jI0N027X4UM1LbcouQEKMMuzh63xiR4d6ZLSzFpeX2kVpZo4KdRnEIrDuaVph
PmgLnRdL0M4nvnvsawfYvp7EHMbTNAaZd2hmU+VB2eChlJQTegUZIqQn99vH3VJ3
Jw8WZCWK7+5jzTaEA1bAI2XOLtDynDl7NkgJk+oXnoVM4xEc6gFWqIFloVZh+2on
nEYvrkbPs2hjYKYDFqDLtGUe9F58O9AMX+eCSMsjljKc+fhJMaZGYQeofghD9gSh
1vqLglaX/1Rh6fR9qnfRx0Mi3ET+ISWVmPhkDbfES3FtAnK/vfSXopE5xVm66PVH
QHm/Rorafq/sm38tgYpw/FYTtBfrv7ptJW/slEgAAqvfNT4C4o1P8skLLjc4HhS2
4Q3VhSbHSIgPWFzkLIJYTfTw+FDR70NADwxgltyuzUYSjIrJUCnv+HDABr4NRgX6
hlSkqsT6usUdqEcCAmqhC/jFFADWzE3LX43jjOR9iEUnqja6j7gvoDzMgaTt28Av
BrH+PqK9849EkqROUDf8vkrBFIvhZWzJ9JVcx2hIsTT82gFf2ASM2/+BH0DfJNsK
bpCHIu8eACWAWIUcGtWAvbPOsyefbDnvZc/7z1szJCSiXWDrL5SYU7m8dWoZ586L
fAbPJBrkIGx31KwLshEHyVNt9BmxFLaP3ye7Sk0w07f0wr18WpLVf+PVD/VMHfl3
N0CAk+QBqCEcslRsRkhjNRIF42XQqUA0tmVp2cGJSq+tPQM0Tvr9A2/p+hMqMF9O
9OaBiqaw4R2nbNIZJujDV+lfJPcBhv5WMq/CC8ttVEiQzyVaV0UGBn87UADGNo9i
d7tGKOmJXYgFTOJq+qexyzxx1vZm5Lp1IEDZBx1U+keA/K8q/mgyifzv3UfXZxlU
PsCLbg2AZKyqLizGGQJ8WAy1LoW7qpJoDm6iRi87XgfOiiiVWICj9lhqabKNENu/
cju6NrPmp+GfwLRB9/5O59Kei7t3mhfAZC8hrJ6xrgx/Rlh4iBQ9YNcw+pPuWRkl
XZy1QSht4OAAYk4kyw83kSffWIlI12Jgjan+L/6YGzr4azi6sCeN/RO2kmWx8vRn
NgNMYuq0a52mB2kvIMKlr/sTwqAt94uD0BeLVyU+Qx1ZZz9pT9scP9g+MvtntYnq
NfW9CLCFqb3a2UmGpHQAEK8DPRBYTiXSoQq+AGUCLVzI2GTUdGLTXpCB/yHx0RrI
07fc97ctWC2/EwrQLTt9xrVXDlHiPqxYPgZN19YxxZXA8BhWGqdG+fmdlUElV9fp
A389OKl2S8EIlFIsydZzGDvenwXaT+nKSNet3Hc5jALsFY+bHDY1im7G44Qd9o0j
pxzTwggoYmvAw3bNyk0ynOUGpkt+MtP4i4FkP73X4jiCvLlNEPwQe8VD/5j8Z+1s
xVM7psoELD8Msd09P2n6YuDVEWBMdGkCu6noh/yj2uMXnL5xBmCqesGEX8dglgW+
oVB3jpAmDDzvOIVy3SW6jW2QxzVJxBwBRVtRlz6TXkZjXVdUaYlfW4Kq3H9NEtEH
VnBGq7G6nX9krcKfHlfWhC3WR4Xw0yakT8a+uMni5PAsNJ165H8b2yFBPhr11MOq
XeR/5C+JM3yWedoj1juCVQuivSGxs4CTkcKskPW07plKpXKZM/eWYpFLg+iqwjEB
1uruoIkgthjkqDbkK5Fe9BeUyxpZ9CeUXSxCR5mCp42fVT0IAwK4gxZfbZqmUjJJ
Um4RUuR7k6l3P8uyXlWTLM42fHfvPFRqqvPpWJBqyq8UHsJOurrqBej5wrMDbvaN
8u1XXNdms++GD2yc6Ic0oVkAGDUNlRLKscUn8+QLHAvgzbLgTNfP9wEyI2cqMGR3
bJov3PiFQaBXEr7pk4oBc/qucJnYrEGNq6RfLULmTZCNEZywAIYzn6TdD3fUvgrv
9b1OTPwoifTR8pdY9cqT89yv/1xVgnlipfjQhPlKUNkzg/09fgNct5U8OdGTGNf1
yHZdR9vUclvTZPkAPXVX63sO6Z7u6+5vWkugbW2e0iM9hwqhJKpZG/ytnkP+5XM6
p2P9BCoO2/SzpxEN8tQ8wbFT4nHO2ex3niqk/414ij5MG+UtgECSCpmMdxVoiejS
InaCuZQpcB1RrALVuQpH2AQ+DZdKd/UPIe+FM/MUplWZjDkxtXWr/CaUGJd2NmNJ
/d1frD7XrDSSW8Jakq3IXiDIcL0APa5XfZQY0l8jHtasFZsWHQw4p7+cKtTmF9p6
L6kEeAg5JGq3rft4OzC/JaVD42Yw3hkbiJUuYzTYTOqV5HNWuNp6+9V9zKWaIQky
fl7kqNg0YiF56/jKrRcWj2g15kRjUtVYtkY7vcWD/hXETYBkmtAxTYgKq7qEhdsZ
4ZtqtjvRdj2JdurtB3667F9leTism8gaEi9v7EpT7tHzTX+Xe05xun+Hb0G/e5ST
JkPhe3c+WvJ1lCR7U8gQSIYVHSTmtB+xID59BVIHxvfFT+H4vfIhz+Vsuw/mTELP
fGWWAbRRJ0Sme2RHihuYPn2lmrLhjX+XBLe090pVEmbI18T4ZpOp2zAnHA9sXu9w
B+U0hfw0XI20RJHMM7eXOMFXSrhHf7Q3JU91FWfvBZUap/a34nX7O5pm3TTPqeRt
cP31CJ5xGLjvMaS26Zdy7pOGB9hKL9Jj4OM+79YZCo7BmPUXlBTwHyFAkaBDxTnv
B3Bb8+yUA9QFlJZNigkOIKYnN4jR/LBlGAGlW9+Ao5sKM0tIwcVIQsI85fMrzOxK
VpvuDcN5LiIYQmpUwqpffj8wTtXuN6lWXD5sn3B/3kBFuEem6j+4ITjbdUokUrEx
+zGjatojGp1kx7Uqa33vVEkk14MGE2YLOVSAPxrxeACB2PTglsNjPJRdmuXmWcUO
4sYjfzVqk9c0o2q3/v653dyJ5RE+juMnDZkSNzzDAjWxB+khMTEd14R6QlJk/1aI
A7qFLAqT0E6cdzqD2tC7Wu80jXMSu8XmiTWcZEaJ2DoBXTy+Dm/LyCuuDtMNpDTK
mV7OQrHZPLvQMxEGly5RlGxgMQeyTlU6T9DfK+eSa503rRPFqN1i++h2qvbMHqW/
qaC79hLm09V7TpHHab4amrqqFzZIEOFdOhli9Ft3EK36voEe8LPZI57EHmv8rqN5
tHb/rLWAE69iKgF7gIhetCci6ubrULdXvlNP5iqK1XRRrb1z5Z9h3XJzIIlJz25Z
R1lB+ns/V7WzvsXvztSfe6L74Izp+A1qDHm5IlRpv/vutFlr1QKT5l+qWcT2+SDW
LOR7OMM0cLwLgKRF9uu2pLmeZ4sUpUt3gxkVsLCP854+VFFVsBKwxXFz/8UnQ1yk
D4vbK4PxY3tQeH1s40Ket78qU+d+Nh3TEvnW0t66ACAz8DLoenbtu0REE+WPGGIq
rZ48nAXVB5AazK2QQzWaUOelZefipJz9c64PCL5V2rWl66XTYtzVk0vq79ByrEVv
lAVcPMEThc27VD/z36u+PsbipPL+QMxF5fiucBeorcIbVYb3eyMTM3y5oLO/0kiQ
6tFrice59sK0/ji8B5W8kETIbvm7SNUBSpZRIN8Kt3t0lNOSXeIOPduX8EMcxGRR
p/r5ifP7UOHGd6KGszJamX3I+JjM8RFd49HcmlwitWPMma8890NHS4B6oiAMSh0L
kkwWOumIwOK9awvZt1xu3OlEU/+E9a+YOG3pOEwNt+faz2MDfMb+0jM6wfoa7nd8
8q1JF8KoV62vjlEyt9zXVAh8ziNjdKGKTOnsrffu4hcdoAzKNQl26dcf0Dp2ghHs
ZbSxJ8G9LSMFDlXDzlDbOg1LpWhIfemG/IVCUsOSXepgXFIsz8QFd8IAGovFQ4dX
ZBrMLUPdW082f7Hn+dcZa10u6tH1hvslI0PB8XjIMEQpkqiZOaCFQngc9kwsYrRq
S3oqIAmmlbORr5s9a1qa1oKtYYB/+GgJhYcSID0/QsB6nhtmLK6yywdR8otiFfc9
OWTqtl1jzZY5u5rUIApt6CNTa7+xqncQ/vXhatG0bsfC9F39aKJdb6ee6kje5j6c
DYTEgIEpudlxcrh5SmaSIFP5IVlG1DLHw6ouhy+EvUVO126f2ih/TtmfeqPgLkqS
jJmnDNFdXtpcFjzOrYUNhZmDdlcBg0Zqu1AN05GxPSrO1+FxArw/WFu7RJMuNcnu
WluBrIIQCtL2ue06tJ3KANlT4thZ8GiJ69ZYMlOejlmXmMQyKH/boa0kBmYSrAI5
eSWwadmkkqHguSiwQXptEeP6gk2APL40nYiYydbE0hk9Q6OkY3fe8QB8d6UXKhTR
LlUIbIpVlnp/fqMYx9FNZOXl4Kc6p9qX7xE5wGSdcNH1Pq54sRu4pbmbyPS+wHsJ
qhpDiTw8O0IjYl3Qc98KfbajwblPOBYweO7Epcf1nYYJy/2idg4VwwAdCZynhLAd
VcIm8aucQZYM5gBAskBh9vM2nIprYw7Wo4kLwTvKnDzF5i3Nn9wVKjUXwRWQbCp9
SfYuq0ONxxfyst30Nc3D3GpYqTJXqoqfg9qCAFDXr2UL+v+v9LEyf2f+Vjp+WfrY
ztfPOjTBm8areNLTxalygJsJXr7w0bKCklV+30cQCJHkDxdYZEkTwr1574/mC7bt
wI9YW7aogKOFfXBlp4/A/fmSVLCqTc/l5piD3SJ9nRJDV3glMeJdGQK742np6TDq
HyCcSoQ1LMP0KeBOM5zAZqGI+NnIqCVk4K9MSOUUe8YPTJj9Zo8BMoHl5eZ/ixE2
Y9YSE5gm496u32X0KPYxVnUQzCljqO1FawL1cj7eLIvn1VciYC0KqwxlEldUfXOz
HEx9C/ZsLoOfcQdbudOknmt0ARGzDB7xLVXDfkWAmfQfILg0XAMZfAMGdiZgoQ9V
bJQa6+/h+8eqIPpUXyey82bKLLgppfgvELvyJMfj4cufoxf15Iw+LiSjvcASrX/Z
a+VMnUNTbo1GWRJr63avloA0gdrATr3H6SydhT51sOM9EaAof84UtO2QiTpfw6wO
t9R3dO0fQrQnPoy129xEzL385jPM/Xcc/P73PjAo6Q3UX8KxSeus48QLfsXilCz/
DD1v0pRA1v5iCUEjtr/rRCp67h5rCDZs8r3w58tid3jSmC3OWisEVXzYslmhw9TT
j9arvE1O6jJR3lpPO4I1u3e4ZpnW1mfd/UBCxzepIpHoYAxoGZIWBtOcauLnS94U
n2Rr0nQKZ3QXSRS1Pb2XMGL8pD4/wbaajrqCyFfxXvp8UXp5w1qJzFLjXrGdMa3P
nVuoicV8Umw/hopYWiEOp+LaSISzqPIYpAHL02I/1QA20bEk+mOhCgNTm9UegfWr
UnCUTan5z56e2mrGHQShJL73SheRqFQzS0TmKnoqh4nCFj2KC6Amf/MJh4z2LB81
qab+xMt+XvNMG2TX6whb0fuAeB/LjTbmwbaURPS5JpKQ/LOwYASfBfU8uQbRkX/c
9B/+EmDNhcbR74z6uHgAcB+hJaybHTJyXLKErdu9R3A2jmwEtjvAaNJE6TZC8SeE
5FgrHYjLrKu+kG2eYGmTN9uDBIWzq/WlqUyN/X+vCyziZ6fYdpDKVCv3E2SpcX1H
0Fi7/lpkqgm7KjkWpU3ATGLmAnLThNmZFFZ5HamA3whe6Ir1FJGGCzlkW86xIYPC
vSo+WgfYeo/YIbZWMpRyQ2E2rb7JBPmUm78pkSeZEBjwGBCTzDzPl2ZRqeSu05Z7
n4OfszRG134c2tCoQBJXSqgeKpvyIgcb/E6IsuVZ6kr0XsRU93oc9u7yxle3bjaN
uS3n2E1F8FLVrbRpw435Kd9THDoOLpcgLuXs4UAA6VsfV/V06yoXSvWuzu8qJaVN
bgKWwD50qqlg4oG7Z1UDtQ==
`pragma protect end_protected

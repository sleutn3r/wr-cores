// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q0Eo232eAvg73RUTAJbfDREMzqLzgU5TcO5eoCESfDjZKNLMh7Az3tdeuA4+0eJd
BV5AILKziXyMAMRm3L9cVeUFgyDEZ6eGhkU73B7C62NjQoGvl5SrH/RM1Qa/Xub5
1kyT6kdceknHHaQmQMROPwGHPtZ7xJKSGGBXwT9KMTg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10720)
0Of4pQc4xyEBZQJe+lCfyTxFfH7TtgkRYLUTnKAzvOKUC7+YPQfnH5g03JuM9bd/
QAgrju7JH6gZCTUXLeHq0MHhR4pWDnzRW36MzYGs3dR2PFMPurXvcKVF4jfrNN+c
h2I/MfuUlZvUGpDYbQxEOtqTH/KUoKDogE4+P6pZEP+7NoujSQrOfvchqRaG2yPw
ZF3WMS7WCm0IjLq4uKkVmz7FQcqSDkdSGA2HLgMMDxw7pLPDms2Rq5QA1t9jGfN3
sdD5r2Jt49CMt3sy4zEsIV/fPYCatDzPv3XO1mbs770vtC4bvYbMGErM6IXpEPNX
/p0EnKM7jExsYBrFS4/RBDTz705qhK3klDdoaPVCrGoIjQlPc+RyeC148d88Uj/E
lSum3l0kKUajJuHdNA9Xr+knXTZDlMQUqZ9ivQTwUmsOxqqntgpEUv9lu4deRkmC
3qU+dtvjSBFraL4OVGzmo2E8dkTBcbnd6o9VojMZti5As1N2beXz8rTcLk5M/Xig
9725Xbw5MdDbex9scM7V0fdCs13sioHBcExQ1i3KSo0ewRphOeBOQq/jCgKzxUUa
Mq3Tm2XFAV/SzEU1PkGY1IlmkndxwUIe3/wEaVpIcecg3DsYUaMrXot7RWRlqBhC
KlpvsU56MWkMeu3LaJxkNZFYY8kEmMZQvrFgF3iAbwP80wOA2728y0+G6SlY14gD
Y+g2YVLDw//fkTpCm6BMBo/FQ9hNwxW4u5gJqB77yeE2voOjCx+GlWdeT1UzDNtY
m9q1HARtfNcNaqIA2+pYV42cFuR0ZRIjdYyLf6XrA1g1atWcq0uIVDSm/i21Mgog
Friuaibr6oLtmtkK8iOTrKAQejFSnz5PJwcG5InVrcExzX8Ozdo3vlxEua8YQSq1
0l0p7qVJDbj/mmIxBC05RfvMRmtHkG+vPuuHPVnWHHkKxiT0kYaMGEkWmkm9nEKY
fkmoN0crMfhktp3T8h7jcO18dI42vU0opZ8Zu90TtohXQkCtn5v23ohgv7ykX04g
QIHWSTvi8x9rqeyPT9Ggh4Ja0k9pY5PLdTg6/4O1jd9/CORJAqJTGAgeRrddWTen
aodA7LbJYg5BB4N4Y/IY0/TCrZ42pRApemi1xZkyxxAGvv383bhPrvMG28ZusIac
smJl/i7NtW0RfREvq6ms81eoHjBJTTcTJ7xZ8uqGBUB37RbH8NXWxfWn6QFmkdNR
L7YIxKXzVWbcSZxyhG6l5OexLNwDmqDcpFO6OM0lmdp+KEqZlBCmxuaayJNN46cJ
HTP5WzGQj+AJC/30P/gOgQm91NVi4ID8iqjigT+EUpK5rnp0TtyVJ+OQBSk/iaZj
ThEIHuBo2roqEAx6KJ9WUEPDtDccS48u5edhK/yexq5370t8YrK5JZj6/hUJMTop
d7YgCRKo1TchPVMiY79fd3p5q3kAGv7DdmjbtXFyQsDa9BM2Ge9ya7A7dB0uTLfa
2SMsY0hERki9bGI1s7dF5ftwlJ92JbJKAbX6e/bLIY3Apc4HY4qxRo0Se5kZ7xD3
u1y7tH9+X7LV9ixYLvvqChOEhHocuuWC8Y9jwm0r4UEADkD4VMfVTUflaVdCWccY
oGHnfZOyJsMCeMCZB6oqSZp+IwNx60H6H8zdveX9+CnuNChQNadqpRUYgL+/1k3D
zGHdlGFnyyV+KKFXVh4fU0vV0vm6sEo6KWxRIR4SMKnBIoLUFMhCKc5nN+gLLhRk
7Gw2GExcBrMxnrvP87GbsWTYGuSqBbMYRTtT7X35PLsfU4vO/Mywqou4DSHAWD1d
3wJyC/pDKRb99ZEoGGpn/3x8Mm/FMRVosjnpiVRH5wsAX39l5v0+QQw1zbuZ/IaO
4deg1UmclbF67E26/spGkkO/+a09GZsMK08fpfmj8ZNglTMYKZxdSSfB9hbmp7St
0Ymn1TID7tFiqwtcu2BOjDW9Cd6XasRpdoOib5ZJED1w6FHxsPPxlqs3uHuK80+W
wWKpfvAur3KUCF5rUG5V7/MIeSeBn6krvXfpF0xdrSvovm0wqHzoZ8CgJLuG12jA
rO54IzRV/wA8r3hUFYZ27VHLuRDDTSLDkUjzIrMDwhurM4noo0WbiN/0xzFLe2QU
Mp5pAMSIfHBKMDalk7mOHNrum2SQ5OCZb0IDFjD918VJ3di/KXgPL/o3PCPs3yfw
x2t062EmHggZDclKER2iEgHS7sfTcq3IOFIMolkrI6zrxe5pLm7dn06WqMyIPn2u
F6f9lEm///0EQghxAR/mlCJvO9aesctWTkdwSgnjpmKX3OjrVcG/k3yevbW4J8BE
v1cchgv8AuWxGgxe5OLZo7B9eXDvXGDn5QTuOjOaUcFX+UhTYjSQ5RN4QbrB2N0x
TkN0t8Ip/yC6D9wK5kPtHSMlIxa8GB2XX/qz4sCvtx91a3LQx6dBeHHMZwWUgajT
l0buDbU/XPLsEyfTgS9t9940rdvlIUpNM8UErTtJwvxfVa5DMtpoHHofWsYn9GHW
pGHNdu99AQTGmrfYEPPVD9nuIRFbcsFl4JGYj6RO8JpZVGnGup0pIDeM8Xb/lonK
OX3+FCGyXEIb5FPAy8vEG4DHkjQL39jQD8JlyWlHEBxqPeTWouwcTO8qSfqfjR68
EnOEjlQEkfjTjDhHuz2aUFZ19EXzrLAN5wi0DcfOvicv/JkmFDjk69Z4YFBFkgB3
5MAwsEJFhAg9iWhabrhvmdewpAVB4kLOawZCFIvo0HRM+7j8autU7+2XN9dFZXPd
zuwl95SUIg8BO6doKtpf/56DEviAWsXNmGcab9WbvFj0p3n8PmlbWym0HgnQYO0H
yMQ7Q/qLuwiBLxB8CTU3tGTgfF0lZtkg13gkQ5FdRk16TLYF2eCO+ZwGJztfF0Np
7CHKUUrUyZ5vGj6MgZlnrGX1k1dmyDmzOiaIU/RHZsIH1WJ6ILcjWo5uOq8Y7eVh
Xjle1DRY44vWy2yNl2KGdv8038JRtWV1fH0xUh/3FCLU3dMXLFp5+TroojQAtpL9
D4UASSW0F0aUnh+8w8MmdBh8t4qNU+CqSkIPOvmHDPMtXwmScBOd06Ds7MwBt8zr
cpuJD8AUOEq5ZPsGbTkx8SjCerLUODhNXOimMCmaXTGeRALDNnPdhCQ0K0xCiHIA
qa5fQeLeKDDsF1kDzZ2xmM4rESLtHOH84EIW015gvLaVMl0YMfiB/ta5GxoT/JsP
0JmfAZqnclnYIBZen92DiERYbnTcvwWQVkyjFPt7ALPsuiUitxskLuPc9o8TQnCZ
Rg1WnbAjiQLcZvNZoM/NMara1KZin9ei5BmDEK/J6cyfuZstTeznsDxbSR1+QYWD
d6rLhgTAz0Cd/p8nAX4qjleVaRDFQ3FFSjt/p6J3LZ6bBgUWXGsHGix/pdlS32kW
DLxtRmlJORE/ItCrdkmIW9LEHQ6shWBx+heI+K76C2El4tpcCUcVet7ZP2ci3Ube
QCJvBKa890fM6O7ERvNN4cFGACVNx8EnCApWeC9jD6SS3V8FQrzk4B8QvAJJUuTU
KBnFhptDBsnxtKGx2sgDCBZAKDnjIta5k2hdqhh2vnJ6MXQ64XLOXYg12T1R9vSU
1dnERqHBvBFTHmqxSB/JWv1seUTfyIvDUj5tRDNbFL3nD1OKZe+1+AXevxjQv4qz
2wHK4edwqgZgjBVbnoOLH7e3lEFh6yf8EUoVDRG/Pd73wECyHzI46dllt5kvU7o7
bN3DkCmozrrhWXJIGISJoPlKWbuckqwK8PrNzWnZzdz4VIjs/dhCDcgGSp7xZs5a
bQnjU0WSrMyoJ9tK84+EouWhnnHQ87HEjkgCEu7s3YAAf4nXc5+N4u+B5+dlf/+R
wqHaf147vhQRrO6dYo8l9wc7geuhgQOrul35ZJdWx2R1mhFrHYf9ePI26PtS1CVM
CQq97jxYgd8oLbZChlaowBaDpQBfQgFPBGO2v76dnf/ricAZGSUK3N7P2kNFwXCI
oGe1UqMdncMPW/y9zHKHp8DBxDuYMlCV/YKYsUZMdSAMn2Ew3xTIzB67boGbkEQ3
Bsq1ZIdNfrNScjvwywgDZc45jDMllZz44gpJlMaHwxS9B1sV0IJ+AjtO6RHubkkC
AcpD8fy8XvIcToTpfcfWoy2KcDZZGGSMrbJ5zsiwH2tzAYws/xEq3xcNBzZPaLw9
+ddCYsooYPFhdXCqXWapABl60siT7JRmM2d0/Ox+Exyn+3ipXDkb0SUAmWnMOds7
bp7m7v9Ye5eDvaSfDom8T2a9lmDs0dXt3cR/LX5EViRGAPHlkjoW1t4LFhIG010b
OdxnairB01PhabtV0MxI/KM1PvwE24MhEnab6PVAYDYc019jpa9hKkXeEgprGGfv
aqixs3clh3spZAUIaXq4nB+XLeQMzbdR4nwIY1424EpySstZE7nH4v30q8QyDaB3
gbqO8Ix3H/RQLarpImxnvT1kDgPdauqM60kjhaZf+rWhq9RWL4l3eVxQvpkQovaj
8sF6/Jw2WGabtmX3skkDvGutmCrMI9Oyi1qw+a6oS0VTzPYXBtm6yVkkVk5LNFx/
XdIpQI+BtxFldrrF5t3PHMoF1PT7DgobBj+KJs4cLyOOGeQQhXreYLuTcBo1u7S3
SXK+wB7Hu95+Iv2V/t645Dbp39UJHCd+MLrsnR5wiDTeeJFt12rqvn+PXs9Rt6AP
xPxo5S+/LCaiZl0fMOuUPOgApIvr84lBqJJ+F58c4kZO529FTf3s/0rbASXpchZU
tey+EIkau1dqtx6/19mg5+O9lXPf3e45CKuUt4gTWjpfBwkgnCFE2cib3xRi3F34
l/VEvCMGoJkmAmrPef7FYNLNDVpyTX+/b8+f+gVUOYhq/OqRtvLUIhBSbnSeoM8v
X0EuQ9NRi11VuHvbpPFNKHtgrPnzaGEW7tL6UGciyLPLM7ZNsLFPZRUe9wABXO8z
r6jjwtPpYMSwrsm4oEAwnZdTZQHOy6kDBiUdqzsHxlqGNWOlEKk473BrVvdoyGUT
8xTPteaVnnXfCaI3wbRMkJn69XvXtn0K5WgjVBQfvtEy0PVyoDTcOH20102+D1Iy
ur4AkwHtx2q5NiLI28YhhkmbYfiABRieubfO5Hs/pMfRMTp1SHa4oIXDoHgeC63k
oFbVgBJ0BS+EJlN4elPgJzjVP6Jz9T57DnDOC3kI6Hsur3OVeeO3CYr/ccne2oPB
Dx3lzFtgBuqub0KH3UOrnzwbdAKKpAzIw27BCsaF0kArISDwvIXm7vXrdeSXDKN4
DOgNopwTwEzOA1HX9iGmhIgYSQsmoACsyfqzRBeKRQoF2NyH7u0mwQNZLBQWjq7K
sTVXmTpXw6qYqsw8pDMyausD/UaG5w+oEYdFV3gOilHEAPvCMwlahTE8a522FEIT
Pw6HLlVNmr9me8qANImiiEAFi5wt18thyPON+A8mN9v0EW4sW6M2+p4g/CfthVso
oKf6H1rw8slUgqomvbVF1Tvow4MIALoudqIJPRsy8li8gXQqLSuzBHgMkCQilU6D
ugAqpRQhYAm6LXoAxtBO2MlTb4ikdeDiz1gcRbzFXw0O3U/27IcZR046ieRDB3s3
/w02xGVFb1PO7qYj+9CzKhJmdy4h5u4I0NELqIWWZM+uCLtcbcQk6oKRxgVirthe
fMu/22ZBqtaAEtDyutgT+uc3LwkA8ZWJzOCrH/pYgay7lYBZwNMNRr9nhgiwobBf
TH4V9xM/bJi7XHjidE4LEMOI1MrGrBaLCZ2uK/AJlkunUUszmKsrTmLvuXch73EO
nttkQPVpHzG+xGBIaFyKCtxiRqo+gfWAgWwvXtknoTFdtItozDuCXlQBKQhvNQ2V
lmr6ILcrW2k43FDdAiPWuVAzCtBD33mWVUWhFYhvRjgJKHZ10DQo0tg8Y8GyZzt6
aMzL1Qu9ZieGqAeODxuuWbay+INktytVjX1YZOWWUyUcMkv7Hwi9RBD4fY/3McVD
ZUYc1mEWCK5EghowjG8vI5XlY1KI0BFgLDt6MuI/gvN6wGGLljbKeocN2kx18nP8
ygn2HPEHbd6LXU+K0ovNANsErMfBAaobN2MQTzNymgxwPiouaXWbWym/gCHoLNmA
C3GRIM6IAq86xHPzyvHsr9mWvUFz60Z2rGLLWp+/YIxabwcVY+e2aRDel1St5PVM
HdXC3eWda04EptyXj1XnxfOlH3Sw30MiAs+totFldpHFoQqOHK24r0aTKCenae4J
p2tdAPNKHtosNrZHM4K04Sawq7jwgcEYtUADkS8Y91h72E3n7wFb+wQTIIAiikPV
CQEOHREWJuN0uMyfU6L3EzExOP5w/SkClDzH/Gw3Oow0h6HVSzH+DoKc2sFMWRrN
fUGQuchwcJFKyaLrAMw15iI7vGYFrLWihraJENTllXxua2E5fxp2DDVEtFK2z2bk
kEtyB50hEMR1ZOgJAZbmfbagwfTFuiV6vLVvAg+3U+02u/CKkNXHtXoVTVLlYEVt
L0VLRtuIpn7IhhA/Mmzfy4fkwO+aDaih3avt5uWqolsX9nKWEVs1g1/OkJlS8w+3
72SjyBYVRVdULnmFQxluKOsVj4uEnTpWKFr5cm4ltfm3wuW3lmrQTQPBO/0Fi/Qy
Cx1AnbRGjpGxPxAbEIUDf27YrEXAT/tNJdEGdVfNN2xYoTOB5WgpjGxEh7OpZbxC
9zCEcI1hMzrzPN4hJud0faR/d0beZvzvIUe4FYM5IFKcGHqrer0puAxBJaPmCk7b
IGee5vQz6jUj2dqc9P5R/m/+8LYv36ZB8r2yukrSOp74cTlt146FYqtOX/myjYlw
PFuABnuIT2yJXy/b6vckjiSOScny2U7C1H8XVufzQrz1ovs9EtjHr4Ij1qX72l5e
HQtIDtAEeQpPRYvNq11T0M3MeDwfYJEz49AKQZOewkUHSYT2ROKTcAqXT7bH2jl0
RBEjkymeKxtrh/1jCBbldveeUK23yc6b1lDWscHVWlIIL+Ze5ORC0mDS84f2l8Yq
exIghGXAl/jblwZfls3miF7zL/29OAsvS3S/TJ3i635/fhLyeezVi0yJLrefML4A
mUDAjl4AJ7VljUIZ2KbO+Hw58LMpLgA0NSp/rwdVsd9n0d71/NXofeVeJWt8lcsP
hR8VDQy/ZuFPJzqcmJRZYdJj1bbuhE7JuWWAMrF9hlHw8Elj5cP5iOvZbD29ARQp
tv7rOiqMBXYKfj3NsONh8kO85XTgvFssxIqYUWGdX6vVA88TgfgWjVQqQxgMSI+k
IclE888VSX0TotzdnByJVvjAYCFWQ6ShJmMI7DtQjGBRO2gTrVAWh9kP/eQqCI1l
ERKaxXxnhVFMZSH0/2tIpA03u4CcjxChkcNlbG6wIn4np0H73gN7YyYO3J6hM+zJ
faMY5XxFUyjFAJmupT2GP2vT5DQqRJYRrizXK41N+qhfWJyiNdzY1+pOIWqMkMtQ
nYNgPeufqdm5hy9ZVRfuJGr6PgocrPzLjA2Ha73f6zaUgKs/jYc7mwVQAVCep6eS
qgNdvQElQ1LVuXRyX7eUR7OgV9I1UqCjsxTtEadNU/uLdrcLaenDX4w01RJjtKqV
6M0kZgynAzq48Dl+Y2J3K8DKThVE4tPCOFWhQ1eevNgRq/R5Iq6uAcPnplYLs7dk
1bJH4rt9iiP9XzyQFilsieT4db78UgS15lRRa9mCbmO8dJWgzA7I6hMYBebsPnLU
KXGkDwNJjPB0iGRpw3S2V9zB4QIehB/1LDgPiM3BbwxeH9FVdVWYztX6TwlKxbIW
N8S1X5Ywfgg8z5M/XIrO/xE9QQ8X8LtJ+lKVDwo/GvU9w3TVDVoTBVEu11f76I7c
5qoGCp2P/a2UiyWl1+mw/FKKDk9TAVOAQ7TU1/H4+Z4AGrXaluGd6ftxXuOKIaWU
BCaWXDLfZsF0tKRFy3kA2SWp9WTPTfy247dty96uvaWRvaK49g+jvaj/tNKkEQsT
DSEBlCc+kn2DuYxaatuWdBnDDgef8ZWDjM9XU896446MN1cuB7BVnNrZlmwtUWXD
JU2RPKfdkvnc/ZufeeccXmJMaZr0lLJEciBdwjR+lBp3kC3XRJSJjX/A2JJPuIqT
DUPD1beii7j43RikZveNHUljyzrLiZoNmoxJ82+Vh1LPAoIPKQLTT8UxPRxzRxzf
4r5H1RZMDOx00DcJbHzLXww4nJzj1LGhim67K70FtA9JKYgOq1XDttVrYIeKgCfl
IEoBzwbatjLOjnPCLgdA5zmc66Gb/ozK7eD0IahepIYHhlBm4YqQKVuUJivJRnwh
K6rd6WWAKuz8j6ilzgy0Ix8lNxtSK/wK761fGMkVDHeYZmYhYPb5k3uqA8WIAw1K
udgY32VOhnWI7K1ciBkYg+XUGGL/vGE9mZTeprHYaQrGFGS/SqUoAJZC+3TPpsOC
DF3Y0dEH49NaSf162r1Hzd2+9BPGT3LyvBae+Wvo2p1nNpGteSRicYv2dqM1NXxs
rxrvXZRhTzoptvoi36uulF/zQVCDCFlEfZKu20JrB5SRj2zNoPcFYCc/DWFqcoX6
4liRIs4jYrKWCL7lNbTQCTB7NsQ84063VtRHqkxhMaOUMyPyiFzta/7ubrDruchP
sXw2X3xvurcEsIlegztVxt0bqXUEejts6i7pvmU+QsEkoD38102O4+Qudtb2R6nk
Pd2sBA5STIHv00899vI/r5u6sNM8DtmbJDBTIeLCM23pApY/093rXVvT6XPs8zOL
kHHd5lO2PFIIBPSG2cl62lzUIlix95lFmLJ3kJdt0QPdL37zImwnGzpJi7OdZ88U
8vD2NViniU6a5KaAudK++HrBHjn86ZPB7oslWXziXQRfBB/09E4gUaaGAEQDs9qf
rJOD4p+MnCr6EHJ0ibJjeYMzQ4cwChjWCTcDWiW5wLP84MfQ4FEYs9yItDzbGnwQ
bCyCHdDQdaSOt+HNsCPjr8aN3HcS3CzGMeGb8x/4+f+T1kpk2XVx7WGIQDO9+CJE
0tiU3yEyfkr/9wuqBZuKga+vA89taaM9bVJwvj1HmFy0qFJa0lBzmfxoIN2uMhlU
Od/5bh+4HI8/ttTw55wfHaibNDPjdi2pzDfQLcgL6S1LsrKsdvm085GU0S6jZ3/b
15+bCdsUFB00QjuGeOBrfwJh1w0MAEKMhtFEGmOMnOz1XbuoRkGaG+uVKIccGV4W
S8kkQhh0Iy6V3r8PDzlA3kWAYYzyILx3rB0gx2Mup7GD98Ne9wRt1UvjHIuU8dwo
pYkq+7h3HOBgvq8VMKWs41Wg0H3J8cY3IKHyr9YlT71ec8YCd/H65UafBNYYdI+1
e/p6Q4czVE9+Rut+BN3nLwjiwd0KcS5pzi2lDhmX4Aouey30Jm6QEo2YDUglOu+a
b/0LPuzbF/b5ku1ol+BDxVI+RXzap0afLU7E0Qx1VIvBYUDuZa0hGwKcd9B3tHVO
L6Ozud0MmDNLIl1koY+Q5O0cf8SXXTqokZXit+nzpB1QfBbVTEvEetCsi3Ct7IyE
PjzjpveLdM2P3kH0unyxe6oBbwgaasyBevodsg0IwA5p7a7ONOy3harQM+8OqKQ8
3IktQwynSdpg34xWeR1aQtCA48sSTjLqZqZzEU30MyVp8ALraANg4n2tDdF+rgBI
wvD5+Ii9G39bFZk7srSd6+q6t4RvFRwG4T48UWkL7Cj62/zOEhEioARgic+bR9oS
XtDMtz2HwPkVYPvLO7lViy9cEIbbN9wKQFUD6pMOlw7Fm+1YhahkBAQFtbDx6+8S
/P+0PhsNqnrQ/UYKzpgY7ZsdHJoCDzw5Zb9KxCabnDetIhGT5P1DcBoV3bPG0jhf
tI3X5Y8Rq7MD80kBNyDtCzpob0Q10smke1gpdKjtyFA1mmPpTECsH130/7qLjvK/
6waZM+zoMyodi4Ul4KenO9qyH8tX8vGcHDwlmZIlwzytdosU4L0P2p22ubzv+API
A+1rwvUyimF1XdS6XmUC7zENiu5K0HzSprs2tTT3mdr0mrSL0CrSB/C3Opri3zaI
kbEoM7ZbWdYHsIdNE987wHPlfyXV3J9iBDfYsClN+PZvmfz4JjuSFen5MZTZ5oqw
ZAG0O8Td3ROA2HWeChpTmcNB2vME7IsBT2Ke8YcYRlAXlIN7rG51M7m/tSLHR1X6
evDU77nVhUtmoDPD99G0EpGrGQzHz+SMy56WZ/pstKCuXrIGsxvrHnFwt9Em/Bb8
XCmo52qM2nWfNK+TgxCgVbV38jGoFWCyAxiHI7G6LkOGM0rax996O+73FHsRNXf9
GEyp4mv6HFT+DUEeSPpmYuxDTWzd7n1bMuU1Mw2ijTTCekiRslZUbjdrVsJZev47
LHpHsLA9LIAhOLMQwaHIs67diKblH7ev76x3JHo+lGFLNJEDXeb4bUCuM2AHdUR6
Wdfng7frhs2zEK3IgfhugVpWPJV6YfVaQ094h7AtXOwk/5NUTUlI9VY9zcISU1Og
RKoVPYRNYdrwt7C4Bkh3eNP/EszEevBfwSb5pWf7lVurgylK5jpl3HeROHaZzvcm
IFhoOWKPg7hPNae+eAjpuS8xeUgv74qLugIRiH9N8lA9w0lhmwKp/h1PAjkza22g
1eg8ETK53oSH6nZgQ7/Ys0GcD0Ek68ebyVy+REiNx0MFKqbNOWceOZxX5MM5OTJn
TE1TnzdpwH0LmSL6p3+cLvprLiML6f5nHcK4/nfQoHmQMJa52RCxRCrNciO1F4lo
pkFZyloskPJV326Hw/vkHijeoGbTmS6bnc8ryB8IwqbjiaqcQ4MUPuOj3fAKTbGT
A9AvG9pxKogbk3AOn86e+mJKpqcEiU6BhwfM4KxIxpDwQYOvwrakGX+kEuHAhvsI
Fi9lDRvDBkZLQXbkB3oCG7xaJ98agyl2fLqhipUhQVADnuq7r2JdXLgnTY6JSs9E
qMh19oGrZGwO3nIzzenFXajf8/GV7qbnGiIozhwcMUtofp2sfzyPlvbNwseGf4Z/
u5TST8ca9pGnVfZfT+wfjxZOYuPOoo/yEy69OFHiMWXt2eWwGdkpePrKA2CZhbZz
vzw7xY/wbVQK0BzY5u2cRIiptM97kzsDI1ymwmyr+ziAT5Wo0ZPysn2WGssn9/Ub
Z2tWQgQO0+QvLaw2qQOMeG4Kc3CrtphZ6B8AkujvNaLPeQIkCKnAAa3vzVUNJlM8
Lac6+R1O92DRDewMvypPzKAVbUSlqQe4eNoQxP8kpsFn0rG7RgvDOdDWhRzmAmPR
ZtIPrWlo6bOW5WdBs2GA6ktGkiNJMGzt9y0sZb9r8BUvy9YAK8PdkS95O9kSK7r8
vWVlFexq/zICy7lXfgxvdne7YowZUqVCKXmBn7nS9asrualOxZRN6lIKTL8TFf/9
Halk7ULNarQO0iiAMGiXBLerIoz1VlwqNQjV4wa/X2h9KqHxZZSd6rODe9RkhOwM
M/ciRE9LobGVCCBGiOe1Siy/r9Xh0u7tZPLyLf+Yl4jO2VYghZ7p/hUE1XqStkI4
38X+8q2szoGkNqzYJcE2G6fkl9Lqtnwifjoot/Q35R70PzOdB9mm6b6mp4eXJ3EK
3KlkifsGluOZJIuUmFZPAnBHfJ6Dk+ASotSwjz8xcjHsyzXVBid11G84rN7IesBp
ADND6JW8OHKSHbVnftEadMNn7Urp0NAxPFBFpSwSbJeNA/rcZhtevWTnQoF/q/5n
lCjrQXqSB5Uai7cXZn8lnYFHsEUqCV3bXGQzRhk+97dLM0G2Ma3N4EIYNo58qdym
jes7sIpR7APiX3kJH8JEQbL6SeoWy2+22vm6JdZcK2LtW6Q0WwIBTXIrUYs+CmNU
kfhKPX6vo0x84vg9CE+mfxJvAdqcRY+wUfwFK9eXBjR+DJCCgi1Q/gjJbVfKPEmu
RkQ7t5oWiMhfFbIL3OKnKsSiZcxE6BgHt1AxOHSpdNfVz8mlJq00fPXB2f34tsaw
U8THBZxpObo10lOX3xvw0Ryr25fx28sDfme1jgnuLN81J/AAX0hWYNHoXnymmKn9
p4MYvMlhttunoCkBFqR6ThD/TzZjAl+BQmW8u/Twe2l6F9pYBdXcIc8wOThZdfqS
OMgIaRCVZx8I2tszi9UdN+Pm+haHc5gGFimO1+WfL96Rs/+pRvZoyyxOSX9Qaw/z
RpR+/x8y7u5KJlOl9rTZgfpGzbzkusULQAPvqFrKyPSQYFsaQVQ5ywLeCmRFrDer
M48hJfL15ft2OvSlJD+a7xwMSoFzWNHr8FyBdTTNjP9Uw4rGg7SVFGKtpD8SoDP7
nlvKjqD5dwK6C6yqtcZucIODT/PDCJqyEsYgIVTTRbFUsi/TKWUY7Krcxx024Cdx
41VvuWY+cXrsocVVU3kYmJScklm3smVZTQDrK5yEyALWFFbd79TdbU0hpdA4GwwE
o6Vfn+89g+DAe7LXwiOgemvKfPGMafoX9RT7/1nLmc4LGpe2jf6vf0h3AgJB+Eo2
/NaEOfFr2W+paO/pPwpYxGYQl5FAU2fJuszvM0JVR2GeH10ZzL6sknWiiHjW3ebr
g8h/kC9pv9uxu08B5R1uLRUe0Uq/14MdC6ha7/uCDq1Hi5XjNPYGRMBAYxfQkjWq
4tbQjqUHgSNFjxoSoEK+ldWfOX+f+C25MZ5G3go+QnX7h/8LjehTPTjsarldCzGr
qwW5OKMCMbMhgTJPWBqyNJdW1ykMq31zMF7FJvMQhxMiP8HKvX9JbsI4o4TLzZSp
vHfeU8VT/ptvAwHiguvk7qaewig9bhW+6eh/4pr/IOZWmVC3kJOjzSuUNdl/bGdD
GqY+/Laas7mBEe3SMokLFfYVy/66zfftLzNicIAUwE5ASOgsE2/+JxYWTkFxblkC
eQJRW3aQa9pZvnTxbaVzCkSIKu6BP1nGxi+uvMmVt5Bor6326482bmkv4Ywigjy7
v9W9FqbzBxRRdJthE6ieM3BCalnIlyD4zBA5mwHlmqgQ9TOOZ40g8IsUVf/a+dCo
uqR+qsT2X0F8c10TOmwiX2iyIhwmyQxpwkwODmSjmCaF0AmWpDaO88bttkC9WenC
WUFcc+SKpHYR++dwnmdINIZeHkRPz7+HWk96UUIQOtevl0VsiuNEleaxzmLT2eDI
RCZZUD0ZZONJ4gBZLIsM7m1zG4DO9M4dv2bJmbi1gPQ0gJ3GKc/ffVYg0oHQeACF
FxRSVIqW/kTCfUnym1aZoi1acSUljmWpyNQTqNn8peDmhTlmvFG7+Zg90CfEA8Mx
Ga+MQOarv+6or9LX7BCa+bzpGX4NUgbw8I+aJ47Wz2WOLX3zKFoRxnnmBgOjaIRt
hm0dV2IpRzRpS1iVwDYNarNHIqUPL6rNkeE2SsVuMlZ1yJ42jnvR8WehJD/vc2kR
e1KJEmMxRu5Yonxh5rB4SXjT1DKXWwjllDiyq/+CruwDmoJHY+qz7d7KozadO1fs
59z+7wlzfvMRPnPLiAII/QQIsPXKHXvSmzdSc0GrVDky++Xmf9nVG63BiTvlougu
bIBMqPITTtvUChuivEsuvQSwvPcv2BpuZvrU0TS8vrHZoAKxhLbWvukvyGJedJmE
tD7uk01mZA1GK4uzvaN7QqjeZwqLh1QaM9UyPvTU/g/HAtiKo6qqP6AehqLSG4Yl
f6A1i6nqZsokucxXrpUmhSAvtAKHr4PxaGiNKqAusAjRmH9xC/rZmroccLfqNcMa
c4gqqD8kriIDzn92MtGHdvlKtpcl17t0b4ap85UuNkWQz7T9ZS/N7uJQfVEzvNSx
N2xyuSpJ2USQOeK3uZ91ieupmesONXF3Pne3yDRnWhfNeO4ZbZWZZ3XrkC7Fb4ON
QMaZ8XQt/wKvYy6cCzxv7Ody9MdR30tVTQQSTbuV6IhtBrw2IpJbThaQI9D4dD37
N38LS/VuXUNF7EN2vgIjD7hzU3jqiBYIz+EE1LDTsA66OG0VcB7cYm19cEYMYcEj
AwAVtwxQKeNOuWZZ29ndzlMUAj0J8xYmn3e1SRQl+nQQ9E2RnRWnEM4Ivt2t9XNj
fwr3TM270Fhgz5g/rIJdAaAMT1Krv2utQZ9Xul6eqk8BBVH1AzlNQv/JX97GkM8d
VWL20my8CX2SeLQAV96a++ED8ifTjBcWRxekj/WnODCfGG6U40NzEsv6qe7YykUm
7eoQSyjuC7UpaLuq45bmmpaw6YQaPQcLm2T4OvcOwHdi5h5fJSeJmu7r4vqv/4n5
onH7wy4DmSDrH2Bzj6GhhV+b6ePgmDnn9VgKdZexvmTd06FQcE7nTrloHc+V5nH8
ICsjrr6Xx58zUm1jJOrlV7TZBtx7SFhEghKd9QiAfqpwefQcUcs2Ug98nmSjKmiX
KvVNg/EZF8fSyzc6ohUq8g==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MEoimOcIvEqdXr72XnOHYDbeoPmFdxmKuKr4PqIDaNjf4OSPS3zWQoz6LJlYonk3
LLLgIeYE/5HWmGmFM2Cif4UJPRNDm0tfnncaFoHbeOIasEVAgVf2qHyOibVzeKoO
ULGP+WQsWTjlygWFmyGAm/BrEMp2XBPhDXiurCLfZPE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 103472)
mlbvLia6v30OWst9eolXGjrGMSH5omPA1Zl7vjemeI+b1C3/TdFZPIR8LDQqXojg
2oxSC4OH1glwn2D+C5CY9IQM/PulfVHZ9kBJgMmjEpRD1NWWv9Mto7v6h9EbgfTu
CxULSDa88iSJCJmM7MXV+SY8fte7tgKW6Jfp0hXyk9oqk62FyLZXXva5MsuOd7BN
1toiERmkGe2gUmeT6zlzn65NPI3yNITSxN5+KcCu9KvexlMcPPHurCMUzKOS/YbL
J5mWGmiJhatodF3lYeBqyDGGw3l26y/ZGoSV0bjylfJVyRW5vQ1ZDGhIqnRKfFXM
xreQlIWHyrCDvaAcgIzW/S9KyQ9fG6bb7f2mMbvF0QiXCh4uByNGR2bsX88lTyxr
m+yJU6FGjLnYPLVahbo2R9BIidBDDM6IBmmp+nnqh+xS6wxqnnXR7P67KLVUhju9
XlvSYwawG5DN3gysG+pPGGki+riAX095uKZQVrMqDfYThm4MmM2EiaOY5gu8wKcg
6I0h0EyvGXCnDJ2T5TwWkna4JCiSHQTMGR/e3i++4HbfR4lFZiPR5lN3nU5EAgth
dJOIw5YgzXgto0YNH/Bt2DVsZR8bWV1wPpWIjsAEVjA7BkHh/hUaPlEQWnzmGUta
Vt3k3Dz0ASkxq5DcNj4s9hYbJzxj7/ZkH5ZF8SwEJmg8VtY52TIk+047hI3xcHYr
95w/EcBHb6WswC5gttdpqWZazu/7iffsx0pCjrRPoH82qjJpcWyu+UmrHdXIwopO
0oLrtXCjRP+6P0yKFn2ky3SOeukBR0eMTwpXlHYFMPkGqsfRl8i/YvoC+YWdrziH
vMACWaHMD8ZThrZ0cBqUKwM4W76WQUPFm10/Fl3PsB/rSQOjREPtiRdsqst735Gp
itWyQEyjNlIXlFXnkIVshe2bl8tLw8yrdC6XHRs4XHVGLS5RgkdbRyPw7ii8Nja4
scqqEbYjW8HmoO6Fu/MXOZuWw1FlnSy47v7SoVyZZ/3mGgmcoVRA/8KPCDJYXHA9
ElWHqkLD0duN4eXRMCYJ/+vz6yi+tLTOcWOG7Lj7WTmi2uKljUWnWy4QGa3NQPVN
PtLr7lQDrmcZFQcTzZhLMetED71eLUn+VIkcf3KIm5WuY0rCkbG+DowoFAI2OJeD
R8lw72ggLbX50Ce3KCTR0dwm+15zO7aEWN1ShbSabpPpZDGYRlZZKenZvCKUGNCF
O+k0fJp1VvYdIkt3wXdbh5YpC2cUHx8nqatEqBDoYPClGtSAxbaW6O1JE9ObZkZO
WtmvFCVah793Zl2ALSiXQ0AJkf4auKiibnWYtIypUdK+hyKZgMALjEKKLsOZSDzL
tQccZzMoSrtXXhra0RRO63TQK9LZ2WPZArQvdJrYtIFmDjO7+p7xESa4NzkvzZ6H
JlzJ7ePr5HSKgNzu7Sr/CP5a31XyNmiGE7A36r02k35f1wJM1cR0WA8cPzIcCX9U
bS64eaBOAH+scNdia1VKJVtTa9pU6fyHjuEiJk7JlmWjsqn2F9UzmC8qMIjiCAtO
0G5vTKp3DCegqjDkW+OVmxulT8aYc7feqTeRW/Ly6381yHiPR38wfKNswSr5gqLo
542Y2rOojTjyoe8RHJ3nuHMGTvIxq42fOLu8FT0SJjnquymSHD67QPiN0Jrk/bEd
6JAkagwkkUPfB3S3RLarqsYwXleznOF1iR7Dy4LTOCxtEC42/WnajRsbxudGXpbc
X2XarnU0bzvLcR8YyGCf8glKF/PTVXacTChJkmFZYT44SZLmvl0LP/gKjix7f6v2
R6aX4BYrvtBu5+Q12+UVIX40DZNtuOnT7b4hqgTkkIaDG8qf6ZUWYL7G4Cg9NcNX
Q/QSf3gt3jGypYE8xB/gpqXsPjD3BJlEkNrDRMlOMsFWPA4eSiB8FEYmBrV8Yxqe
a45BMORuIRhJiQh6iS/vTlMQ/2zLU0bErYIDkUv4rPJrnVhPCA4gZSdzOvycOIl/
S8l+I6XQhOnzQu08KZ4O3zQNyszL75gK392VOGN6my7vf+lzavguoUKqEAwmL7RZ
VvC/EEYLf2GotO9smo+CpEhQSyuJQ20i3818FZmyrFThFMAkdTdlC37xbN6B3Ld8
OlDhxL66q/eNIvROfahUuU/a/NLe46GFueBtP+Mi1u9fXArGl2OqeFlM9UgWAjfn
dBNgM1pdtNxi2feNdZPH1WODCHoP08PKn0O0THwb0XvcxG5Rt0w/kLOD504p5pyS
bub+ZnCgXv2oKSxY4IkYZCw/lcWZqY6spa627eS44K2qYuk2/uYyj4EaJIZdlnAq
wkWHQsF7u3QKJIOgCXg1Y0JwwcNG6EdW1A0HF7kRWTcmglZLojj4EdZ5PjkkWaXY
pckJRlYWpzq7PB0uwcvM3zcD3xJxHphcxvjdJ1DAYZQ8C538f5/POQ8EEp0FfgQS
EhKeuc+JzhzBcCsToYpeZQhvzvSXy/7tcRb3PpmiQeGb+x4QJciap/Ru5+od8f4Y
BfLsnLtwxE2kZrY5bxdwGHoE6QHhGs7iHQaZDBxQcqpNhdLIkGVL4He5lcsgXhKl
bawwC+Weu2DfibRIEZEY5GOGxw6T/fgc+xGs861nhiBJ23RKTWin2bJXCM3GScpz
ZGuqnmJSs/QUA7HEP7YhobtTGLz1YTiFiPLdHf8rTTqOoPws4utuBXQU/qvySj5v
cchKA78SBe1Er87FDMUms/eINq9LdEA5v93JZO3P8NW6NuwA/9jQ/eXDAya9kOe6
wDQMVp/fh6/hsO5Fm9GtFNVGvRsPJafOY0Nj6QnH5xM3XQewUzH7PvJJ9JNOGVRS
6uc5BxXJBpolrjChB8MhsfT9TV7Ib49luCoeZxrc3HgRk9G2Ey0UvfTz2xRzDsI5
PphNJP3TmGjylXn8cPV2B0X+/JoZZ8sg12DYFvdoyk2SG2gIXTqxs9NNfFaVg/dC
0T+9VQeQRL4i4/ZadxQu1WLaoLHra8D27wqe/04zTOPuT/qUE3TKOVt8TrhOG5Ft
BVzAqjrX1DW+OxJtD8xF+MSVa7GQFwWI3xvcSAtRhLxHb6LCGV1Di9v1MQ0p7sKC
yJAWeICUce+Y30V555mSd+Myf1zw1lcT8rBncbLUC+9zshafCCOQFcXx4u4oIvyX
DkyXOOFqzKRhnfvMgUOWlewdRmjFzYN+zn6pmhXVztrE9br/DgkpMAknYdBQ9ukZ
ijn6okSL2uOJTL9n0X7a+BSDeaxILrk3XMKvmUQkA74wcKXa/NPN2ks4IlRLiQx6
hvIgi/r9xjBsuzLBH9oY2l1sr5GT11qDt6hVieWfN6GyAAu00tCv+ihToFnX6RHQ
5Rt/fuhz2yA0lCN3lkJssX7JTuLBhJwbFMRRC2hugDPE2Fr8fKCY4dQnj0oG8WZ9
ZmGg4P7JvwuN3qdAzhdThMTksVFBUuq5DzyojvdYAkYTCRZoeX2lzW9Wq3DcVo0z
FNpIaIR0rawyl22boWzRzItAdDyGd2vatmfdX/Zj78vke+Zl4noURDvAmx7oljko
Q04sbJZqK580JL7YwOdyKuyfXfEeVoY/44EH9H1jfQoYOlKSk/WZfqZq+f4ZKWw4
Jsxte1lSIEJDzR64htxXWPMfhubnS1y2cG7Y3sZmQNytM8UfKYHJOIHRdTKbc6nt
kmUqmXYwuOS0H088xVMWIo6uRsNOlLosVOuH9kSJ3kZUR7Akf4RzAP4O2ya8HXCv
v0JNitqxLqUqdC+T+5xrPkKRjq/HsOkdoc5IXbbqC1Duptvxz84qkNZAOQuhzzcG
Lmo1EcezKA+/YCwY+Daa6ecgKwqwezYqqCZb1mq/M+ibMU+QhMYSSPh0N/lfeb9R
bxS804boOYDY+YmogTTqPfrCH8bc3Gw9uMsbRk0d6E0kJ6AGllG+8C0TDoq6Zyln
2hllMpF+FImHRln9zbX+Xbodx8n7fvVHxr6ZRN52lOisPxHuWFepNOsuOfUg8XP7
3PJjHZ9OGx/Ro83DfISQZU7o+tuLd4PHElniOPJoSXjmMnDl1ko26hYc1kMa75EY
9QNxsnwnFb95fViIVCDdW0WM6LIdBbXz1XqIIY8zdrYUDrnB8ibErDc+yJHOSqA3
o5GoI70rXY95zTRrlWd9ttYVG7umr9J9w7FsVmee88sqZAjJ8DVu8X50rtMLQolO
yPGvmwZozdgk3brsv87kMRGaKz/uvvt5yrwba3NF9KPkqNm+ZDyWEOVI/mzynnCJ
HqgxwDAgrbmgBqxjOXYGNjcgHiJsX3RIts0esC5KJ5+xhVa/jQJtbcBhwSyHNBrq
Ew5tcbUPGh4M01e6th9REzhbMss6NhT+95s948ric7YK+vtC07WmDbHCXBAVZVpA
HKoDVOZb0tJALbbJCq2wmGwD0Sr6HO2JW1btIiJ/tnVuJG2PisvqDfIUf/Dmu6ib
HCUd7EqWix4qS5qLtDWQAIGSMnjf0DMqeh3iPemVvkP40ObkJUgFfXllejY/xh3z
6xwQBBuo8zZ/1Z67QxXDx3V+ruW4vftcOU4uh6QU6gJSWRsX46uB5OFuj4bgfPv0
CAFVyiB1a/1Bq6hw0DpjX/PstljknictL9wWO4eLQvb4IHC9km5FKOTBO4fO8uLI
i80vViDiAUpZ5m47mYYBfEpswpwkuDCTGwiw52d8+GBzohd9NvzCAKb0Pc8Huzcd
5WBR1xVeKNX5m736sjk4KzqU/Lz0zMwBlW6hIpb7jIHA5DQVfi3evlqA4IM8rSVe
PYp20gu99gl5DNOiWg7Bn+2j/DhE01kcsDrJE/PN1eQ5F/rxIchZ5aBo3nos9M8s
53lCVQ+CInzI3wMjRUaSm2OzBAHQacp3IDl/fJMfvVbfoLvTMGOeOTTJRePMmq28
ODSqkXUo4tesCEp9Dz+Icz1cfVh4NG6jJ2jTOpUJ4FDUUhB8A+4HWVTXS0iYiWXp
6FXBcOr9UygPEjq0O92ViuWXOF760ACRzIOOcgJG8kg9rZiuABGp1YYpM1Vwj0UC
fZg5VAcNgsD5Q9LEoo6daWmX2Ulmqr5hJW/9YvyORqzHuAv/OonYS+C447HKhMk2
n4DB921NjLP8A3w3vl+gzxJGaqFMqvCs4VpPAe+v16rd0eNWSk2WYMhtgaaAY5Yf
Dn2fsGuPKHSDjsk0iPGC0mIuQf6iSrwJYjiq1v2Tmb2kmtOYpjba/e7YublXE2Uj
pJyPtvlaYYBUmlNQd2sB0whDb2eW+XxvuaTyXNajxmX4seRx+zQlgEQm2DzCE4Of
b6Ic3MQExsB7R29Tn22dGabiWcw5XdQ2X1i4MyF8Qm5JhLcOIP4FEDfES05064tV
VzxE4YqIobJbxfcbWTyA69hHETEux97SkRgmiVEsLLMo9eiVzbOBsEkkH7jv6wro
CqTFhL4BnNfD5LLZwg/D+Me2Xgrgc2it/yMvgfHGpf5OFQjmBucr4yPxJo0oH9MI
fP5MvpvYZ7iLuYZl20Y3GCSH5s5PRqODvwfkfCqF0NAs4v4IQbr1/sg0BScCObiV
K1Pf5iQQGOhaQUS3LJ5oehAzUs62WhtJmwjMc/8+3HpSEGntSskEyTM+ol6+BX+U
W84ilsnhrnYs5O9e9TIZXyLPd2zpuiqbffotfGK/tCamWP8Nn76t4antSkKes6xQ
x2U+yxy0+K/fqhASfazkUIQKWm+lCd2VyfqqPtsY745gfGlDQXVjsHAV2VS4E+mb
ypnEpZGCrunBypOJiFlwv55ut+gNviA4JQ+VvjMKRb2ELMUc0l+bTLQw1qf64+YQ
iOw9e14Tm/WzUU7idKzeoGVXZWgVQjYHbFuPl9Uv1eqS58+CLuoiRFCfBd5T/MTu
mxNzJn0Nhp7s9NqSWvFjkbC5MHk9wDh6fDS7iwpAdvdQH6021Wn2Fr/scaNRhoIH
TwIzp1wx71TAzauI8LGaHZPCmlj+5/4IFvtoOnyx4mdvVG/ySDSAksAA3dhwXpwz
jI70108Admvksq03u1jDvSrriheH9zdmUdJnmCUZ1cd+8/66d5Op4svYm+aoK6SN
ByzbYtYqdrZ7eHV46KUB+w1PqIvZwyJh2qUgDzcgQPgFv1t/kwo3bJ+jp7wHogSa
SG5uyzjvxm+bu9n2aXgtYqKtQD0VzacPc9nBnoZQSgnKwzrJbRZv8xTahXziBVyj
dEujh6maoc7X3Mr6VzFJs7jzX6BCFNcYp95Wk6W4HyTES1te89zdyT4pxuYxPOkE
Igq4EVQvL+mNONDYgj5m3r8QVydMqgXwPu22I0Te6gkJO64NolJE3ClxEjRWoLmL
JfTAjeULwMCtgSnt0vuHBYNaS9YUXL+xQux7hy9XpcY57WmctMIDy4VizLBIXHjl
56kHQurkCI9275IQcAyfeznk/g4xtNZ1ruftz8JzEnvQSDfl1CFatH9aqBXjnSNQ
WsSuLEvFihkalhskDnkCJa3c0dJEBnhdJfCG7Kyyx9oNiq9MHVh9ywIMx8dSyHBM
Ho3gj+k6oysoFHtJzSlvY2qmu6OUMQXg4X1aJeje0VIE1vpekh5dVcLqVwK45lJ+
ZfOL8/yXAiNLLRRDqeTJI5Xh7zeyEaiv0IwpX8+wRLZmxUMhtwC14dO4qixvBoop
HkYJSogJ9VhzpQOjXuHZtLvvePF0N3uiTr1yv95Gwa5ifjblmLMz8GpzRqTFBJOG
w0N3i7RblwOQCMELsUl5p5JtJ7nAlwfkkPF0PuEibLM8d4BXM7WlXLHL5YtCbnAM
NdcqnWgpAq8eYJKcqvQUxz+uSon42br17bIzK+ekOSCzUi4mf/WOs1uSxb99gtcn
06ibofrDtcd0mvcxBbwBKxeqwj7KM1Hh8o5E3PZBEhh+RkWGQBkZq29N7wt3LsPU
MBFBnub7N3dPL5xCVIXKvBqFxL6wRYLAZTVCDiuE4zO/AKstz9r62NNqeVEXJLWO
mdCHOzC7qcsYzU3+kllDwQ5hEAUzpxcQK43wrTQq2qt4PyqiVykJqbSweMJl29Py
qG3QQlmiWdUkPbbTA0ipw8CchozTc5O3JlFLblK1/Y87obSJTqgc9cYUGeFfgLNz
F7elKo9bT7aXUB8wXMNtKJuyeOKXaaX3i2MjnmArdSWtzkUM8H/VOMEsVe6qwEeM
qylrJk1b0rnSTjcewAfdiI12uxBp9eggGTTTNVOOlFYKmur3gZUItL575cCKDJS/
cjSwefjW6z6bROq7++bxJvzYXBmwGdnFdYn/v/maJEhgfAGMHcVhoQsojfWeQnU0
owvhgh3Qt91uKIBkRpt0cSCxkjH0RLv2wLyh/0YDVLFqgQH/rvayRjOTeRC1uguj
RxmaHQZN8ZvwgBZN06aDO5B7YOdJpp4x0/WX51HYZ4LFWAPDLv303fdjzvzz+c/u
I7p+LOdzpB5NjJXS9L0L2loPGeBEr3sXJ10zTvQ+ClEXbZZoma01/JQYFZAEbkhp
r10BiMBN3zaW8Nb3MBVVLxcKRpf6d3XdhCmbqK+JMIdAIIFkZpMNSpV8nkHt/WxD
3orpKjX21cKcJifAcff11x/yoyAtH2L0DDj4RjPfg2F6D3GLwb0pUu5hG4HpnM7l
Jli6lysWJe3E2Rl2b1ASlO/Zm9GPy6g0bWX4RPpwWmgKIlyBgxisi7QDo4BVbugo
X53Tm2yfh2XH8/5LcESUiKpiCbhfjb/IG/X2qJanDZr1K4LhgD7rGlFf/gnVdtdE
aint3iqSg2JqSdTS/qLuepiAV57jpYPbugnKRSumGvvT2DyOlAOZCvaEcpLVnZ3u
Ry1iTTR1E+iOD/RglR3eRtniDa/4aa3qU3KSPB0sXtPni1va0/G7HwLD2e6i1POT
hjR6bcZGXah5UgeBx2TMw8/+EBOFBu4JnZ3Vq57hPfmzT4n+wLK5L9hxuU7XUaTy
rWciu4dPnLTEtMJZBXkxKqi2mglUQL40Jetw7cpyken6L02rw2G6OZdZhVXz09AU
+K0dLx8mDdaddv4c4GdbvqEbDfLsYlo+wMzHdyGETgKQuSuoQRuGoWIdVPpl/ifV
OrN2N0De3S91uJr/WccGJ/56uHKyAHa7IYuYMyWdkjgkhy+oVvEOT3ICEAWOqr/G
UUJJp66BmeNaEV6hFQuOha8tVbVeO8yczey+zV4cm0PmsS7uvgU7QFZX/FlKrRmI
/L21FP0Hja4QEwYnov2D502aI7SmW6MKWdMXbOk+2oEV/2LZCMIMG5eY/9vS9yh3
LidcV/TOz3ZiKvdwmi7yeGs6cCc0RKRc1fC6wx4kkgPgBLcwk4aHvGuy07VvojVc
0BHwI4694oAiFsmZ/ip6oIkbiioNmxLHJH5JL6ClljrJyFVd74WQRCjuLMNAs60m
NlrNrh9y+XxDYq91a0OjAiVNwlOX253ObzOLCkdI40KCJtPEERKsCv0FvJSCbJFU
nXtO2djpSKaBd8OYeLvNLUfxtY/f014zL+7/6VHiJ8SsaGepyovjOYnsPFCPoMoj
4BQSw9h3BT2LFqYwS0pptsWoeaScoLanCEwDH7A7T83Vu7GSIrdUPaqaxdMpyAZR
X3XVL92bz6hApChYNIbIm1zmXSJTPGiW1xbcvoSSF79VHWnx2mg3TwmOYZZToS48
cLyCuWmZ87nvZf7SckTSHvZxM71gyJ39OKshiOz1H+jg0SWXVj+PPXqe1imaahrH
OMdUhQwcTSTMjlr0w23l6vo+mKCO0bNWpaJuQYu8T4+lczmTOE/HGhvbi7OK+8DP
U2eX7pGKVeqUVEXyDZfaHk3Jzg37am2T33cYWQlv5HtQrvEo/ESk7hg1tfjFXetf
PJkJG6QwBSkLaQTtwBx3+TgthkLljoxOYBtTq6qvTWDS5F2/xMTes48y3fSavHy8
2Hov8SrDGh/LEAm8fpriGx7xEa4pEEsjyVA95vYSz0tawAilYN8qlfihlIivuwyE
+tw1Sq8u4nxUlmeq3FZxk53/1Pwjvk7D1okKp9z+l7u4iDbltn65ioGBohkuQqqV
9GdJ+H+imV4nusMjrbJoCukxY/7WlFTH/gR2qh7LEkr/TRXRaBZSjFUiaq+qWAm7
pDl45ARh/KFAiZ2QmgLFqEmZ7H8NYdnvKFhB54QDT/UQr/kvNAik/B5Z1T7wVK5o
1vUsWbDYYTNbTF9XOAiJfYj5vwKUX5Lf/xPeb0xfzCJS/80DpsYM+8wVZeD6LPxd
J4scj31yAGPB/rT2PHUSdzEnfToWz3dISOO0QPd4lAnVKdyIJhBTQejAvahMWZ7/
bcNcfHQSE9em0uSzm4ujg7UhRXTymola+5/Wt5/iE75BeE1IY8YpbZ97HGCM94gt
AjBLsmBzihGekcROq6sKc0UuUMeHkP7WpQfm5EAhL78ZiRFmSEX/yH7FpPMJsyRU
RRlxhSVi/+HqLsJqOIxPNJNXu1uw9EuzTIhE03Y13nSO3aUv3Pu8nx5jD1D4XfwA
3Cdsh+CD+qzxzXlgmY0l0bCpKa3pM9zw9W12uX2C9W50OeYvwSCwlUTxbRkDtBHb
RrS10S6QrZkkvL0tDLDDf1Ae4Ng9XCciF6EkPhQNcWLtq6Owqt4DR34i4ERH/nZ9
Tx1qjvZIBj0My1UfQuq7Xl7JyCqhc+1OmzCN1rR+EaqD1hzlCKCjQIT/Su7VtdCj
KCqAegAoTbdEfZcdZX74BgLCoN6q0c2hYQxY6p8Fq6h0bCep9+85SjruICy6AoBg
ysNZ/ag2TYBWkm2N3Hi0YzUdOhebinmZp87318jsF3t7qpVqNZosxEzzEVjzcqCR
ioPTTIeZFTDXKJGlEdQ8jGUbfXS3c6QaZWaLbHjUnqj9d6ZQ05HTwB/LjXmi06SV
hahhyucOYbjx8VIK1bJu3SRQGcQzpcS7Ydhta7X942RE1hWKlmrO7WqdP7E2TNgs
umB3xlvltJLa2Rm5vaVmEyey6ZhVMX9OUFT0B0StLoTEAjKhRUyt8+AKMzQcBwBx
WRhC8bGjasJLVktgrD97Q3duWTa6liNdw3kzmJrItm5wkvMiuTJokK+Wx6fWoDCl
eF7LwFXwAgReeN/APij3UaDsz6aVKGr8gDg8X++KW3txVYGg+cuJJYNAP/YkfZns
uNwKri8IBs1PMYhzrjxkui9Y9iadp/1dNVFZYJJ6rqUrOu+t+pDF3p6B4rubegTX
9ytSwyFtYq6Dz+ulmte8ATCymKKZ92Rgzhwl2l1rnjsWRN1achgHVSkoISeaUP8/
g2OEeG2NGB9qCQg+B+wo7X/BneddnvAhNY4DXKrMP8Gh96eFl+fBvFA/m+vbx5Rm
Vl77SY2FUD7moulV7x9eyHLyIELKmT7FG4cSbrnch1M2P6FfA4X0pPnL+pogeZUV
clNprAL8aY/86VENbcDeV0gvqBiza/bUnrKe/0if0Qnraf81JZI0z3hmCCn3xRMa
opBN0sxmQvEDvfcvN3LXSiDIY7WQE6Rp4Wlxmo9i6lVsSVM7SDznu2PInYV7cHk1
utnScvkCQ+c9fbK8PFxRBxIGeZuotrFtp/gbimk+F4pR7te4gwnq0cWRu+VkxiJy
NGqgtVvASamHwUmjO6wVQNpjJejtTj02scDJ1PqpoFz404Y0vqJ/Qh6F11FqyeTk
NcALNZtIgURhFiaHfovMDO1aNN91YROS0JeNJV/1QdS08pHIBV3pCCu7dQmkvZIT
02Cws/Zw4Cx59njcyFTK103b8Xj6OcVcgL4fiTs/6sri7ERyqQyegm6MdA8i/bgb
RHavXqatA8Z5AkvxR0EXmwOdBDmqTOwcujJyyR85dE943AOAKWKsTt4Yf89/nKcy
mGVkJGVf420pc3BKWl35XU6Hd/IE1ln93qg4D6mbg9y46gkGpYRbivsFknxyocIi
7l/BkTGlZ3/PPUHEYRPXgQxNFgimag1T+qB54yZXy7QUnaJsl42urYvJrQ8l+NAx
YNhVzy5gA/vC0CBzydtB9iYqTwt1t73yZGwPx+0Kvf2mSaqnrOif8o1vgQXrMrIn
HVD8Q/VZtt8a+vUT5FiQKUcwN5nAoF45WnnPuXYUTzWjPGLV6WNrFseuDnZgy1up
c+8aqJsGyLusQAg2Becc0aDP5y+kTUas0/do7qR4yGBLAqlg/wDSDsGglzfc+m0C
zZlqhTnAHFeVVXH9MXbOKux+/dKx7zMCY7puYiCgRPGkKnwj3z9EvKBA6g57YoIU
wCHJ4m9yv4xIc9bTd/fypz3UaITANI0E99iGraiC4JCyIU5pB+Mb/eup8GQATtto
0/UQZS0N1Gx1sxS+ubYwXGyABzTku6z+hnoEV98KwT2tpzMnNhNE/cacYyfqqQ5D
0rfQ6VP7qXvmrHVP++JxAgUq7JiUHsRUYj1+zed/UThcVMUZowdhQEM1KfGlj+Hq
FfJQUJdFNNTvD83cZS1VgloctFXWUu0SuKxF0SyCkgGAmrE5iG22LUTLzPsiHROT
2B4/Xdt134MRag6vNPoUbDJv92wN2ImDpKUkKwDbvt3ACudGwtjYnHR6l5GwKiHb
Bnpci8atxRA2KFs5mz3MP8jFe/HGGEtbwDvEuqo3yuRJPcmZ0XC/f0x7AxWorJXX
ViCsVj44z/BvpdSn/xOvroGLZ3ynaLXJ1CJN9YGb5J5XmSOqgvOG0Zk8iMW5cnir
sGVEyvd5eDkJ+nD0U4KIzSeHskPS+26lRmio8XDkFA8WNZ7FM0GckXUI3MX1cruC
abxD6bkUEPLTqdqncKWqWn9/FktTQ0OXJKv7DX2xBDOxwYuQ0TMTonFYTEoyW3iJ
Vzvh2nQ2gtCgK0RbJnrFCU6YA5wBcblRd7o1/LOth/Vl2x089Ye8qYjIUovn28Vy
Pg4loWQUXcy/SeK75WTD05WJ3ysdqRNujTuFXcidEcoWY16gu1z8d1cqODClwqfE
NYJ6I+u1F+zqXykkvCgD2Bam5cFApo9rRJEw2hAnLnn7AFRzGhwJ+Vq1WwgOsdMU
92qoF3F4hM0BdmGZORRbmtjr2UPJwLqtK7toouE5xA1SIPsWMQ0Wzv40K+XmBDb3
aLzpaXs72DMMRFnpG3He7gAzf4DUMw9RFank40TlAxG4NSCdb1ipSsz322qF7IZM
QpT8DcFaqnueAAlqQAwNXFD5sxBhyhGNey71fZ5tLL6CUB3aK1RPzOFKYA4xhst3
y+sOTCy5ibL3d/B/1SAOR3QvKWWKqA+GdgW+64cHZ6YKBVPvjkaZhwhv3HzoNAyD
+pu4thRafWtebnjzLgC74ooBV1n+8CyXWc37Lb9jGoELJCyiodssPMhDyxTzXclA
s1tiHk3SK+/4SAn9JxKC/WDW5LqVOtwB8n0YuDE3TDnKxp0BRQQLx5CRUK0jzQZw
c6QcGqImzeDBlWP8iYwTtye1O54D1BHemzVNSI/EpaQwsmGZ3bZZvEys/nssTiOT
PRXKcXrRPdsFijcIEv7/NB35dFuL/S1LcZCiRfNV8i+xb7jZDrMHwe/t7ivAlj++
hTqc3cWei7XySqLFNufisJYNRUOfzeP5dVuyZFS46AdSscHoJfyD5oS2B6lkT1v8
92F468UOQAi1v6FwBdsGHZztzV6D7l/BBcUgAa0GrIMUc/WvtIKd6Pygw0EIQJfU
CPCj4ORkuWbev4erinDlehURfIBxwn9g0ZRX+9I6qUW67R+sw1ZvVb83c9+GNltJ
SafGhvmD02KravFisJhmrw5itNWqgqW6Njd2gmyncjbs8+MgtrZNMspwamuStt2Z
cLmnYvlcnZT9SKkZ5qjK2YbM4ni/Hhg30r65wnKvcyNNY/juk1lhl6ZMCXx/udMV
53a8IHGj+WipoK9FHZ+d6QJnTtBfEy/Jy+2wSv0XybPYORoGNDm6OEolQKpyRSwq
AG0IMdnOcMmJF1UCXHAmLYbyWfluKJHVLSnSzlZ07ASXQuLRwV01tlVdbrtHVo18
jX/QZE86ggyvmD3dXuB1eLBt8EvunM4X60PvuvicthSXSdJ+lf5fr/SA9UkaeFxO
TRIgGisetPlCSfWMyUnGHWIalwLPLPJ5cWfxhE1UzeEqk+V4lkzNp7Mj30h6TYzX
Yt5G63E+5GMR0fDYQ3LNFE/SeIrp7OskG/uJIqhNH/PJ6mHgp9YjQA8gs3yJ6fmS
41TZr8s1EbrkaCcojnbPlHw0xujZabruOGsD7AXkhhoWN9rHB7m0Awt6ItuQ1zOe
b3CSSOjGJNpG0KfXOHx9Eti8INM6+6DaJVlySU8Kwo81nhvOljSwyK23ls4vTHsi
6/j2PB7c32WB+UkOdi5QO+lzUE8URx7geUr8esLv5JmYGnk/wuz2jCi/rAPHGOIX
b8Vt/fjga134D3jbtGdk7tdYYTgYiruhvk0hhmnSC8d+1rWmTXMbFX5t4u3mJleG
Ozr8dJUnJqCACoxfic98D+T4N5IbjEQL66K/1S8xva1/rCeKi58H3wamRKoHAB1f
cINDOjeyTjpnTt3U72swY6pmUlC8wAo2/Xll1vr2V+Oqt9lvmdet6xqM6PXpn/qo
wA+oPdby7JOmh60eZMWyUf8lbIT6Maw79x9ZvYq4ZCM38+ZgHSU0q4HGjGAE1nHM
AiK5NnAj5viPx+YtxApgPuKRF1wqI5ja/L8jRTumulLZ1Nr8VN4bVEyGoDV00r15
iQJC+OFdtdId2sT5OWDncpRDlT/krkCvz+8L8/SSpjHGHG6KH79hPINTHXgnFBlj
0BjymXH5FOuicBX4g/D4sICQ0rh3HJ2r/XBoWz8/yT/CpXVtOGbkJk43g76jdIVy
YQMRBf1GymNqhLiiJcI7W0gp2dARaokRGw/eD6kh98wQWBN/KSCwoig0nAtAH8Xa
DBSgxjT3P+//pn3xr0ewIXnd/3Bpr2lKLXRXwly/32P6VFfxXIlBZG9TIXZOMcjf
ZCwaE6h6NBEsbSK/SVLT/iS45/6/DkUa6sYeyr72OWw7mO3hVLEGvB0lJTgD8VXE
yDmMDySxwOuAOE8FKrPKoaEtKhG6dMr6AEzL2NKwyH7c/5MUDCCIKqepKU/QOVVX
7DKE7obxO8xzmfXHb2O0XzrxmQvCOyMtLBALK6Iy+X5DBMO4Nbz71jdjlwoJs5j/
HdElokm+vrsNAbzOFqbmR6uzTQ3nYwpUYmjYsTN5tGqrUjpSz7iGz2HtGdf9rjZv
0JChq4/xQvQ4jSb+Gs3cuSOJWLGOx3ukh328T1Ex8dxdFQBIGm2r47xVfwS7VYOD
s2yNxcI9g8afpzkWuKdvMzt5XN5IeW4wtrEFaT9mPfJC0J2IC+2CnF/uoknJ5kby
ASZxyLBsdeBwvCvbhkDt7w3RcmYtgY87j/3vJpSWDZ1PRtt56u6Z1riKGFFS47jk
0bTTDkAzQpgPz9ma0lVHaOxi7ipbEm9Qt8lIBwyVvxgAaH/8O/Y7LB5ql1sD2E8r
GO28lc8+osdVJ1r9s3ft7itm2hK3FRCHAT5dkbHFmw96dFlT768VTMiDdhH6YY7s
sSYL4I+P52VaSV6XgdsCS/fv5iPDvue/nR+BdeP2KE5P4C6tlDgw8qQjul63dpJE
wanSxyhgZJOESfdqVfG1O80sYae63tSV4rnjrP/elUeyIO4fC2JWZVxd1knd/fHr
x4C/aiYbsogMszkanjVsEmiWQ6zNxrzIBGld0Fbkw0uabha9EG65JmT+N/Wg5vPP
lH5NXX+xIOdKrBDMcb2KoVj+ZotMXvllmWFW734Y0g2Orl0VAe/bqMo7YTTTqCQI
GpjzI4uLaUJMxXX1i/SOAZ0iXnkATj2MgTwo3AQ58SMdkSTfrgj8km3w6bHB5zZ4
Ecd2saf7vy0hlhJWe0jBLKHBPnMJkvMSu40ValBxPaQCQScCfbSV9bmoM8B8LUhv
EVaHaE2uR/Bz0b9vKJWuOSc5lxfGfedxPtZCmhv4jIU9ybZY3PR0Gsw/ArG8FLcv
F2F4YUxD9S+yki8xYBh3BGunN1sb4RR9+cSGsN0tA+IRRYFdrRZSXAcoue2PPcbh
dsbYVTUMerIr9oZaj7k/ECr6369LKqMNLi/nvzWvkG5NouMevvjXg7NI308ytfGr
6rXZqpFyEWWAHnKmrGX/hkyQyXUUbQ+8qO5AnijtWgqbpdS1UOYsOI2nP+jbuyWm
VxWtjZkuNUvAxN0Rlc3T5iltlktgT0N/vb8a5JCM5g4fhmYAEioUH6Nlnm2uq+88
1JmU6IVgUE2g5knjUqU4z1PaUjKJJLg5DHio9kPJRi5TMOuzJUja8YzOcwDCV9K4
VEyGAZEizZqnqnEkvCAK3Uy5+pfEgUkPsackJ/md8xR0sgogkC2FO80JRNNbHD57
haxxXOfKEBd5UmkNY89IBBSLt4w+Q9/xVvY23IW9IxoIy9Rzy3HouEudMhMRzK+X
Tf9y2aHSIt77Y8FWKJJ82tWWB79JnCNQfx8GAkaUspKLZjVkIUwgJQqx5wp9RlBb
1VTJbdoO3IglcrlzI3rPxexXRfhjfK01irlIC8B/79X58xAQzC9KH6uQoo/7j3Se
9IylPU4CnoiwssYb88xKp95O6A5pYssYRMWHZtX21zdNYB8mnp8na/W55zoEgUU4
iKQeC5k01A84AHuJeod4tzaSIgIhC7flUKRmOB0aB2f607SiNDNZEmnn447jQ/bt
aJLyItPQzU5/T5xp/58mgUjnfQKVBrt5iL4ydkQIdUKb7PJuElBhLR2R/nM2hJ+p
zZrWuglHHIUzsV53pKhKs8vQNhzklefRpEOnMIrBhvhNxaEHACY/DNIcYxDa4lE3
zuiX4vr8UyZMDL+Rp0esZAQE7yAZoJDphq5zA84cLcu5rMIXV0Pj5s/anFdGbzwy
dbxtbL94jENcrA81vxvptguPMu1Q/+rK8TJ4k+wdV1ZrqbxGOGDRT1x2fQLYyJaO
Kj6HIEmq5xOk6cEldbr+LSxrcm9Mxbc8akGuUxIahxg7CuEsHLnzATl1ke7GEbEl
nwUiLkAxedJGZq9acHjCiI4ETeODDkVRECSpSMftBMLBoxd9Gch+7GqrqX+PtJTf
wQ9SqI29kqNbJfs7PSMqCwyE819XV7JdicciSd/kkKwyDLcHgv/r4XVttoHeRzNW
LqUlq7jB9owYLWDHLlxIaRE/64GLLI3lMLRasmTo/nGgu8cLEqVnh2JpXOw2u35t
fiQpskVkPM0gwUMFM+OBC2Occ8x4OpCP1nUanty84uIIadNZRVrA9KGjWr0wkipe
GHjOshS5F19j8xmMg9RFy3IufyFj0UFPLYjoPWTCkBCm32K0R52ErZW4s9TOfRUG
VONfGWb56Z6A+LLyU7pLy4CPu718/O/67nydtMCGJlT/2CGWbe6LfmO4POtGpVTl
MOBEirSWSBACeZgAkYPBH8f+jXkyHfvT+2oQgxHjeAGq9ig3370MvYC8RZ3WLgpe
8zFaLhvbNQLZT19X2AUpx6Lv0LFrbJ/0ATIseobdUDGmd8e/mCJ1T4p7VuB84Uh7
sWAJlmtC72TbsH2YJw48mSQFoO+aj0gsjAdDkRc2HuoscAPA6ntJPNQAj0kWPxrH
JjPQ4Km3umbA3o+kPqtBe0Yj8vN1iKA56JcJFdZbZ8R90rElVlu7tdXmelPTGF4i
Q7tYlLN4HUZi9HBGfep7b682j+FZQP29zWkFYXOccn+DwP0uWz43GEtVWQmVR2Qd
2hdTZcoHAC6Ew4rOG9Y4zZPMznok5eVjtI/XGh/5nrKLbOD/TS13dDdXKxP954B1
G7Sr2ag0p3aicULEfuoIw8pdb8PzltDUspL2H8Fc92g9dAYGBVOsfTJ1TcU5zhmv
Phwr3JDZwInmGytyTC+GttnJNl0J1ojs+OAhW6tlB5JywGXW51W8MriPAgq9UuTw
DjxjbG8VEs3h42hz7neqDtUM2H91mzrMQIo5YQYvbo9jsBkrO+NjJZ8AinigZFxh
GjGzvqzg5W6O/n1cYuB5efcNiMXP7aa8KsAZBhqOF5YL7d64H7o0VEh5OM+sOj9T
p8jlqGKCpnUv1lY1f8mMWn9l/egeaRtd62RnWL+TzZ4qULUAOPZrHe8AOWQrBnV4
AzCbFKmYEq0n91wr3/dgmj63ljP+yJnmwcrAytMJau0LCNCeWpFMVwhaOQbmONrs
s/41g1B6D+DVdc/c+puHUM7n8YpB19ilF7B1yt13zlqa09xMsoTwR7PO5vh5cMDF
Mmpm3AbVBUzoX2FlPoH1i60LFrJ8sE7EUW//uSzJ4bRAi+njk+CQyGktoo06zQ+M
i4AEw/sHDIFUjdxpQbfhB5wikaMgs45LNsBlWFU6ocwGvx+Mf1waS92lOgViooMe
ECu2eqs0ztWLVkBMmIhxhQAi/fgqOp4SfrTaW7es2SQD9Z6OXH8cdjP15ksqkFie
x9QkUYuiAX6Egofp1lN+QzfcymaorEOrmNx/5Eyk3zlCfs8dcpvoYDkClDyWj+8N
IsHI/Vl/sIkSyI5XgoPtbV3J7pzbHJCq94+rwNs3HHR4CjviaPiAG4gcdnnaFDD5
ngVzjSpxNQ6Pk6D5t6dkiFY3/j80j6Ue0rj25VWPQBSalfHilQ6/qeFD21EDScSU
U2ZFZA37Dxz9pqzGf4r6aZs/K2zXCRHxFdgeZ0EcWOzRw6kgltyJzFdnmyxFWo72
3ZtZUMu20RjiYiiSBEcJ40lipjPsqA3o/5hg6kcwogBV6bMAH7JeUVPBKJRbrr5o
HTfPM7sZib7es7fLhtHhpHz2uEdFACUjIJ5mCHNMrfQ4yuExbfM6eIsGsnBKdrHd
ARqjRyHS2mvurZn1RoN7FnkHDi1gY/hU9EUb7Pm+FcMjW0p3ESE6aBRDxfPmmkRA
Ja3yBBTyAjxRL8z5uWd59xNypudU2XN6+0E5b1DjAXLyrQIeFp/rpnKCCSXOuDjv
pv3/ScK644gWGdlEnDbEPqJZJTWkDat1CTWbGD0eHmtsCIB7GIEzkqNdnOhusmZj
ofbLPUFx4W8QOua5QBJpwLmtQ7liH2bhRGoUyNK7HvO8aXNrOsQDCQLmAiAt1M+s
9KY2dnzyBakbUoWlEVWTdP6n4VaI9pfXmF44SL33Ax5XtV8uQNRZKKHcY2pyh58i
/FwVmwj1qIuSje+MIVOlNYc7AjjfUNqO8fBpbq4pV8+wqRtSs82hkiQ2PPCnfDu/
g9THFSUvf/6HFpiwFXb1/cqdWv5SqE32KmscDqbUohR2vtnJ3ytfK/PSg7hBwd9I
mtYkegIMP4d8k99bwTBhmjy0UpBEOFtblzNn/SpojfC7V+f5vdye6scByw09o1w4
pvzpn6oOptlL4gfCckAaD9eEInsq1NLG03lK2mWEWbKvJ1up7UXpofvQaY17fIgS
+5vUdd9fBjXTL0HW/L+UhefnJK8S9B8pMK/9IQBDZ0ZBB5q+sAZyM75gVhRQNTRl
YydRmjMyjt7DsTJMMFHSZ3gqNqNOwR6RrbOj69oywyplZHl4idAFd9XUDDRJ0gpO
WUYO5Gq2gqg/CPJY+px5XGmsSRC7HxVRsgKI5jmr3lRoIFdF1DLoL17u0VcXJ9Gn
P112Rx8pQVJ9KVCdUN+Ci7HZ2zLoXtW9zXanc0SRGCzOFaU2FQe3nS2FlibIPlmw
6mCBlAen1+EYlKFW00rrJVR/6M5MgfMex6D1D60nX1MMcumYB1Ja472XuHlvcdfI
EwAK04P9Ncyx0yt6PZlPgGSD/rLee6NbbnJTzcJEUSos8aiAJrRyqj7/7SMhieyr
5oD8AY+YuuPDUu3MCD0EHRVKidIvoaUVQfhBXK6c9JiPCQmPqzebO6MyjEVQaLmZ
RCW9hV87lydfuSBzxuoxZgYCAxNg5U75S0iAUd0OxsGqEnFWBbhP2i1slEYILSCT
hKzPZRxegNDsOKpTcfmmPH/N8qfhccaNn8dtQ5fli/lfftlT5Km3dAFMjw3Y/N+A
oMOaktSpW54lhdKxDIpERQcIZuIxKb+9Ai+h03n25pztfRiI5BxbseoeoORWoUdQ
zv8NRHDLIQxlX+i2nIVXXT6yVBKNZs3JnHOyRPMSnixgg96VhGAaFcMCzy3naUJU
F4pMGLP5dVQBtGZN0eg+8AIQVUganEoS0xpj+F5KjncOsSW/bcBHj6zdHZKBeMxF
zE5qyfp/t82BJPG/1d5HSceEu01r7fDPPR5Xo2zwRwUi+KbIelDLvakPr/GX3BWI
PATsiIyMa+WMAY/spksif+e3zkHDaNPttSS4lfWp5Gmf6+ucfx8O0ehm+lyWKK+R
llHy2t3o6mrMAfwrbHTJgg4NDUU8sRkgy470+aUdcIxtMqnERKeUHRPNLowrTGrW
3sEiagfYseAI5U2Fr6IaZMTD5wbvXSpJ98il9M7i7AwGl4AX/MNh01c/MlHV36Tl
zyHtvhlJtYupbJXpcqpDWUT3n3WBrN/D2NQyPqMSimKpVv3gyNJ7WC2b36Fibk8K
m6jSjdUooehs6u3E2gwIX7s8PyHvCoGb30RWTWo1M7aku7KId+BrzUs/YKf9Ra6K
fLtXPF6ePUyQI4moFWJcu7L/U7DWy7kzdGqldXA1MyNEQQvAGJKtiWiSqMTCk/O/
A18SimNyp0rPYAY3gpMO/c4MEIHy1NwYp2PQCZdqmDV79ds5CZ6qN6T77yROQxgs
0HtqW8NejI4rydHEyUUgS+6P2gKQ0ziINklqNzJ9JWOZXD7VqoyfzTgFD2B9bbyF
P9s0+cNPpQnhV980UDXkKB1zUi+lFSuqw6Pwo6Adk30XsDO1l/1MrKEonWy4pLCG
EAytsrYCae4IlW/K2arBmU73GFDMsEBgdIKCyU4+ijurL8iS0ndHGmwWFqbo8ffp
f5oTdwJROuIZU1yM/9gO4DtFwkyhrkMq0QUqd81Qndd7InwMZmkeszo3jAhi1a2s
Plvh+1Sr2rOkujmkqlCGS12ZkzaAk8dN+kSUCUkety1R9HZQtGictf657i3Cm0ks
YQoNdJ6JZtjPZDTOCEuCqC/CfNYfiGKeTyavi2WqakOIIQhLSFrQv8KKgCqmvHWZ
mEoarePMOvtu0Q3dM5Bo6OH/UdYhWn9YoN6bIypVg8fmtc+mfAeDpCKNT5t//CDv
gn5m6ZbHjAX4rxwIpMWEqpnXntHiPuvpZcgf3h3AymZik2rk33M5M0c4l2owHl/W
tkfdjqT5Ros08egzExnXdlIvnVSj4N2+kxSKLEv1RLoPahDn8PTUWg+RXTzsgCl2
KYsXkH6036RW7LCo0Cyl3YhJdazgafBhMMLPa41uib/RMjd97dpy9m/pPfyoD2mG
sucnuxHKj/uI/AEkNq7XrLpcH10NOSoh0XpbXV0mHrEGKJUJ1SMfuXG3mASBPriP
TiXfBu8RB/+UC3hIFdG8WGhvjSpD7622lnlontfj6IsGeZn/wRjtrSUUC3v1rkWr
pgWNdAZjyhrf34YgJmk9fjbqRFxg8gTcxKHehLmrtwlXxGX+gjzmwtH7iAltK2fG
HWA0EveQL01HpY8aLNMi/n1qqwysLF2hvCkrs5sYIsI7UxKtYz41j7Wq8ieJRXn0
WpDKEA4IToCixb62t11sVrU8HXJS6ysXN/q/1D2B6ZBiehpsZX5wlVWDfexCK88X
QYPQRQgag77XWfYV9ieUO4eHj+HLg7M2yWJEaS4W5Kw7OSpynS2yTDswDzyChwwG
1vOruHMWmYeO/vE8RS5HbQLPB3LMP+XJSfInOK9ekKmHDT5ggK6pr4xnqYi6aDIC
uldz/6aYuaaSe9R4B8/M6FIKFdjYs6E9FFPv5L92i+BNl+vXBxr6RV5HqVkbjMKM
O6onHUVHohjgfYPQfDjcxxy3pZ34ajBNWjTL4iFQWoIRe2TD/5FU3zTH+8tg9YhV
GTv3KmaeSoCEbj5/xdMn4QX8LeOfb2zQNcgqrBeJylO9A2StB34SRphsZVze280u
RY75Ewa84Cvh+qxFUt7ZcDy/4XZ1hm/eBsofBVL3A0s9YiPUy8xg1OThi12EWTE/
pnV8iThiD7gQBSoTJsDNz9KOodOJzySWqmM3iD/1KUTIpCQ2YMSvbdxFfFQLRXaC
0w4qsnzvObEh4/tvyTGiJkrccs/jji0LzYxXbKRHkqrjgVQwZyn9G/qwvvks0ML9
LkXJWAjrQeTNHHD+QqmabB0w1oP9WPwIK61hheAwkfJiaOlbw0gS5juj5xOCjPVW
cUu8PeULtSLAfNtVKBkfRWVTDRk62o8Qzsw+cGbK/9KBouCX0nQSqu8Y1mMQQhcM
eNHq0/F71PQRBbB28BjTMFoeyxqSRhTGCIHrbzP9Xs7/WFr3HdZyfqPRIU/ptjsP
pwX81uwPWEDn39z4Ckt+ygX/HnOqphtGqxgGZJqAetjC4Tbr7PxCRf96glGJ+GMN
J8Ife5PxMq3aktlCperle+VPziNlCqjgGciRx0bd8h2CEhKwGmtO/O+YVdPSx8jj
xbAo2k7TB2CmSDj2e7kETHGJjKcHofdrU97a1XdvE/mBZnbD5bCwLm/l+REpBFS2
4Eai+TEDar/yBGm6Pz6XzzhHhmBuksNFFgzn7DCrnMtAymV2XEMpTBLe2MZwRpDr
Jkhr4QelpeNtnZSmBBOpxCM1wtPGCYbeiww7njOZ4pUs/RfUDF7XF3fxHfYu9iCQ
z/mHnSv6JellgMclWGSB5nLlJHWu94grMzKa47VjhcwPupXDiTjJaknlTe0gPvrh
hfRPYvPvd2kk8fM8A+WZpUktPvpVLn/StGptU+lrXQW27YKKpx4mBO+Z6OY/b+Rp
BDq8/vCl5GFsHZpw1g8hWg0Yom/fLvmXbzWFwWk5k7EeQCRr7THlewEoDfon8GSu
aYM+op02o7JAGVfm5l59edTTgVzyWbLLa3IChMDApP8KCBGSmS+QNTNPk/NFYPMP
vn84DpvMYch5SmYJtZDbJ9f1Qx8UKTSyzV4o5iP/PZUI1xHIpkmL89dXrSHbPOep
VDgvBNrNRU5u6Xo8JxlwzwPDMC7GwXhqZzZD97wyz4mjzSU8nldbvncGGcLVuxxw
LC/5RAyq5lc0jxVAZ55r61Qbqmo5rheE91L5NuOpc8Or2O3lyaX/H54pL2nAO7qj
/QVCcIK4rp88AbV9p2C1I/LFVTa4WJAzj/i4E0aYuS1Y48t5U5YhbQ2LE8R5GTU5
rCu1hEbrZOho8/74zEKIg59uID72hQgj4vBAIj8tCCjStBJXFWLPLFMQdHw4xTEF
0uJ5bM2k779RHf/MnE1PcE+snvmEYpCCtBDrtwcaboSnlLBLaqG50NzrtwAxfNZr
wqgkMT1fF6eKTV736Aw5DaivIcZRBMJCfkUc9aYmZ9u3bXQd97uySjC76dErA+Tk
2yOEYn03qyj7Fwe9S2MYlZ7e7WgrfxxIN7y1eT5SObr8IUtPCM6bs1zMtFqZLy3+
+82c0eyWcjh3xQ6LDO+PEYKgCiDkqSB1gTwO7LlQ9H2qsXGANwJSsytdVI2geZt3
b4r6qWemfGDBIw3HPfgI6wuLPWsXo04NM5TnvEt4Gano/iKVSjaT/QFceDo0jYff
FnH1niJa+ATNa6hcUREqCpHNB/3SNjQhh0bL+Hjjzja9VYoNFrLTsBDKFwXDo7N1
/7+8zoQWCEG2PTk12qApuG+MSETh/yLDHbpUwoIUyBkOVUtgPL+FP/M08K4GHE9V
WG+FdwtDFqkTLa8TEcTW8P1C3VvbgAcODegvf1WS4iME+BIl+kW4dimI5zQ8B59+
TNYch3zN5S1wKd6q8CnIvC6Y0mf1RY3uwnZ3tWDTtz3iZPneKCT/T6frE/quffyR
MJcmZt84WB0+hQeoDj2hLwQve/0f/woPtpODFEhTl40FJ1FsWacYvzHZTtCQwX4g
CsWl2pEkT7TSHdSqeFuX8cWzDhVKAZrgOtC9b2+HJY4r2PRd0Gc+t85/4j/F49IP
4LH2fe5seMOXGLOcgU3+oZYCa3s1TeXhL5u/6Otmqe12W84rEXmiTzf+3yaOXMbz
AAC0oTO8e9SCU77GEOsyiw+Q2HuXo03YT9+axE+Y78d+Lpb1InT0OaJCObEzdVbH
7l+aC77d+GbNkNJW6K2c7T6iSxf9obQuihPCaZWKQ+HSP9cgf4aP3wNLhviRkbCg
b3Kp92kwsPD/Q2v+LPXJFTZxvj9WuF081xi9qay0YnfZ7IEDp54ZHJ/uWLveXwqT
9vc4EeikZJUr+U5dxtFOrc+U9GG0uoanKZO3lpT/AsGS+MN7T768PkN1Phu1ySZa
Z9Fzx/anXWGOdYJOH1SsWIlW9ZqJSg/SNLmjintouju1eoj4ArszQFXRUb+zgSCI
Oqjfzyvum98R9O+pxTwChEBPQ340nhWMe8yswIDceoLxa7ivaYuZ4ra5FZUS11Vc
6AI/JHnCv58LnoGwkQcjjifyvhOLdwQnfuw08pHAnFsst/7YjZN4IHYrhAyE+QAn
aoHGw3jE/C2Ml3B6sTdp3JsHtMukqg4KKr00jKh1ah8P3f9T7F/OSnAD5TIhRrfG
BWm+dJGRsQC+ooMdX4kpWDx20jDXh/sc/LYSDJRb5mx9LodoYnD9JZQQDpMBZGIX
QdQzCdotivCJDFJQONl1RtFZENH1A0e51MyTutuFy12CurQwOjqVCSQAUmXxcrEe
rq3ar1DaaDmKNu19yG6iwbjDxoTI2oV5yGChxNhcF/S4Hs2/4zqgl+pqbb/IvPTZ
iejFwzQfovXuJYjesF+6OHT2fAUPwhAgv0WFf+yuZlLO1Yk1QXIXWzN7iq81wZr9
4eJveWOpIKQL8WfScNjhoN91QgYPyBzLf9z2sqK3WDJoFENEZbFC5oGXKCx8B4oD
rmzpfDCIksbdDB390gLh6kqzi+ziIkYtHR/PU9GuRR7KjHOXxjaYc5mcFeqKbae1
hZgY1veux/ySnZRjpu9BWLL4cnvDF8lTtb/DV+1b+s01lInLEvJDgHXEaXp+fNlN
fYFGxnD1YdySoikrQIF367qhkvpmhqanGpdmrWZBTT2V2RlwlT4iSTVXhafIZFyG
XQZyiWJkwoNMl8Fk16dzL7nYZ26btGHe4MSKBLSVwS6HM/iiJg7IsMQRO1T9haz2
hxkd0cPtL7T0FoKMKC9ef0EqalgxoxxZmRsZqCT284EeBqnLH+VDpMP9RT2tjUzT
E0lhLLwW68OPmsR0z46+T4AiUrZjTPkp/Ueqa/pCjdIwnfKoCCTGet5xUlbBxN7/
Qf7+SYAZjimp8NoYN7ABcDmJUKyBO+opWvf0Qd6dGkjwWkG4dN8xNDhuNEYfkH9i
TAf7sO2bP105pek0fS5/24PbhgbOdSXH0HoB9i5r2RAvUj9t3Gb1Mvm2kC+4Tnal
+JOzDGNzl6Pu1mXO35t9707yARZ6K+r4bfszfKBdhdkr5yv7VNt3uA409mmAkX7s
IopWMzuI2IoEf5wAvM5D7o9m9r3cpp5jD/H15BQX8O08azThWXkStOUM5s2ugHSY
sZciEqSArEURbDVjlDvlm96oOecbqwft1GqgiCNa/9quUjhwH0t9uRjpsoiOOHux
ghc58Vi1NGa+08ZpH9LUs+Dy7qmAPRkv2EeNbH0+cDki0z4V1Y2gCH+9CkBNRBDl
We1Y9srTIHhoyJHpmXtRDgtUnPTEq+J9sHqXl+DysXNlLRFGNt1cjPCz9tVAD+Qw
ZvB94NGgEv+N4lAr3Kj9bya8k/p863TPKwZ3PAzOVhaY2J4VCgdqEBn9BLdatZTp
eOU4J5g5nxEUgV8uq7JWF5xnheOTmIdVFt0e2nehFrAmEIApQtBNaFi/lMwm/Gvt
Nn8VPEU4LxUPyyefTbbc6ucZjXsiztIs3/nlj/sYeQ3EOnsx2Qydb/POe3SVtWzW
qf89ezZmcEWvQ8KkY9FkFUghhAiW6M43B1y+IOtEcOHx9BZH3ylwgXT42zjz2fk+
SBrZS/0C9R5eY0qgPYBKQl8/0L66Rg1crMEd7kLAJji5jFgzNYs7xEszN7b9POoF
QN7ChMCKNhDprVMafRLwDgw7paY5UQF3t4s8vVglDZCtibEbNRDbFyv12jWMOY0j
T92l9xZovaXpZkJBWiPRJmD9lEWpSe71hUnTT2SlmypEEHzkiLFf4qKhyTv4FMra
GyCRgRRKqZPn2dEHLERzXEzOs1bhxfmvw0tqgbuMhGRg39ZXK75Dt2kmRMYJztc1
op8nSGpMNAczFEuzaE1qeS3kM8v2Sfa/Xh2+hW4RVLzgulruNo2zsbxLcE0X+z1L
rsRt6lGadSnOQyewfQiWwFq47HDjFBUd41Jq8c46sEjhZTbgVrs68t3xIYaR1yo0
Xl+ZYrIvT1QW9B5jrHFxy8wey0O8ugyXwy0neYLLWMLi9o27cHMGYbLFaK38KP0W
pFP3ITuDIpTNNlLILBfxCAntJGU5YpEz58U+qZknsGE0MQThEqP9dHY24ixgVC8K
3ISAfz4SCodLBuEXtE7Bgp4EKOzUgpx3DcPwdQdxPF9+5gFqOJR2FhXUasK8IUlJ
M83lu73j8dGGwPkLyPu12Ngh9DPvwgnFZodQ5oMImSH/SYref3JznakUvqeaIGkU
RiHtEcYCHxNmoMg+CWcpZPVRS4FIMmLWSb1oeynGgu90Ppwmcyq2OdrXZgZmR/rl
uLd1neLTYdZneMIJ6dbsFG72R65D596Dj9HshCRU+Geof7tl440TabNCB6PdXkVD
Auq1aK9Rw6ncyfzrjG99MhZSI48QsUVpcAhMe39uHh5vm3UvQi4UuHiY7jlLNpzP
C6oMIKtoxhb49wNKFyxrZx7x4CddUFZoecXP/uvCNg4f5z9RzUqpvJ0bcdL6zsfQ
W5WUr+TvoV/ZLjY1PegReaZmtyKu0fF7I5l/DLastLcYl6GLibVrLQnYONH3f99Y
yks7pGAijRMJQxN8DKbu5KpnjIh3D63C97w4k1i9gc/eJ+kmvL1uaq7GLwXmVzDX
zMeU2LWq+uW/ll4k9DfUprhlUtxqG5lIj+NwbqrmgOO1hTuUEE1GZcIY2Q9DxK5o
WPvQ6obBmIhm40FAdb05KoOEbEEWC9G9y6506dpnesGu5imRXQE+rNfofLkFEBc7
LtJFRI7FnrR72iSBU3i/JK8RtgquHtLPCvJVuFDazjnpnmjr+zFaVy4r5SeJHU3I
t9bTE+MQtNEbClSVpXVCuMJEUpBgMeAlycafKa+n0SBvIz78KEnGS2gcN93miEQT
fJ5fM7n6rPxjJ6xxc+b9ugp6gi0SH3zQxcmdPFrHkARV1tfciyJJg6bjuRT5RGZv
FexMhChlbdRsxLfI83NPpFKEHgG71SBzj9t+qD1OqWzcEtlRaNXGPdVzb0+x5VLn
FLNjp5Dgu66YZHiEiy5pfVne1ZNae2o+p6FIzXfsEmkRddYnnxiLhKwV8Cv5x7P6
wQs8Vj/WdZ+V5BHOZrtwC6OJhxq6o8uxzwtpCDlFKDbZI/SxfBlJVygXgcAnBOJm
y6ljU3s/7BIO91oYYiM7EQZAAgPHVVGAniz7vXEoBN7t7Q8sYqFgARh+q7IJ7BvD
L6oaSQkonAJXdCcn8jFiza2h7Lp27KiQ5BiFLR2ktP+ek9RCyrYU/nUfGeCdr6vn
DNWLnPIp0kzhDs25G491QVwavZ0tmQ+x4/GE4ozQNWhvYAYMvyNBV+gp5QSCkOYQ
y7grhsau595UwFfzqjrsgdS659p9f9GsqzoYtZPFpK0rqDNXpGSvM4tkDlGZP8/6
LkpAyrEAk+yDnl+LlUxPwZeCMUniL5vXyPtP5pUQuOrPskcZ1UmpOxeXeXnxwNry
UMZx9uqhofeMW9r6L/eE2de/slo68inbq4pfXuCZNBrEmAn90WMm8fiAW/0CUlfC
bnm+yi/ILwsexUlfRqdg+NDWI2A3kCupeuejGwpw+ZmhrgmoFf4HnPj5NvuhlFC9
wgvVZpJPABa0Nzg9j9vfIyzfaP2AEE8uOPbP0V3T18WoLBQBSvk0sDbUJswNCTwu
PDOm7tWfCYtUnk7k4YMOGlxfDc2vt9IJGSD1FAkvJAOKdlnRtf69nt5FFD62J3lr
70K2YX2No8iop7385C3oWtOp9SjhN0RgSVZ59AUmnv0Xb34XXXxahe44ZERLWpdU
MWho6Tewro21UsSOOFotsjjVvtKXeXazTKaO58P9UjmoBi2iLPGKblt7dih7LAld
3xYuNOzrzj8ZAcBcyDU5e25XlpKSbwTCE7kwJAqubno+EBHYJwxSWV4uuUC00f4W
BuDRzNXIHCyHJ1AafQIOVLXeJoug83Cs8wZ9zsvSXGu5V9oy3WEAxOFe/HRB8dBr
Ez2xcdmGmTVGdZFTSbPfUGfNutX1A9q1uniVP7RJhFChttdqVdce7Q1VR3ufrsXt
mTLMggjZUtx+WZIL0nemEM1yxTjM8Wz9MQBx+0oGS2F0rzKfmh93aFtvCIpnscWC
BMEjDqt2Y7A68R7I4zMc8sFa6hkI/KOSXmejreFBprH7bYBkudXFbCNPkvNMgAbu
7fbgFlUChmJvgSG/f5tYOUZwu0izui+7C2e1bx35aVp8QgOmYMP1vbIYeBKHzztV
9mYGBdn2oMrqi9IfAhWNSkRz21pCpRTbTyg24ehtmYAJbrSOTPgBm4c7wuCLOrw7
6eA4fNYXklbnw+i1XhG7M9FMOTLOXoM/2Ql2CdIgY6xB0day9UCbhZacEtaR3R8d
Z0cAyTRNjgSCDA4tiqyKN+gDZrNw+2KocEMEw2VLAvSrO3C35Rr42HOuHfC8JA27
FfJwDuFS/fAlTW76KITjoWxq1sr77N7huLYpzGT2a9XT8olTCDpoV7VZ5k2GLLq1
14VGzfn88ReJCOTemP16aYrMBY0s9mwqHpq+JQX4cfWJnB85ZZn5hz9iSW9yCxUF
u1HfJpdJ92jtuYCZRyg5xsR/oo0jGqXT6Up3F35WJluR7B9SJSVQEKVuQERqcH77
Jc1JLjtCxZGAykivD8jMIztF7K3/lmO2h90B1nzSA5I2arobGUBorKKUiGidJYgj
td2RVArc68iWHQX+TC4TOg5MwbXTRLOI4Wltpao6Fs+Mt+9NwSxgHzo/5KYi/Vul
bNsfw7tjxVOkWhnK4/yCicYuKS8WHXlcxSBSRpRCQZZ16ps8l6xJdfrmPW7eQk2p
e/wnEKQPYtf3dmUC4G7ThZeHJuOd/4+RVR6DHuafuqyLSXYv216yDyaPlOdK4Xuc
S6i58DGlyqJY5cSmbrSHIRahGXCfZlhQVzG2fEIVFcZ3Qn74MBi3ZZnKbJqt1o26
DHDK1wyhd8aImVUDH2MGdJOIKLTaZpr5UK3ZKf+Wi6QNB+WWpCH0tPFv4pPcxLjf
ZfgCG6yl0b+qOXcLn4ywrHPTjIOHw7PxBAOryvxdJbNIQ87GrOUMKEbIUWodF3DR
PEqpdsWu427YPeK5ztnbZHPADXliuLmUmHPV6jOx19W3p8WouGImGFzsPcRF9zSL
Sf9TLMUL4dM40DLD+mMux/fE6JIHWlUHWR/Bf8MMxX0eLHCsVm5/JPnbw2OGsJBm
vBpXffMWp6pi5FYwbXKok5raapzsjwPSJL8PXZOihzCAVsRqqIHpCIpSZ5oOLnbD
vUe2oGo6Xs3LvF8Rv/VpyOj5Db22GZbwI+zs8c4aEIICJ6It1BXoLgYRdZCarkkx
7D0Be0bHoYA3lf/80E8axW9Z7lfUTriZKKL8fu5aOXXdfcLTiaZ4FXvgQfuK2Qgs
cL87GUEE5iYSt9RbKcVXJTh/7D9NR3dT+R2Fx96/zl+HTBaVEgPDS+UBege6ChF7
MwClnf42XKjLoTy0EYgH8ZhsqVhGv/o6suce7EkDCQYKyiAWdmuO4UFx8pP+M01I
y9sgCfiJGgPsjgXD4oebr5usP+JBKBLezklMS62JEztVjDc3HgCGPy4SK4uzPKI+
t06YXlz38sMQoGUQ1Cy+z05NX06dl/p+Qup2d8mTbokLk7za2ZzPYVbGewtV9GVm
UACARWYbh7h5/2cM+og0AMiJNGPd3RuEXiyueUuto2Vpn/mc+6shtQsYnyJ+cvIg
f5fFGtfuEEslf6cgqdv9b1oYI2x+6S5Km/DIby0dKLAU3+yabu1hRp0w7IhToLQ1
4RLMfpmpSTBjz2xWhPRuTlX7rDtpk20/MDSIgtqNuF2rf/++2dZ0l71DPiW1Hzm5
yH1u0ZBimXgyhiXH2yS/7jkmL3BS7Z39N5lc058x9VUObXkc504bZleeNaroBdmQ
jY6y7dfPBiMjcVmt7v0J+vBrKQlgWvxQTTdawB17xlMve73r6s4r0NHFibcsoB1t
r3uT+y0CiYSYX0LNln/R1NEYIr8QLaBveRdcUAGP5rGi5Pe/gxfE655VLCEJszt+
1bMidJpdX5wCNabj4W9HddNmP2iji0xqcI+CUyKSfOjSRoBd582w+xWVD7eCTMYD
32mVAR6oZXFwiTudKMGjL5sMmJim+Vb8869AEEL0i5y0uMUmPMrb/dGYX101OwNM
fPZy+dEEbdhD4BTiTUiEDGAJqhvMbVy4iXysXVdD6MeQP79g3veTBpcPEYVr4fkn
ck1Jl9WEpNBfbnqgQX3l0ABnOjsYQKOWvAUtqUINB/JCOuEcLVuVSjkJQJ3yTqd3
2Dv0ZuclOXW69+ey1KuXhGsZEU9xuOSedowD447O1MM6BwLoziPvrQwbp4c0agQ0
LLCpVAsUf8LKHMt+zZ4ogShyWiy7+1E9ZRK9ys1YSgFPV07jSde8M3WETrW3+bTV
smTaXvTcC/VUayBL1hHxl9L6uEv72eM7fcNd9x4RLl6QAUvZZo37BPrYVaHe4kUq
XBmkkFcUvWmiQ+Jticbuaaty6Ldwh07IxSlwtAUQ3INjtdXwy8dTCx8RZPmr0m2R
J+il2MHuqEXPrP9mFYEQuexX4Yid/EottvnZvLVb94GbxiyTi72YiWhwBwpuLiNC
CSQnIXo78Dz3USGAUEV1FYVa2y/ZjkCqxum5duFr9UzwE80r47fxunc6S7cbn81A
T1ACggvF0oXkwHiLTZf9qUO8B3eINI821nFwPoZbJENEPQIRSjbAzDZs+hlofB0U
+/mrzJ9Nv3g+1UqaPOeH0qr9Rh2Y+wFr0tNWHJfu19Cricv9jV79eMLUDC+AZT5d
fKopfndsLbouBm+BdmSdgJBi+nhu6mijVst1jsM0vm4BRuymNp9uQpbSlBBlQHMy
DHaFiwQnqRr63b5jiiHnfrjRC0SMvGHpVAWY+1WYmUJLaq00in8djn8zUngiW9t5
0i57SG+NsvCJm0Jk5x/EEy356rBkG/mtsk0F7qNl+YWDWCTPNIvsMLcg7Ko3xsJA
elZ5YIbbWzEZyv+rG0t+sCf6/kDO6BnFX3vKt8tjbc3B8mDks1mE7sWRylc8sBY7
89V8yTahZVw+ZJ7eP05g/aSbCFtpQQ+Dx7ehVDmtJ61zWSosd4zVcKX/xZlLpjbA
6ondUBzU5+bb3wjWCGtySpnex20YbadVUFq6WFXJ1S3c5ebc6Q71yqgznwkHXzpc
cidX5Uzhn6lat2p082ngpthCEs9bkMhQSx0L8LLHUJ0aFSwrDIdedA4NgghC95tG
ZPulZ6vlB6H6j7sXX7i5DbSCQoyc3QL5CVoDTVwANAzgVt/b9a+KcKIEwZPqoqgw
ZMv7GB8n3bWpHVPZPMCB6HrIrC0TvoR6bdhlTb3tqLsFbTT7CrMaNI2Hb5LXplqY
GtJpR0eqwyU2ld2q1nR5ReaHoCROZZbreiSSxhNlvgLb3Ifw4EaE8oOdsb7t4bxU
lwrZG1jGGgRz2wbANEMuQF7/mBEZLZ/07hHChN5kTTo542VJGetDskXNjdxRca0r
9Xk2EQJglAgUMtKXRCHjRAStp0bvoNVpg74ZfHlGDe+hcmM7DOUgL/5PMO6UzN+x
cIoAoEA5PHXDQYA2/NdIxGbDYJa3ejiATmmLWFvJztpPZ2IKxcSYLm5sndvGK5Ty
kZFvcM4qabqUwXlu7pvAZ49P56/3T8lLYkjmuNG1bc82sEL0AoIWSzOMNUwgkbn5
qIpVC+nmsKVA+8/Z4583lH4sA7dp9M+umxKg7XM3HfQzMpBhtDBW+GWd7Pouj2do
r/+qDj/85CGaECgNP+40KUSDDY6wZesFI2m7nZigz7It73+pOrqJGehvEQDgQXdu
26OettM1oUYBRmiamqPrkK+IQVftwy2c45YD/GFRDJob3h9GRemJtx73+m6o89Yo
2+qWGeOoi05OyxtXqa7IfcDVS/GkXZvJgSI9pjbmFiAnuzqgAvkzk4iFJj05u5Ol
3mr/DCktq5gZ+EO9fVppN3WB76fVDtQVEKpVToLE2w3yUM90awK44X+MVnNy9Psa
rNuHSed/S/fpgR4ZC/QgxAwilM1UOFyhewsBv7LAP/k4MJTw3AtQdf42JM9J6bU4
CvqEmis8yMUF9ojb5IXavbYRFLoddmhBypr5UnFevn31gThb4QKLQ0fcdH+w7l/X
L2rCTl731l/3UIvtOQFaO+UO9ThZYRoQ6uOl5V3VUKbMmbzJSIoul6+8AKHwsUHB
A+bYhCY5PoFvzHeHWnV7BFJpibQEfh6dPzvpR0IDb9rCtpN4tD94audJZLY+KBOj
82yMni07GNawi9zLHT2WNdzrK9P6QgnIoRNz8xAVZdoCAxFpaqwnH0y+Q7lu0wUu
YkaQG4SF3o3bXMFvHya/XyGE3QYMElAFBWWAKKFzbInMnSj5jAGlRp08a0wyo/oM
ulFNqUSkfg8ePFdVwht/0IGT34Y2T6m2FMjSlmaEX+y/9jQvLoSjvSMF7apocHn+
1jGMmDDB+qzC9wSaCQBD0sTOfKWy5aRfe2XAzAl8kFmtIOANzRcXaixr2KZDoc+U
IdmA8ikNxUa+JHyiTr+jknz/9NuFAckodjlIbWs+v/cY+GtTttulGHZEHhinbVcJ
WMgeFBDbJ6WaFNtSdlBgYZAsu5j8CuCWMNBsmtJbNBbFAvyH2PeaT1fIf+fFottP
p+S0FxE4qoxFHfTZTTdwhYIQu7as54083kEns2PZesum+XknBTEA9DPkiAaKbb1G
EH1MWC4p0O4Ag4bkLRhCM1oTVlGPcR/LDSdU2VsBpBpC0JDecYqvO/C/dAXjEN1W
6LFYH1RApfXbqnBNnepmF+GFjQcAUvG65I8jNTfcmr5AYn7bfXaAj7g74JwXUyC5
x+thPtjFfzsZ3yOfXYNh4V2uVasnfG/DbSLbVqmXeR+6UGqWN9yVAMRwjIFen3Ja
y/YhWOSGRoXsZTNEgf7wGNgROoi6KiwqgxZkgefNZmNB5TkS0RX/vmRY4c/T3cTv
aptQLnS7W3HPoTT1CDlje4F2tI2VRzt2HUtMwZ4p+oxkNUepSobo2ZIIZsHnZeOt
OHZdjdgutcDbI3g/eajBVbDMRMHKazDnSacltJVyrOKjTcmme0XXIlrtY2z9eeN/
43Ox/fTe4WAct8O0k8iifjWQvJp7KJTilADxy1NENLKymV4DsTpdZspSvKRIVBQR
C3IjS0Pla5qgIHEwH0Wl8HNeQcwRhDp3LEpZjYoYYbYIeQ8cBmY7zPAbZ8Mfi4cw
DWHD+q6gkCsjld904jGZ3BtdYMAiRatOHFsndF5y5jLIkODu4Sk8UpIuf/nE27kw
o6aqi3rZ9BKeIl+f+99GbxoeQR//xV67XWXEuQhu614TyOxzGmdhnXY36e/AfN50
AEqAQMPC9I2AJbZV3HpIn7csDhGS0yYEoYMBiN/vx3MAGPLIKDtq6YLiHQyA5ivL
u6quDk1M0z5FB7AJqnBrQoCEEYfw2fg0h+jnrrAUsejfk5w6FMcAA6nmW/cj2qFm
7zdqLzqOj06kW8Bik7z6cHFh9bJ7OTehBtUgN64vryyPPSkt6MdqIqxq7SxTOAVx
6GCw+MHQ5dfdWI23CFJkxjgOCQkCl7wyWqIXW4yHpSHV7z18lrgwzRnmL0hGTd3N
siXwyl8GNWipaw94QFCLfPDjEEWnLBNBmOYS2LLcK1RbeTwW97W5k4eBoluA5D0Y
Ttklw/hthKegBruq+ACVionPciBoudTueyNPTQFIF7AXSTm/k3noS+nLuDhIQfAf
5tet3j0/DyFCQrsgCkQjAUqPTMhpiu0r3uld1/NszuDhObSKyVYT9lBtjNwQLk2H
vxvPaPCLoC3xtAXh8glyVS1eHNLZhb2dCdhuaNnev6nCe+qmQXBWkftItzeB3P2y
Nf7bpa7NZNewowXsyiBcvW7mZGuCubMDcwMorvRdgYWG2nF/lJz2W8L6zlZZmujR
JNtOeoQOQ1BPnVmeuzhllxN7zL5RMvEqg027HzDkX4MPTMtibeE0OeEaziHNICC0
mXfQyDtfySoWJFSAwFGjX6bPE1uo8r2Zag6V/qbtb8wR1C/VPriIxd6jjQ96Df4W
CpIFo2xju+KSpWYCFL3H4rz9bJnV04yNKxwY+qzMxuzPia8IamF9FusKg53qkhdw
ZSUumpkf3JTnYx/FdctuQytd37xLq6dV06fcEvRgTnmvbBcLhmkZSYdIY2CfyohX
Avc+ft4oAK4pzb272V4GU/Y6QnctFmI/nqkz4SfJarE5uw4CAAIiiyMn7zc/dXDr
yIs6S2wjFBE39T9/lXjTVqBnCRmdvuZ+qnY3ctsw7yiKu2c7PX7vtNsUAeLaMM0v
O+YIz0hYOy5x5lwVE6OYf5odAXvqJLHg1/N86vNFHa8YYRJM76qEcQwDzqy30tOh
EhGUMEXsKwWCG5EO/Oo+EdKM8lHtBBaZk7O0ZSoUwdRoMnlNhXXx3yu1cp0i5Dhc
Fh3FRv70i0D8MClU9AuNdhIWEo2QnSb6eJTb9Sdf/H672acG1hm/FboV7BlMinB0
oUJ3xSPino5U/yGFSH256dICB2ocmPH78SBdVvgw+jcOyE0wD/dfCz/yKJSJeURS
D/7lUNVN4Pjn8dnOl19Tk1oScPPEELBAX51iRMkugkFy94VvpAOJU2bejHvIIocp
10ZLkGaKe8hyrPqVE8qoYt8YVk7dQ7qSr+P94ugqJeg4q5z+bfcKdMLzEzCVBy2N
tcL7AdcANS4QkpCBm+XlEwkq1GvEkZybKv5ZUOamexR+9vyKt97q8a0lHcjl3tLs
yIQPfT34XyHkZk9+GgOCsInrCqqF04CFNI/ThfZB8+8eylu4wPdtaBbSZlomxonm
e0hlaAQPShY14tsCBS3FmkSyYxmNLNyP0Jgdbs7rwsnx1NptdWbZsr39fCcHAzKJ
du951bqgX4oGtPmRi46/LC6lwC9TrNo0UP0Hwh51pT7/tMO023TRCx7i6uZQZD20
k3LKuXNUZr3Sq0zejAqTD+HmlJ04qiOJKTPPpH0Z2fUE9qdajy0CsNVRF/XtS4Pp
XrDt8lE12iTeWh43MDkDPY8MgF1Gt8XOBncka5cXGXnOQvptK66XSEWBPsEvbcPG
oIUfuRHrU+iwE7LBXkwetB0CAF3y6+2ijgRSAg1xj/KgZRACvj01wGvhQ6oN9ekH
aenW2EN558ZLmJs8UwfVqCDGAEgRqxFGYXs1I7jEX7frEGw5fZr4qMUPQvXMIErW
tYWB8n/KR31XNid1EUfgAShyrZHzAvtNCSZpmDfKbjrmftY1hX/e5d+CGTAUUMTF
wV4fb2kOErnpvzMTKyz4UNDSfD536P5NjiCc9X91cQ0eN1xqXKiyA3d/QC14vJxk
oXWIwrTFLz4DlHFQkQNesiMxL8u5AwZ+ultxKyAK70dcwNEW+yiSxloMce4XkOhZ
kwD5vgDo8727fPcF+5uuDopwQhCoVDJTHiS15AhH2eggG/eo/dyAWk9m9k8iRJe7
k7a+s8YNsW5Fa3WYV29ifOCb5PLmHJtlRpg9d5rIKUTi2+LFRLCDH/Bjtl4e6RPk
eRKEy8pu2jixoPWQizwIJYW4xVvu1zXW298/X52tB+YmR0xdd+Jg9jueAKxEzcw5
N0tmocHcQZ7HLAvLSgOf/GnIlxycJPIg9Hab2he7IPEjOjHsjewoTDM7nlNxGsDF
4bBKAFF5X8YSSxxm5j5yp6vjEv4xyCzZlWDHc54N7PX57qecfbJBpMdpnJnEGewT
OOUzODzlv9CF+S/cAqMcFqP4g7AEvZNMDT0SWh04P3ioG/f/K5PMJ05WGqraycFz
R+iJ3VVRJFbwsvsnK5ZlG4KTLbxT8XDTCpmiftOLiGaF/XW/Bq3f4qaTdq7HhNxa
P9Tku7lXE9veLLvTOBGOS462i0UhkSd9cJL7sv7sHb+RHAAGfDmGihBVgeET1beb
HEksZ2+93SkLeRS3RPgPY4zKTm+mhsSF9dZ2xIrrugWlm+Tf4sr0jFSBMoeTgDuu
G0OFrC5WAfgmHVkoncEkXZgUiszm6td5Dj4BYvOOQN1LswQ1K1BNHrk/9yociAJB
pagEcFBo4n2slmTHyQW5gKnEFXdEIdgQnMqBU05bEZDxGNq3I2h+8/plkC3U2m2x
3TP87fCcwkig3Z0c5legAJoeXc0TeDi5p/T3e0S6ZABRA9/akcdNjXeMeKxjEGXd
SWYSvaerCOYG97+Pk+cpwH1EwdabuK97snYzGyrV3PdN9oy9U4iwGB1Ud7NT4sss
+D68fhDPTVgDO1ka6wl1iOqROEgoHYN1bgpW6dCPjibOrHxDncVEhBj4SYHjMHpY
RmQ+O0XAhj7pC7QkI8Vjk7AfzHRtVVvaNg6pI9hi9Yfs8c9pWw37RuOiiatutw+y
SVYzV/Ngp+U+Qs0cebhEEOS74q4dYAzY4pVH79qVxodg6M5cDSL+8LRmtpXJSyKb
VY/h2ZsE3b8PbGogL+2sG7aammQVmW+8FiYxoRGRg2gPDtl2aUpDnkWWmkZWdIyz
w26uxxRZXwOgIGH5y/FfxJeNCAX8RYJpF1mAwltc4Ijh17uPh+vuNnae6EiR0t/V
ogKm2YyQUAHeSmZqFXfJYqvBJIXO9dPz579hiesQ5p1YuWwe1ae9kcT4hJKJiADX
aRhBcBVLhUsaYo7bafQdfdGADf0R1aGRHNli70AZAcP8vgOD7FRB4egETa0ByhKr
HBdyEG8JROZ06XxbDW7fZSoHIR63vorsDtZ15bxyQazFEl5kaYaUy84sv0QxOVH/
OnbOPLl0ZDa9yNadSWxKfuR1yjXyUYerZGvnFoNbOlnh7ChlzT9mR6r/FejQXAPB
gQx7yuRggtw4ivv3HAufCD5v/9CFx8OmfjjGdgMx45OPnUcFcKqetJJaH7GbjrZQ
CaAz7HT8GKeUC12KzV2Xb0L9gy7tJ6JkAosterXl8BX1cK2v0M9e2fnBaYNamfUM
+DLa+rbLesZZg3eSkUgRnVnxG7veHmXLD2l3WlEESsJHHwMQCdDos19ksY70iInG
WemZRycot4dduB9B5yotNpQNPqIkWPSHCzTurUxyUkW4zy4fPzdD9TZrSf2hk7b0
gWfqGpa6NpElfCt9RLbareng35bkhUlfm7UFZ+VkdbfSLpmKDsyK8kIrpfS/Kkxx
IFZ1XDL+NlGU8KIAoDt9CEi3hmkvlYb8e5uhKEWrMUdyltkxo++PNxkyAlXa0NpD
OSBDDnooW5igKwtfPnsRdcqqT0F1Caluyo57Q27iuCwIyS9NGtm9/NQT6KUTDvcv
V5hYwP0LIHpb/EgXoq7w2CyMCeNvIaipAha0W7af1wAcPlJUV1kTQcgrrH6wenbB
4lDd6bByESjbjtULbfRJkcswemNgTREFIEPqbkDigbhWbbqqz0ahBsDPnNijcas2
86KDm+JErjzfU12S69jwdmKKFKkOOQU+heRseWtRM248tDJL1JckX91WY8ipS3PL
HuPJ/iKNWycG5jxk+Wh3t9gemtsmboyfIAAZxPoQUvYSacOxbavck6xyBZQSXISl
9+/e6Tsuy1tyaPDAooxLl9NE2CQcdsufW7ZrD0tiQFrPtsWYyVndjGpTOXBNAVcw
GxiNemVUk3QtVupGlJ9tu/mQLcWHeICE8plkarXl2MtRGNnjDWWXvnJVGRmheLPo
mZgtAL7mj1j+HSc8QlXbz/5WWYivEYJPOmXdXKer295StO8Es6Vk3UBFoK+HfjJs
5SU4lnhi+p608MgVzmLKDpxYwd8llKkpmWsXtSn96NRguulusVa5X8sZb3q02LKt
Okk113xI6KmYxb0Ae25dFFdCoCRf3X/Bel4tMr7ndpYfo4FiYRiYJsNyGEfqeaTy
l3Z9wWdVqI8YAuGbt4duHQBNJyZP4c8CUhL9yp5OcliwxPlRt7E/4XE6RGIjHmI2
bBM1ffze10ipLJLejYZXPCX8V7YxQSfdSS1/lUGMMoeilcBDhNPKcP5IKQR2L4gI
a7X2EoSHgOmBvmR+ndGCkrbfvV2oDChyn0rH32ZRejxjzAOHNmHXKFYx+a1TBgoi
xQPkgt+e/fW6sZYMwjOT4J9eZspN14p6yIvptI8uC0c1VWbK3eitYINH4iUBJtnF
YkuQto41g16biU578ntsof5JCfAkipsVLuXhcKryeTM9pVqZcfcN3ucx83i6tW/b
gc5FEW2jQw95cf3cFm+eK/SpWjhDXz+A1VxPzEPIZRinSgCFYyodUSR9Yzs/VEoM
ZBOaJJOnjDdgYeRZJd4mkVKFQFAdI1hhU8ecRDCThYf90pemuLlecWp+O40NAEo3
tUM92WXk4uIbjt554h/2vi88KuTM8aFuopSVi0NdpQu8JdEX/IrqPsLceXPTItez
vOCGS7ivRln2jSIZmQEnR6CvgGkNHqejVNr6/lIExdWaIERLhE9EE2PVQWJunVc5
UzWkToLtyk72aIxi9CfAt0OQjhW7ww3JY9u9sr7SxWMpL8qG7ispW+/vdFaHs/QG
DZRQZrPdd4qpJynsCcBWL0ZViU3rCQOnpd8L7w+orYFRxMq2Dn6z0R4se244xTik
wfuBrOxAOhNHVpOjVKlmyBnVKbKPDh24IH4kWWlvV9/MvVZYyCikzmXqU/0/Ad9s
OJRHmWIMlbzJ6wCNFgpmx83MRll/RSPsV4177qtw1phCtgvSPFkXzG57V3oqIuRf
RXn9ar1MckntouTaxy0WnRwKLOVqwqdr8b6uLVabtvttcs2Kt11oz2GpeSv0l/K/
FexbiFK2Ulz3IQyuZG87MvRt+0Gto5/37lPNEoXCe21hk9SVZeBLOrcotJaZddj2
KFqyNeghddir+U/+oK31cTpnkoDlGLCCnkbEpiUsYWMDS/Dqnf/V4Bff3ombTuSd
6ww1Avmqj0M2gCSHp5ri0Hv2jOKz0Lfd7/vp/6ve6KtpqU/+m+kr4eOHlPCc9r84
KrvUslCssNJUdZniGxE1IfvkODkTpcV0qdBIzvZFgmMaSVFgO4Vv4e6Wqzin3enT
8NI5/Zlj69Yz6O29aGyq7mLEZS2bRB7uChfGHqyx8yi185u24qwLqzvBtu+dASX+
qlyUYOQOqfs6qpXvxGBQuQoL+HobVJg0A/rGevaiVjgejSdPUzBhubZWFKGN+v06
IXIeDQVZIzq4Pip2R5+R/A/UUD95X/opaRSnZ1i4pAKf2t6nNNLHfyFAV4Xn9QGV
jCqaCOyMCaRyJysqLI5DPy7ZhvaROBjI5Bi9uHQzJkj8QkLudGMDlx4PmaQga/53
f9WeBYVgWZWmo10v/vA3VfXP5zQbb2Lttgd34Pg+vTd1SWlXXTsrPDxEUDqGuunk
Jn9G4/3xgUhcCN+gR3OtyEVfCOe0GyxLYh/3LVrRaBjhOSVBArQjljtZoO7s/B6N
L3IzK5ZHCvJ4yRX+SkWGTO1FtSLCH8jrv672n5Aym8JA4T4nqAFca26c5Gt/ZCpn
ZwcyTIkr0sXsI0vLnPyFcQoOrsoJMpA1urf6UgCXXWKem4yGqhEhxXXxLKWatyca
4kSn6SPHIhNLHXh9ljhbnwRJwG/gRlqx/cdVmcjut0hNWlN4dTdgEX8kxdlwxh4Z
8aU30t31cxEaKbgVMRJ8IAsZ5z/Q+EFvcrb7cbT3zzrrMd/ZqvR2OSNNoHlO+CkQ
MOZvCkQzsgPwkeE2FV0wayPUt6+clB4pWrdSWAIdSBFmN9obtsbJkhujiEzGDMyJ
PIU4sFThmfpVT2tqmm/zlPNsYWrPrXOS4rkNOypcmmr0VUW3KtqXEGZTbqrKI8qB
af5qhaA5zfiv9ukvh+mpqcKc283A1XbzmoGTaKDA6QxRGzv/H1Rfkle4vMWzX3YX
RmQIgUdA2X495vqQ0bu8zpDw7RbSkpxq0vG7pXdkeYj+uFtf33GSF0uuiBajqRXE
Hgq774z6oPKzyOQfN9ua4MZPpRzNZG3x9XqqpjsBsE8W2hcRTL6whcgx/R9fL4Dl
sLxQQ/gEHyH4O+i5jFN/7KvWzNplASzgJu+tis2DNnS0dLIjsvckAN+JEHxFvkOk
VjqevLF32RFbi1Rdki527JGOESC7WX4ru0kKU96UZ0EltLKNI9KaJtPz8PUEwBMY
biHx9uS7DQ6S0+c0Ii44P7ltWCXdLYsTK/AjmObmPbv3qtV8bFV9BrC7W2hXACSo
+AsEJx+PmtlHBmfp2tRQ5nCE3EfaJ+hznlg8kJS817ZM4bvHhvu+fCQ6YrMGUJNl
PK8+gCqOF+m6PWrbbBgJ/syr6+Ysp/EqN3Qm1QjitLEdkQZ84X1p6GY0C+Hulcun
qWsqaXSnZWNvMks56k0kD8Fh+kYcpYpa7pN0BdukpPmoRHQm1rSFbGI3n28W8xUD
LDhNARi08QFVCVB4co72xvyQeNGR6OZCN7mpy947EVCjnIzwfO0WBgv+lHF/hsC6
EPoKTQLVfIv1NHEKFquDUeA9Lks6gwbj6KijTasVVkUcwGF13EvdwKM5AIE5zC33
xVRryDlqvoBeiCmIUN8bZljUcPCdM0gLykVfX0OViNb32dPm1/SCqKOPGNsqgWGB
/X1BmP3KL0J/+5B9jlqbzhyfrsVNEbgBQXByVFummHMYgp6TFUvtCPDmbvYZVTy+
UzrvLLHDgTl2ejUrBcTgo08GhuEE91apQwQQBnNDgQcI59NU81cBW1KbF37KhLIi
rzhxTSYoLFR0UgL2E9g/6JqftK6sbOOrz9Ol4D3pObvEDc3scy3NrT0l22AsJzS0
KzxvX/knKmDBg+1dOCpRX9RQqOscA2fYSq8j1MXjFXa+ueOuouyZosbgigkubRs9
8FPKd7B0sttZv0a7fo5rbyAkeLrbXJgu/1qJGYqimJ7Xfqpk5+O2zwjlvaX8JrnV
n22pl7sJUTa2k4rnuya95TGoRu2uuF5Kl5kImPahHBLMSJdPHJw7h20CFXvkXEOs
Zv0P/TtysRX07GbuFQ2UH3HA7uL6exXBsyYkeZYePJpSrpp9p2G13smCLI8F1nTr
EEhZuOoSItl4U6zZTVp7JlB97IQyBVqDow7zXFFNUNsjzddvAcb4pg63h1Y9lvjF
H+eTpvMYU2z0zI7QZ5CxmWKzmlTlJhNh6w2AQtH+8+WRXnlbskigvQO3kfeiYKQy
okotfSkkXivc9pncRQ1YOCwFATIFvhIQvo8Q5nj0RfjBaORH/LY48I4BzUbaodk9
SaVeMmHOMaX8sB7cUSru+8DTG84FIpVScrml+kqOxhcfiOIJcmd4g9At4e8fp+/z
fRa14hVq3+wji12JFXCbz54TSScLYNxYW8oFNcqYvZTEVh5pCizLR9thxTStl5NL
39MJzkVw8T2LetguGjmQi5GU09pEZxlVXmit5DpjK4Bwf4QU4M/zPnbn0ARxRfpH
pH4MVvN6BpREhq2KzIwdppEfrOjFfdtBciVzfKPtSbYXFBeaWFUWvPuuWoktkS0X
d8dpMeH0jivQ4PWbusvP0QNNgO45E0KdR3oRwRBhsxPINoSsJxyXH+rdcMMGcXyn
rmIQXSSk4md/AXcJf6IjhlJTo8Req2Ed1D4fkxWMZhhwKKAjqni4p3p8CzH30lli
pXSwySJeL/I6/61OxTS0U1OVUv4guXnsDw9Hh3PcLRsXRVylV+U6KxQZevNO+w8F
Vk0a2RFuWvEEn9e+3l8zpOjRy/LP++s07hAhulGMgsE2B6TN+0qrSYwMb/eOxRBP
Lw0qH9B407GoNvC7iyTdw11u+UIYuLONUd5ZjJKjR2JN8QOds/cTLKrDemWRey4S
z9KlmfLm1B5Fh2O0RjAF6rVnid/JXVFyCLFdjiGTukPBDuzjafzk0e++ya6xHRI4
WQ1vZu6ckp/ytm47O5KPNFigt/PBPRiwu1x7lJrhYrTuxKypMMl5RdJGjLmXa17Q
hK/wcYkGFjg099Q3nhiS1uXKt1IQfOpEYjjsZTzQOFgnXWEMiACtDv8QkIzyzlQf
FgTnNUWlQNUTs/9srfCDJMxwMdSvozDDNnZaDXRx8+gXomugZOFVy1T3GrOq4urR
zbV0S7P7jN75xYEpHbbbkeFmQFs30BAFOaUWbuHKX1XNTGs5Ip3kflW3N5LiydJ9
IbEfpWaplRQPaz95jtIxK0PoNYmn/VoqRw5EH2JB/isylw7kW/Wu/jUYtdVz8VDK
9P8PvfNSPnKL9AHjGhYd/hleW1KLm0cCpjnqjWebR7/9FatDf9WunVWlev56ozRg
M8hikexYMkxrI6rcqzot0Bapu1wGAI8bBFOV7F5RE9arkzRP5XE+GvtiPyEAJO+y
y9tvh07U06Tq8KIp70Y3x75JJx4dWzzcgKX5Neme2Ai883XcX1MR1RsfzDq3Bji1
ZXZ0IkCXMAAMK0s2MC17aQ6VXO70I4iNm3D+yYLNzOXyc9z5b56BeTh2SpyCB+2w
+QzG3M5D4rLpwFCre+uZSVev6cOleCchEJQwqLreYvwrg0Fq8pJWDVRvuDr0bGXX
i/IEdH1b+JNMkziRkRWBw3jko1KvBbcpugJZa/jwDmCHdhTqPAUWtZzg9FDO+0nG
Rs5GFPCeO0u+Sluvhh1lLVdNcnsKjVxF+B9AMYF+kauk6qdjpR0liXWjMIFUGLyO
7ddPMYxLNj2NuEfR8BUeinV1o7uWxmjoD6pv9dSuRQZbmrwvFzaPofb0MXuCqi0K
wG/lfPe/wWwaPAB6OlnDmwZs23RTmASNqG6J2d1gx1nVh1lPCdt4fn+yJU2gwktg
VOzVrX0Jo1oufbNUww1sFK9NjlD2FdJL0y9JlaIHECwC5+UbnO8333+FgC9h0xe/
5jHTsHwZCrU3Cy35kdJ36dzAJuNA8ElRblUE3uq7zOr2GaH75pO3nCSaxxMuALo9
TuD6jlD7SuZpBubuw8PDFBJP2PJqf7xO2F5UW7p05zSufOP3mb4ivvOT2TdOHkzQ
RJhNs3s7lThS1ftYyfKgDnfJjjimH8h221j9dvzRjPvIyjA+yY5sqGjVxo7C5BAe
VJBhXV4exaci+vlx2nEDX+G4sffYuhSiTx8xKZVzXffSW0ixbWmXakD/eyqJCT9E
rX0s4B+WMsi7pjgX1EO5TzqS22eEQm10JyV5ac+mxGw3F494Zi1yOnQWPfPU9tlp
w97lR4Qa16iag8ShlQ1HOkfO+3rGus8Gu/FNqU28SKkqe4EZaftDtJ7flIF2KmWZ
WcwYuH/dyHLeWxipBzGSVDqYKKPtZ5lrYBMghlVL4hLUSvMa0JKoYuM7rD3imvp2
3NtOan9Ldp116dvjjxlQDbxYC4aq9D4XEERNYNUmFeF4KHcFF3WJz707+JLf0vWD
3tUL8YZvm9d/XfO5WVNQQS0nVuwXqyG2k7r7L10O3nqU94c00PS8vjybg3TC1Bql
lRp8Cm+j8CgGCbHdLC3HWNqBIytL7PC8rsE6i70ZViySsCZS8VbREBOCbo/3vHgB
hOoHxDmpWs7z5zcCz3ozk20VPIX3jvjoChdxvKUGwoXuINxzrI2vRNUCTdItWGVJ
/YWDvWj4Y/n9LR4HpYVH5gNY3f8HRJmqHxIEGVM/SXnUSQSXRx1V+s59JKyHlTlk
PcsUeY+85FF8DuPv5gpHBHlDYF+WzfrDp9KLolec32FqLaC0d/0Xk7ffo9ii7xQQ
F7+jNA2G5ytbBf7XeFS32+yA5vPUKoTIUk6jxYLEDfTPXcV8EQ6AGATEY4sQWr5y
IswRgqTILAF1cwEbY1VRp3KH/ETpVNonPgAaeIpKKaE1Cd5eUWdGk9trLRdKoJNe
Gw1iQUwwf/nEgsu67v5vbQ+QxQzuYE2cSOpu8Kcb2LOD/fMJw2Xo0mIz5UdP4hLu
6636Yo+KrAEIeLjJE76mlT9p5Y2I2idsVJooWREtk3xvrguQhmygrwJvJOMO5qXh
+FpHKlhwoiszUc1jo6zZIA7ZBJqagBVUk1t/c1xLKWtuIlD4KcfNjJJXjdf6/Dbw
dSE3WmQIz6qjoZXf5w3csn3sJgguVOpUrSFPptO/4Hd4NInPKGbVS6xyvljTpZ4r
TCfJghUELpSzs32DDet2umoihX6TzMIfjTArd7knZR7G0WdIz5YKfirQ2+z2hhoU
9A/LwuZz5N1UN2abTARitYEmw87FyETPjrdTH1jSW1d4YiVdOan5U/Y5sWoW0+sI
/qJxYhoQGBuRzne1pej9l+kRCHOdLUOjQFIVt7IIsQicSnGFDJwBpCsqxd/TvLt/
AC0tTpVva49VZF1AG2Nc62ACz84u2Jf0IthvlNjce8TmQKQHfyy1nD+qVNWZqAmN
IWu0em3YIJLGjR8UKiiRnJQvvxalrJVmwHI5Yao/gCKiVvB/+zrP0GBZRRmeIAnJ
tVgdDi64WCVgEirIBFK4yM+co8RTNNnn1O0jHezOaRx1+GYltSBkPmxB4ARg5HkU
Me0EZDbdDaMpKMlmkT+MMJ35GbM/HE2F2iQVXcmcJQJx6YtaiFG+SObAoIofqMOq
90flox7JMNM1NANHrR4V1y87kUvUKt3rYpYam2zOFGzSzp7Xict/+DMabaySE0yv
0dk5JjqdR+VeT+MuId+rFhJviHcmWRmiY327cFimUMWsATyMdS9rsxYYZ7kHrzlQ
cjGvFq64BXAVBtp9uvWmkwRXgAvzAEKBY+AngYlnnSOFLQkvTGhnwtcE2rZcPpus
LKbouGmi8URHrEb8EFHiUsFb114Ewdskbp8uVsNi21RTfRJA4e3W0AkqBiLXiUea
ouLLblQjaUsqYOliZ6MLM4hOBxSFBWSEhdHvl4fkU5oy7rA0XaSlc+Wls1Er5EaR
yTWcTX2N8iKd1HmAcCd50fqKz6S4A58zWLrJoXa7j+QrSRaWH+RBEnGTqI3Jo3NA
Pa2HN2nknvCdw2iuacy6QwfFfJXcnQYuVKL3Pfg0+tF2EwySnf7H8SPIOY6U1tcd
Mk+RfqLHDI5xlWCKb2tA/toYHCXA8D6mk/omqR6v66LHlgCDtF3kFcdPNis/OKEp
qkepBS0cJtkup+XMBo6RYWKFS9YYWR031DwEwSlprpIJWE/AKIlwhhXNe/N4GTv6
kSAC0j5y2PdxrGADHQIVSKVXI2qdAANVih/USy/3pBPTeI0zOZsGxSp72Y56ZN38
U8ZVmVbtkCwN186neQ1mn0bGSW+yGnUg4K8cV3oIcM8yfHzyJobmMKC9xxWIMES0
efnPmwRvnX5YqxYfmSU0aukJIvm9Pj+GNgjcAEztvBHKD9DvRXvOw4g2F7kXCbph
BU5GAKQBjWFqUuZmbnwjld0jXwK+bsKpP23B6kzlQeilUL0yGKAzczdn6SwGwRfp
pFfRfcw/C/JzDKwj6pTf7FoDhKjl9rxIVZBj79NLZi+MgyysyaspKtl9paIGktec
vqSZ4xUNgVQBbwuuY403RI8hmydy89bHtEphg/AVdtWDfpU4gwx6T+ofLVzruIE1
5fetznul/g4VRegEgLWhoVSra2RoJxqkm5QIycfaUZsng9IGk0rsdBjT0yMYV9Kw
KgmR0fx1jpDcCiiDynGC2QkpYAizbgXdI7yXNm6OG+f/sI9LNbe1snptDfqv6GtO
ARLnzxgk7RJDxgbIZC/8RHugEt8WAUI2u6Mm7xURYM/er9BSSd7kH8EaE3bX/aFQ
O3S/pNDvHqtoWMrN2uHQwbJChfyoJKD2TfsogThkFWilPef+lUC+CENq8IjvaR30
CUNt4nLcOwg7aUR6hKVcSwEw+tbKCFCmN8t3/MHuP4K6sRg0NFricMwb4NFO21XL
w9i3XkLrNF7wVRyUxeSVtD3ehDioGr7a0elsSwEPLpZTPiENZXnG+7Fygc2gMCLL
/4VNY69S9mxYsMyPb7eeFrbw/BgUqCFkB3ME7GiaC5p5Q2p6zLYnxntNEM1x2gvC
JFfe+q3q56UDJqkSQd2h0IwMZVBpUBENLrk58swCyGfG2Or30PsrgN+ZvInsFl+8
s5eVPzpZDMb6WnjdZl5jpzMgm3j/IJyMHgZHsSwP6ke84yVhDlnPKVA9f9U9obzf
mWvT6BpxOwVjDV+FT3IjHPSfz76MeBuSWoQIy4+a/JyHFcPY1maDJgBs2gEaqTmx
D8M1LmDQlFLTsV/+mOBj+mCMUaorki7eLiP+1czSSkCkgYiDE5O3gak97G0GxpLo
ZyrVV+vBkHODE/UTkNER5OPypNn6R2oLlFClF61IKfJdfHk5RZQ90HtZsgnJ288Q
K3Opkd3i0h8H2tc91y6UrjHaWkeJTBy/kWGe0/EaiDfYj7mUw5byO5SBXMfvHmw7
dMgQB8M8QgQklXtOLru/JoKh4QfEZb1PU/v3yi45t3WGRIZKWE5kWpxaosNACSKU
l42bRhbkfeUEPsQ5cWsQvw5pOyLNhP4GftjBiQU3MS1vgPdhRF420BlaOrKs2APq
KVlq8iNq7Z3WP8kjzQquKebktoRFKIHmSNyZfHKnV/i7wZe6l32FklM6Iwol+Txz
/rdQpw/EUFybL1KJSVeTNMXeKTmj5cXtQB5fGUrG1+5ZZUAJYPpe6YlgU84HFpQH
uZltrwzzzpv4JibbI88Ib/os5a+DO07rHYh9dL1mdyOHdyfrIlEIbqWouA2lTEIY
l//QyU12AzC49tJITOIyiaFFnC7KLkCgVrsCrWNyLXe4qd8f/j9yxcmNeZioCiWD
IkwZOK9mqmJWuc2ZlulHj5KYWiyhW48dDjBvFpMlzBrKIRQkyzuRmB5Cy9DV7JR+
MsMFkLd+wmcvw+DgndxagRZWVPAWwemoXqDS/RgdZ/58zSXbNBLAHqYbaXNhMJWr
J/eJXYQ3Ky4Pxx6lWPVxigYrjwyPBFfqgxNfIf19aTuAiJoMtNeADFLq1XijonGX
aKSsvG0MoNJE4NsdknJl7sdwujMwZUXQUNpWOFDKgUCPKtk7Pd5sN8I5Mm7cbzY7
+Iy0rxu8TgGD+Pp5rBZYm7EiMuKz08Ra/LcUBSMPfW3bqlMN7n4y2hm1CirpUByg
55vXjEHGvI8Wn0XPuL46SLGWZmQBEwjIAQ4XCMHuLgmwwTge16ebaAU775P4rQOn
lLhDJWVhCMEfwaeDQ9SdK8ibaMbSPM6+4VUOMuk41NQdz9XniU+TU2vE6No+jQEY
LhAEp5UeSwJN1h2m6H9Svjgpy01O+sIcFW7bnErXDhJMbgVPMXf7NLm6kEyYQ/bS
0X6z0QU1euXACcIYCgvwnVKAerU72UsxtT58xsUmzvJXT2DUuTxSFcWHXtfcPTx5
+3eFAASUyrBrtePmi4QG4jseF8WfQXAGLDtw/ljJBNB6/4FYKCdaw6xqSzX/q3hk
lQndS7a2ebZfx40n7JjYK8Fz4DzyovpXNcT/3SsbmFtjxoDHDmp/C5FQdK1L1Xon
G4DZLPxi9oTLmg3XNaRnOxyoz5gjZtzzc2Rd+sreMaaaW+RtVxwcEE6lV09Jwbxv
w0Iyi96U+m2LCBoEBtYEjRo6U5uzCJ81jPMMA8y4LtOnTyyyw0J85nNtCODm7Na/
Tn4XtHg5v4LkIH5wg6AteHAq5bMRGG7a4F730X/SyHXbpEAufM4Pg6vAeWGrXjLu
KHvy4fC0e82FxFDp4ruj981+HuIROao7lURBU+zyXVnpQ5B4IeFV8L4tR6w0YUuA
opHGUuputMwS7y7MDA1rX9S0xY0qOluWWV8XnCZO47gZMJ8dGq31JMftWJM9ooDM
eH2s1WyzGtjErqZEjYGsJe5M3DkcDyGbHhCOteM8vE7QxUfjKkXANHtt3vUHNjqw
IsInXWIY+80yiaisc0BiutQGN0pYj9vwmxLfFhVye/TlUs4gvFn5YUpXzHhvWKeA
8xGpIGrkrqpqWCRJKweMDRl+qrYPoD/F0Ww0D7fXJoirqpnnQadumzJ7hBQr90hj
og4fyZRpuUq75yapDNPyWdgHUg6bakz4lUH82JwUObRbASclVqFrtqi/OmJdhQz9
O+wom2Mc1r94U+uMzt4J7JAXe2r+xwvldkWVM0aV1Hm8zl7DBZuPO8ZhVUOpDJsZ
e1xuew0weKS59KIHZ9ECFTGEGf/+zIQRM6TbZSlWYMgDv5I9/qEtZ6GpsU8S5CZO
QXV03ByB3bTzuIkDnpRRatZtFlG++FW/hyOuVkIeNCdcJ/q9jMHHvlhhjKPCk2oD
b0QKsCYoUFmfKIz4VJ9s6fCdd4zjlEMI+BqbLokZ7IiD6z7CddrrOOwmNw4gwZX2
RXqKCr5Kug6p4o5MMrKLiJDJ43oh+Kh7skLYWHFGuT0S7nV6M9ZJ8IUF/txoe/to
CYzVH6lRkmHqH5IVXsjVNqe8HXnpTQIHpIpDN13P6NxdmptazyIKTLhYLdKJcdKd
7HO3B65JQnuh5ekAHv7jIXHS2kd1H2GSl/Q0VRlKiH94zgctGJC+Z4QC/TrA/PER
FXM0Fk/uU5KVsGs8kmclAtTSrdn5clxpkYon+eu+UzvpHYLDfOZRUVanp0KvU81n
zYrAcsAk3kcUXAtyh9PhbwQTtpAJJlpUnZj8aDlZN4UheCpYKzCVHOkiZe9stVtV
sSWyD0DMt/JhbkMrynT8g1omVfZsxqENWF/UF/JJiFMZUcXGW2Wqj/Y6JfjVfKns
VHGlH1rswrdAs1HHftUeyliNDU27C32occr16oqZquIv9jKw+TB4qaRcgly9dT3+
S06v2rjQZpBJgbNA8SG0Wafuz8zikh0hC3hBtcFEMo/SHpL+9feARezGeSoCQ1Xj
xZkNPsIn2yJjL92WhZKLPa2ZHk9T40RaY0hk8oEltl2rTe3Q2TMp3/LT0jOeLoQc
J8OQPUojGQcB3oAPQXNv7gGUXcBf/XVwjngbugHt/l+aWBaV8QosNG25nzOINxtY
kFxEYCEH5bkLu2lUhGJDD+zm/fKEVv3tks3qeU3Zr94fd+x+VAF1ByHrZ9phJGRO
m0F7YBVh3ierxmXxaAxilDCbbAiu+0yiOgLQ9TINy3McFlKdIdikUXv/B9cHKz1C
x+Hpdq0UH/KOI5jXQGXUuL7tRtzkMFrz845XzSI06RkX1ewP4seCxezBVsz0Lt3/
mVMTSBs6W3iu5X8dkBlqMimI+KDnMMFXOoXgUbQjelIqmR/+5iXrR1zgrI0+yUuq
qMIjoZHGZL0BgrHRFvCQ7vbgTOz2PcWZrWOjdajbe7wMUJcraYvP+mprxT+b59Jw
Pig3PpjvLoAFPUvoMPp/CDqiciQKUA9d3PGohA97pMomE5oNralDNgg7Y6ovbrxb
BnGARe7x0DRySgtP4M4DJajmz9KxireYSaYl8wFTy6Osv2LTgCQhNShQ0icIVw5f
doLnUiQTZztn8UkYnkmWAJd0/vzFewUcGN+8nhRRVJJY4Jk4ZFI9ui2PnyPH2qMX
fxLQNeizpPOJqoFGf/xnZV/HAyZlvvhdLHmiR5K9IaSgvfkEIjaXfEKtHcXCQAbA
q3bcR743LuVWPje2ToC/CEOPOWGkLTJ5vOgyP6yN2Y4cnRvJpx7njydLicTCWlzf
oXAXoPPG+J4jYxRClLRrtI8YuJQn6g1tWkPMJSgkzfAJ3KplwX4270KYx8KABEKS
oxe6u4005oqz+U088qZL9NkyZDcX7/zNAUzmxqgnXK8Y/zxbqa7nqYRTSV/8jlsy
B/JbHyWj+1Yx4mf5X6u8EeaEL/H6Ct1b6E95BX1QXCdRBBiuqClclm7Cg47vG6sY
Hb3IIDilqTWfR3ZV63YFMS4iMWi2tbB0icaJKOfEGaoqQVB/ivSO8ktdT2eQhzGQ
D3fEU6WqdT6SjcMGOU7XAOpGxUtxVnBOcKsPa8N3Tgm1J+G05+gtjTQ4q2M+AdQz
7EwknezgS2fceC6s32xLr57olW/dw+ObE3q/rIKZcJp9dpQ2FTfL3+1XvSOsOm9n
WSNfvmHqI5Fral6vkwY5yzyPjB8hZ9mlX3BxUlPGbt/MNIUELhbt499DQg2hb814
aF0gR0NFihS4xBtBBBk5kJOkLWy+/PyVB/9pju7izo38JrFHixlcLj13TY0t0EHj
AvlGVoUZoPXFT/2WxuSDGuYrv95C4LITxrTnGsuJimHtjxv2L05DNOSiBqZLMMTs
YW/7RzHaw7aGMCXdnQRvnF8IwMT/jMk5p2ZOWAhierPXnhZQMX/vtrNWrB2c1n5c
dcRQ8RmakyB7w/fe7YpgUDVkjT5kRyQqHGZg346KnavUOuBxd4O1YEpdKyEJIZN1
n9j4v4Jf6YdC6z2mJdy+9MlvwDawCgEMrImdO4FrwsFy5+hkdtcYJROv/zB6UCK3
NRB7I8AoOka5TRGA+G0HRoV8WEXBwimkNWWH8DSSqJ+2ZAER0e7TFcEZir+Awp/d
ZHnRnxOF8VE6wBOuNkffbrtOl0mkVRUHK6wrqHEgLIfHKHPLKPjhwMYw8gWpWdur
d22uXGrA48V16EAExTLJoz5tJHxSG3xnu7PD8CoG+pWMbrOO59hslHEt//sO9BiF
Z7E2yXSMD4Y5YC8t5hAPr2V0PTt+L7EZZPyia3aUduCtBgm+Ks7BsKKdp0DX1VFd
73SGSdsRgFRln6Ggxx2TK6S51xYOh8meK+y8jDkyaDl1ONg9L6csPzn27VfSKg7o
U19lnRuPGaLtfd7mmcLDpAzU9mjFOizYAGDHaWL8DmkzeNHU2JVUr2p51AFMtM2B
MEyKFKuLRoOJKbokj8Ka2QHnP3ovD1fBxNU8mnUsa9a9zDoMY1wp7YfTPtreo2pT
sdYEfe6v6FuyW4r6URbGL0MGlLzWA68/BFGOq0GV5rhXgLnhxKnSjJkaUrq5kJcy
CXb3MsNuLE/jnHIaoVq4hO5t/PDLhLOP/PeU/vHmzdiM7n1h9tGMU5O+fqZtMDTF
7CYrTEGGjv37I5Ipyf4VEwWv67eoVdABH3UPmy93+jV9iXPnojLwzwgkzIWOO3ck
/yFKSX1wYVSKKO+EQ0Jc6rs6DB57uVMIBEJZD7R9xaZ1YH8Opl6fR1Vpa2ywl92x
VvhG9KpsWHUEqiY7cg760dseC4OrD5b9UDZpxGaIFF3HxPvSKXR32Xr/fpuY1y3G
IWfiQxRJrxjSvnsXkRRmCKUoBG3XukpfQEQtJeFZbaI6yCqyRFd3SBZjx5UxoL79
Xdp5HzXEXzOYHN7f3xbiEmF/LYo76scq/OQXcC854/BiY1VrSjPR70S+hNRI+8R2
dmNR/PdUx896spsWUMiVAXhZI35tbuR7Q2xgTvgphnIvWJnUiqByZnWWX+6VOivK
EN/Ivg2sTODzr3+31dkdag/jJkqac6GEpSCTxgJo/5Bl3G7ZILUhC/sUZ3PkcfUk
EDEzUVQ/hU3P59k93V0/PWmrI52BU2I62gGKMKgzVqX969ONwTLgas3iTc0OmdoN
JLlRf5WoEt7IgxWnRFN2Oi09NQfAE6cgwYVV6IhHhxyQEolodBTeQ3dKSX5ACxOf
Ox4DJ9prefl3OGJZ4psQ3UYCzCdwAALRc86IbkmYKx7i00VFKaSZz9KqOFZ03iLq
DBNjpgG+IAM0d/LJPLmQhRXqmsgz4EnFt0jGcJ6sQwDxLLJU2LVSiIsypWxI/J5S
MrU5EqrbxzM03PPjiQzK1UVcrT/2HMGgMd0sVMQL1vCW72tehYymwfNo8gN8BFlb
NtOVd8muMgNPYoGQzfDB7r3oSjU9vUSMEzs2uM9Bc93+kH120M5WLo6EIYQgInHX
7ZHH6goOxaY1S/HsN8Qsl58EaJqjJFBroa30ywSGmyD8VlYtb/Ng/4AhuGWEfZbj
1xO7DR3IHvZVGR2Hd+hQiSdwcRFwFTjm3KDnITbzhPDMSgPrrjZSAKC3A9KHjngk
L5HCIEwk3SpYVDHQrAvkIgXYs6o1qsJ7xzw1OV8t7XqNJoFMfW1oclkZBxf5r4wa
tRSLLSs06CHmhdFyrXZ3I/6gr5bsnR4jC6ploNiJ475QFRl8Fu85xZt3OIc2deYi
evH7kTqgEPt/cDG6A07OYwvXgM6ghxyMmVUyI/KRqerpPveLAAO9BSa273BpXnPS
qqJ90Y49TcZc0slI3kOAMxfUqiCI9DmnbLc1gvM++pVAXnJULsc9zOxzy90kaIkl
ws9Jey451BdNjqoY+5zQKaDWO+GgZIV39zeg+xRyJA5FiBK4jJoT2Kv7r3THrlv1
sk6VIesk8ULP6c8yGPyTqms/1oi37gmNgBof2o8PbCGeKdvJeZQ28p2VRe34EvjL
w4e3bt5mve5IdCAQd896ACJ/mKZSO3D9q3+NNM8t85Qo5KU0oRP6TvGY5PJ+jSkz
qz2+9urlk+uh/mUclNu4bYO0IsKSMSBy52EHmlbkXEJfnx6emmcp9v9syBZOBWM7
wv5/bUfIfrwlYNhTapGh9fKKaMHHVAeMDceMtwqLAt422bsJl2w/l6oBlAiQs/m9
MNUX8sjopefMEAmqxxLDeg6wa+T1QLzylxCFrPMz8tDkzxXktCNKb+NqRcxXYfPk
zaCsGOOUxDzcDO/3Yohw6EvEfzwtMEHbBXEh5fkn+x859knBhCUvf73Kp4eFtQ2D
dZes6/y9LwJUvnjZN4Tvo+Wv2F7+TT8BFJQhOADx7ljP+hiVGuJY6Gv7Baudmpmn
4kg3dRY10oClCEQodpNELlNhnlNaT21eyKpL0c72oUqh6CLxkXZd4dhvowM6PHz/
V2L95pxvX1QVnt354f2Ytko6CSMnFU/LKGwEF0M/Gb00bn/WzxWiXKNBGq3x0UKD
KYEaS5NP3XtabQUWUgFJnySwITHoQXPKHcGm7NmBVwEeLiGMTW3/L+b0AFqycN3j
lwqFfX3kxwk/+BjJhnDRWzu0Vl4xAEfprjUUWvg53oIEaYKnu5jt885TlwawqSm2
SE5EebR4e+xSzTfqKAfXSoqsH67j0ESJUBWQCcgismQze4FG/3nYO7X0Tzm8yaxo
g32ugpInQsTruy6fxn7SYiUkbzMqOyCFdshttMhE/Qp4kwhWIjXJQ+Dh9libqJS/
cUHvNscFqwMdDrNCaLMtvFO1TSg9cw5sw5bQ64QZl264YoeQ/J25xMOUujlHCEE4
dI/qfnL+9aCQT5hb3blfSHdBychwjn+EFb3a68x2IY9Abpey+QdZSqXcsqWk7WLC
FQKNcTVyF45PSUHq0WlBHJXXSnoq2QV3DVQcbaX/cVTuVioi0MRNcRCHm4nZGDnj
YNoXEucvpSPUtu9tNcBP0W5ogl7SDnD9/S3WUYXgbcrEUuhobAGWy8EfBsaq5J3q
+fB1yjPYTS/MMF0ZnkrCA69A4wBoxWx2V1GDvFQ5G5BvQX5fqNUccjm8vcFpDYFC
eR7QThCwHd2khOSCw3+gzd0ubjVAbaC1weqLEBRGdxD5S+iTHyG4NooX6PgWR52j
+wZVFZ+D+iTXUcE2hD5tzuTyqBOva68+tQlZOPgkbvkUrtpAHXL+EyvSrZ7+wGcr
dps4c/iuZxcoQPnVn5b6qVfAyyFgTseASFwV0FObRJ7VxYBTlxU/8PBsgnRsx9Kh
lMUBIt4+IRZeYhh25eokjwTFmnGOUcikrQ0Au7/iXIRtyWJbeyn2cRcj0pdAkQUQ
wN8obHh1xUv5wqoyMo8I6Jn5iTDnxAkbT+7bY8one3P7zYV1jFJGqBNEUYkBjULn
NY2+ODRgzNqzlrhv8aK3hPrpQ6aIyhEd+rcf2L+eiyvWRAInhag53Rup2IakUGa/
iX/i2hepYKYDvgFk/xw30XeH8d8RzYvzO0oR0oMxD695qPYyo6Z4tSEnwgJnMShi
MUH412AaZGcJlLGSf1DuYexa5wttFX2zNjTTnnbUmAIWwB2q1x5BSPhpa/Lfgyr3
buEX//b6lAMCJeioy8hlrREvZ5Sfz/WCUgDczZ4JIDRfepxznC65yJSxN84yTaGR
7Pv66oDTDVcuQjzkk8bNDu9wxw8MQvKsTdSqOzBdQ5CXgYq9u0Y9pvvMv9HOlcOW
RXHFWWswgyccqi6wjD3iNkrirxmlH6lpGpkGv81J9kOz0U7cQwrJNHCTHxJEfoNF
Nkzz5VV+uiqSTyQtPYW800YWtpOaD2+IGJe0/wvWmtIrRitiVYpBu9HQlZIxMHlU
qmkeUI2oZyxiiHgUyhgGWMAtBw9n5tnd+KmR+jVitTeYy+RtxPDwXxxXWBeVBESw
GjeLspVeOwWGLO+cRCo4PjOQop2CV+yMyAN2EdpWLHpQyzmYsCOP8qUsVRvjReHf
B86tY3ERl4fbq/GcZNf/OJgZJMRlQ9KZRJTq5NwCWcHJQvbAhc8GAI6ShndEq4dr
WYkavKcV0crnPVTv8Uk46aO6a3FM9I2yBF2V2pmitzW4FUqh54Tyf0EO5dr5RIV4
BYTK/0ZVkz6lZ3ofyns0oa3EPo47Dk0oeVAPzMZjFlG8k9qBUJXrS9mlbFZKZP7Q
lpgbQJGhwxYLUKgp7Xr+Fo62y0iI4arwrRLHwi/7wEm4nE1jn0wUyzDaEybXccOL
i3/op+LeNKWluAJwQJAbIS9l94ewtHFPFbys8Py8OcrPXYDZNefhrKiofPCBFxDG
wxpUi9vmDpwAnzm1BiLbvxUtOBGMmlxCSdtgmI0IVh0DevOsy8IJhCKENpAm130T
xVT1VVp01R8yfSWpNN4AJrnNqagRo8EvmTvG2liG0JB/Lp14R1HHYurVy24OcJAP
s238MAquKvT1tQDg1xAbnqfZSC0N9+FLyMRJSrcLvoOyd7TNYeFgk/oiwD4O86Xf
ebsmoRcbn/yqKKLqcStbBOULeapIzHqmy/l1njqY/ezdz+RN9+XKqcSFD9KKZB27
ooRdCsH6jiN4zgzDa22mqJ38xVl9v9xXgy4/MS5b10qQ60wtVck2BkPP1LqUAMRA
d50xyPe8CpQ2MAquW/9f4GxzYirolQYSa5WpbdB3VUONiixHzFviA4ybekmmPq+I
fahroW/XUPGdFnXZx0K4Dlb4ib02gUBiq/viDHDWVYofEzJrIckBQLi8TQ65J74/
MOK8YPNHPMFyrFMrQs7EV/ch9Mzge2rzqK9uGUU558Haza+v96Ymwxg7VC59tiI5
UqGS17UkOYpz28kh8DUNVtnoBbSXDST2BNxLXYhVcvVMBAUufw8vMwY7BVxL7Vev
WkQaA6Vm0iyaVooNgMiZhVbNzPmhduZTz07LRYdzC61/aMDLhrRGD18aoqUdypNA
l9r61UrN5iO/Yy4X7pX90AoyMDaS7Tto7BWkqTdKpwWIlLEsWUQoON46qxcLiFgW
UKYau5xEWYmA0J3hec59f7bCyENms8rnvWT6d1cC3q+/1jAWtQZL1CUdoiD9sIR7
F65xuGsNvxkzWB0yIUrTv2gEy/Vjpxpcz5hYe4POwutwoLeye+XvJpgX0kVFmrTZ
HV/LJo6CBW+sJFmvnvpNc4ofLpp5LvvL008CkvrE9NihI55qp2zcOadmGAvFNDX9
vj+OZ+DMZTRR87lOGRwBtLKJAsr1/o/lkuTXH6haMBHUHu596ly2Tm8qmWdUj6XC
hQtnzBBK+nKgJMHEP+cRZpvKk7M6fR8/Q9JeSHInbDXS269syGVJJc71LNPFtZsJ
qX+3I/qL6c7Zbs7fAmOzFL+SgCrRNrawcbPIAKJ/87jWrNoJSc9xH+VITFIGp7l1
qGhPi9KAjdajISkztU+XBfPOC+8vkSsTvS5Uns4w2TjMPZesNur6/vVHaRWFNIEK
BkIehqCbL+/7TUrtHxCpKIMT8xULNxEfKiTVQKZiG8DW7dZPBOZPT3LTHzHx/W2A
LkqTOzOKZIgy1N30gmuGh5s+5BCpCfpsF5l/riSFOw19NyezUnpG79q14Ggd2CMT
NMD6hElpoZateEZzBefaFNpA6mdIest1KT54gw/wT8nGZdmMOYlrVKb+mJvnf5eH
wAzxK8pbFpmIDawXvshsxlqls+Q1XlJfyDuSjvEA3Lg8CqgUhYq4/GStGrwbDIYC
SXb0sTbPMHh3OVkSEKXRBd7KvDZF/2pK/oGy1xuTYf1/y25MMca3uo6SNw1g8N+v
Xf28LifX1HscacMayjN6qcNYJ7K+sSJUUvFNdSnn4p9HdKaACp0gbQdbn5vCYZ9J
KHvNnI6ZTcgISO3dDq/c/E/rvo3B3tyGD8s1/EhbGeOQaKeQ1xIbjkNx/hFGvKZy
BBOPTb1Oe3O2O9gdg+47Cxu2nAhOcphIJ+UNOxO5dHwLftp26uMwExPg8pkvcdYp
de5XMF+Qny++dh2w/0zPKO2kHXOce66XzAkGVGl6T/6dgMiJUNo1hsC1jaDnyOfr
O0kORLH73hcxe0OJGjfpXyHd2C2VWZ0TcIYaVeyIaDvcQV+L7/i/9uhecY5OnSA6
FTN9ERKOkhTbB4GK8/ZAyNOe+yFSTUzWUaySU1kNQC7I8rW0iy0gf/JmrmN+uXe8
UNuwusb47aSuGPNpROZNuCN1qKWpB6/pxCqNuUR25M8VDI1+dZ1G0N1xJ3vJIn5E
8eWgm8OnwPDb7GJ64KCAmhiDSjwZ/2k4NXKcEPv1Gb6kbuPh42i+z6XXhDg3rNbs
vUUVI19FsFtbzuLHb+8EraSStQmQZIIx6RudG5f4PIBx/wH+jhJ/IQ2m1zOBVEor
gbTesa1Kin2o4P4iOul9AdIG7d+lK1wUAYHgoBGF5Y1xdlgK7+uuzg42EzrCPRyV
tSYeHhig0ZjebsptbXWlqsulpkkySY4A/+1+43M27aYxuMeOdDRlLSpo4/DVB1Y/
jTO2DNDivlW5qUQngKUXzT2IVEVa2hmxslZf5uPKYxCO1Tx0/oqpQ5b22o7Jefwz
sBdbLT89YQPWWDQmWA/H1YshCrF6k4Z0x2nLzggEA2akL+5oYccd4DoJNC0THrdv
Akv2pq9xG7FxThXMOL11c0MiMenTQh48wzWaS8KyMxxXSRTsQsko6dMgqMz7CsEf
j7WTXpgsx/4DvrAgm6ifohYpFIx17N0O7gXi4IHevanw5PJ2gEe23sI2yLL8S33N
0aXsBB8lryLjr91Fn1aKrwjzjy7OV1SreWZ9/y0cmImLo4LaOWIMOwoW/bMUwewj
O01NdTQvHQuUaPvUCDXJGMwnf/PffdsorW2q04U5RaoG5vMbh54HnbsEm4IapL31
vab+EznSymmdLAh8Rr4LHMUm2VvKbFfBDIpcQwojHrYedaTAXp+kImGiebuOguxq
2E8A9P3MR5BxF2RWESvf2UaFi96enedyKRkgmX3aSatdoq/Ne3Be453nz1Q/EhrP
wzbzRWk7s5y3c7VgLE+jHUiE7DZ7Xzbtg6GB0JCKg8FKDurR8dtZLQ77lCyk8bWT
xjmeh1W08RSQJeOk7LhUy1mKtt5s4FGSksf0iiXq8vCYmc/6K7nm9optIda+hmRk
6Nz4nW+JEera6/dc1Fa0QyVcAHULgsQNgeUIluuxzc77E86hensoyZgFxoP5oHRf
pcOqJN5d5643hqfdtVE7mgUtJVWezDKvjmUF7f9FhuQvGek2vU7/ViXyO/jeTEd/
hhhYpMwfSu46sapXxsQFmWxY8J+3RHJc/BWIoJrTcyiUeA1ib/W96lUfLZHidSDA
gLROUtBaC23aP57Wn6nT43iRieF2nIWRvcqr9pof6lfFOkOWtMcSVHisBlDyDeEW
qCKQZcMTFX7JQJs3vLMzN3J3zFicgcFOL6WXLSv2KDsy76NCo5usutgJLlnLzS4Z
FtW/BBtHfM9Bn+Jfz7DdPWDqZTfKtL5UvRyrLlDW57xNHgEKvx45zuWDonYunwvu
QkDQwmGrQd05hxruT/xham75Fc7s2Z1csC1WzSn23o+tziJV1inovOIBO85+yGE4
8cq5hhRxtpk1+lehZb2MbbIP+1r7+VpFlzXjkqsD+FvQwaLMlYUcz+4ndnOl/8sT
Alg4CooHxhdKouIvoxkNauAIny03p7n4HoXc5z6kb07rvtnh5k2uelLK4EXBOrdE
v2xtod5r87cDvHdsM3+Zv6ezhGQ5U5iUgghKGocToayFiWeDISUFAhcricSM7SbQ
RJpXXX++f8PxDyVm0kXNF+4xkTF5edxYWLSRxIVZVJZiIfn6KSXISZkS4ICg7RkL
+gRz//6hVXdZhXagF8+8gcRm5w640Cn8BB5/lQUy/MuUKASjKAs+6ihC+HnSnI8V
1JTr+72LcnfhcsrjEE4sL7dYaxjgGvzpo+ixYKoywUgHoiOQSpXF5/TV1u8wtFKG
KYvyu9fmA9+QfENtJiCrwPJCfDUdhiL9E/PSaNUZ9a6FV+Eo7pjVBl2STLN22GYS
72AdAzr97esSeQT/zWpKJooQgw6zJRooUl081rMiWIJKFHw5zTDO/3e2Prge+OlJ
Rfm6UBpAsM/AiKLzfz6UQdxlHMzvJ8A73VpdSc06OPnVFMOhIs1pN5shocKMqjyX
on1fYSt4QIkJ8utIxhZBcZPFG04MbXzrWL+YWgwe4+BnchdA6cYSC3kZjfQUci+d
CNplgqDIx+3o8VqHWhlKiUTN1A/7EkJ6I6aaqwwddzogpF0szNMf4NgUYXXykWda
QXc7ELKwRHSBAf5GWUK5l1Zodnl1dtgY7uq8lMnQMiAdS5zW2lMoclqMPI1cAzAC
0XCa8hjsJJdhmNS9zrx0wP8t6GUDHc9rUmpBcs1LfHujh6wKqdbiw2ulKU0A2bLE
f6v/1qhdTYwF0dQe9NNR7EA9zuVmPtft7iKI+VA3BFlCvvbj9vCUmIoojwj/LHCV
kL+yWZJBnJcA1NUslNElQsr7h+auSsQbpNtjWVbNVEjS3Mbqoii7ac3lGLrXHEfH
subYXV+BtNS6qM1lheOuTft22+BfLJ/1632+fOIIT70tKcraULBKttFm3LgI3g7W
XxMBe9cwgwkicvz9Fxlhz63pScJn3sR3OPvRQVX2KFx1nICH83BA2B3off7cJBSZ
O8N5fuK2CM9ihCBKj3BAItirOuzayAmGXnt7gss/NeFeXvQIuwpndY5r4WYsub7P
v4cNSEk+U10DPPeIOhsq7XfrTGF1dpFIko0HbbCQoBWh/fU5XYaNELK3lgDhBgML
7X0VCB45bKnwjTYpNswahl1ecT81HyKwVmKYTiIVk9CoDlbqyhld3YMpo3KCOpo0
WTW9rerxefqVWr0Nz2Gsll/h4O3g6r8am8io4WwLjz8UEsNNgxCKhtrnmCEpfN0B
D0rB/x2frbaWaMWSltIyQ9yCE7BYWW1gsCsQ3qOuRjlEfqxvD1v5ZMoexnG6GgSY
mc8Yyb97X+S/yS3GBbiExiGBl/JEZF9dTAdK+x59seWjsnxoq0tmaVfr8J7TjDHA
m9Hu+b+MrVRYB5qScg45HbrHBojty4Fm0d/wfy5X2WVnGW6GJdvTAo0esrHDjJlZ
J7X/nQvgh5lLf5fqtVAbzm5jx/tozoTFfY0YC6l+vDwBqroPfkc4mQ80AOyskwbP
DxJcRT2+D3A8ZMJ8H2MBPvLid7EhrUmEK0L0vTQvCqbn09PtnNEgrn7B2HBwvKao
9jouIcqwKnMj926chudCmhoUihbrhxn892urVT2UTQsHL14FtVWBNGYYleDurz2A
3RP5E+qRMnAjVfBrL3QhVeGfvY21KIcbvGnnRXVOa5bSYjjSxpuhfQArYedzL84+
pZ19CS5aCMazzlKKFgCyRxtAqMFvx/mZm1XaceePT16/e2QnR7DBd7crn9Tplk+u
T09wWvtYo8uqHnk1d7reiVQzFzcbG0m4wZmy9QPGEmjmPfs+k3Mkt5t2LDoYMGM1
MC2CMPKEB6EHCXy6+90VX9+hInsiQag1Nk4x1ogy3a/+xVZtZ+jt3QH4+/eRsaJh
6g8+hje7VUJ0LPD4nRQ1WBobYGaMuD7e5x3NuxQzywMGcwelqqMX0bxr0j3kyi+v
0v/jYlsE5qHE07XzyEfqaXLybsLrSBZXJ2XyaRAxZk6r0rGijJFLVfatYMxw4lrM
MTAQeYr/O3/4d2id3JNzfxNxxpylgEggsSOEqL1zPWLb1GKk4RTld5bEUvf0IJsg
hKGGvXJrAV8Pj5gCX+82EWsbZHu8QC43aZ9TvEJb+b64vYfl5WhGeGucHfInFTvv
t9TigsOfpB1RtaunOngLoQHy/KmZAFqNzhCysAUlfA8sLAUKDSWlC2BIgOYCWCHH
QW5X/qT2mijHZ0eYwEomMip4/08kUYj4EIcHmVg0eHSvIP1kjYZ6P1POHy7CV5Ea
DKAIdfKorEDbMbxYzl6vPy7H6gsSsX6KvxrKXAsDHl/dk+x8XD3aNoeCpdCZLLJX
nmmw2EssVSP3focfF7yuWvyCXwD/tMLTX+VANIJKazoDwXurxQL/EkAySJg2Cu9z
dxzElAPJbfelVBHUoLejzuztm8ggXaDvgb51ScoGFM7fjridjIOUT7ljalm0GbGY
S9DqM2f3Ip/ucsmdp2/J+cO9SjHCxpcJrG87e2+pdfGqVWZu8BTcjyYMrJQrF2ua
fLXDva1VUAJ61KC5olPjlkgAXyxd3kluRHZ4s+7M+gXcLQ+wVPll2zSqZ1KrbvlQ
jzuWZN8FoCVM9Z0GegfDd3GW1m8WJ/NaDOzUzbVC+5ePGru5LWIMTOc/ZIQz8D8u
M/Z7rwwSddaqW9x+dMMyR6JS+UwodPuvCv/iGsax8513RTla4xC1UvgBC8POP7IU
mSjAvSCOw3jqTFjdbgMKVzTyd53FK6lnJmR+zgw+m9NIzbAsDSPvMTT8meTp1TKK
yVQP/CmRAn/q9aJhKd79EpxruVApf04DHMq/iquwrv1HIEbx/zPrXgFghMhDipC3
zm66EMt7z+R3Eh/g6hg0rTSz+oEAgsezQsZB21Dgd/NBceg4kwDkeDITvqEu+wsR
FBlThP+v1TUu58Cg9KPQGIYv/dwBDu0qovbDh/ULM9sMSosg+Dns6pSQSJN0vRco
Q4tI264nOFr6gWfelmXzv0C1FV6POKFfPggW6pwsoIy/f6fbbA9pfHR2ssxMLh41
dOS+EQchTWAzG+PoGrLKA/+INNUl/ZxxtZtbS1S6qFM4XXDLiCr25c9d8kFvgpEf
dCHHelC2gSbq/nuzfWHU+pEEu6FWI/gmiiP4R/kFthO1UR4w/liXKJaPR4jJYZG1
KGL7CPwWmLb9YG06QV+AuMgGBRgjvkSk02Oiq4vsSBjoG+02oerwJe4rMs9jprtO
fPjGIre2b6lR8ikTHw7ruJWnuFF703Gc8vn7ZQ7U9F3jDOfWunz2yp+G/bfN39rS
9GKSkcXR40xDi2BWvK5fa4f/0U/vsMeIW1sDRzootWZAb6Zh2yu20i/yjqM6mXYG
GfnNEBnBrBFIQ+dz2zvF3bN/aKeBRjAgQFe6jQLXz5urIbhEaJv7QydfTgMinohu
MvocLt2wu236nJXu9v/B/vAQeHMLwPSre9tYpk3eCOkyx38qdQKeBxAAsxPLryjp
sCo4ljm0ZCLw6q6bOAqG0wtNWVnkREAIw5Qn8yiyB3jZG4ztzEaFUE3dPlwCjzf6
E4RuI//QdEs+SqZRU/kM5Ub836KblIZgP6MZ43lSW/DoWtXYOPwQDF+OVJgorHUv
hwgnwm75hflMIHa+722RtirTwNmLzMwpJX1YtBVfj8nK+xoHjem5bpbxUaoLQNsB
7WsPrzid8PMdMVR3z+Qj1bseTgajaNHreKWDUm7VpLoTDt+17uBj8jL9QqUVuWkj
2+Q8VJg6osrAN34IEsZO89dVFaOf/Uo0wpM5MRQIIUjVqKjinpmFnvmsRYZcDBFJ
s6/lvdBKXWxudAwTfRrkFvrkqSTjwobts3iEW+Arnhlf6woOprVKbpuY1Y7XGIiR
MmDgHdWdm98z/c0Jf7XRxjvBTZtbedKrVAC9SA/+hx04wnPG2AVfCHhsfhUlZCy1
0NPEEfkqqNt8dtgZCudfsE3FmdT6LkNr46gMRpwM2jkp4g2d8dNA3TJ8MZO4NVKV
CUjsVzd84/irkZ/ENaZpAbs9/f0s75Ap+xDi976011Ii2d7NAVKJVn7eWeYTyMWZ
OU91GUekY96Df1+MN3dwejxYBxZUkTqCJwzWJjN86WlPQ6u3k+Wb7P0C08Hhcwoq
R092JwfJ0++GanlKCMWkKFv1kiHvRCoYz156VJajLWH6Ptwmo3SHy/2hVCbIM7hE
9CaUnBNlH2/zdz40HyMl8oyvC4/S/hkyeEwFgEOr+5cB98JRCjblBI9KgIdc2NHj
Y49d496K+3HlqUqVa/F5vmjy6D0vxxbLnycDEors8uDUJpzKv7RySAJtEG2Qmr5x
b5+H+gQRD9A9emC7ctOVuYtkeqVxi+ryYpNUoOoJ/lSV0cllOqIbmb6qagjdERkv
Ym7cZ/DYyzT0uCaPSbwFMVNTHSQi/8dLDiYDgOhwa54qbkxD1mqlcOdQE8qoE5w3
0y10wB5yHu7vV8WNCY+nmPpagoAZW6HqCum7TU0b/M1dfKpzFEYlF9vkQR/R0d7x
Vx3Hbg/Yf+f/KP7LAt7D7cOqbMFgT+K8Rn2Vb9pbJEbqo62+3UNLPGDvmBrUTp0j
SLOfqRpA8SCoMTLnzAPUBQPUMlVjP9rzFV23CMTC7GrCK0e9pTlxGB83nZjtXK+3
kB0X5TQpyuVWhvVWOvu7GUOnUqagy1MBDmazB8YuIdxOs+28rniX2OLK2PiBm0AV
G+vskc3wT52bkppNluUeNkn6GlBLTO3UN9AaEi/K/YxGWEkMyV1MEGiV0E/Swf0Z
l5Z6fQ2hnMrmITFwGB0sOLPf00AR+C0MCY5KG3PQzfAxzEOFbkyT/I8Oxa2l2jps
/Pb9kOb6XsRle9lEVhQVBmLEhjz9TijClC9yoDR/j3YxAYQAqus6P1GsHQetSi9F
Gd08S6DI/PsXVJGKa0ze7d23++k5bvqI8XPpuLbo+Rka2FR/EHdHjmAiVxxodTeh
f1qzd9QXv0bdXajrLCNOeWzTMfSoLFhNWC3gEJDngWLTjOoK64QYDSSo88uFcP57
+hoSDIGbA0uHf303ADoFRFRceskKFkNtTBwGR5aVe8BZrUX+2Rp0hhSKzplI2STz
WUV4UaUOdTvXvAf7SUfP2g++CnGXvSFhCrzkVLv0idSEnlZAb2M+WTxlwZIFbccH
wMFwOQm0tgnLRCyzORgJ2PYWwOmQM+gcbeKwpxAhyhbKgp3GCK2QeroTTCIznhzm
3hQkBKLEK8W3EOT03Vyugb5NkrAHLt5/RqLuvVmWUQcZeFOKdtPMNz7sPEDktce8
BMWAPLX1aorQnfuW12RpeTsJGlSbZX1ZiPXQznjMIdYhSDuxqYbd0egvdi1L1ARC
s2AF7GAFkLoHuzbW/pEbxpsYDa7roGio0VOzPeg6HsNJ+Wkahsbog2DX0jIYglB5
CrgKS89krmxUmYUKSYPCHlWim5gpdA8uN1qxCxkF0EMJZUfOx49T7xosO2kL4fK4
rwblUG0WQtN3SNCzZBoj2TeAzaRWXe0T3xzHjipTjU4xVSh02Iw42+/H5bmYOATb
pviNe6lhfETGtg3F/eQbMxI9fQ7/5yHeU5qjdx+irwUotqL+DvD98Tq6R8kAgIN4
4a0qpLXHWWwhngVhXPEYhIOp81Qxov1a8F9GCXtd12xXx8cDuRyKDaUOvcMTbzNA
GM/BVhjRVwVnmPER90ZOTdjoWpjh6kx9ZjEox6IYkhcujaRXpxtJxZim6S8cDfm4
0iOlZuqI8/Nqs8giMaMTnJp3rLLAPBpHwnsytVStyjmMy4BbS4a0suBaFOs5doey
p413GHAzpJukVs2JFvHba1B8DkhahrWskOspWVAkHixNSah3ZVbRO0+XuKi4tSwI
T7iCg1ebo3Dl5V1Viwjsl4LjerfdgeuuFuCVfgyUyaJ2WuCt8/oIMyMbq5eD5is1
0ZvfnfYhULtrEGPkNmOKLnYDFZ/Qbpv1rKmqoVgv45T6/E6l5c/XvgF2nrgzBZHa
jamP/rYbiLefXlY3KKVrqoEQ0DCu3XeIt+3zdrV8blj7cNVJOlR3IqPAvOzSNte6
nScMYFYqPRqVcZ7QoaeB6JciDEptk/x6mWrtSHajxa5AIpVXlhd6xUxRKzOSPrEE
9vbvA4h/xfiLYmgELkGGrM/1Te2FclTGsWHSiqLi911tMiDFVfPZpAWPYdvKiPxt
ZXSRj4g4R7qJWpSmDuthvxGjihzbmkhCrPr7SoRZEpOGhZEDCPc6SqHI+IKgBB8J
RTWLSU9RNgd6F3NOs64WJ/95aoInoV257Uj5/sgF6bVZzre+GtCYJ/YP2+VJ9tyV
WSUw41sJK/YbacxUZ+OQu38IdRUMsTOKedrZTSMzGaR/CSKJNoywkw1USCfJZs1B
d0Mbpn//MExZM9xckUlwz3YH/rMJ50HHatpCzuJ7/ButrSsuNYgkHsBMeQYb9B36
l1pcWqiYDdSeXkTlTsUrsxm6EtUF++dV+Bcef+f4lTXLtZGXoPKOoXI9CFJuIUv/
GccRiE7cuq/MfkepdD4NXcauEKSu9z9H5lYA34BmAX3ROmRyqA4RkD5HAe2Swlhe
C4t5FX0ABMVINT5fVyeoxmwAgfd0+6YdEVoqd3y3Nfxm80l9TFG6QikLyEX449bT
3l9txqH2Fgc32bxx+GzIlDelaJO1/+sryQ+DotpX0VnmLL8CSGpwVDh3X7smBpsY
LhOAaJeGf5/+YNzN0J+F6tRLwbbemZwdrdphHZn6Pk8vq5vLzTu59aLUZPKjZaaP
tBzevyluUJPcIy12mIXoxdGsQ+1zwtrwBNwINz7TRmb7rBUh71Ffeva/1SPuJ/9p
daCFfw5J6E1t3LsKkebPBIV3xKLqouwKkUY0OZfKE8rzSpvR//Zik3hxIoCQ7pAq
jQp738Cl/Fe9LJuRPpjhN8oWoXcvuq4ZBjvSyTjBvs6h5/la2crv8WRVScdZ/AQp
ZgwPvFSgBV0wmPOKVqmMlxc6YW38Vp4+u4wccWq2RuB86txDH4jtNeY3KBmP5CjH
gPvKtGO9SHO0MXJFYfX9YnTojlG3Z6I/IHxqjFSiegvkJrAVees1vJJMiBb47zF9
i/eA+XaPEEFtGNIpqKYIlsH4YlhoWRa5sguLNPlXWABmaoYILt9inYuL+9Rnavex
cm4knIN5+ESBejqwOqxXYkxaxBrvpP+k9byley+5OAVuKUJj3ZoZ2OwVyr+KRkes
ly5UPORuAdcsDaawczjMAYJvkiYSzxLpDlTYFPsQD/ujE9ZQg5NzAnHBiJmLfDja
W9GKvUKbKPNC0BQEBOABSg0DJRxdU6ROBa0JV6pM3V4zEXiGawBOhDLzqgSxrmLg
8h/8m4/JTdTs7MIuIfp7O9qERRewE+alRDjlEChlbz/0CJc+7GAluOou+N/LWTFL
br66uT1oj75csop4XFKZuTcsB2z20tSCUFIVUEcykYq7oClSUfmoViKEmUtFGTto
+D88FlgNfHajqyuvIz/Cvk085i37va8Lk5zIpgkjkheZK8pJO1QZyUbGVurq58JJ
+Sp3o+IdG8ml4n1nxQ7XOwtY1meSzcNKxDkKeCSzTiu4mjM34M/xBeufuf1gqg9y
38ve2M0R4YlqXdQvGUa2V7cXQnhqNquKmi9AvQX3gk1ZGu7U7qtUh8ui+ZggWcPM
zP3SPwjTjlKVQr0ImG5Uv1HyQp7ulL9+q4JRG4Bc6p9dCml5BwfBRv5SXRknbhfd
V1aRR7HtC/OlsNeRtnC/nAr5ToBDopEZWdrJIQsbOWwSCcQwG/WuGy9X7v0PWCpk
bvRxm73xrMKlHLn/+ocHWilvhCLqaQPZeakZ9klzuOJFNmsAhKb8QV3/4BfQCL50
bjy07YMCTdHi2wOovk+ONwFujPWFkjvss27lfSLhIbvbr63ITKD16HDPIM+1dbiG
ee/lX3Fe9/j+nwsBn119t/rlsSMZOCKRRxcHkQn/WoRYDvddvUmyhQP84bwgpXz9
2auXxEAC2tFW+2USMSWpFJC50e+2zcgnBrhjbK5wtimfGMWYt9wcC/nggj5vghRb
+FDsdN8d7R9aPe6Ishi5LMXa3zsFc9IAg79RhV1GYYwJP0Lgy7LFP9DymfZOtZ89
Bkv/hzKADkOOkaZePGxVRKXjkBhhfGzo/xP53LoIorp1M7EL8nf+BBALn8088lKk
ryw5NYYtI95bBFN4wPOdSyMTvEknYY37gOMN7zhVdMayw1VQMLhA2OBo6XrR0L1F
1o5PnmQnWily0M4tS5iJTA3BOfl2MZ6cMXzGyuNd/jUd/xEa1ct3JzcLS708QRuZ
O5OT0C2d0Om9SqdDzvJcRwNkNLgSdl/4I3gwV1KzWMm0rlh/0KjnJk1smWaeTc5h
fEGKqWLbS/IdwrqXIhMtnBgsW65spSUdUlcpOLZO9mTIoCTLmS39q2Dxgu+u+hM6
i2AMz2d8Z/77oY4r5JddDN3uZWg/6n5cVSuO47Z0c/wgaYqOjgXgsaQBuwydoAKn
Kij15gIA/Pv7joR46LEz13C10m1/CAqKI8cCBUQK86VIIp2irCdhL8Pxj/1/s+qW
uHsH28I6K25Tb3jPViQ/XU9Au8IxT80AMRqga8MJkisPlMO7wQgFyH2OaUY1v2Gv
XQ9KRvXayj0jYNrhZDSXpR1wMMA0rb0MlbyvkbWEF+mMFzdj0xfwgscxgYt0PPd3
D7dZ7kx7XURxE/05flZjE53y6tKnnDnngeIOWRJReCtA5d0KhShzhZxueqymjAl/
OSv4LQh0MkcQSB+3XONTCX50OFWvvHo1C8hkOzcOcQ0FZfHgzQ+d97Dp75tGgoik
AvFJBLUHdtyDvkr4vldLTNX9Tv7ZKC2MHs86+/8sDFUZ+7FlKOp/kt0hlCY7DT2z
d20FnJ9BlP+XXlYpiuJxcaYSitXG4ki+z7+LX5M6RHV0ryv7KXsa+mooe1MQaLWs
8ysmSA6XRJlqmQHYh4I6dxOmuIUlz7HRyI6BXFu8Hlo7RX/5LKxMJYlgrvoVCdb0
v5UCC6MpCyhekxGUAOWWTNrkz2utWpSS0eo0VKuFUsBI0p0W+7JGJAJv6bxoxLkN
rimW/noGF9j6XdBmn4ycaY4UGHrowJA7+6bJ3a53UGtd5aTM0A2QPAQvUtiNC16r
8Fy+WhTYssQJSVVPEnmNpKL85aqafUsDe3xuUD2swwuACATy32Vrx7DA4Z4XEgDM
gcjosM4E0puQRuwUADKRUuRg41KSoqwKnUJNKpFz58/mVC+8rB+4fBeMXcCKgHYi
R9K8HWEbP0wvXw37n2fjSpWyFy0huYMFT2DfQPgxWVbNDPjjyxIIjoUCyAdVNCKc
DQ8zLsuzaJp+U1OkxkleJDwtOGGLu1eTt8MiUtlHJzw3EbVL70RG1IM+A3uR3hj8
2pPyUE4knCpN/wJQ9oJYcGqc5cHiihRmlw7Kb0CrPepaAGYwJHzc0Qg6klgaQCrI
lIDXYFPkSl2kZ49zI1yJx0p+fT4fGVgxekcE+gkphEjgt1RLfC3XLm7PPliIA/Ru
Dr0nzqGal5Uf1faoxzR5q/+L8K6vBf1MKq6u/ipfqBbeW5r+bxxWSFHye5oQ4D6r
Yof+xPdgpWO/rq2ODVUGzC1VW0F83LnI/uS4NeFu1ruu6gA2G3TuxuEzgrmbKSFd
Lo6+dJrrCZiMJbJhBwMCZptTthpJkyURQKjwAAbHs2XyjhYUnnr3S8ByUreRIOUP
FFa8yk2n2sS4QFQh/5rnnf9bBoxeTUjWBcgb/krTLrqKH6Ycw0LGMmyZZK1Hjtvp
T/t6rg9zwbhKxGRstTdMrFehzmzmLkd3FlWhWMgbjJsanV9Kc8uOGeMnIQfdxkTY
PxmyWYxh+zN6G7Jkybci7NoLTUKvhk7MZDxEetx24dLmEj/CabJr9ds3uN5ZwUvZ
reN7nyOODwjMhSdrh1H7fiSlfW6vnLylUQ8+tivn5WwYZU6F46vVzEQE7vK7EzDb
ITW1GTI+xuVlmMwkB3ai5lezVwuVRjEDAM3pNFkWSmLy7l0vq68nnUyDCmf73cq5
gwHZA1h3yoFfSFsvc9QCYFuAJABhPa4cSY3hF/U65bSegnrS+QUsdJ37ifuyXbK2
EVtDKo3shd8s+TqgRMdRN5Z6yow/AX49BCCrF/rjBRDHSBIP40pVUGawYfbWxAce
hZeS7Cvy/JdKbsnvoaf4AFMWDHx7ojf0F3ygnJa6k6agwC3d4VfLFAfQGtiOsugM
o/XI8zPf02KxdbiEpg1qAC1MAVdr2epEnS/L9KCP3sNQylH/n4sdBWiQA/+DiGVV
iEpqeLFx+umtPaiD5tcVYW+ISWZUEHly2mgilVLNYKI1Z5Gww3ruTmN0tlV4ieBy
AwcPwOEIHD3YGYAli6pQoKNpk4/1PYwuRYBTnwoUf2MveoXMLxvzlJspTbme6yqr
K8z94wgAIbwprFcyYDsF34oOhpaTrqR+S3ArrA2Mz8hOGaghscyEZM5V9vpKwOal
qDI7bH8EDnqsvAvUYfVcEOLhADRSiFJyRKJra4/F7VpfjHuEYA7iH1YxSlm3y3iN
lYZh4kUtzNhh4qRKOegwgMhbOg2upgHovDOnc4qfXg6UagzyOXobWlr6zZxtDyWT
CZSUaH1iXpn1v5dyCFD1JDVzTvjAXtVfK2rjQwUPRThZLNx37JvDQ3bw8Fm8Txf/
+v1lAj+jNZ3CAAy90lqpWBkZT6QiKemyULTSTg20YkYhqMTrMS8CfGdVwxt3U9V/
ffeBTerChHU7LDyXImmCXbd0kZ1oMAwZwY9Mljm4QDn8n9ixYE4/t2azb39oNl8g
rSQjlS+jcGHD23LRcqDL4/B6FN59tmUUwjwxKD82qT2IqxE1kQYUJWBmlyXSvLQh
GZ+w0As+4MGJRHx2m8KhwJwbdv+DdcuCyi5Ne4QDeSvjOVCQXHSM/yWOVW3NrnIQ
Yb+FIVajuKdPeBzq03/7xCTydtmEp5V1cspRp2Te/ssIlYzRvNmpdSaHS2arh11E
kgr7gXkDJbyILgmKiMU7C1S5e2KvoeD8L9ENJwtIsX9+i6FdgZGj6FYvZuo/Zl6V
P6QaT2xCOCkujrLKINfsHFO9yN57B9SM93mSoAwdQjUz/DlqGwhpew3+GVFsgq66
fcyXxYDL6uVzPnNieHvU4LwPPNwAWRDmqfLdTG7qP9fwuA4A5klIP6AJJhvhsx7h
n7/wlBLuMgFJvZugDc/T1M1ktsxHZl+jD+f15b2fMEdOFyvDCxnj34PV9ehDoTwZ
GMU4XRRV18azGcqPVz4Bvedoq4dK3WCVoVBhcxorAhJq4308bqLkQKYvrAattEGi
bViGzVN9BYyDiEbDWPvhZ/ROaLCFAv1URFlGS8PFyZEsBsBwaTxod8G96dQmbkgR
TxoIl4pW0pdaMIA2yVdZpWbh9/RhxIzfOmKEZS5+1E0nS6asTzTVp9ThpgQYuLx3
6R4/Y70wo62XtQNeRw/gYnzmYXq5VmfKBZme5MDkdIZ9TlzfIVpRYnuc8Zx902eD
/89cakEHGJeET0dsSpZmEBUh5+2+mK/MmDY/yOWixsLWMLVGE7VUvBgeBbXrvQU+
Oz63OSuIhx+Ba6o6Pkv92ke+ZqEiQoYgcoewoORQMXzNJ7WJLXsdFV+9YZSCKJ3D
nzm9tp5MdPzjXc0de+eJVVQgrb4symCMVcM7I3GeDU3c3WKy4sKHhbl/kGZ1Wrhp
VUeWTtiWOLY3m/8wiFics53kFtLFTENIDU7VxZ+Q/PMc4DasiRxZVmIftDso1Gf0
EWBXuVFuOsaSGJs4eCywH9/UFpIXq1yzetb4M+gYVFcw0dSN/j7/7sE4Ei5ns1Rj
2ssKP1h1T4EseNANWO/a4+CeiPdSTHGq/xiEy70utxAPRot69qwJref1HG2VK133
NXOGM+7x0+jCigKV0D9hglY5qt/9THukgb1QFbcdqnY1GAYPjCxco7NFDR4TUHMy
+4Ax6SildMLZQHbImaS54IprmukMwxyCFDwB4BLM3tUql7/7tXE5qb42h2j8mhnh
LeoThd2CyQVv0cQYOMWQ19z6BUACa6gmjPG0628jchXZzjpAgzPvs7pA7+Of3i8u
rlqYlkTjwtzhM1n+OrAzfhf2KpKz3s8kQVrtufe2vnOOgvwMPsqhreY+Hm29PmTk
aMbgGYafC9bUTRuXVA0N2bj5jbvrfUxdBt5HtnnY5AneQiBdSmLSU7OkoDNiXGEI
utMx4hLI4bDGjv5DTtM0z08PZSPlygs0KsACTdzbndE4cNQUr5QS6wy6/kcJTB9J
1xvp/zU5SKs6iTTNf7TfzIS2A7gqzlxASDHBUgq2ODWWBoJmP7x5G76WrHGEoReX
UKE7au/6nsXNjE48NpbCa230ujFdy24OAXAibzJYh02yRkbQQuOaleOcfOCkXrQY
sY24vV27fDfdd8AFB3b2mKndcHluxtTLvCZezcNWWMRZydknlg9H9cYrIByNTss8
BF6Dsw0GyUwUIYw9nZQs7Lo4zCfBefk9rsIEM4tpwuDiPopYkBC/oqNoqbfRCd5t
lnT8D/zuWt9hb1imzJQaAGFOyoveGmkOm5gj2blD4aouP3peHl1o5rlh09T3OaD7
C9OaN927VyuvmKDaz0WO1vkAZxf1Id4ZbXG8MaVsQibqECkWp1MC8ZF+rcvm30X1
lKN9jHfcxy2icrztQ4jl1r73SPl7hYJYRGPpmJi6MidKUUeylNcY1mKev6Es1ROj
xQH1s3oob1dOtPxqTWBrZaQsFJlRVRm/J6AC9XCpD1lXvai97Oncn/LgzCa4cLQp
nyGarMRAksuDp6g7/OY0kN53xAyunBOE+Kfrs/VQ/AZYnBncFKfN2EUxfjU6CUq3
qAS5iPAG96CovUKMdvyYK8yPmUhxePXxddWLwuYd2qHogpM58qhAkukJ0eo5tBv2
7TxSk64dKrNVy2e778Qq9r7/riN1GXRE0Uu9vMqhAh5x1IxhohDbDCN+wNZ0se3q
oHxqEAX5ohJpcd4c0LiDucT3etQt4flnyIg03GMKDBHZxKj/8Ug9W7p/csrFKSrC
JcMQMkpCmXPrQPfXXYE/vs2CAfLAgNXdpZ43Y+01w8tiCiOUh1bmztpCegKHKMrC
FCucz6AIIyZlaK35ke/XlihC3rxo8RP528cItiGCjCTvHb7JNLnHufdkof8mo9wS
Mrnh+S39HmNnurVwpSibs7jie+CoV7arTILu5ZeaqspRzwmLv/KKBCaS+8cohfBn
d0VZArImjl+SG75ZyBfL2NOwKOQW6K3gPiPPclEpM+/ISKLq2OyGXH1n9dbvtcB0
EbemKqOA+G/+GAK4HaI7trWh9Nv3xq8znJnXgcJkukDolkGDqh9rUlFNi7bCAK81
kOo7TCC7RvyW1HmhxbxwVkA7bJ6rCD+u/Ja9Gli6KdjC6ucQNn7kMaWFy4yaWErP
equDRD5SYdNqPDNrfwxF3xtrnhENUqAaOSXdZcRIiXPvNCGdvj1UYmr7Jw47BBeN
NpNX9rURDvScvwOP1+5fGbNrHUKAqRXG2T8AtvxIgoJ9uX5Kyjs9VaYxnMWNOoeu
/9Tji2vYXJZWktzY8CcB0AthfXC0Z0taVAYb3TqgpFDzxWZVqhupDv4gsrQQjNmd
G8mBaEgVk4rYJYp6zmYWFRbFVtFhKtthcgGPl9+8hE2AH5yfBA8lzWwevcksZxDV
7YppP+2a+sIUTRGF3Zd03zfvT9yY9zmktV6UeHySw2SM4j9QaApvp/qTpmb6FWVr
qEnuewFf9AXrLm7RHl6i2GNci903Igu9NIBmbAnDEjh2NhsDLQoxMGOxdyyfe4iJ
AmQkywJ7x4w3IGbtXkkAXBgdaeNcfz/bBUA/qi1OzSlNHtZOf+l2p6Cw5FiKexzi
PxyFotHjVdkZHTmOKMdO5pl/V+Az4Y72aGMV6jxBDJLecepr1Xo9xO/x+2uFzUD6
x1ZH/0wi2ENiuTQo3AU75PmIQNat/getPxwTgEpAsTqCFcDVZvi1yidIuEitpJqn
S/isV2qurN7b4ippFQ1XnWKXbPZLCWZSQjnoi5vVE1C0RykD7JVc3g27IFe/1dDo
838hGFRvSFq6oJC7V6po8/TxMK9KHyAs4+V1IG8xs2bFCMLcCOIVsNNKMddWqMjS
G5FBVBZmSyixhRIvbzbVY1P97OHGRT3WqCdF/jFC9DdbDRTjBfAwDJp4uDneDq7L
qisT1zu52RdFmeIrbpU2fmGRWWpJSMSSwMPwkV4WYH0A7JOtpgpKPyhlM32WwIVM
Fa71LwEHADUJWUxYJPlBn4ZZ3yUHIGmkYpQ9mdQeD+HqR5/m8J77DO5umpuwcP7I
0jO5xGFepEseTGN6LHgqG1s5RrLavGMglGqFXVxdXbsgiCN3t9tO33SGWf5ij4w3
stRSwjb+Qhz0T+OLP4kV/pJNgWI7HcJAFLq3xbbHhd5oBObnhJ0Q85uPBCj7YNJa
ZOZ4nx76dpizdCZtAbl1uz3bvb1WARgchrpMw1SmOe8Sa5pGm541Wsh5FCpiHZOc
eEGSJyPmwxxO2sqFZGrpJcrLNIoXz6bjIrCQ2/Mnbe6NUeJVcIdWxFBw0X6v9H7H
cWa/Eg26Seo6eg5nsXXcMC6lSv+V6wlsU1ZhRUHbMz46xrwZi3U6ZdH0VDdzSQyh
e9owxrzxsIWJ2MvSyiUQ7uMZmYPS/q0RUvDcWygA8Ey6KPW7g0PVoP49F0OmCV7f
xVExukY7IT3w4axdjVV+jPOtoEpOWR8msFPPahhE0tYOEGphlDT2+ZyRq7mQeyvN
n5PRf+3GenL9g9qtQhPkzPEvaScY1NRuuezBRTomh97rIOZwKtpmi22VWRyWqus1
9fhVbECGjgRu2pFxwxOGRf2aOWuur8JIrgjPvpgwgnduvQzAY275PVontT4r7/3P
gd8prdNDjZ7iMOnOqNKPTxCfCpE1T+m9oGXfA1tQwd3njrGZsQDObbjJM0+BigQi
aTFQIe/A69UqIKvO0rt/Ug2NEfWhaeNSZBkovlugcQprt0Yo1b1eSdjAAWt8xZdT
H4uz6JGKCEZcaMir2A2mAWXV85wN2pbYv8uzzrlAylMRYc4M4C5aZvpY/mP7eVy4
jNrUvjRNS0S2PeQ2oEgA0258wpCL8JZ2IKvMF/lsssTBRY4NIP/yPOqXojxJ1OrY
2tVDc4gR0oxTsShcKVyryUIrcVekgZjZFDLPXh7sn0440pQ0xVNMbRyTes6wt8Wv
Muzqio/Vc2I4R49OWKyplBcmX2Lp9Ulplj91heZBfsyVzk5JZqRV6Nz2P2hTbx7y
u0rExk/dtMvLcHSqwkgDvlOoUxbLXdJZbj33/ogr5AMocjJxFJzZIShxvUCxnxef
nEsqt33Xz1DiRT71P9HrK/84jns60dOKEf5hFHgk+nWE82/CkHFf/bYPRX8BjB3f
Bi515TVNVYUI36uAByuK6x8BEo9lMKAzwpiSr1yBF/COPxmSkeE/m5bsnEvtgMK9
koynf5wwgC0zFTmCZ5/hfRXyfhH6eNdaVS74Gze6fBczT+tWS42vpohpATbkDYjy
crbHjr0H9Yh+cNKLu+M6ZzZa52SXXGO9HYkvDz+rb0ICsnojaTOSD2Iv+yMAwGu9
xaCGEKl7uoGkxVfiZZDzb/G0YfG7mleOej9C1+q7Zss1lCbz3z364okjpPPXNgnd
2qF3tx/fVbWj2UWN7KT/+xxYWqiVXkQdz93mpPcA9Vg9FIJH5b/ydvVjQarPeF/q
wychKlgkp+2RSzm7HjUjAqTEUJ3oT1OJ1kcphx4BKIZzNj3KcmRVVVLmKVpIG8oe
8dfTHrxsOpnKoFnj3dhJLy/gdLVpCRNrIyEPTPE5goHQGl3dp7s2eI2+a3OV1EMo
TaXhs7ry5jfVOULQeWw0x0jthMr+h2DJzTL4WmJ9YQWIZ2+lP/+WIwNiwffRM1iN
itG1cv4GBSUGHW3KcDQfynqaA8YgFzpHZSt/bhMIokkR3+seqHMaRYvbAKLBqtBh
wQBWDZSB8xeSr34CDQhUErofUib9RVEoeBzgXor0IGqD4M4cEOBocAuyxhom+v1k
UBYI9gmjeIq2A1HkutAfK2lMTLLthU2eUaTlY4yuhBPeWoGTPlOntjpVcvMWrQTD
W1Z9ewvef3riAHKv/S9jX6EykXp0pzRVJttpEZUiqk9OtkLFSmioy3SjkljODRfA
WzYTNW4XwYjmbLIep7/ytlutrGLYIH1gdQzGrfYCPcOFQ4F6Lf3ZousOc/i8PBzT
A0UQRq5x8/i0BSASaZB9Eq8g/KR+8WT1+KN82rfz7NS6g1uzQdv3FYRbbhMzTtHh
zI2eazLF/pDvSWx76JsxdB3IOIwpkBKlgFykwfb92Ca3dNjQ1JXgmOYQXUqih9xS
J0R+kRcCJICRN5NfX5IDaL7duQCdLSSe+DPYGf/5ZWxkULFPhufsbty/kHvPLZ7C
DN8HLxj3P9AzxWEASsWQNxpKO8/U5fTHfg859X6MklEdFnvhLuJm4csMqv+lBb2n
eUP1Ff6FuB3bK4FCGeiAcZHPCuv3rYVL+BVhVP2KXUsc+TgYPSAUJ7PFLvugEgqH
aG6EqIN+j+P9d+SL/JL+NJ7rn6bmYx5f+iabOfdVBFX8DeFvQxiwJkn6S/pHKA+y
3vjnDoLVNdntbly1CH1Er0sy9tGYpx+CxQJCG0V2ZWySZQiY3n/6IaOJ1WJQjNvZ
XerhMKKL3JfNJJTUQIgCVCARo0PJlF3092WgtGhTe7dQcclBcY0kqYDca0saU/K1
UERgKI2w5HPuAQgJj+LazKuQNS6JqwV7vBv0n0IHOAmbb/XQmtk84Tx0JYlUk+dS
HOnmybERBjyjWoic1QqHjJQ9LZYaxjtmdM3X9j/PJ315KqmBmpPs5rFtNbpVNTB6
g5FWjiamZ1/IdI5o8QyqGWVMPvE6q2CY5shPHuKrb9RYf4ihpwJ+TTC0gAX6o0yh
nnp8zpcm7dAz6jGLPrptnQvA2yA9DJKFYvaXsgYHURX8SEWFso0GhLKGnxtGl6Ce
kq8ReGR/0JQ43OIsUZJwYzckiwrhulMZ4SP+QzOyiVPDscCmdZw4q+Y0ehQsAtTt
fbWeugUlLWq+qk8jP4vVvgcKD5/EQwR4GzSsqaFfx3xpXSL6NDQ9u84O05mrzBDd
1HfAzrjh8aGjuvxV4x/3SGwO0p9nBhNG5Auk8TNh2Nu4RO0YpBBNV3oB0kbIsDNu
1yn1NTIc3LY+49TeWcgo9gJeF3uKFivZ7UkaInVMgV8rAJ0qqOrtqKEYI+i2cfkr
zc0pGbmTtQGDRZuUMXUk9uccu95oclVfnmpbd3FHXGhFBx96VqQuMg8Ni8ZN3RJx
KCbSFmT1Zb2oAwmGlOHhdKr9U18yLpZVs8U1ipfQgAo5qpa1JnBuZ2ibKLeMXnpt
lEjh7mXzeySinPfB9tIavXSNWxl06uMJJlTdWYxB2pxRQIvuEo/MPUXsGT9elE0m
Kr311PSLXGfvP37+c+jn+s9bJhWaWUBTSm3Gjna2AK31vtQNFB2Wo2012L1Q2sOY
ih29+P9bPcf6HeQhd4Q+MDPZj2oXupFvHsR9CcPpah1q0t0lTm+tbfXi4QpIdIAS
xB8/8T8ujosiry/ofGUnPyF0MQhLhB/muspolrCGBvUNxbUa+XOGjV2mwErFPIGe
bnqRDRLbFRVOJpn8Sgg3P1GwOKz6SyjgvZyEETB5qMZfo6FXlWbCanCHGoiK/qaU
Xrh3ugfq1mWrtyNNjQGHas5OUS0viuSN4H6jEaL9PM5vHOLt+HfiEX7SQqDQ8rXD
FdlKzSFSNBEK64QCjgfpngDNiU4RIhBCuiWhfX9wUH5SsDuiLRQq7MFGvOaK5eDL
9BGSu6jXqcaNuwZKH96D57BIMWodXvXV7Nv4qluef97FNwrrdPu7CDRmBfJ7B6H5
FmECxtKs/TEyXVsY3rlb/zMJQwmfbimX6e88fd48e4aers0F5p8zKvhoMpCvTol1
hD7KAClz/IonKKUlkauH0VTbAHosMGTufgB0AMbMIJdwukwgHlmXBR7FLrkiATBl
PuAie9HJ40k2/zT9Bj/NGjlhvYnQhbtVNN01Gf7ppGNQ9C4/IfqyV7pxGzgc4bXY
ohma5pVsQ5jV02yV4Dg98XR17XvRcvE6q+kkaY4M1EBrDJMQ9NGfNq32rqJpDyYb
XqsS2/3xux26zk+LyYcd67VqrMTH3euBWRJeuppCfHowJo4T88ryMXtkrrU8Pl+i
uaA7RY5V7UYLLeaU7gzO2/nX8uOHYpu2VtaA2jQJBlFdEN/ouEwgPMWZxO1wH5x5
aT3bB+Vevq4p1fwC6IZpb4rLgo3FJDhCDZOf1eUIVVdfi1QzItDTaVJwwCLBX415
ohxxsSP4UO4uFHGinYylUUyoN2DXkw42P/JJUC2KeOykxdwpLTW1niqwhnHQmuk0
fBuVtDyfdDU+SL2kC/c1KjhJh2VmN+xYXajPnOJXNbiuPXWBSnfGVeazfUPdjEGU
VJT6/p3YTPJ/GjpUkVeuQxcNWaRS6fI0L6VP8YVFuOWW0OjRR2i57nMUMzposkHj
N34FLgbkYM1WGDJyAvTiAgy9WIgGfnv7RDm9HNC9EtPRjr+dt9LA8Nke8BI4kEwU
jLg7cNC79r4f4N1vLFU6Xd6/rotOfkxZy49lNAl/lensxIPqdbOwqGT/lKWjb/P2
0J0hf1kqcAsPA9QjCx0UnPZArJefAba8BXzJCK/R0cknH3CVrdEI6f49mh7/CAe6
DdCJtTiJDBRSmfLGNoyl5UuU9ce5adi4tikWYFUXOeLIfBOQs0O+z3JtCvdby88/
J0cEPYPsYlKgT+6l0D5aOu0uRvmMyej/yVqAjnit62UcsNus1XP6Pn/8CoYxnxB2
aTHbU9SXY6WSa/cM39P4ZJQxAqX95KeULhJycYnok8vbLO5qfzcL5FnxNg/0+lTS
6G0x6uteMLYWBESZ/TYLktfkuwoG6Li3rFPOhq38LVpUBL0dGTDNMUuvsTp58rxy
0s1Gss7/8fXd2R0Fq0BmsBOA/3uJS4SfTEgU1YYP0DbRyv4/rZBOf2fImXnz4CoJ
GnI+6CynlwbDYb8URq7ctc1iqF6qg5KqvSkpGZ1K6dF21VTSNmYSTWZYRpfqUlLT
Z/ud10KS9dkgw2H2xXNmm4h4NU6PDpci2nnSLF5negpprNTPpwwtUrvEJALZcluV
rmL7YQ2IZTxD2eZiSRvBve3WgjCgLtUg56RS08K+8r4AjCmXrVwp3w7tMd3U9iJH
uS3lZW4W4MvkkHQ71SFhIx5T/6zBdWp8O8HaiqZgQf/Xg5okEWYrceAMViFI88MW
90FaXZww15PCFf3nPhDKsdpNVLIKc4ZwYXTKZ6ZPZT9lW98xkhCqY7Q23nkieFvE
XdysvUJce4LrkhKyDwveGmlrrpijMqlFsiTWYuaCt18kjiA4oikF+Wn3EsyHf20D
dk4njH0EE2ugufOKVdQ/6OaekxXVMiDEQM8jX5iQbcA5Z7bNNjhmnKANJo++lKZL
cOJKA07aeVUL8ZtLtbAEIWxCKu1k0Jcyp+Hx2DV4xO7OQqr1dpjOU5+PCF066u7z
o5zMGQmCyiLWdsmbakUbGcLvEErqv4Kl7nhdZNAmGPbrxZFY36cmsgUV8u5J8Cz/
3x9i7Em9U8i9n/4pBardlJql3eaTvM/2Pb8aiOx+/OVt6noN+GsYKXCz90Q+Rqts
jAHEP5Lf3tKlv+/yMQPaW2ExMpcrysTFcyH9EiU1+qVArzKY00PSB8evi6WV47J2
iDj01AcfRgH4qEBm+2rkFBEEGq5FZqlSCXThgEf5xn/cWkHXjmx3JIKMJzJGeufL
RNH0QD8JHy0wmsFHt1wdWOHnWU/aGzTNJmR6EXD4YfQPwr/Pz6P3wKA5DzWATli0
Itk+d/0D/7LEeWqo033lUaw+1a8tq+VneC/MzvAae086N+rmLZg3Ggcsxqb+EOtK
mcc6ScLFrPJp0vJy6BKML5H27ANzPdliYhGLZ5F7DuDy/4xYImbGsp7/b3XuflWz
VBU91Ooz1OcVtkraShZ3+KQPtDpmjNsrC6+gh3u1rPmlZR7vJ+W01duIA6wkXPZM
MAa47PP3sRtET8MVUnBo655Xvk7+2FH7j+R+YwMU/pUUjEHekThvP/9WJEVMonj2
72hn0oAcQ2cPOUsCfVEx0U6uDFD8nvr9Tjt813lYykqKnxG3RpqYKg0ZBfD57kvq
xMJ5hraBkK9WY9yOqCauchUdHgxY+t8PgocmfRgOp1gnhDCc8HCHTkSy0bLZsp8l
MqcT3oKx1/KvC5Gazp+yR3S5RAFWzSJyh8KWtRqC+O31B/xqH1SJxAMIsOvnotyi
HFbdqLU7k7VHmvDd/1VVVA++Xnt9yHeE+zl/8T46n+hg91wBaRwsiYJEo6yVrgbc
TcekZApyBejWsYJL/gT+opDGqbbEpSRHkjcsf8cCQx6gF48T4/dB/KA3uF2InOVQ
iEJTfjOEqslqmvSw8YeI8tBi8ydKmxrY5E1vX/n0R/nPJKlOX+Xrt9dyLYeCjx5U
hRZP0ljwmwvGyrzSsgUduxe/vTHhNmDT3QSHUnAbz8zi8Jq6gK4ye0I4R/t4mVst
AyCe4hrPC3O2xiuXM9yej7Ovgt+JIEBXAPIFV1JNXjpO0y/llew4NUKrfPtq7Cc1
Rg+ISo+e7psv8f8jP8M1cXUpiL/qUL08TCga/+btzuF74X+96B2ZlLDoGmFiD6yG
kvl1YIsgZmi80aIQIyubByfyvAXxNoHGeKQFSVogj+RJgqXd930EyaLjjTos+5TR
IWczwWH953uJcjYh6OpIViUypLQLyGvAdyVXWRwGM3rqwC2vWxgTSC6BQdLjlWe+
3HbZ5x8ViMjjayWHdSYOoYV5S/Ny5mnX+YSZgewiR3Zqw48BPY1sgZRV887uPa03
ORIOoXuSKYWGkXkwqOPwPg9gRhwzewlcXAyvwclTSpRXry5uDvP7jyWNNWkxPDBS
QduuRZxX/71xOmtkmV/Ryv7InOSYx2StotwUhNgVT3wtYrfNJPU+dwyc0sssCQBQ
m2ExUM3ll0tin+3GommS5rZXXm/UALuhX2dPaUgOsrcIHbYApZIrsiIa5QdfFy3u
kuwukok+y/20KB+xtQpFOBtPrNLDBq2farmVhBnyrdyM7yvanAFi9bPxxAbTOyYe
z+RNXgx0hgm5V5mSib/FzS/+152vqizdH2uxaecm5TLBSf3jRF78ns0z9JijejT5
W8Jud20k0kXw74B/2qdxfB7n94+LrFLeGLWcHaspn21wvdYEEEDcYvNx8CHadBeH
AcRYDp3xInVRr6vAk+iIWrCFVcfwnLPCJ4woCqtj4Hd7FlT3Y/ansxp9dD8+VH2V
glPvasqY5rAim5+Keg7vg47FsAHH4D/2nyERLlKAAHysGYju+qsLSunc4BOKemml
u9j+uCDAMk/s9snmKuBk1t10kwmUbm4hPwCrUZHsaYjJA+IGXWTaOPcoDHujiLvo
CE9d0O6Lv3rdxQG9TWaY/Cg8ZYhhppqvIDve9IKC4q0dVUyqYrMeMvxhtMEB0cCi
OSGOid1YdWCQRhjXUO75zVpZHwcF0EMeyEu6+mGZ4I0EqmblLUM6GlVui2A3d0Ts
Tcfjr+uQN5JQqZW1Vr8OOskwDYEddHDUgUHZ5sr5Q19ZqU3RgRj/kDc2Zle1GEyS
knezxRRJ+dfm4FSfKqoyuijDEHMnzgYzVcr3IMuomavcc7Rs0mUpbc81h9Kw+84g
eR1l9/Z1YqAZdteFLAmYuyx/tQ47SUJQdr2QSSiSCRvk24WCEsySIu12pAs0lyO9
QRVD40/uoaYJWhXX8JEmyNkDB0nhuhXsWKPhMz7Aev5rVidtPz4CqOASsPjDSTKG
tBlhGr1rh+s8ongwU3iI4OgmKA9GjFnlnPXQzaTfYHjCTBWc6jr6IEzHuRbofVZ3
CRM47uAF+c0OcTjB2PSSZJYGcofMxwPnEYYGne0m4f+gBUoAPgiO9iZhpJPvM4kf
wfxalCNSJ0xas1KWOmPfxa9MG30GKAdkYFubOIGTZNqfjC+Va3eTqNlw4P3mUEMI
Qpf40AFFZsHuv+/iCQ1WGqpazYKEnObJHDUo9P/Yi3Ey2dNHTbVZWXXaiBESeJd+
69Y11FhXvc50Ehv+zc6lxmP//KC4G396p6OHWxkm2R+FSVS6Mqwx2dZfa4nSJy45
EQ2iD/NBH8xLfPxdv6jZGuAWFSHd4/JaNploMGLkztKkvhwbLEd4xtTx+UioyZOm
sZFZQzoFP6aJpZxTn853FR25Xfmt62Fn+xqSr6Jv3KGKIdswSYqMx2l5/k28KmNI
oRwTjPV7gWGnWX62NAciCMzidHpChmJ49vvSd7DO51n2r6XzbjNCsSviYCw2nuBb
yQ3v/abDQDJQwRQe5MOPgjwYVcpAdoepVnwcJn4DOEUpiS+/6J8D7s8f78EoyXNV
NQtWQA3lxR9qcpVi0ERAPx+Yh/BpbIJunqNctkli2yY8XV/dnyvMxpc/U44tMIqA
wJIfo1YrrSs5LyH4pr4DcQ68wmAhMrGtT1yoGWOSIT0xqzEoaT+gmafjGEh6fKRv
0b2WBwrHRbsOWbjGmOwjpz3vLIZM+TxBTJcVblbjLGhkwKlPTYZ4nSubVOVNUoTK
CfsuPrf+DJYyS8QOyAUlo1Bh4ozp8Wya4vCz+mx3Mj9WS/c43A4CkZUrchodTtGU
vlr9L8Ys/TwV5BaCVteGTRueBab6SUJf55tANUuiR+jYt5ZOV1t8hJ8bGGImwzDH
o9BtSX8vDlPyGCJxaOOsY9ndtiC32e0DySsQg9XnwpHnJOEbtp7LbmcLM3DifBgi
kg4trmyqDqw9UVbIqmSPvzc4zf8zrVeF79x+G/MCqQS138upbnbpbjZE5jWtvYCf
KihhQoCQO6fSb4nwV40Y6xcvT4s5UXOAGJkzcJ7HfclbntzGEgZKaM/qIwWblf7Z
Z9jy3J6YOYnv2EUgk9SQfes8QyTxadPf+j84pkGzzSCrksFePdnKKkw/lvnz8CwH
TP+sR8p+sn/pYnTuleBPOj+6uC4Z/leX7NXjBgp1VJHb4Vcbn28HCRZi7WjCLFf8
HOF0EhlsxJyyrGZEXrROBfLWkUOHuIDo8pZOHBBmYcFkDtTxGavLCcZai7NGKHDy
W6wtrD9R05UKpDgQME6om9pxnjK7CLf8K1Yzh3D9HMlvhX/Wt9v3dNZM/tmqEXM5
61kxoAxRJHt9agBTPGSMa/Uxv9y82YGxoRMe8eeZLKZz5Ffyyaj+mVcwFROUCOf1
C66id97RZ5Jkfrq1thGMVw1mcCtqzjha6RIlEiL9+2WGN0N7mhyVjaxsaoMUYJDy
UL/4Ex8KWBy/mN59Njhdzxu7X6llFXKhcisl5cz+dQfZRCY1/X6obmH0uTz5C1aq
zTjI7jLNp8HEV8Kj2ZwdwXhU5iaDtGbDu+3tgtVlmTwM6wsbB3k1GpkGVQ2YL8fI
pV+bx7cDnfblRbMCQMIO1Sg5KwDkQoXB1r38/Cb3OjX7vxsCpCk3i4sbu8qGXOt3
TJ2O4Io3bx5gUnfyv60jGeRAV4FQq5KS4fbPC+rGvxSUywOaXeJ9V3osOZEXenLW
t8ixZvaIoMDGjpToAd4WEs0hUjJCtGYAwqKyJ36GcGiyAtt8LlqGlWAq81I1F2ai
tCQlh8L55/NfmqDZS/ZWl8gukp+paSd8BM9+tOieiXmQCIlKXOmj9KhLnXNuXqv4
Ta7ijMfqZPyYbTYX5j9aL/uErQ4w6E8gjFdgHoQbytP7v83VO9xptU4lXhZlDl1D
ynXec3DGcv8mIpoLgxN9rcKx++z5P+2RxYzSUtHRu42iEYJU3QnYSckt0LkPh0IP
SRiRSzyxSrRxNiEbyR/CL654Zdqp5htB6dJn8lxmGE3+LSPZJxUD3IIRBiIN7WpC
9L2CL3+I+GzYMiAghpXsUOUoqvfnDf3a8OriTJ4UUDo+hLwiKSHDd6qvNAlYLBYI
zbSEGCGD20b8BVAmVtw3+pc/edkvmjZBjzvUk7e0qUokABn6Wo2MIcYSVpCbAInO
oCtSqWW0jtEHFhgbTZGCwYnxIVilHzPleLUw7DGUdSpPoGsQ6NlCFiCu6t4ybgq2
babVIWiikvIrjgitA9Cg6t17YWeBghZHmEc4o9Ya+YWMt6oYm2Euc4DCvxmCo4oe
xD9fgRFCpVtScraJKd/Q74b+J5fci8t/v+plA+jfpEup+G44XtxfAW1dRot9ekJZ
kf0Qea6ofAXmrK4DURzOjSjDTOL4NcXob/ufEIoahx6GjJMa7xsQifgSrfZNVanh
ycoogmXsvjL7zPm4OPtHRRMs3Onad8ta+vGiDIdf8qcNH0kCZcyCOnz2HG55dNHv
/whRijN8M60MrApR/gUy+86tLlGtBK5ojtGZt0xmYCxStUH9CBbrK8CpMO2/or2E
ULWGuNzxnsA/Uis1VL08FeS4WsyS3x7Hsn0yr+UkOU9YVVVZERM8Qal3P7mXtoYt
2lIua6lcHZw+ECvtqzpAI8bcuagxE/TKSxR9uQKz+o4Frdr71eyrWnms2Qsy+qRc
YZrK4LEpFHXiBlakhM71pTgvm7Ccfpm07HaB1OL5X4S91VGBnuc7b2Wq52NN9jsP
Og1eiRzyiI5MOe1lDgFRrSED0hEn/6jWNJzhM9Z3Y42FUrdRwtNEWRSvLA1XTsWX
g//3651JNkv7dtaOSvukNtj6JH2vUz30Cm6KhkqVOxXbf6P6pCa9n6biwg6h3w93
6fuEYjXgT3mtjluz+lB/DIiQTjLlJjHChzXE04dXd97SiUzmKoD5XVhnJsrrLkA/
Fx5x+PxzTNbSh7qDQT5+DYFEM6PLWJ+TYqpxVQsGhEwaHW3DKhPPIUAf0Uv9Rv44
6+IYI3QYHSqk5Q/ASlzvts2q41t3BcooZi8uLbWlcdT5xTJsV6ro87hcJqS1iaFw
i4jHITOJ8+zkETx0vQU7re8S+3YZmBI2pHN5TivlG0amEgo80BcBKoXMwk4bk1ce
sVK5+GEw90pwH8qtfdIvv1FNQAxAalixBQMqqtIuODGo6XUgRmY8tEEB535sznzJ
2b2vFSYSB6otfDaGJwXVdcFinJIxYbp0TA4sFVyTndB6kADFMhrpPMYrXUrORA2f
XTPCD3ya/FFAcF9WPWu/AiPSBIFAMpgicPWduRmT9JG8u7XpeRolP5RI3lskSu5k
VR1MDI/Dm0CbNMB4ygGKtl9w7hrUmHjHA0PiffJj0qv/WzbpoarYAmV36RZ9GGV/
OgEJXYFkpEuxVSH/fYBWElVNak8dp4X6U4VvR49uXAPgJWyI80+nmPkzVts1POop
xMCENTsFYM8RaVTdUKRtMNH6n3i58vSjkcwhFo1OQpNokUVSw+xQLmM26rsMJqfj
we2dAWEH8FWqORtS4N4e4mBvScCYc9PMFcarm/C/B4RyrBLnTx+lmwrwTvxmUpKx
3fTvHycRCpRfbCqpjLiGFzNSwO30AFXPOCah+TuFUMyFjc+CGCOeXAylN67OYFOY
PhNDyiRKN2vwFA7Y4k3afnDGuRhvMQ6MW/yBpTV+J5YtZUKFdtM1/NDh/wmE+rTM
jkxRHup03HK6I5jpgeU22hZYq54GYNNADX5UEYKB+rBca6WLw/wzNTfZj7YWIvWv
k0Ew+55unoMuW/0aFgpx0hcYgOjKhhnHSnwMstSgHEGHn6h6nhR1CLyXFmo9bLmZ
+zWu0jcPjQcQfTU04yEGg47i1OMKZsMUX3w5pptWhzHRN3TjGcz2sf/OFx3YOvtc
sIe+E5lFxY7roUujUKZUPZmAmy7alYZwbpWB9rffnhIoYI/JTPQbkN6cnIdIkZgl
ATyGF+a89NE+5g4zyY65FHwYk+KAbPOKAMg6YygFuHxyJHNpZBYnKec7LNOlcVUs
mpEaA3up8kdfYcc7Lf5jcfx1jNHl+mLGeV0zHxk82+smdQwS2jFgfefu6oOBp66k
LDEhy7DvESaSZ3ef9+g0zby0hcONTAS9B1gRTpZ0bQcXMItP2YFJB0kByfMxonLj
dyJBYY/lx5hHgG61Ahf7/BL99ZN54aaIgm1njfnM93kcRRiIzFjAo56ES0qyuiYm
KAtIsIT7yyBlTXVqtBXzE4dKiGjT88g+1szofNiuesmzJPrdEXyvoNRZP38anp+p
WTy5CKTzuOhNlSg+DFOvrsPAPH2foVoOYhCjhccBScbkDJuYSF5CYP3YNvnCm64Y
4uvWvaTUtd/KRWkxOqLt64KKkW0uzIL2Qx1tpEiHIOKPkMxQ0I2uWq90DJt77teF
sk/ifxOibg0s7OYpsaXG3fUmNtnlz0Sh91I2wM/449ojiExJhUQU+Gd0WZotahae
LM42JIBU5FFu2pf0Dqj3wpn7/n8cjvvUE/Zu0f35dZUBadNHNXjy3OqlTVGR5ATd
9mPz4EZy3iaYrGRVzp87gEqzH0lC1Kngg/spSFhOj2w+jvyoqGkVTXTzJbqiTo2O
ysEsIoZCBJbzCl/7FfDIFl0oWaQ6vFRL2SJaB6w+TNlct6jY8mRV3caTenbYMMBP
Z12Kc6YOP1Bu3ebD2TY/yW2+nFZh5nMCJTO53K0kfnsvUxTL484Cui1IMa46UtEf
MO1F0uOCiZYsUk+duvWPvtdg5JI6Ya3mtUPdl0KrTeRhrJcWd9+ITorZxhStSlOe
zvJhPTwLMidkCqAVPk/Q0Zl3X0qjSaHRW6V7j/y0Nmu2xF7lMlI/96z8o2RsxrBT
QBpwMRedSjlPX9ipKSK+eLDQk1zZaocMGl/TisncSd+A2c+TdRBSJCG7PnZu8DOU
uzq0ggo3yudM+NUR/tc3Zu4AoQOZl8IIo8cELuKGpvDLWvMw4ZrlRavHr0EWaAIt
+DzWmHeW5ReAkCok5TBSwz91+AP+/YTSKTBv5OZF00vFeuhJt6/Pz+0D32WlZVe/
oMyo/O6TNj9t9VaPWXhg84MuGx7xq6BdmxNZl2o5a33TdclgsnS6Oy8bHfzDNkGe
TNSHNbbIHfhGTJ8b081R5dZa1APgZs7ZMnv2bPyz/+Zt3AqnEV6wljzd058jzLBS
RnvOgo4/rjIsmausoDii6tovAH3IRCcbHVXb/0K3tV9zUSLDAk5xkcNoy5gp+GBY
6bi5Dr8q8Xho3JPESnsDDDEu28wAaf7O4g1QFJXX5kQ6j+Tdw181bDXC6f/09iAP
iB7rUppyadRrPd62YJgKV/EvPR+QN9J838wLkaZuJnsJPpJ7LQQ5m02bkz9VCLTt
lo+B8E6xwuWV7A40/084oxlUG0pGruu3EW48uG56qywnnxK5u0T9Gr+Ted6zR0Ai
GeoF9pwdaaHq8/AT8EqN2cbnuKFvD/frqyn+dosBsDTBy7l8MRIwmhlNh5MU5doL
/C0EbPd+QWJIZraXT+b7/3soLKsMBsaWFBX88/auDxYWnK8e5jbLmkpabh+STG2k
xmvGZ3Ju4ZGM6O0VbOVtx2EbkVXBcCtfpIvedzVKjFqy9QOIDGLmTNsNEq4b3533
4aS78d4X3tO+4ZQWVVn+tcVgBrIPjbK2MqWKnf7nZ7swbdvKafgW0TbxkXvHpKUs
VRm8u9VrJ4lsxBTPCa3/PA255ZbnRpvhOz6qNL6ocnWUWYz2ttAtot2igYspiO98
dxZjXJklEcQOUSHmar8sh/iQ9O9Lbj8uIOLArC4sjoWEsbBn2HmfpxnQW8HxYZ1e
wKK6wjdUADzQ7rdt+PK31q0KEKx53YjQeq1ZJRASc87JiQdvolJQvh6erevwVz1o
94FXaDpLgrD3RlI5iKzUuCyFXje98xfItxtmisW5l5yR8CfJo/4sBpFDbzhh1mAH
DFVh3Gda8HV2I0AhEsxbq+qwtqTRKM/SZXSJu0wbk8bsNKqbqiaepmzgRl+6IrfP
pxL/v98F5tGuPs9DMehy68TlJd9Fy4qWw/3rEa3GMK8zDiSIcCmYhoEjx8qCrCUU
kT8xlmYFA7RYLaHNxU434r7ommL//DyCzfhycawd5A0QHEoMkgZ9xQ4kIiLUSo5C
P1EU9f8d0yYLJLFEmRUKsSXCsxBYzHTCjYevM9N0slOjzm+A++70XfA1AxyCeIKT
dxE3hzSjgEocL6YpCM9kakhse2fp2yhcLUToHYaRocSCH1qLiIUGWaokk0nx4OyU
ajLfjHsVhO/oYDazZPzXpVdpavAdOv2kBA+5x6Ew4FaENTGuwRgUe5XoC7wVjzlt
Pvk9AYCrgTyg83EpkW3BxxI+85helxcvPUzCO8PMjHeN1h1E2hTAOqdQfOJbkMRH
SPp2ZyxLOy2974CU+VUY6Yo8Mqa7ZaeCRSPcTg7xooVsuag1P6G0IrCjRjZRF5zj
elyTo7oHBAZWx9z4rmlqiyxe1IjduI0LD0K2lH3W7Zg9zvXgtMXMkx2dMsweiY8Q
3h4kghTa1Z0b4AhimlB22tlnOtYQ9zjpU1W9D1fALGX0EcCu0+lyTq96J2niKi9X
KfnQloIIfyZAJTVv8noauqLkoCgOz99dP0SHNbS40Zb6k3cOp75LSbRtACjFmniF
/Iki/gpKMfrVhrP7/SU+iWHCuPMswV48HR5YzWv5AgbkCBQ0WkpnMxiaWVxw2bcL
aWvWSnOnAGktjPMovLJUXuRNAI+n63YRiyze4cXjI51NppqpoWPi45zGN99loVA2
XvIVG/FpYDHw5P6rWKkHgeNz8fZLyT2LDZOjinp4L/7X5hjrql/4rMhkDKn2/Tm8
OPlFmDyvbj/91OM+DCirG5l02l3ibPvm8GzZFCTEhzNZOkpioaKKvp9amDlWEDZY
o0ZFXkzWVc7rvH2zlc0LEdBqHFIvj9zzlapq4KHZzchAo06zC1cOdNjqcVWoUOUb
dT5DIDHckb0WbMburWNhSS1B44o2OadhQ0bjFpg4J51UiXiFdV/HJNc2EtnJtoBx
eWQuTlx5xap/2Mlc2tsqEzJ0AX50zT7GV3POAueZiVuee9uUeFFucv5C5n4H25fy
Owe++EHI72F99QdGOalHWeixzwS30MvxQfWRkXqQMtFJdw6d+WFBuenuCGPHQzyV
hfhWRdAjnXApOlKYcuWlM4uw9PgKhI7fY6mgU4ub0bhEK82vGRqpKtXiMOabh7ph
hQz/PmhV+8otV7GGyTrLKFLbtj31LcGlNrWnNkELK5qYxEaEWldED3Knd0HSp/25
DW1QSJMLmDXI4t/0U+gMbC+Q/F/AA1toOfnzCvA641HW6M6zWOlwPA5DnHNHfqXF
Xl8gXP7eoCaQ/Ow1id8BB9Hw2ML2ZlbbU9tJnbirirWYjUr0LblVouD/glsVgryP
UdsTslYOPZhbkGaSVn/mW7NFG0MYopvnKlBouAL+BOz4n9jj/1Hl5fmbQVgF8occ
f0Y6ANRa4n4m+SoB9Yj086383Qz6mNWgN8RXpN97SI311JbC2uUH0JU4bw7M8tcj
uBn2pvR83XvM8rwvmqTWLDD/HoYKdMqItVvbWqRHDlpZbyyNolCRi5TgOhQp1yT3
xOAtmunbUSr/H5yYjaT6AK80bL2YI6+A290L/l/ej5eG9ORCq+mRemvYLKktjEua
a/mXZuTHMbhNg8AYeeVr+d++rWH7z3CZlQoU2Bes3Suc0PIZXC5UU4/oF0ArFvlD
axkQUTumtRW5juWQ+lZVsgAhrQL4g37ZvEuArJMXTBSTJfv5KeqrRYFxFlt0Imdg
magfkh5f23mGHz2WD96k/D3PA5sjG7ovetRUWxiPyoM7Dne2nlCuz39OSgVbK2o4
XeXpmK6e/PB/jqCI6UJticvU5DRwTrXEpmc7H0GpZhq/AU/RmV9E0gYtffVeBJJB
rnV/QEUSsLKLWnacOoo+Na/N2S/MrODEPnqhtsaouhmUnQGA2ZRAoOcHJ5i/1Uv8
txzt04TNoJ8DX8+6u7PFhhVVdxOPfKPIcASj9IGiaUMdZqoz6AFYBqMSMlFV+Kni
lfOWiDSrZS7s4svg3A85zDHDgGOJX5zxmU/3H3aN+RvafejiAzZ7kIkvSQ3wv2KI
jdKQ0WTP0+9PJj9sPAau35EzAp459Pt10BOMvH5vbBAPntm0imWVYYjNjljhDshv
wl1F5wJxHis1Tv09ZFmsxlIK3cTqmLlpr+gQhD5HfG0QJzDUSa78RRLkPMJ+XIVV
DTsqxNosUrs8gEwMXlUsJEYn6UUdfRUFgtG4KL5+CoABj3bc9B485ALeka4HDkog
jSXti3+KCXUlm0VXjy1vomSGicIsE5ic2XyQyQUM9j4iocYwZKyIM8hlSxeErrAP
qnUnToouk5WqQu18LfbV8LyX65tP3GQ4XDiUM4pvJaX9Y5fipqyklSymTF/ZWKYa
Ngl3XpP73Fa/StYF8V0mF0F5IlB2xQTifEIm6ehr1CztsJ+VqF/6A5sL6E5kLtRC
WBBjZnlnOg6mcqH+8hPbF7KRaVGjeNvRyKgFOhaQwqnUxIH57urTAeNjtxiVUjzE
h3YgWES9mtW2FMVZ+SX68n/t7r8Zad2Lv99N1LWgif1VloBhEEGf+UGQP9q3l17G
PI4FRLjcbCE3tzfYkvwSSewVoiruYcjD5+4XoQb7ZgaKcYLhxVQR4eDkos3Ic61f
9aro9OpNho4zA3BYtmuZWf7K5A4M4LwE/ldjrPSVGSU6+xY8lwdVr5AZPMhR16vN
NFkqjrywrHHZo4AN7JcprGVhRX8Ro/01FLi+wwdx3t36TqL2+Mi1+U254e4oZpJJ
U51Z+ETrKOpJnQDkg5TC4KAaz4JsSnRDMgroBh9zcyqCSWmQ7CEGQklPUnogwrLg
/kKAYkZDcWp3WUR2+2r91S0GfzanMyeLg3oFAQqxPH2PaWifhTyEGKTPBewCFBJt
0e23Poe1gWTnNCuXKz8QS/dd09Ssp8eb3J7p89AtVlGa6/b3SxI/0MlupKpSqptc
QJvJb6IOYMqn9SrI7JKGUVyWdKUFPzCd8jAofEzHE5VzwBVDWRLP7N9Rawyx3IXE
UWjEjc72LUR0QIlBqW5drASjCbz2kbGv+b2nyq07lDYp0mhRf6z3PxVYbuoU5PhD
vn6q9OirSYjppj/MLiBvRvVbiM7d+Mi0mPt2UzivvtMEt8y6qVN6qKL2v68IxNWM
+7OM4kb9UtdoGloOAvHHK1ZiOOZeLo2XtA321bpT3rDOPXz+TKPIck9tz67OWqrr
w2xNtGQQw9rtLQSl9XUVDQFF0W1GMK4duoOt5TguMMWfEyDdB7i7ZvqJyP1HhCKE
lJX44+EWRDr719OHlrvVFVIDqAJFBKlRS+4poRct28v+l5Ge7QwlIyMmBJx1o2yq
bAr5NkfrbL40KTg/UygzqvnducV1678WvO79y3kc65ajYZy/6itR9WEkYqJ9y/Sp
qppuhA6PyRMjuChzZovGdH2SMUhztQWo0h9/H6bAN9YjThDwokaARoAD6Nd7iwhr
blj88qBzEdlB+k0byE+aRbKpymEoWcLT2leLi4kubOOG0Exz8fzyCA/QHbgQD5Tm
4NBbbUbQ/B/3W7NSpzRmylzsHomtLZXA23paN1Fmtkwr5yb9WTALhzgihmWkCmUA
rSFz//O/b3k6n/iHcT5X2aklI7ECSg1iZCSlYPtDW1HX/53IV8lnnzvhDORFo10N
MckhkW/MtXW0k7Jf3O0Oi3qa4SY2qtkiyNh32OTmmj+zce7iQsdEy50aytuU84Nb
fjYmDwVFWuaoQQG8Zy+FibB5hNeqPPINE0P4M7/HatXTDiBHRF50uZZFGX8JXMuf
h/6N5dos9WtEeWJC1eVwRH/yyiw7XhNj5fnFHPu8IrAiJY5O3cQWXIXrvN3MDLeZ
02KzNMBFZQIRzF6FonPwk2a0lxCFXDW7Q6RRcCvblFxTUQ0EDEVRH3Wsap8TdKXM
fptZ6BxKag1vhKTTguk8G1AEmKTV5L6380yHaldJHOOjEtWVpvowdBmSDa0cJ0Ui
k9yVbL70G14MHWNQterazN3M8RSb50vEHNEwh1TiqxEStQicVKhaoVw5PM10CZnd
7pttc9igTefiCBIOlXJyxVCvqk2wKCalidfP4H8XgenXL5i/JzuRXd7NhEaQzhGk
z9lveoMMJbouMdC63fSWS7p/S7ZKL/NDePUA1VDhqezcT6cSLclZy58x7da6h+oh
RRfgdXBzmrFLAHiKKQNoTAKvKg3H91bEry2sLMQUhISzqnu7myXhv23S57hZxyaa
tTjfLpFhCToymIQXEluYkq/Mc9q5WThieUivceoKHfdQHt4Hvhj+7LWT6/Z5shiV
OkTgGiwa3ChWKpQItjvICqWYjBs4mf5q6WKZ7D0UV7XBWlk3SQU+twXiMctsw/2h
Zeo1INq4xmQIS0qIJglThRrRgjii+aWPLooAoA6MrnDTNGcpT7RCNOsaQ6ZMH35u
7uhCWQJb08RU2Tc8r1tdrRJ4z4/gIavxLJV93+FMY7l8WdCyjeLGk994hVPZ5pry
CnZQhLm4Quvx/78u4w+9QeToWHbbZAAHFzutW6ZAxHrKr3oW1Xh7rRJC3a1Dhnfw
BVSul45LhI3GuMiNnjW2Jf2xmUcT+1/uFgWh0OZdx4WK/QYNTokkhm4hGUCj9ZkH
SrYgEcVdeCAwmZRj/p9RV4OuquR3e1vMJLz57r45FGkJgvXatlIB7o/K870isUtU
IeEM5qeEGc2PGi4WFsqZJqszkntBNuS1WGEnDsTnaXuLa1vzse20Xh9+nxgTssmy
+cX2rnveuBgpcpYs7d7a9/XAt2YV0+PO6mqV1Jie76zwElClR872t9NwtgQiTVxM
nG3VuSPvCBujwk36Zm++LHiaK7GAea8nxxNJemRWkPySF6y/Z2AgbFysrp50EkTc
DkxpivUw15lEMkR4pcdXYECf9nYhphR33AW1538pZCZIk+dD8DuwJVc2qahVdQ0K
o4BK04v8j9KDGwwD4a7msWvHi3KYDt5XEcXyVQD7TKwCyrWN+oCo8cd4d9sAFiDU
f+Mq/4hEXBDbj8MenBB5kedkc31FZhlw/ax78vp/K7bp30/gnjdoF4WKHvXyKx8/
KSVmBgIn2IXTAyysp8lk4pQwfzqRJMHQWf2GFy0De7+Qg5MunBg0/YI/bSvVaANc
CiMp+gjESitzX1c6uQY4cFDyIPOB5FNiuZ+3FjqYt/VYnqRhpLqSDecgN3dUBOH6
ZttwMyAvK5uq+5Z6zQ2g5sctUz+fFLO50JAzOZkQnUkm5tIN/Z2kukKcxxfB4eq6
/8toZIAElL5esl/h/QY2QDUNJoqcYOaPc+/H49/Uap1rrqPPv77/c2LvJb3RiEcK
ra5XKUItEnDOaxU3Jt5ZU4s34pmh7TpacXELYlNMcNpzF9lu4cwDJwe4SABV6Q7e
DyKzvhUDh0jmojeimoOvSgiGZv9v4s2GaEbretOxGg148Y6KO5kCmKkQG6zFNW0V
4QMs465yPmpH4XoapwLTVHSmQ60px1KefID5mNzKKwFLIegIb2OcA5WErWWneo9f
4qwFK3Y/uVWrDuucx3ppFoL4Zxx4XOrsXDD8KW2Oae7rMY2wwnyUee7geN07zgQ/
X9cw75ImgeyfcFUwgff8yA9PcNhD+34zwos2xHCrwAoGvr/Ux+GZC2ax0sV72hVx
3FsJOv5JHzw530kQUDK8WvuNwf/7xoGIQP+6oaHQZpJrm9PHERBI2gWPDLbBm2QQ
EErvcPCnutr4eEMbXXgg2IkuQnPZNME2mBP2mINfixPpU94uah57/rH413uYd5rk
DA40i0mGKGNirOqfnmy48IlcmcKbwhjw4dvwKd0MK7pFENJVFJW4hVLuALF3/XNq
ciffoRVqyOF/1EYSFasgtEmuSxngVESe6dz5BCl9h5pffjPZ3eTFAk0E+eBo/Rte
7eM7zCrUmWSOw7kpFnf5G8GbhEZUYsXuo/lIpMpHytgDHyanp37H1R9Z5Lbv4kwA
4yy7VYl4SgjrIJkEv7o/McFeLZqvKAaoXI7bqnObtyk/R7gd+jpRDx5y51nMdx0e
4GdGH5fHoUp0ZPJPpt4fkmQ4X1Vn1ESN+YY8wjqD631yfDl0UcLWZ4cOL8sO28a9
dHb9JXOpKU0Ktn7Rv2xZ+vjkyIUm2PieiEP9Ze0WtN5eQ/KprLWQ5stau4rOGJkf
QwfB5wWQVRqsRqSW761i0JfUQ/V+9w8BqUYxHasgs7hZAmV8ngEnRY5iz98ulAA4
vY1HfaBrfTAhPqEqXb8Y9aFVXakV3kGUGW5+5nJKX6XxF7YxBLq3Ycouj6VhUhYq
+wNquXaDtJzcYo95gcpFg+0rOSQOYm9nYxCwA6s5D0eaw22Pi4G5TV5KRpXA/pGH
4/Bra0UMSOnZO07RsMbjaGN5nDNyDISUW8H/oZX2VjFDIAYDML4LnPDU5NlPlNYi
IB5VI8A0x9auYWLrlV2daglZxb2XtK4+8uGyjkiG39KTxRDYadj1L1qTw0J3I/c2
wq5lgicgFZkMkvvtsKOggxLZkOL9wJ66k1mCL2oXdGcWigYZduTU5e/rOWoLZ85j
NO2C1DaEtsuyXN8+/tfmDe/huEKzWLyP5+Jh6SDPlili+FWSkIZX0VOWTwmMm/m1
BGatovepbQ5Im1diPKw9h2g9YsSw1ankWwTUCU1wJniY3ypJO6f1rIitpQeGCh9M
S4ChemLZkVdMkf1bT+aMNKDJ0JeOrFy9raWFGJuj5S8otRHAIquNhn9BLK4DKEMv
rMWPlY5hXWoou6eu4Q/xOXTfYq781NJywXp7UVf7PLCCcvQsWECKR9UwZj/rTAhS
sXP4r9VCxBGMIb1VID6vwi58kfrQ4TVifTSmoE5KxrcLkuT43e+4corB7liR85b7
7axcZnatFo3CEa8jr/X9gc85X9VUC7xDHzPmIjYmp+EK0AVZYRoOdQyGuKHaDVo8
Yhhz9OwJQ8FvZFGf3TXp5GJVEX+xjN/lXPrdlfX12pirK6uERVDLAbpmS4SefMVM
LgGFl0Pu2Z5QIf7hvAnAui9QbnIzPK1rP4k1lbsXoN/iaE6JKCPPz3xYhbh6P3Ep
vKT40OhYwyDkda9daygo9kUoF8l4pvkFb1+s/KVeKg3aORarbrq8YBcXTJajTToT
2GVknopskIbXUCmKufeqjLLIJ9j2a5/kSVp79ehikbBoKcefvGplNRiMHzgMQ3ly
aKGbJ8awvUeDizQks9CUuT0AffE1Kbis6QQsVk2uokjiFlOuDHvZOoDVeDZdVlS9
LR1r7CS/Zqe2YqyTquqFYimzdYzNHHK5xDoyEOOvB75FT//V5SKqFcWzwzEF3H8f
EnKcnEvngLDodvgsDvenlCAMD9ZpWzLEgcfh6DrmjL9HmJfoy2MRB0qjbT4e6p/0
/FhGGb0yYIPvsUslZgCqMfY0AzRiYP4iW8RVMn2v4uSqZq+wc8S4Uj4C7vG/RJi7
o1EhRjOZneFf+L/pwr2jJq6q3nIfvjZqozra4w1/dB9jFdP9Kg19q4sX7ge9q/Dc
1mQ4pGr+JQcCrrAnhuEsEHhPSQqssd0rp/RCIlpzxsPHYKhEQWxtOIa3B0qPT8x4
ZI3IljPfsp8HyB4Tp+0GH3XGbLmKVcU1GVJD8ZDw79xervfq/q5VX9zS+Db/GSza
G7SFg/9BErw42wyR7IyAFCZ8F5IbuTt/i50jCDKNfISogU7diUdZ5xlcn4zzMK5j
O6qoHP7fLDCIIxJcybLRHM1N0g/+3efunnUpyeXBADdUejTpBH7CO1BXaQ1ZKxSK
cS4w2EmJGPjIbz42+UYbgE9StQ2mMtGUyl703PQN9u9HcJr/VDmLCFZtFsS/XAkC
BQ8kruve3ywvHHjV6KnkSwobpPZhthocxdLLwWVHDFgth1vdfOPttwCcvNsTjXvd
X0f20TvWfLU1ojiP3BRxolR+tAk0P5WIsVnu9qihNaFWx7VFEt7JQcbSYsyPJf56
S5lj/x7jV+jL9L/sW0dQeQF9UrmEaFOQ8zNa/1VzyHwp2Tv4SkV0kDk0JmkBBWjT
+P2Jo1JtcXcJuobVnQRUJPzVNhfyrFmaDWSaEshSbX0D1SkjXsHVqvldpoYNDZ6Z
smvaTHuPUFVMq01miSpfL7iBdsX9jpZGbgo3RSH7pKag0ofH7Y5nGZnKhE5i7OLo
TFgXxv9TmQv7nt7fYJ9qWWZO2CpH7s+tdU+I4W0PmGEED3EtedxpMmLLCsFfaZz4
H/rD4HxAljLkND8f+Td0UYOLz0SMI1QbJqVoyR52n4KSQ3Hg50JsA8l6OVS/SqzT
7a9lBZzYd4/tJ5w7EAGvprh7eMPwNIbDUNFjYhUm/lCPXbi0G9T2WU/0zY0raYUA
BJPpPBni1ANCbJs6dJaqyUSUZQbBETIakAo3D5YxL+gdSnJ83/DP3hyQdze67XcE
k4NNXcfe0SJhQNtv1ZVH6trHh/blqbdMxNPU/GSpw+H+pYvKeE/YOITGYdRVcI0m
JCZlO0zSoNkN2eHs22pI21sodLTQWQvmbg64+MXCfOCC5d249nj0CqxH0wsInnMo
EmDazSOi/3k9t/57D0YaUi17WyQhPqVshBkfE0CsiNNnYZ/q3d2fatP1g5V7wDr1
FoiaSN34dNV3m8fJL15HGXkoO+GztucSmib0Hea/R3DvGRNAtCMhkgZu7wbcokX5
qLU+XhbhckR5xSIPx/QC3fZyE6oAEbRfmS7ELJdQMa3q5UCPYAp0jIMQJ70oSR3d
EC4PrIwnwKH1dJfekfa8EXRK/2AMpk/hBro8a1mw8CMgDTZo/cVwGATIRazvLOGi
hqPWw2qP7ENSDLlWE8+ULWrAzPNek5Bd881e5eMN8F1ms+5NT9xrOjGSw2BUHXwN
zAtS0RRHJhV9RhDfK+frV93D3NsLuUchMDHhPWlM6nsGLVw8skx2yShdtaCX+YbR
h77T7GB6wXmCTFnnvoza6ygbu+uD4B8u4isRQZq/wOWUwpdiFD25mELBUDxdPGvV
PntwC4netOUMJXLyU0rsXzwiG3PDcOB+5DneyWjzVaKqngbTxSeAyevLmtBoU71K
1sqisAzm3DbYE8GQtWcQ85xztbhHOoBENm5Q/xlZOD4Tm09YOQOm9YHrzZUeVjJb
MWUdL+b15xU4ISCnnVm3JugLS5booqA1xIRfAQqvrlp/d/b022CyT4hOooHHNtUp
n5RunSi3z+IbPwvHhku7C/1g+y/for+VAGbD/cs7shFLy/B41LNzSzWhV0fbqxxe
X8H8WltQudWKZWZJazZ4lcbyGyyTZponRkwbcY/Uy2MAhOQLchYHoJHWRk7whE+I
DX1/HUJ2rwOrfpOrVF6dq1hHWWEIjmcPlqRMcnD50oaXevqn92iq5i8tcjW4TDsD
dWsR5NfXScUTNraiEaXOoV/IJtYnoA+702W8IXQ0sd0ECahM4z1u9LH3ZJyAvM7L
E2GWD7WEXWzPf8V76IJjk6mXVh2TchrT3AwKCg/p50ZZseiLhI3SyqhoQKSWdCou
JiFoWvUpvRxsnbZMpClj3uzYtcyf/SoWBaaA7E7l7882BY4DsI223wmAYvxSGRn4
wVnSFdrkaUcH8cSxyd3atzPB/Lvt2vLPtAXlCot7BOEJNQU4AtRykT9DFugx48hS
VtFXsiMnaL4w+aiL64JWwYnRQvHtr+ARkOJDtwe3rZ1rciQrG/Cc4YptcElLbtGP
e3gxlLHR0Ei9cGHDpwVDhx69Q+WXZ3jEQxjkjNrivcVLTmT4rE+jIx2sfVqNq+30
V4oztCnwmLWRI9HQTtCI/GNf1UCalkqQesJe38igdAjxEITV87IQvK/5W0Bb6fMJ
hOOyiLNxMOhCjJLmKpVk3sP6UQcx8iNnlFYHa3tqJ7HMXV2MxI14+N/FShS6IJcX
pbrzfIiWRqnwiq/OM8Rw0+lkPHlfYGyfJPeSnvsTF9yP4a9NMxgSP4Mui7znBSW+
9BOZ7KdGP/AsVy6RS1wizhQPNd8c12z+bZfSKHA5CaeNUT+2ptdAWgckFg1Lbm5R
iyg4DjMjofI16no3O/svHNq8cnonYD+jwlfMB/kSz7mZUO7IC7s7j890Ix3kf/4V
M2gcejrejH8c0tej9MlRJpQD7M707GQuRTBTwotQsqr43xJ67lFxFpP1K9ncB7Dx
1vn43F4VkPa2LEL9eSJyf3kWUGBpqGhD64LXDUgjUzlMs/BH342UXtwhR8wlYvaI
VWxdk5BMDkTof8b8or7hfg9LNvXhC8H8MNwUb8uarc/KG3bf4FXnkZVUV2n/kQ5S
pKYKXGrRj8k6Zo1chUeRT17dGD6LZms0pOxG/Y5d3QbEO7t8ox0DiDDUBTg8tLs/
+e8eak2kQ5x8BZAVhoOG7HQ3lFUX/cQlhxgAUWoe6Y7syXb3vSP74wU7H5i7hUuV
VkZlaSSp3+1VoEs7jdWqBO21w/2i2jEsgMyfq7CDQvQFpfQ6V8qavBp1PKFrc5zI
Qm7MSyXMG5LOsceXmwI4yVodgSJbh4e3szzYFoOsuG1MVux860OqD7mWz4ZSje+k
84bze+negZK+Y/rEdoHKELyh0GHWhqqHVLoufM6C4ma2i5x5aRLrlGPPMLrBzhC1
Ta66f5zpEgKCsOlqCuZZL8ts5x0KhixzIIeFuWfDBXWPjohgxcaAifdhEOw20A2Y
yC+kVlFvbYroG830Yrw9xXrN0e0kzxaVMS7pBrQLEEn+YfSSfzdmt7BeS+RSeHjj
FtrR3bJglsnwImJRdAJxgZqDQAOt+YCutz1Wm6w+Ut8O694/l3JCHEEurrmErBdR
ljJTjmBDCdBtRYFR6KVZOghRYbFQMfPIbsRo1ZQ1tUd1ASKOPqGy0iUY8/1Tt1P/
oVxqdhNTm0fgVr0LFZDSaorr2JUeGIEkxUjWPpbbVnI7xr1eofUcoMAOHVAvvp2g
WOGwW24aL7/0EkpTzPs8LOqYkVp2ftv8pn+zMbZr53EgPZ9qg5afVXDyXL8FX1NY
eBxRirVvwLVZYrKRvS1eQ/VPbOzTouKJZxgrkxzpHWEjymtK/ZkzFckoKMvylbsu
iXVFcSGWCG7Aiacc9bBVOFMpyt5Ou4P1/ylQ51HCUDjYsaPNiu1BQdCnKid4YQS5
s+dgL3RIXfO0QBkyb4F6bmX+kH9KJthCc4kDDnZ67QU0qyrP7JIidsamc6srwwCy
mnsX1xqcMtW+DBsOWtR/8B/AmCCiO4G+H6C0E5PLwp42OSbjDeBHj1gQSy9deRdT
E9jRA5gXcW5c1T7n8tq7KDewKlpK2iaGfUV+EsnBDECg3Kmzt2HgxduTUUCHv0YF
00xryaCBiMg+6f3u9KIQAwtYybLYKGcCjzNRLuJI+iYc2A1e7H0UYTWHyCO7ncy3
xybKUham/ustmBbkAqCuPl3/CeUeKpObI/Brcun42Wd5zHiIU+jI02ytjt2Bum0x
36Q7J6hxaFOgySsscv7sqfJbJbf9tBvwVWjDPL9W06UD97ayz/R4ClI6k0ZVSxZc
fK4pQSE0g1NpYNH266mnHSBNmBDpOQhI6bh7em+IxrrO5/5l+HCcXpJFij3Er6O6
srxasOyP7+rAUC/3OM7PGoe0E48lCLvyrWtlq3ZkCBGM29pMmkvDR/3v1mFKJVBb
8FAogM1b+kOyL3pAQZzutyxUUoh2LR9m/mH7aIKKvjKSa+PTn6ziNOmwNYYNP9w0
8RPkxvjybed6e8tqUb4GH0MJM4Stu+x7aud+4PCeU9NJuqNrx6JxOaAANndIUj3j
LWWkj7VjfvJswjf7DOg1AvPtGtRgpz0SPT2Zx+0D1GuHij4tP5Xur37C7s+nuNUb
u+m/dBucy8vohhy+fxuiJzj29GbR1dLmJbGP3QTMmL3aqL+PitjKvRsfc0620PHq
c45jCA8d4TCh9O2xgbYbzS/NEQzUq/6tmyuvq8qQSrXpGchPRp747S7CKsxt9H7u
msFkb7XAi6pNFRCPsaBLNZ+QYDX9OvzVZgK/PJogF+DMXlgStUvC7x5fRzeCUrTT
I+8UVWtd1dQFBdR1UptliPGIiWdeMbp94z3j1EErEf1vn8TOFPBV4hUVl1t7MTUI
YX9HiHQhkCU8x+ebuyIbqbxC32sA35xt7H+oq2/0CBbjCz+l4BVMB7urz0eS/C7U
oZkpGzHa/eYyWZkEqMnno9w0Q62RvZNe6c2r2FZ0W4q8LlQS8ML84zm6NnZGwyiF
SvGqO3bf+sJ6kEBkNR04zL5oqDJpa19Uj6UJ0OZi0eMyI22f9npLeqAwHw5af/Zc
S4fsOP5jBhiNiPu4uMviQUcr3zwyA8GtiNHWXhTAE2lNdFVkpkm1MaUa3cQXpBOu
vSAopjopGzWdXcpNuBQ8c1FJNHI1pM5da5fNhIrp5SldJrxYIQBHZM2347RdqdNK
cxG9ADx5OVdo5qQFV1jnGV8W77xn6a7AgYXCnEPVgYw3LDJykrOprE9V5j9SmcN3
olDVQeeLbc/1vtMIUtUkIK13OL/PiRHpa5LVNUZ2a/why+dAb6fY6G6lAlupmCjD
nOlQdv7Od4RxjeGghqOwh+01skCuVPqNjSECxUHLl3aYN0s+DFV3sNMG3fD/OooE
whMadQPK5ydGLWqho4UAW+NzsfVSQMtfYujAHlucgXEed30aipA7NbD9PqeUWUR/
Lvz/oZ+vJ8IhyODxZ0gzp+1pRIC6PGvEe3rn9o5D6TmszNAZhoCPA9J7WGv7N89s
8MUeHJrEgHYtF+/SDFEl0E+DOQgqJp5KL8IThe838zosVyJjmXJ29s5yuigvO3/g
1qewAwTrdm4DZeL+YYYfUhmIA6b6w+j03JtUpZHS74W1srAqmpp6H5hMAvriTrml
YCdce5NvcsvKjE2hUvl32N5BoGWSm8BCcKy1HUXhnYARr5wYLORrTomJuVz+hQiZ
PETdY1NVar5L9UGNjvlHAGybOXyAE77mTJxr0XD9KpbnLps+ELmnyyOMn14T3pUO
SMRtLA5m0vsbbyxmltIQRyeo8fSadSRuSce9Uba84hsSEbis0uB5fv3FoRWsPA1N
PdfWOIlgEo9APW/qrtzKVKXERQZ8mVXkEWPQ4b3GYPgT1Hh65V/PfII6ILVX5B/g
PsMd7y0E30f5xwM/he4Ik08M0J2+Ds0dbSJ5SDzaANyqoMAgN1teDH6n8mGCns8H
cDX2Fd/IQxBMjWoQNNdK5UUXn5l1C25Dt5iWml4uFo2vxsTAg/9ZnP3HMv1Fif5E
8GHMxHzDYIR4wzT/7Qvpw5uBkD1Dfo8RfYfOKa7JS4+dPcNsIC2VDTw1o7dDkApy
h8ZE8moeq09j5wfPynRKRJFYRFxWu69/BHPzQzEMC5Lx3ELDYYnbDbswEsgPZDgk
lVFSxOhpES1n2BNSav5ivaeR16qoupjy7peyfDA/8r2NNzGJLeasu7X0FOATNOBD
6EcxHW15ipNA5Y5YQ0W1D1X4vUc/ocyKjM7wn0bN1FDTfVrANFjgCPE/s12v3YHk
ZVlXOpM55t4Stv2dHM74FU2tDzG7LqjPEb7ka0tidvv0QWiYSIdZaO7ufZiFhS3X
zycHHe0YKgUEiKglktkmD0/+WWmRGqgDKrgLUbX3uIMNSt7ty3cePGGofOKtP1wF
Ef6QAf5/nbVhwGiRjhw64f7i0/bp9bXwH0UIb9UcFB5jhAyi4BXaBr6dtCTMPYew
7SR++PJlvEzvQkDh83GbXXPMqsgH9NCtDLyygZkwXpiMPH3SYt43ecuOtuBGPgHm
fdpVpnRcao1kW0BXB5CF+ge8VxK32gjgufWzKr7UMnqJg5o8BcVZ8qJErxRFtwKW
Lk4AK86bmuAIKae7eYWNjpUda9v5E5si3Y68QaVV5L/Letg3yY2aRXYprdgw9trv
7+y51ieJb0mMC6gghwr+EXLLYH9kTbxs3+nIBFdGXfNI2Xu9zblirmVcPj1a0G/S
W7+Ye572K/cO0zdba5EeSYCMvSuN5jKRfzyEDp8pWInXNWrsZGnTvphQMckZkhqi
LiiKrcmp4TCqnrD96R4iR4PyipULF5zEGI/iGXeK8hNNgjPvYdkaPnj3cIHLcX21
5mpz/JyiWCEEOFEpCQt4QexoG5fag0io5pGdPXuzkiguBraJUSqVu+vhWY2jOhCZ
LO2Z0bQyRTTLdf23fGVef7lVRL461pmklc4qc5of/fl02+iyiv+Di+v5rAzoATLJ
4gxUdH73xm5oNJ88Mkk37jvlQkk2EXbM8ZRTUKr/pLgVuygH1zdYpJ8HjjzifXZw
nrXFl+vx9VdF7OszRYTK4RZvhqQ2r/1wZuQy/zohMC2g0Za6y/CQzh2QHHKqjA5K
gzt1eY7rSYZaPSoMEeDCfDNHbkJ98+B569eueCyFJfhVU0mxCVfg8zbesPpdzTbB
tLB13WyiivzVu24yCTD0VWYbh+8h9lQqpR+dzgvxLlCj2bJ4LjiHe8kQwqvrjw6K
uDE6z12x8bNloHRmsJgn+jlCETR9TvJppHLV351O1Y+pPqBOYN3kfYZbv3ksn/pR
ACu2FOeqQoYljknT2oyOuiyuWebsoc80f55uqlmKedB/TcMehJmSu9wLLj0UpwOu
vxUnvxppmM0dutH1C5TdUtar3QhWibceU9ntXe66XVlk4pkIRTtFCv5DBJ50WeQi
KrLtmXgXOtkb6X6NtGFbp5ioXQyYddOL21HcWyNq2GSea293zktj/W9cL4nzOFtC
45yLkSXP4tV5A0B7k4ji17LXdohy0MARVLIhghLb40edLgiGfrOkmnBHvNGgUxhZ
bG1LyXe22hlaancHgdTRYuJf14F7gQkCNaDfjIr84CKW758UykrEZk8+pqZmODs2
MFCjY4/aqsYdi3+R02lRLr1TA8piTJNNSa0gywLL03iwD+Yxq03VHUDMIhP5/yhb
X6LvWvQz9bFpOBV0KcMyz7M9j6qbP8ZVGNzbFkkpiRA2LmIdJuhk1NlN+qDDzjXT
zHO+/ihgQWKWUmGA85U5muWAJPpbnW4ikPLYrmWHN0NLFLJGyGxZwbLHC/coNtyw
diQJk9PlVpdgZV4P9Jr0WvJZCI9FifbhMNa6UVvrGlPlyeadcWPLlfx8tYTsDs47
TxEmzk/so9VQtAUMI7skWMGBJqdh5vW8mxLIa5emNPJDmPJKaNFnLMD/z7WJUo+M
GEO4lx54z8P3kMb/f+h+525YUol7OZk34A+PNcN2kaH8Q3OQ6pzPpxXGMAv5qagC
YtfEh1p3dgdaxw+hFRbGnCoQ6++nC2IpvnNKvARcgRngrHbfm+1ph3cN1Ngc7FV1
DMzKO16DuXbqooud/Fi0KCDIhuD+saP+t/3FuCmiSfNa7trvIINogMNw//fpW+c/
TMihJg8isGyTlkPG41ZFSbq3J7Zx7kCj4ATn9ccoOWQlY850C1yNAqWyGLwtd3zq
RJs/7k61HH9yNEjh5mIWhGZR5rXevt78s6GdvY7pk9BhAQoO/t7J61klkhJu1kF1
5Xw8K26f8eLXtjIE5QWKBZNfP2TFh4OssFWt34JrZuca3PHyiYtCK+pfnCfYTLdh
wSTp0MjY5KwB/7xEgx436KrGLxCOg1DJLtZzQ0vxwfybB8J4SFpTCBY8KbwwEOOZ
PjEgdmhukWydCRhqovU3Vo5Vnzbw/ehUU0FCz9bfhXhQYqjxYbcRwzdURJ5D2Isk
dbLXgN6fI+gdJm2QaTHBE59cj24rY+tw/tvFtTOtAATwov/10/OlvRMYSPstT7+D
aLje+pPTCO5njG4DcoK+0ty7QnSTb+qmjFv38S9lSYlipYFAXR1Qy6i+0ktO65/W
8AO74u7DC+HEYSHS2d9+GRqXUKRK+DibUTl4Xi1+x1hhj3KNnTjQpZj8GPbilEGr
vw47P2EOb9X77ddMizwc9+khiD675oLQ1OXX6P4c7ub3lStoMotA7d3Gqa7sG5c6
FvxAL0G6GzQ8y3kLd9Qge+eZCQhckPwsVcrGEvMV10SAuRu9eq85JAwEZvhd1c3t
1+eXu4shq09VxKBY8jO+GKBBkwXmsP50GukewF5blvcRfmEVcYeFWw3+G5Iml9ZX
CYMvOIs4qRxHRgpul7HDd7j6fKDBmGEDo8m4cIMyRGComr/pzT5PFt8VTSR8oyBh
nabI2JOpgjsMUXrXyPF8Y2zsaQf/iOENj0gagxUfq3JPZD+4CiXll9U256jhXlaF
r1UySeY/OIOFN+TUJEUQpaVDX6Y9cgWyIOlC/ZvYxqbU5bUvGt8IXqnph8bp1Xlu
YcqrTcNO9Opqt2NCemFhwM7OGX/+jTL52c3ODjdjqZLY4xoIhPX+S6lZshEill1+
sy3PPVCFzMMSHIl02fnpUe58Oo/jJqXLJil07MUQGQprjvGVIAMYOtxRcGneFZW9
99Q/6MCyJ9QfyuVs0UnYAuNeZSNs2Sdt5T/dbnDxJzLJdC96PRH6Wdqh72tn9bjX
47wbXMCdh/hcA2D6l1BPXy72coQjd52ufvoZ0524lrGsV/2M+USL+e7z9ItA/uMf
TqlbcZj7ON03sxQvz3CL9MvrcR2G01Vil2WLaxkQs147pC3m7kTyATYS90CspEhG
ONrTmsEsRrVKtZseoY8jlqEblLTWwmbyR31Q6BKX+I8+vpie0ny+vamh8jHPnsMO
0f76rszyEzPpCwkE76EMMvNPcnZzLju+LnL+sMl29DMV3RqcsuSwIirT4CMFki1F
V2YoiigSSsr4UmENNn38s6BIjas9R7j44FEYBT33uraaBJ0Mby8YFMFMMiQ1cE64
QSzfaWBr2RanaLjBKd+Kp3A7UTmCMWWQ7RA1c7dZoZvbAtSXsRZ5ZDbpBBOE8Xbg
sRNuLSe1xcHQMfRktSP+P3dIVzGEA/2apuVqg1s/Nvw4urqZhGl6VRLE9+StKnLG
DFoKY3vACF31mXlQT0WfzMGj2r76CC+5KOXiNP8zCR9EAQK5lrIQHDm5ll5UOMsT
InX/Lr1TflRspwleEpWXgfMQKLLZ41Jul2A2KlTnxS7z3W4lwn8Yvfyb1a3ZE75G
CTob+sB0dlUcxxAeSTNuqqWxfvqd7agNQDFEH+SOa0vu1N7OI4nP77k+jzom5Meu
PJLBT8b4Gba+DZ4MyiDFgUCTlY897ghPQ0iuX3ALWYckK1wSuRkla0yu7P7l0/fk
w5kkukpFFY5wyjP2G/BjKBG1Ur4+MSCokupqdsFT/CO2ixIhtRogNPjK88lWnghf
jN2oSs02EMXT3YE/cxWGaPMbOcWDbx0SWGTcwM7lB+TI72t+oFm7aeJwAk12Mhl6
ilts6YrXrepj0IAcSBEuqZmEqULo83M8BlpOWfQg6kbb8wTFcsuUcDVlSj7gq5Xi
n8MgKZ5HENZkw4VGAT350KxLR7MmIvjUvy5MbwY34PEplATt6LdaYA8jSgGBasIQ
1+oPY6XGCY2a0iYcfFMUKcYPYIbaHX1AekqqfeMsUOKX+2cMEzkc9p+N6e0ai2aO
nIBDPHQoypN9Yf54vHc3ywKAriZRIJEXANVyZ9gr6v82JQwE7OKN8jBOtlettyAz
TN9dwybkGMA/605we/u8Icr4rHnLOvuaT9z3QgbqmQhzSWPRkdgNhUmDExvuPipC
pyJz4RycDJ556LQtH1VDgAzXSaIBQT6ybCLotGvdV6fm0D8iB7Hf2Gn4p45ws+/w
4Dwk9H+VM7YE0s1jztwvp1esEi6Be4iRVN3/qrgDPEPPL8NaHrIXWEx82Z7/8p0Q
4br83jT+EjmwfdrxOCy+FyghgjSSmdsUuRLh8y//c4FhotTZq22f7QiF9Nnxb4Il
eW3fHVk6dOW/TDGs2N26jCQO1E5mZKqgQRe9hLPyh/Hzr5JdmPHfshDwPG6iFEeC
saDdUO9wIXA5D7YmfGaZ9WM5/ALQckpd2E2ABHZM1KzNOhULsgj/+IpgO4fIREbk
4M2N30RcBNkP1iefBCK6PqS7+QMSBexPff4CW4Vu/Q9PSe0+vCbqd/xVOQjxVHS7
zZokphLHwctV/rV/DWpnBXixiSd/yAh+pvfA6fgJu4zjQ0nQTAmFsMlQrazCNRn1
MexDfNKdccjGMibCa9uHlE9HSOhmYVcy/1RbtMTTxCoyp21Hg4+15RVhXUaGgav6
FB/llV58hCo8KxjxfceJllb13CXQ200Lki8/7ClWVa7iADJ/TEWzSy6nY1Jw+Lhm
yQ2shaD82JxVc3gF8mMdGmG2X79FBkKA+tcU0SXPV1cC7jnPOsa6sYpD98mWqMK0
WYxWs8wr2tWZ4tdFk+xbVKa0EYSO/H23wIYiBcHgkmMskttB2VAJhkeGTf290R05
h56W0OJ/RbtJ8QGXxX2MZhA0XbgQb2yJ2R++/i737wORPgmtJvzWkUy72gMea5YK
++eMqsOTtSnDrpq2HwKZZmYV9lQf5zhj/iZCPhYb8if6Ej87VQZpiyEMQIk8aTjJ
4R6OHZtbc3N6pkIwvakMZ1eQySyV7dRG/FK/MWxEgbDiynWSwNlX8dzxZcgudoKq
//Vc3kWx0qPDlaEIIz/sVtpBvtW1f57qObKCIKbImL3hXIgNxbyk9htfiGQLA9jO
A1z/M0jXbBl94tFGt05oopPdB1bxDFBdEPlW13BtaxxspyXoqJZ43YRBtYzq7lwn
L+ZmFLYVwrxOzDdUAiW+/MREk5iEAu/pRwSsJNSwm25QuoaeJONlpwoAzGxscXV2
WaXvf67jbEa6FSuUeSF1RsVp1CfaN4Wig1Ju5eJ7tABF8Sdu6/NLFtkEDRBvNgK5
/bfrLje3LH7O76qfUFO6RHPmdSh05K6mkrj4vRtFwzetZr/2WPxhD3sLE3D+MLlv
0N5ZrI6gRPZ58Aa7E1Y37mBZhHqhdkHns0aDqx1c6xtfdkA32LwCDoSZkjXSDMeV
oYH0mta1Lp/2pPH/fjST0GK1G/vNniqP1JMslpeIiVGrCxIUjnXRog1X7kR2AftF
jEElLqM0KI5lyWJnli5dGJvqiDO/lTGfBnQE41T2iJsqeUhoizz57aSxLbNZg89V
cTq3u+YBlswSQAQF2Cer74bBnhLKe9uNR35Md9ETmxApJlK6EHEqwYrl6c1B7dp0
ZZEoI+rtV4neZ3vpHR7EHIJLaGJDaQFZw4cK2MtoqzL8e5bxGCPqQo8twmi8dJz9
PSThbQvYKcNQY5GQkIcIwU/TrNoyUXhRxucAsFJCzyUqEQYdTzyWAcm9VpA2y0ld
eEpfxMhPEYR6ycA3PYaRJ+9IGLjBeB+6s1P95cjLscwmQECDR2cvkZlW0bV296Xw
GoLA4ErNu9Ijf2H7/Alh7wMBssFpMgx4rhZvN1d6j8HRWbfSqar0x1Ad7Z5S8t7/
tUmycMyGFOmLrdhzxn6vA+OXm0A/l5NGgO5hPIWlAELULH067x2nnXLBIdt0cAo8
OljPm/INTguUxzqPK/jp4FOwL5ubTZOZxohd1qP9ZP8c5X0v7khL9iqYPd33xQMv
OOVJiNyq2Nq/cal1+HQGLy88p977+GwHRWptFGXON2s+Uw/4nN4bHmhxj/aNZvAY
X8gQXMEzLI01xluFKqRNacRD8IDSJobUmKixrUBYEQ2Lft88Z5RbEPXl0nhQiZRB
kr0QJgrxkX5v9eNkaiX/HGuYI2kvLJs7+HJe7CI+Ot6zcEaJmmDzzPBdTolOWjjs
yMVE61KqINW9/Fj+uuyNHd3IPticjDYLn0B5VCq06r9kXdiEXcKvZ9hh7Xe2OcPd
H3BUWm1L6TUaY3na1sUAbGrq8YQcxjKBS7Nye59lg5iCn00v/4s1R6DzniBjzFli
8rY+zLOiWEWkEDk+T6FLmM5w10RRijqSwtEPv2YlzwKSyCu09ul5+3T3xkjwf55M
pCRT5HiYqcCo+j+OgTP9sCg4H+G9hCRmTTi1c7WHTkrFZY3Xxdh4zBG3JMI57PyT
YCHkIh3sABTwtzI8L+6y+MNASMMQ39jFdy+4+YxmOuR+06HwPSAWoOzyyynMaKIx
o6mKNNG1DiiJJflzjHnbq4lpKTUv+Gwd36Vxp7aWMsYZ9lq2csKgh0mYpU51/qRr
vLwBgbaG+AIFoKfHyf0c4N9Z+4ezhIf8xpCIhgFKSGeOqYk46Q2AvThgyQX83x85
pzS5Rt39LzLXjbuXDdkQ9dtFgRFbyNKRQuEjEvDViE0sKozhQ7NC6kGk25DIY4se
pUcJ1jrsSjBbcUCQDuJ/nEByLm5zLQiKzrQaDUNR7GW1rYdqQWpFq6U5eJ94Lo8l
x6wqyh6C0mpKQGuKvYBMn33KQlY5LIkkIObs6a8UIjXw/INsVBnbCLgwWgalhjtG
EFN2MnvPY+uPsweR5DxXZJ4MBBfWoFEyFPlTiMYC8xAsG0p9oWCodbmjXNTaVeJy
uCoqBSAR/OSL/fVh7hnAo8NciUDyqmXoonZJPSQhMYgn2nI2LMMJujW+kVLCjuA8
OGzhEzBPe+7LiTNDxv93n0t2XNuHJ4l/FZ5KsOXWdaevlCPYJ/K6tfDwZlLFgZV0
342HzRYAylT5bjQyjbYCXrAwJ7XCn8PLpD8jYdMCmJvwEd74cXJN8v1pPbBn8wcg
EJEurtfuY18koCkuZhLQPbDR/hP1looj+zuJ8a5orUMrWAAGETWQA2e22iDCl+44
xR0Ep/tlTieeSiCth2Ef9BpEivfwt4lKLI9MEkZQG8oFUM9oOZLgia5sGMyMHga8
kvt6xVpiBkQzQQNt8zZFBCY746ifNskFOMkA/szhRSCMrao82rAIKIfuRYhh80dM
HreFNCu8BYXN2SNnK6N+B9LYuxtmqXKVdOb8VA23C/9DKYoX8GXV6NSZjirzwQ+G
NOefWu5LplssjQ7M8f/ArkYhcjmLVcFLstRfQjVeq4PRy3Whec4vAAqg8x1aDQT/
vSep4vPQ5e+wqqpHjhX8F2ExN8JgYUwyzX/QWS+w/u+fdi80zXd18zkC65R176NS
LoNVLGpe9SyYMg7kmijrndR6kDCpM8DIVsUATQvjhcfMymwgOR9bAc1VhMZqgfPw
1pvD8URFKUMFg/McgJZ+bpmOWFGH9vGk1uCZWnMC0h6DIOm8GVdw/bK1IcYAYqdd
A6AZYZMiiZA/0Lg7im+WVqAGYBq/hYeLpCQz1TSNUMADD4QevnogVDgAVmRT3UUR
1GvWmvQCC3X4kZfGNnDzCIw6e3wlcqIgpkw/Ro01kTs2I+Xa2bqHyovqVBdkLxOI
jQohayTmsqyzvtxYRaYRWcdmeAn1/jcQ3D9+jHFKlSYs54Y8jyVfxzmzcCIYQ70p
VnmgT6fzFicQPS9xPeLEwPDxrEqpZBOqjWJ0FLbWfbnyYU+X3O0qa1I1L58X9FEV
qZb9A2FOFCMN3pOyNtMeJHpxMMazlJZRPPRURzfA63hqmw3iPxDkn30UJU72F3cx
EFOcFnn4q2CYXS/2JaQa3qqIYIriJSH3E231PGU9166tYD+4QPB/dVx25HaAbfTL
6Vc8FaQaLfqBA8e75k4X4dRRBJCtl8nuNQc9cfLEwuWUysDBDBo/n5yYGoSfFvSR
JSjbhxDpqxzo0xoaQwA8zDx4kC/2iA7G0knefGTyc5NdZwqPGXQcITc6qNOjTamh
/sFrnge8u7wvT2lby0eWxa171UQDu+m2MkF2H+aLouKBX+y8mZ1VMdE/uFBjDZ6d
/8Nsn1iJVfW3POlRI5huRfiAXoM0/tHgoEGGSdwhC3w45TBmQyBfouDo6FjcwRd3
V8UlR573s0zoX+ua/W5vHwACi2xHdTM3fu9LB8YPagwg/nqNMmhlIII8IvqN/Ucn
jB9lBLjVpJgRUTdJcqmwpe0xjSgTbcTHFkpTTM+ZdbU70Ja1IQeXVZENuV043gaw
/9Qrujr254biRWSG3RbOsirw6jPg2pXUTgVjgN1jd2OtBHAqi5+WjtLtmQFO+Srb
aWRnE1ZHdRiGjFTfweOF6qv9IO14Vv9YauH4HtAWv/XeiURf4rqn5jpznipSAa7G
fu91fGWBm0iZpOKcBXPndmGsh4PtcSMNJ7X+tenX+7GEzIg3rL6xpSK98BHbOC/2
nKbnQpycX2XOBtuf3bnN/QguXw3ykiVvCsoIClIQUR2WX+a9TKE6p9n5lkozApQT
+fnpb+YBAhS1yKBon/E8+2VS2JQg1k5DBI+19BJFH6i9yyfmxUm4tpQPriBy5E9P
nVUOKV30t5M1+TqNdnt0zzoHrEAbLX7Mybz6IfXKVVoKRRz1NucUn39Y1/HqP4dP
p26E5xSpCy1CUx7wJWnXfm7YD4WYv9RznCxt7nOuut4FIOPunzekUThRSehkaiOl
sZOnjbf1/En6NUc34zRulcKTcG3zAQjOeb+q7JAmhoCLdHtV9XluKe0zQqUUyXSI
AviBxSYiexcQwMVOdAAFXXccXGDPvJScwVoSfkWwbka2VaiZz6sRHTVkS412SV6E
HFEGCoiS6+GJna2r+V/2DxG7zRfOFX8A8U8pQ8VpAFeH0CHUBt5BQsroJDnTCnl6
o5p/0SCx8wto5gIGZNdqU9/31a+E/4kKAW5Vc/qlZrBeObcXns1pzuxF3ya10yor
ac+ZLDCpJH73gSnSSwEOM6ZqqUP1m4vNfPqg46JVZjE5pPFyPbxtIhrnYUIKJBky
q0b8dxfOa1U0lLQpBWgSnOmp0+5M6HO9bZ5FFEzkOZzje0kr7dr+7f+bedg41g91
ROTQ9ZRXBnYUN3Wuba1i6EyEAMBB10VEeB/PTInvy/3Bt2qbncoeOdriiwuRQzJg
5iCkVfiSn++x72H22OxZMW48e8OsMWOjbbpABVGljItP+7Btsd3DgZwXI8hAYr4v
7lp90voEcOukiioAWsccenJczQwKBax/wCu38iIr0EhluSOaR9WByuka0HNRXJFy
nbtiINVzo3nE7IT45kxOM7mlzF73YHmzr8TY++MXolyJy8V3toteML65W+kuK1qY
CUhIWDfiAEyCSRIJWiJD6sac4bEUfSI9AYjxZ7buUq/VOVv6EYIxf9yf+vL0kA7v
13ZlZ9L6RHi2pRm0rcx8gQSgbk9Glr7SQiYDElBMTLgV0guPLplLNl7Xv+B3X98t
T9bxc/IjqNg5uzltCq5mqWjqIuxlp2myyGPsN2a/U8DRgA9E4vc0AzfoRst2VrmJ
MogaVTVaRxPV7B2beSpCcFwFbT/raWany7P740R6HI4H35hCc/uUp3RVutXlNNVo
Rp0a3onj0NE/31tHUazkaeeXoaDVvGTcPMZUik86wCKaGU9reEZ+wqgBGMARIKZN
E2fam4XO34kAwUfuqJfgI1+n/NVSCj8L136XIvyoIM7jrzV/VTBBvCCft/2GDQHA
kCpFfuFKEBzzwVDyDAbq5/CEh5jQ5BSZRAPEin1/Fo88ylIOMSqHCSv/fW30+HSd
HRKKJvL91yoI+hNFu4HP8u3jBb7BfNZhbev7thZaNG4k8cQtMH68/Z13/2+iCqxd
bKkvr/mYC6ra0wPq77P/fxQpBjcLwkd487V7zTGKtjKq6jW6FYISvB4FiNACavxY
5VWuTcMYhukGJacsyNFb1iEvkbuCgYPHNZmoPqG/LS28QSrbk+4QzLycV1QBvhXJ
qQMyZXs5jGVkOPqw5yb3vseIWiacEgHkyyENbnr/XBjGsB9rZDFTVbz+krmxpSkc
Nh4LVXijUk9PcSJ81SbuSwEOVbOJYHu5ECvQK64ngxif3Eh3LVPRhudPeKK4fz3i
fXEyGKHewOIuTQjyD4+69LqqRluLA2ypgrCQ5De+Hg2q3PW3zN1SQRhp30KXDrZK
qpp3SPeeP6xPWG+Q58SZCUCMcQrrt+Sv1jqZXdfD/qDwXl5sTflmqm5EaVyRXsNw
WlThDQk5na/yRay3piwmLvQY9+qFCXRLU2aVsOtGs3ogKFv04yIIdzN0bAf7AeNj
1iIAkqzLOTiK34WFtxUN62EGtC+TK4BZf9ZZCnzPSP12yT8t4GTqt4LOi0kguFXI
xxA2oI1L18d4K2dlC15jEpMrEc6sfCN4eJZ75O4/SDf0+opFITa6hc7/oBGgebkw
f/Xje/AVYH823qrx3FsSdPJ/netDQjrGKsSv9cIlq/vsGEwdZ5kKzJK64rute8aZ
RLqKE8TfSlCo+w4P4sVyPcPQ5RjKNmYtD3aI+ws2R5LZgb8NEHpao5p9bGD7FjvM
mW7Lsp/Yai16Mrd5xkd6qkys9AiuB3mcKosotF8wmSoMaOzvEyqK7tVnd1sXFjB3
VeUBKb1fD3bzJvwYat0gV/jfFxKRPDT4JL275OTXT7oyF36dS2u5zPvB4Jw1RCpt
EprpWVKyEcYUaL4hMg0BkNsRvsEYMYFyzsQIO9QH585pAgtlZpUxl3wc+S6DOMsI
UB2ICxMeMs6DxScaNwGatk54Tcl7m9gTJfET8FLvQmHX5Cm8YTRwcecZJTGgPAyj
yZCKeBBoDd8QaIpy1nWc20QU4tfIiwH/r/UiJTWkNfpQzVAHOz6OpVJYiKLjJNr1
t0C4+SiO1inQndsso5KEmFT7xe5vbWHTJf51M/laFQsgbwNqt3M0wJDxU/Zu7g+a
wG3l7CAXOAkx4gcGap2k3agpdgK8RuJJGJcr+AkLs9xujLKdxJiHMJegG9U+uNiK
DyuFFLVenw8P/StTOrhAzrKNsklOnHrjuqAXH6CQL3WSFvIq3CeLL3uOE6yhwmhU
WGbGNleeZd2NI2gltlu9gD66ULstIMsVczLq4CqKXdZ0s5Jh450SvVhlGkl5zTw3
QcEeUwH3xjbl9CWVoHZWnL8lwlUhyVMRmbsi31+wm3u0tgN67ABFy+l2uBwO1N2v
VsxzxGM6B0HUTPK2SWClcrBcEHWEm3TAmRE3v7azEqIL658i/P1/7vvFFDhe9aIa
fZ8SzDyc8MrhV5eJH8LKA13OzSnOmhOHAuLpxig1CCSTpZjiBvRrnIMDgtQG/epF
bJUwP9SwMq+DYJ6sIIoaes91QykPRFBfnFztjHJJGMj3fsBA7GnIbohzgCF4+Q+y
gWjnhIdvZNlWQ1kOkFzJ3/BPK8KNVNQ9cXvyoHCIXcmd5Bq0HMnldmB1ERCpkqUi
xhKJO5Pc7uFqgAL7hWsPHUzqsM5G7tt3Ltjz+O4UjqoPgUeCKsuLZTKSxEYrOhtP
PHOR+F0T4uFlc5RUvSTqkqiqmsrFixRAA6FrsR3DiUIlp1SCud0s3apKKFDTOzWY
jH714YcWAnYBY2uYw6Ccr6bRd9VI07GzdKzipnArd3xoLWHPayykdU9Zq233iH72
mHnKdNHNGKU5nPkvge1+TVFN4NyJUV7SX7sn+ypQD4K/QThsg9Hyja3hq/JKQe4m
g2Tf6sXyyq8UCBwsh7mt/GSZcOXANLGOkvzGvyA7ugAQunJ8/K0EKl4h8rvajzC2
yvHNAE7RfvSnAw0DQ3uZXJowazNLaW7PqDUv0YB7YouK17bsuYtUqJ9vQK4NX9z6
grcDA62c3UE8u3TR0Z/GahINvLtcLltr8J+HKZCzFtAD5dh2caeTJvOB76Y4rG29
T2TCWyxYyBZNJKnzJ8DcrB1hUaO/L5NFwNC6zewdpU75mJkh5ItBHZ9QpF0mWsK2
OMlc/z8yIJZ4kaHqgE5XVk884iRa5qLldNHUsxY8zSLIDIJGW/tFa6KaBBcui7Bc
hDUeN0Qfv4aBQ7/+dzKfdgBqpISH44JgSfhvWCAtmSmPGsnCXp1/08q34lZeUjTc
d3wfKLmmAUkMNrNdudVPJgAimq95dn0q6aNh22ycb+JlMDAyEStBe+OFG9bwMB8Z
dn4dW6Mr2LCq9kPjUBgQdffxFW9djiTH6lBhGeum34DC/mzTuWCz5fHjZKdKDBr8
CUc3H0d1GFW4XkYXbnWmayG6YoqntJL3s079mxOIN3ICQIw62/VXlS49f+1p+j4B
6v6IzYJkQgvKyOeIDIbbIT478xUIn8oA5LjvgFhA5hxj0dbs0xd/RVZR8FJep5rB
V9Kz9FOQIRktwSu/SlD/63beEYHTJeXtgNXnfr9/ivsR5pw8bibXffXB7QFoMx2y
G6/BpPDRfyLKF5cO4Ir6I9qicChsEonxxdTYkgWO4xHeiwjphgmlIOhIrFRczdHz
8QuCX5yYz4fOOSOyOMZsmrbO9gU4IfG1CG2UpturImKp9ehTYl3h2g45UOvnsl8L
pvlVOMq7yvDuPd5FYa7A0oBtrTPQLZ6S/qlmaL6O8c94jxS6SkQd6/kUJvfY35K4
UwWDNidQyH9jed8g7UhTQclJob13+r06c0GhgBGhEWUVqPZSz+YLi41z2ulom4BI
gAUIbNCXagbCX/QRdU2tPo9UrRrGP11j8hOKa39KSKymSZnPRuJi/5f8pGaRoDQH
9VWd+lgNcvnB4Q5pFhcBPY0TuoO6tbrZUoL+sHO/6lGlvtL3jQQC4VLv1Cl7RrqL
9d6epnWDNXnIO90mC0mInYNfwbcJQHCHyj6Jq52WyxmAHMuWZUc3TqTEIfknvvhz
KaRLFsc0Yo5/Ngum+bJFLeaighwuRkdMkkx81H0cGCcBDY7nNQ7MjS6cXV4z81Cv
XxuLX1jMTmMXFreB46DQJrWWG8v1mM7Nt+qmzPgH9+GCaj1IpmbU7WHY+/8EzyoW
LzXGEe2C+e9XQBc8slwqPpM3lVqTOWhQWJw/v6SlSXSRRYKx2gssGzDSRUyJ4hZN
QOBDPWZmTw/gOP48ybLYtwaVTdyWSZvlnRVIneJ6yzeoWGGWM9Ppozawj2v3PKzw
vRyD0osqvuOJ0FWRF7qVgWPmrpCJ9osf1u9RGOe8CqUyUBK8lsIP7IuiOR3k+SjT
yL3czQUJYg+JQ18jSTYPPE+Oc+siuIt5OLdVzWyWJH1ZbeQsUibT4tPR4+x4CdoQ
IGaed3T3T0Orsqd6ahglypKKGJwIi93SiA70bGxO0gK6GGZ2YxYfNVSCSO3VZ39+
l34Rndt99rt4vSMpzcxBhRdiWyIlsuCdw2jXuXWA0cShNNOYoxTShm2s7jnlx4Il
1WptCl2mbXjIHZkgqslgDqMpVidD8gUOBbK2oA+coZ8OlK74L88utbL03gnwJiOx
fXGhaAXTIg+NSD5W6rQQsu3S0ftSk/t4y11ajQ7KB+f7HoO2ZJeHPCFJ7PPzGfsE
Sxsfd2EFbnimSzteF/HzW0OJZIB4dOQM/Xjvi19um406vRa5hYJMWLvI7h44dJJD
DTlMonlwtvoTD3WXPFJKg7n6+Zfv5x2L8oZkFolferOx9nleALgi9B758UNfA0hb
XoHfR81xnRHUibAXgOEmZd3k9ZMujjhHugGoy3T5FOgyiVDedwpTMqBoJLaE/1GZ
YMNy+sfLy+JCR7QXyHjxqaJDtTZryV3ErudFzZe8ttEOqNwIK/ibFIlqcB6ZQwp+
Y/+lSn15BeyIPGB4z0gBgd3BvRVJ6WMjA88fLC2YizgHbUWxsoM8WKQy+AfB59vZ
C60dW0l5vq/kwdNdfzW5zUcAO3uQfyd7Hsl4Drr68C2VKno6juqSVUSDzcma/3Xs
XMcHmmamufIoXjijF2LUvNuHZkZomW0NXwdsoj/WlTtn5KIsAfCN1LuLPxVZdCwv
t1Lfh04IRzaIfye4RXf9bI+E7ljFheBNk27xuPcE6L4ri6PNZiPiTT3oi16JyoAT
Iz1iJPBTZY+0dayYgV2x093xHAZnSc1jiUKhn3jzjoQv7pxeeb8rTOPtkoiSCzMG
wC4QGd1ZbRRXpgcHFp+MNgy9Uo5aXT7hKJDOPFJeiK64vi5Nu/glngozf0xzNl11
NIvFcloImlIThZt2lURlMwpKHOgQ9IAzN4KztEftvPDGX8fPfawKKgvS23ChRMu3
MtAtcOMjqg1Z2Y9gt+7LRT0l+cFKm8QX+t9Wk4wYihNEEGejyfp2Fm9woyEP7Hzz
XOMfikjLIU86q0+QpBXAxocvW+PKUlT3AM0nnl1cUqt04YTATNYvcqs0GWDaJfP5
Ef6+odexnPJlIe47lL84+bnvHx22nk9JXNlOfdYDcSYl6NV7zhkYckFlJlTwZmZ7
JExDP1FYNAuSOZBIC4/s9Kwyx2ms/589TcyqEsZ5MeloCjqn0SMw+xxBYkou0q8E
Am8hb24VSd8F54CaA38AO23MozyhBNzAMyQUxwuoVPu4wtbb3JhUh8WvMepE4Epz
XyE5eH38aT+V3qmgbdrsPZz0qDeqWwIJAqaEEFtOxapoW6/9fj6W9es8guLoUIIU
ZoCEO0DCPFgWkHyv0gVCEExeHMd550kmeOVwtyx9lt16VYmwOMPnPT8rc3rgTij2
H9gJ7t0WyiFGJnL8O8AJPtVaRpy4RNggiAsxI3uaDWqIyWMwfdFqB1Dx9+9sUocd
VS9Q0FLB8YOsWnAsiPb1w3kH5KIwJVFEnm1rp0lMY0Ci/8kY3vKyj7TpTutkxXJC
AuWywZFaexQQl/Acm39WhAINFDfnTZ8nDF1Pok0Bzg+fLdI/MPrjnAvSvcgKme9X
NXSrY1kpU3NwrkSCz2M4tFAdd494JZyKeG2pmZ90qS2uFLCYf/qZpb6PSVQYTy+B
HYGlp4ITEHSiszqWUDKaO7L4YDNr0Crmq/7cXI0VaBV2qNCSoZLFegolIa3549qL
dpDyxT9ECILxb93Ou9JdLpCaIVQ+KVdOda30B6U7sovnzww+HhaodxAFLb04mgGs
/iWXsuqy2sbAmUwI0SVe8WAqY+TuHLvn0R/KHBANXBeVgkvGSxK1MaWkMD/JUjGl
IbceWTkiTdIVVdPFlZkPuTNfr7C2atO5k4qTd6oseP1YLj5ZJuI7Awtbib8EdXDB
6yeyH27g1ZQlbTuMZt3xThgb2jPnJZAMFQCexlF0g5x7HH5i+Sh2Uy4f3wjz1pTD
P7uXyBAfuwJNkr1cfjD3bpdvPolesBDLA0KkticUjlbMHhCpVNrqtD/pGOoIEULM
SQ4CCJe30b++nEfO0rMsVlgfityTUJhgTuNxShLZarm0pmFBreRs7dDEqNCMqMqg
RVRfWwei0G5wdGqOBDuLG8Mr+lIPuRkxkp0n7BjYyvSPjju3hft55cS0Dj0zN1JO
ns4aE3M9x6LD0IKfl7QoorlhQnQFVFEx5e7a7iSpYSF+9ntsnlESN+uxC3QttoZR
WgO5KNjF5Ddd50LqwlFjUQt0zKX2sOEjs9Z1iqyE685XvjMGyjM6Gm0wy3GqphO7
ndKI1aeghqbbZsouIwkYy4NgSmO5RGbOngldM/qODQsMf2+WdRcb2OXEVKARdjL3
BhAKWofREwWrJRpU7MWVfFJ6/EjXl84n6WLqdjKYdQTDddORgVcnBueD6ulReUTU
O1vfIyFqB6+ru5BzyVpyQ/mkhLQFLCD7u+KrImhKphRmNQbl7Kj4bvIBmVdNpS/f
8DAvvG9nlkQ2P4LIYTcxkzyvSjUV4246MH/AKBpA43ypUIht3/E1UvyDUAgGFOzR
f3TO2Kt0gA7rN4VjEjGWe5dY2W80S+KROzOGWe24XcDveS1x3bZqcLa5Bbe+c3m+
eTKcVufPjjszUjjjo1WPbpwzfq2C9ZjzWhAdUx9+FrGzmjECsKoeXqUJ1k3K1+AP
KaKEeiL0U30Ssl9L9GbT3ruBo8DLiQWoVCyf2cAg3sInDVI2EylkttkJ2sByWr2n
aj0OcMSA0DjVeQ6qqDswGHMPPlb1FwgePwa3ysVjjv70pZge0eOzQDTVgC2+InZR
UUSa2s8DK4OK+djekl/QQVkK5xD7A020DUgf8pk7k8ICZReuIMQq+p5XuaulKxap
7Y8uWXyOghwhm4k+weEJWd1cjV5WmCSkCcQLLK0spzt9rFDqOJVA8CLGJ4AJ/fet
2Cxe13uJb22lZItGh/ZBQa2mHrJ+YJwpvrX2NJOncN+tzlGWEMaMmIJ5TfhW340r
jafJ9HMMAV7d0ccAElq1sxwnocgNAiGz7o2mXyoICO2dZXRoUqMCYGp3Sj8POYdK
xGeP3Vpnry7agPL1iL/UzkCwXu/x0bF2mL/0Am6D5w/Yv5uNlwwSAwDC/Jr4TJyk
GwfZrxHF5Nj3UaOmq4mUYoqE8U2yr6XG+RC7QtQo/V1oYOiF6QOR5soKAtbhcMdI
4d9LPaKgle7EBe84supiwfbygMUVpPBZMTVZgRdthPIdxTwAsgs27VWfL0IEwDFB
hwlZq4S3GNYttWYHmt5xT/FgZGGbIcFVQdfSEK3g3j1HfglrozQUdxZiMQVEU9Hl
/NU3Y8QPA8Q6E+V6PEsQtcVS76NVfwPtY/bdRz20MYZjJnQlyzK0WBXNjK2sLEcZ
UoUlkA2tOm7GvREn2TIYBXBKj0vUI2cotrVHJzzpnH54ZnA1K8NkXGUSXwiWed81
4Ez04WNECvFMBMZbWh0yxtPAQ0oO+O//khdyqDPiKUDpFB5msqm3KvvXZIWlGQA1
7bCU5FDE/jbIXGaXM/huoyRpycZACtefkE6iAVdi/Lwq9ANg9Y50Lg6jCEaDVEKV
B0T8Ko4sB9uiAoI6dagK4OmKSoi6KZ7hlkQfBAIshMfOWj1M1FooDrYGpAVBhJ7w
/AwJRYbt8KHGCkwJu2PG4lyJme3V8aUtii2JyzvSONXFR0u/kUBKISiJC8RaLLjx
JaJrqJxhKMJR5OJ0B0mtgF82pFlb633Su+6Y5fl0We4tkdGtCtRJbOUyiUwt5wf3
OWhV4lGMV0VuIz703BUWQdcsj5csmpIL2Tw7l1pUXJyflcrD3xsDLNckv8n5y6So
gm1VkQ76S8KsuftY11ETNoD3tvcDEVCTr3JVVO59S/USRENblliTa7twxPK1tQxB
m2ifRZkeJDyxNt8TqTKtF5PrFDHr6vjX1j76ioezKFfoO/AeWWouqrIOnTJG3GAr
TlPfnx2bCmQxKTWRkFZWDtpMGmBOb2vYvfB0z7YHR00DZ/G4VUpbTHfbBjBIACeJ
aYcVP9KeBs+F5n/vBIdOBD7xeGkZClY5hpKz5PLNC2wj5g5ONWWILajXfqTHIE30
lO1UGZEk4pR1JG0b6buZ2GidDZxFNQfDPXa74wavajsXXLC+WvhDqlhKmIH3hlds
2WjyBYxIMlHrv2A54ocnzApzZ+E+pUZ0IK/H3VT9RTsJ+kuuFC3zAzgE/FsttjnN
2BB17vvHZtCbvX1QAvc9Zko1iM5bGhU4+Yg8pmkjpfVzEtRzBiU20/atXQl2QGiw
hBykS4pN/d4T8l1eACmLtPJiFldemCVLCh00XdE2bGcNbcL3IEH8Gq8N0tqp0QmD
a5z3Dk9u+dDKfdM4G2+hz6qDgjW/H1+iuatiRMwOtZ936dCatiI0QTF1KgqlKtTX
A/9qq7BbZXCAftz0UMxFSMGeWBExaZmVTQe2wvYEgJZiEs515s5C1ZnBo5cS24Df
18E0Cnu0fmKG6yadPlakEPuCDHi8E61pYYvPUspZN5+Mx2LUVQBBwl0pswdrxFtr
Esg+wHg1gfWPlqdKtGelCBIa5IeC+BcOutv9lMU2KjY4/SCDxTzUtOMSf7in3lj3
E/CPWnhXC+qSu/O2uHt0Gf1j1phZ0KbJBTzZIzTtOhHB6gnKdhk5hJszNND+SOEO
jVyt3jnUeK/N3V242BDsl5ciRL02Axui7pkt1BKILSe/rEPZ03+K9sZRxzXnzLHb
hJLB+4M9htujfUxppDDMCWN3GjqOVnWd16kqOvLNaxb7AohYfdX7vjYwDc+WQn62
C5bQ4MCmvCdioVYUcy0GW6lQ9SBi2pDqzNC12oeFs6f0ayTu0phBByG/xJTgxA81
mRJFHXc4qAz8XQYzDj8ubysjni7zaL4AUOpFpkFZhgdgminJq1kwrMMQZx8ZVfYY
DcKNMBDi+mNF4C8XTVDxg6pjKKniiqFF12hAI+TiXGCZ+zijSj2aUrGx2dwg1RtL
RU1k0tyAy9kX7AKNPjHikZoQE0Hx9hruQr/Gng4osCjn1/erGqtrUwoBbZxs9X5k
dyU01ZRmMIJr37SsKtqLoWs91Ae3Y6BXVEidHVV4rbGKEUEW0w16ij0Uy1yxmlcK
VnUqxLiVWt8xGcxLMOxSGzeBqoILGmUgBeXZsVOq+DgEMEqz0fo8IQhO+nszXctf
D02VZfUyV98ort+qQcLU9s8HxkP53NDHAnMa4Igy1cbaSOA+Qq4Mwb6cdZly5ULL
iq8gYf2BSnC92/Ps74TGs8DCpazCbfMVsuUYVfsg5QzewjS6oBP8AY9oOgXK+3da
FkTQayf++3GUxJrnKAniO1ExrNYVUjGbOtd3k+x6TC74Oiz5V7QoYdW1Fgn9J/Nf
lDVreAnxfH1JopJhfjUUYb/Di65nXyzJ4eO/x3yAHVVb9Xx9YsOj2hy9z3SOoyfu
pyNBn0CYi8UAYXqnKHlls8HAosPQEkHzlkmu3EiXGopvNTwll09go+Y4+tenraO1
dHisIdVTyogQPGyO7iIhoZiOUCkmnMmEF4q2+kZkad4kv4QweQMFz5nkk4Tgj85B
xgtZKDGLPsxMkA8eH1ddscnK4zVm9HSqEq8RLPwderU6dTzwlbi30DAbmCfXvkMl
aciNIpB+i5iAWFPOrPoXk1SkClBGyOzamVrxKhEwNvsgFG2RXqoP5wNX79495g20
HIUsK5aattd8EUg+wQwe+01o361vdKW2a6Q3PjpqyMCFhAnONDKhX2FBh6oUFKqX
2Q+B6g9C8puMIuNQPXQ7zODbFrcKASexL/n8yBYPRC9s2I8hcVbM3SysjR+gLiSJ
nKVUNj1jGfsODpNoIu0Ujbsr6KOszikcMXjVSXpuc1V4rSimFq+2a8S7j+UWfjPR
X8XUg2FSwo5qSnWOhuqoCjEd8efP3X0MP+WCQcUiHbrgn3DbPN05un8xU7SZoyYI
XmIdklMs6VtT+Oc236bVaBma/ClQDkFVohYwGphkz6XWS8vE0eUMxeN671N6hEMT
BSwSOvfL4Vlfanx5r52TJpuKjqdoY8lCWHeFD4e/1xZta+5QuiMhEsH7n3eq/v6S
+dn2054WPZy/+wCyRydkNTPkFSXi/kAlcv6+rw/Lrg9UYPmm7jzqRGxtPHp8+Q4m
VVoy5SXyqyXhIdR69Qy4Ily+9mHk+DmMGhMNghLcCOgfl1L0Rmc5ZUmQJIe462Lg
GIXSidmUV0K01fnKQKYaQ+HdwB1+xnbYhdm0iCw/kq5aG0DV0INqU4s0MtTL3D+9
FvZZGQJfMgIVNgnBsZzXuv5sXHz+Wn95F6MZrlpUtBIWNilMoiHK+PaZhux0l6uC
eHGU47WOtSQBM5v3NZN2Dc+dcL/huCCujr0Jmj28VUSFkBSEIbEXZWCwidU6ZDPg
74aiif3K0o8EgWCN3HqrMNZ/bhm/BgVB8x8RhUN0rHrt354kuF65s1hCcaYl7l2A
fdwjMsQi7JwSCLripbL18WMpNCRpBJFPItsxg3mIcEpLrFmHpUvJ8t+dET24tssg
BaJz0V/iLOJQeO0xT/7tQqlPpIgG06SFuK78HmuamqmAjPrHVL8J3wLO0xHpuqT0
BxilhNaTw9lDAvH+yvhmK1gjnq5aBzEpWAOuCNpS6EQNjspTGHPxQ7hwTrg3YCGo
JDnmjZE84POAfmILD6V4PPJ+mvTvE1s6qEaNdF22ZHwtcgfx60KgckE8S/w14pqK
HPZ24imNs9ChJUSk55iE4ofhl1UcGaxzZwzQ9qhxWrdaHQrD8dhB6aRNDArCy2Fb
MILGFfze82Fe2Xpo9HtGZ2/4ABUegMcj/5AGmAzk1m7zLrtRAr8f7KJ2GBc6MQSn
CuQzwPQzdnkoUhx/X5iohWqnslT7wF9cEsi/CUuinR6ByfF9XpuG5WGixZwXAQvb
w1rzGhC6p4Ox/mi6ukaEsJnvykhwB9omg5Hsmm2/oZIjb2eoh2AFNu1Cx9QA/OW1
CosFVjj18zd1NVCer0+OiHU29VFXCSNE4IcOSHHGSNBxdpgR48fJ2dgN06628KXQ
ZjeoeoTWBz5AsWeBXqwSe+l50VEsVUu9UZfAkScDzn8eila63uZig4w5zorMqieE
3aXUaqsA2fknyWH6uRFa8RpDs+mlGy4doxGm7SreZFy8CWqjV6hnhIo6Stk3mIql
2ZjofGa3U323x9DiL62eJwVPbe/7AzdMVjzL8C0BThV2IH4aHOsu9XdMkGotf+ar
hR68raRWcgiFhyyXD5jYCqZZtFpIk8GPo4ujXvrL1oU1ee5mFU5PI5A3FRJe+MGQ
lVmilx2x0rq1av5OfegYh7VcFGWqCuVcpz+KBilntBVvLx+o1upoF6zKdEu8lUri
WTyuhwB6QULMTx5nUCq9tcvtxOdAJY7STbXrKIRppD47z8hqMTI+CHXHo1+slFZX
7XBsKgL0yu5r8AhR/ZgzSbhvSwVZkAOTMnN/qKq7OIGHR0gE3BjNGcBG9KSt8fRj
OSXNedd8lsgRKhxlJ/voDd3IgkyWTaAVgdXJI8btvgB/UDKohOu5JtYsQMR2M+ob
PELz94iqQJpxNPcLwnQ+jM/Wk+Qwy9RwmtJ1vFMJfTfyC7wD5YB1KOacpEmYNOo4
FsEHyOTU1Ir7NbJVfaKBaeiL7dyZVmSuzu+VPm/yS9tYLRRABonLpAYqnyAa+4DL
UfuBlZUayKfCAgU+syk0XNowCsr4sZ7nudRYGc5T3U0PJ0gR9EEq1JeMZTsSItCt
7s+fQ3tVS/nT1QL50lFcEmKlEym2QntuINue7GHKx50+w9KKHJcLXCcKr8wf/kPg
CDhRTcONkhvU1GNclJ7QAGj1MZR+olXSK2d8D6tvKbdXcZn1NPUQag4grOnhfqsF
QsvdMoJyjY6qZlfUftanWyI+6Aofrt2ggXAU1TLvpIymlHBGL8/bEOsstgYUxREv
Ghet74mB3FJfM3Dh9xDImTZsKgFEtNX8Mzg3r3yXNNWRraBjPE61pmPeYaBiO8RM
G5t03aQGKBBsnr+otpVbCMRTsh2TD9x3EXJIfD9w90qtlKrS0/xZgO2rqdx5HeK3
3sLlwPh9seGOjCR3msLNH4kwm/QdNE1cDcwnt8LZXXsKOPJ6NWO3+S82C9ifZKG8
vbw0oW1F1LFcCZKp05YPR0xKMuQfrvGMVGRb9KySr1+6IhmZtNwZktrloadA6bVa
t0hjXK672ZigN6aWJWOmYECIX+HijPGUf1MCglwMibSA8Q1hiNfOSw10QNxhyuWS
P543eA3ZZJEoiCSAXQIXUud47YDTPvm2yB5jNmFRFrW303rUjlkuDYa4egIJY4/B
m+X/guH9QoUHRlr5+HWiftFRymHgaTLuPdyBZioN9GqYvxqL6dsZeqe1AHD7OYwU
n22sOBUXEEO3ijGQOEujg0/HD4ThJlkotzgBkV3HGlsVwVhpA802pw3Vzr+DO5vT
B2oOnsJ2esOcUC98rFyGXu2ongKtIyBD/1Jzy79g7H3nbZ0GSi7IF7tk1zDimcJj
1tXgjry8vHcaYnLpDUCg/Ehk5JyK1ACViUmEAxGj3TEoC/uWr81M7HCB9uBi/IZJ
KhlEhuxr0nB8h+Azt2H8D5JbYz/LMWW8gm8KWhzEEy+hw3ucOErF7tc+oXfuKyDx
+WFjLfddcKTVWeJZL+geGsxRv1rIhBHPXHjNxcFeTx8a67vxMVEWx9DrRC0fdyr3
dqShYbiY9dGamDTklkP5W55bDh8fI1sppmbjCr74h/OoDrGeaFJpN4/PtweLihp2
ClUPne6dDFWmc0K4SaP+liQZy3OI1QPt+1NOdV1rEM1bUfiEalclMJy1iVllUtCk
31eFHD1DWnvkrbzQ03EqnLJ4AINE3EacSNPYI7yWX9AdKIDKiZWSUGzMn6cyYHRM
BCL0GKAp5p+2KQ6+VMUDqxdDSopW+i2UF7luW3R/nOqQrGDtrRAcFCDivizRuPrT
xhhvblIX45UteZC7Kbxm7IvAv1IK5Dw4s09hY+DY/A+qDQ11vjcjeV4cNTVk7zI4
FLag7mlHJugix71rfQgAspT/OTTcegU7pVhfshYv3n5ukQWcAzuCAy36Iv3pDqgG
+WGd9hw9TvK0pvHFQR7tlvFdn1jXmF0V5jZac3eZOctDH7ezCtiHvI5JZeAd84Aj
oOPn72ad346NO+vX/KP84vfVNiLH9PyTNJ0jyXX/2qm0Jruim3QWLHtkosJMALAx
nDbrjwomxVD2hWgvC63PvEXFZ69190iVzZYvNqhhgRdKR5VYvijJwHQyA+axN7vB
SMxe9LGfDiOf49kEOuWFyvxOM7T9irm7CzKBzwQ/zf3Hu5R4/vaN9qYgoZ9+oOW6
4cmoWpYr44l78HshoLszwamT97AKRzIStfOZz+YqkNq6SZQ/c6n233Uc/WGlu5M7
XoOd7Z45S5bgppM9sf6d1/wRKLJG9vWwcJ5vwkvDFi5/JpPdypQnxmRl57Ms/aa7
AvLyN2pRr5hKogcMF/OOB8Zb1i3mZxxIzT6JJAbEVzMoW7qxHNvYVbs3/Neg/Mbu
AXu4EySbYnS5hagWaRUXGJDMDNAWflGXIcOAXMKC+mpN2e4g1RiAdMRRroMgfhz7
Mw3iTFMcU/Y7rEGzZK2RsKHsLpJC/23ZeKRW81+Opfc7stoVvH4nJjzZgOHJDL5e
QCeJpwxET8TVZRnlSfKFHTA5pRF9sds/yWLTQ2CNAMyH5Vk++4UmCaBRxMlNnx5t
H8kNSSHerijrXtNVsGAgdR5IHGojTpj+cmo4KCNARkR2meeOqUa/re5Qi2ctxK6s
4HP7wZQ4S+cIodKstelBEIUjTwHR7bMauHHF5zVDCkqRN6m0CqWHWkSYO7lQ8443
7dWie/5h6NmXfSub4wzfdkRQIRLLKj+tz6sxiS9mu0xUc6kIgfDr6ZupcOO4mX5D
8dYdyHHLYRnZA3irQnvErMl8dLFw7+CTYWCkcrXZIwa6BW4AA06ThKrRB1RKI9Ig
NuBW55kQzw8yx0A7ODrroxRF3ocRe3y2OoDdi/9LVozQb8zXQiUsGhy/7BTIoZME
gZRulnaSPbTLfCvoazDIdyUbKKW0h9esIGwxSyPRs9UcGyqHjf2gBrufPDYxOnxb
WxIGxfarBJeLukc1BEXgra9eOPsea1zuWzEOboUs8FnFpW/tEeVdmQVlnylHEHyC
nc3w9IP8Kd7sVBZqHaJR2lksAzH9AFlvYuBQYsng7HQ7OOq65DcxTx6bFSGuvWfX
M7o82A39K+to7sk73SRRlqElElRId+eYBlGz1KkiiEF7Ers3N1sTdIYhjie/CKBe
x9k6w/KKmJQ6hfpneqDadmKe6y0y0giMmjCntsR33rewJuD1rfWIuO9YyHgJOvcP
GEOBrTOVJA6XYtcGzBfonfpFWiV0sb4TCi1ttCGLcAX25Wsxw97B2N1FEQNauUvH
pNoBROu4uk7B/nEKNdlIByi4fMTjq3qS+XyBuW9KY4FNn8KSkzJC1xtA9sbX/55M
IQSP8pegFptp+Hxj+6AX6to5MA1iyrnD5h0CiG1RQsBjrivSrGcL7Pbk8jVFSFT4
grNd0Rs00/9maPpxz/Ez9xo+4dRWt70pcRCqr/cLd8pQA6MU5Aand3aUrtlieGVr
dHoJ+UhMVIR6NbbVNDNuhUI4jCByy9iKJpPnLG/PrAXqsz+rbKqVYf/CxfEy/6Pi
Iy8bPfdgwo2HQHS3zV6idMlTxnZeiB5JcW/mJHd1UhlbvJKkPjiOyOTxedcu23sx
eOOxxpMvoAmapPM73jDQAWkPh0vfelzVxil3bSbTnGRGtJtqK3FElGLcbyMWhbs3
cRijE5UyOJjVhI91edVmpskjstoBZb4/5re6MkRceJpcSAxiOZD3u8wdLvw3O/SG
VRGufKkWhwkxZj0PHCNhFXOlkwzuJyBXNmZzY1imE9s8rfCPVc0vlKsKQ7IJ5jKe
EQN9sV0UK+bDvPLNtJaO9TFeeeMPqnM7AXoHD0mV/pyHURn39X56FmK82qUnaglW
F+kcxH/6FU/p62isesSjdlqI/t889eb6uoR2bENTg7qfghGFuNS68g12UfhfsA9G
VULjkIrJY9+UNyniKljt5g6LgWWI9jCF+FZP+9TofGqxM2DAz4woVEVEZ/TYcwvD
NKM3WOpRRkoJGr1lhMpxJkAot6Pmb08cIvDuz5A5H3G8XCOixauYEQWd9O6gNkOM
yYSZb92zd0rwMPGGJs0LF3a5+Rwkpq5Gu/NqNAR4QDGCW7Ibv9O39WvCE+fh0NPb
P3eTrFHgLqIElwfK1eTtLJ9h5ezasVs7dqbIPdjKYAqPEYbR/N2nwRw8kpB9rTlr
XAzJAvpEBeT/UQZqcGNLFMtoYJNL1gW0FhO6eLMBnn+ODdG8/wRqIyBMP6RKFNxq
wH4AuOqzUMDJ/bPwQn4pza+okrijKoZPpTuLlzDXQn//sD2dSPIcn+o1PSddeJ5T
grLR7ouTd7x/wRKyycer9FoMYn5EN8ZdK/NLm3gxv+UMsp1nM39saELcy0Dq9RcZ
5+jmXCEw3zm4WcKBghmVawni/C0ig4c2gkt/gHpXIGq1VZySP/Bt0rYUCrCLDguZ
04JIf9sIOVMPKf1vn7iiUm/q38Vhg50J7xNyQ653cA84pMCb36JCt/LuVdL0YebE
uKIBw5/tuRxT6THCMOE/6QtF4w67nsfRvRnLZ5XRncS2EhQzPmQVOM8hCXzibV0V
7/koVN5hvRcuApMgFt4RXZ1ZAobCXW8zjFjhJgKs72H+vTPkuAHkw7osab3uGQ+C
LeC7W9sv68Chglj8G4dPiCOtRal6K4T/2QEB237wzJW13fW2GZwDLjxywoctxjJX
7m4SF7UUWiDRt5uxCEcioPd5T/HQPIeGLUk+qBROZWC4KkOsuUquErWES87lyO3w
hvxJSkkvHJUTj5KjvQioPxncFgpTrGoDQVzfNDi5JjBOHW8rz2cyX3fHWusx1CJ3
3Mc2jcRCm4qnJacjlmZqu/aOHTJL6Lj45cgNCaRgWi22P0C9+18PDvNBywVO3rWS
+C5fnl82+w8oqnlx0cKQaRuNlNBrdN0OUf9vkTapc+CywiG9ZCnigMJdR+qO3jWU
Ah7BTilfsz5tURRp6EEjjewQrZ8bUEDLXyKSCDZoculFD7DdClbLxayN/1faZQSO
0ZJoFAOb43uZVtcaTIWJOVYCV1icmcaJlrZSKlpNGcSkV//s/VHr+BVc/PoNBRWf
MBkLroTp8HQHVOVedkPx8SaO/H1j+653wO/cZaFSwMhMUV+cqm6qy0fGGkmf6Oig
yL0FFs1uieAlWJ6Cb3ZVkYYTboitOwMDHeGUs9owYVNw2jO2mKA4B9/XTz7c+2MS
WErWUjFs/z4lnqwIZtwvODVxFL5RzKzU2DA+OSC/4hf0O3JxwE/YBQeIxJT4Pe2d
2C4j67UjhJM1AT8TRNJdLQd118KX24fpGwA9cN3Smgk39/T5/Ta6+GO2OdBcZ6Oy
vQWJryKUMKBuia904Ln2yUVSiSMT0546arpCQLm5fsoIMd2PaT9ddYRzHvrc02pf
/FGjs0/J0O3rKvoUToRF6fB2voKP0coBLv0mFP4NDvN/LtzPLiPiRroaTw7fNxo+
2tP8FCLZoXO5xjq5WtioRRghMjDqbW0JkBXxP1C+UvkQCSKp+Zb0+liiljbS4vrD
3+Y6ZhWXYhMnDMk+uh/sPU4aB5CSm8agvn3Bl+2SCfZXB0LeLPn9+BuDmGZrteG/
mVsJ4t4Y+7rZfZWRRGXodWewYDSy6suD/jjR2FqSl5UxBsuLyqkAoBvd1UrpXuAh
Fby9XtC2NMIGqi57X9slDpmypD3dg5RJS7hG7ugVLHaQjDXA49zzrKl2ytGvrCNs
R/OMeR8GSvIKQMHUC5tcA5tpCSbV4SfEdnAyrfwV4KmKkvbT6Hd8tt6yLagzE7jS
nfGAx72jrvsWe+gqSkJWFuA00TIN5+L+NoLsXNR67Pe3mmAeT66aQEgDlfjaFXqD
Ss1+02dX9Zk0iqTG6Y3DXe1E/Hluw89lGFGPX2dsnJXBGfU3bclOqFg9LA9hcjNZ
+lxynJiYWlMm05CDinS4hoXDiyq0CT9Wox//s4XZ6ep0n/xjFAB244BMhj0lColX
taiRDINd3G1w3p3ICYMnTI/SEJxvQCCCAiCArAfvTHkWjPnF8XGfIUohVWoFXdJL
7djBgB0f+bzVePamGe1Hhfipo/rQolCOuS0Nb4Ju62dGMQjShMhBvfHnIeG8Dcbe
n5wdyKAcAC2To3G+AQJPtmh9AKAr+WY4pxpGQUKOMMRfotbzQZwsAAmghtlJExcl
T10SNDH1/YP8XQ/pq33i4bKbC2/awU3pX2gxTrgo+X0Ay3w3R6Pj0jSEmSg0ucbt
bn2YOV6/fyWJLODVc3bazj9BDo65+NwNfHp4SOSI6Uv6Ra2RPPEQCJSOEQHfWLpy
Ljoqz9T65W6PopED1zlQDxt8r6FeZqDFpVFB+YDV3/00/DPjvJqPpf1HNiD2lAEG
kZHNK1NThLwS105DQj8JlKtdlunOPrGss6m+0TNbZWcrO9zNPjmEhSCOS24FtHvc
CEIbwh6Bx7U3vPAdR6CnXC1/3zKBRlMcCIJhH2S/qcoFWF8SoorxLxh07oYIDDie
gs41XAOU36WOuEA5FiBW+OnYSv0CmBEDdSfDyxnUI83JJLkbm74FYQGlsIHHxuD8
7JqE6yTwvbsJEG5zfjdWAyLxxPfgoTKWauLzeXU8M477Ixqq/ZnEgJz/9LPT3ggH
TWWkMFWovqy/EDZpF7YQeZ0x72jjx7UOo2tU81UTnmsxORs+5kFz9/TdZCcICa4e
c8DYpWg3sBcUv8e5nUilY+lpnFV4ET2lYeiiemITNbpdC3rON0OCGh85CD4kBHcI
p4tHwn6G7h2gkWXHiBQQqAsWDI/Zxsi3IUHvxJiSgCP5XgNspF5FGI1DcZvou/7/
naqctwH7jWZJaSNG/ILg50qaerQsxVjyy/ul8LTM2UNgvgwJ8QLyX1osUYRSvVvV
lyxxd5yoCaxOFXWqZhQ9/iYjJX9tb2fI2y+8S9tClHq8u782AlGvZ2WMaU055jzC
PZC3zcc1OzQ8sCdUzRWsXhssj7FiSQeJ9DrHrW9ETlZ5zmjYzNoCiG84xanCUqT8
JuuWOBVSE4EV4bTWd4MkLtK4Zkg3b02rLr0HZNj759EPKDqgC8XWAMGxPStBw/qv
ybkWANPK8qU/fXFe2enSWVOTmkLxM73gKLdTNMKqZOGczxDtJEic/aPQUKqAuYRm
JA57XPhCijM6ge0RewFTaoQyK8g3wnNxuY36iURVRI2liKuZcOWJ7Uy5LUMhOWo6
3aTxl1RgyxxQSVA17/LwmsK6S6trMXMkvW2ZP+v84VxqSON9O/7RqKrUrX4qVNoE
1ZSFl64XMcEPfYxYGpJ+MGlCypRo4pDA+MxhRv7EMwsVcV75woCWPU6qmzcBE8er
TGHIfftB7f4RwIFZ8mDw1yOmYhzPrRtlH3BLnm/361tw7gQx3WBLjK1/1EBrIOD1
nUIcI83lHY7+uh+VOo8c3LAPYanoWB+zVpny/SraWJpS0uE0RFxfRcfboVxzBvQ7
QsahWhV+/zPlWK1qXGRLorAQ3Ou7Uzi90fxzZUxf89kB85sLO6IIs78pAAyXl+Z/
TNGRP67CgvpHeJf3cjPdHwn0qySCW8AjWsbNIzCIzaPDlL+sY9noMQGtsWgeHlyw
0hx2mE79Q99L6JG0ufKFyE3dias9W2PpgaJqdqDDzkdznXWMJhkmkTJSJINdgP3d
AawotZbVej6EADzlOxAtQmXFBy3e1jQ/AgzB/B5VGkFTfQxEM5y7V28ZECgUrpDa
nTF92UWWPg3/GNN70GpPkZtMLniNyo6OqxPSz0c36LSQWI1GcL25cnx4OBAX2NBY
sIAIBWNeFTGupjSTAPcXxb95u5kDjEZ2TZWnTvO6gJc/JwAfUWQDaZTu8ccr9f4l
FaetCTzA2ob6xuv3eAoUDxXz7dfzeZ9ugJt9W1HDcUQKVtADPbkAs0IweOVC71wk
WAPNjcRmMCTNGomCW4Aedc2CuR6k2RpWi8Wm8O7uIajw/alRH52AmC5Xj6RhYV+B
MJIFHAj/dpnuOdgvFPm9u8tYMatyIwk1dHTAC02Jfeb1tcqPJx3CGZTflbvUH36S
P1TmLlUzSUDUC4n6pipgHu6PM86tfw2XyT4lNkQLI3Q2262sxXRHcslpYzuCIHSu
Y3yaY/CfRnJzX18goh9jf6TgMgDBjtTXTIf4d61/d/CsFmoYQEDljyO94CeFR5C9
4ksge0q13L6eqPUSuIwQ6HvX9oSMeipG3k0MscKWMIO5+ejbhqwGMNTNmJvPIgV2
Y74oyhPxg3+LbPrnNH3/LAN+CTkM31c4DsinDYVjGOQwvuhNcz/qrJYuw9VCLwsQ
Et4Ocio3xb1K07v6Emnx43Vw3CjOVlZ9i31/pHjOvVV94FYpAibqtg4aNaqxPHt4
mU3x5jrZpNtEtunmvUcFDoqvIvnrxT/bPYZqx0Ycz1jDTNXbK2ivmkBXniDteuo/
77C6zBh0n/og5QfQ7E+2ZRShN4msASzYSkRJIvtkKQlRLbkcZrm1sXitHAzuzGW1
gmljOWLEYgcD2Tosv1edvKdzY7HoqyEC9Os2k/MGH4xtYXX/svS1a4LnHtEycIM8
1+CEeCiOtFMyZptT83TPpw+3frzLYA9zeLSgp5snsh2oDeXIow+7TOeY6cz1QJaE
d0fKHkUK4PkLeiQvhSW55m6wlfqGVYE3nqnE8gYdqCIYMwxJd+piFi5RhNpBrHyw
aZ8u/KvnZz1qybqRTQCPmjYGUszjjCyboQpuNWD7f3X/quJnf9Hm3hvTt1Xpls5W
AIWbS3lC8mJ9XyZzxfXs2XLxUxb5iniTjhBPwoXt53eJIvE7iYzy1GZE+Dtr3IMN
8dVuoNZgP0GzdO2cZppR2SROfMkSG+mArdV7t9zKffxGjVDjK4crbTlSZ1zIhceY
yEiLbd63klDUPOjjhiEJneDc9ze9WveKs4VOxHhfyhu0DA90SW6HK42bYO6gggUK
GOscxUUlFd/q+Lw0PGHd4d04zmmEIW5VmlAnLx7LzYjsgIOPbGYc6EofpWaAsioR
x57UggZSohfdC0wJGdX5UZ6VT/9q6vrLxYjAGzfeV4RgM6BWOhg3jyGyZmqlTjZt
a/uNlAs56b0Sq34b1qx33MY+aW2N04Fv+p7Dm3dxuxyl/yMapqSm6sBzpTdzcKJ5
G1pe/gGQR7Eyw0wzfIPv70yIz/jT7xxxCCh3Y1NFcgJETu+8Z21dIA7FCVaxUxn3
EhYosiYuFt6GnG/WfT6Kbg0/rGICZpvA27mVj8N6iCn/JJMFDZJNDlSQeTiRKDHd
UtyjzJayfAUuXRnk25NBHsMWRvBb/pPxoVIPg9zPoPWRg+DrZeZ2RT0oIiWJJ3uK
6cGQLjF7D0C1mpxEU9K5JYVz04ZmVtuk5fMybGyglXSkksRaoMkziZHLjE/wPGmo
2D4DkAvDG7xXVwsGhhDViu/eqUvJmvBKr1QmgN6RF6dANmj23vnE/YuR0KwNYSus
g8KweQm+W5G9nkKyV+C+cMIW4PR0k+tADBpoOt4xSREpyxc0kPGcFiVHd64i2853
0NJ4wBGfy2jiqll2haYFHX2CyXlMpo+ACK3lb5UlSmVV5iHTsE1ygwKEvFwCENnI
kzjmxFV0e2fd1olhUfQ9aO07ObymWop5xW8VJ6FSXH/WaPdNDdc2v+po7e2ZVHMS
fPoftedvI8ETS+o5bdthL8gtXI10Z+JJiSBIAynSOssy/Anl9P84LUSJVD+tXf/z
9OuV7wE3PCPsyc2nodj5il3FjhSvC6MHU3YWYM5bNxs+mCNCUrNtshTH3pQfe79X
wdT4qgxJmTyhTCdcf8E27W7uZdvvCYJIGKXKBKBOKVBBJG7Z0idp5vUqeiPKlZZ0
39cC+p38AE3wuJgz6ECWU+QK7tDMPrwhUF+H3kZnOo3OSJaXiYw9FcvU+Cjdo7w3
2vj9HFeqnBKHDWunNuOfZyasNavEcMV721saflXkqIlMu/x//Hphp7tiIPIyJ3pt
Kov/6SXcgJTdaoApwVPbYrRQoJbzgtwlJUe6WL3Ui5qDVduENok9y5dF+EQoyhLV
OBnJaIUnyPUslqkYqf0CDBKhVjhWqXILh5GPQotC/xiUtPwJMiiKQHHN2Pgs9rto
Rz8DGR+h3cHL0x9K72k7Hzsp/+tncszFozAb9opp77VYbFklzWIvEa9ilUlyz2U5
tuKitUoUPdw6T77v1YQFmc0t5I6f9P9eDXoIulASeDniMbLmWaF+qa1CrDZwUduU
JkZajzFK1A4nI1LJkX/WSfSNz/GH0Lpdn3nbxhXNcp/m2+wrkV7GUYoIX4imWx1q
zjQL8FNHSprAEpgqXzGsCF46HkhXw1XCxZiE7fs8j9JdjVT2IpcvbF/0hR9J4fNk
ZnufuT81iQg8VyK5ia323nOmlytWeXQxGzWUX2A0I6XR0jZBp5KbizCVFgTqB5vK
eSU/AfcRPa6c7oug9RhjJA31hGgbzejTZV7lVfoVwUQVfl47U8mzbphYht9b/hUu
XVk4rXELtKIvpjpE0apfdVBlHNSBUEYrg9mJ6UlT9GNXZpJ68OxBdYvjv/1RyI6u
pMfd+zY3XfS4LAqQm3osakrOLIFeNggkUrqgsTpFPaqDf2VZn0H1BDUvGPzeToXC
TephDb3dSe2b50xeAZYpsZYUnKGitpTnfzqhPCMZgaTYHiHpEYqpeTKg/Wb0KgRc
+EJIA8O8dFFX8Tlo1WkFtUlSXmVbwGQwJSvQzFAySl9ZnU7SSJX5sk9Xdwyyhtx9
yOYEsDyJJT33HEwQQvGHBnn00PpnJp6OkJwb/FI8zkiPJqLq6ncQLZxP103A45Ez
X7mI8+nhCSeTeFDUpC41YhSxYBB3u4oNKTDFUWntNnIxA58x/ywUl1kXfAZKkARh
4v5DzZlqMCUjVDfZRWUXHhw2W/TDIlfH5ZbfPiKF+V3qvgjcYTADp37W0uzhOWY5
hk1TwH8XbdXOoOGpsah51G/A8acuXr6Oih2ME7UmV0DMpdzgMvSNTXB7KrQxHyxD
niOf5HKqksPQMe0lobO2eCNp//c1MGy4ZNSmEXvWWhzRR1sqTPiPrIMC19J543SG
RqeybS+QZwlek7mgmCgV0W44EmicxzzUFoEIZ9D7sl3EzYCcDC/CZgMc+feNqLQg
ZrE5KcmA/nSW6n67u9i5GulFpm1fK95QdmVCpgZUlJ0lQWyPMl5KIT+3QkQhIqKm
uK5PNSbhRdW6g8hV239smM8rOa4vi/pg+UDXezCeRbirA1eg8y/164Ye2GvPfjty
8wVaQ+jA3Hvs7XUKFk9s7Hd7JmSpKcI38dUpDa0XpoMyX/uf8Mr9PemvnQaEC+Yf
zE8NAEVrwqVkZ+c5Zz5cmUrRdXXvVzQ9I6vnZgg96vhadp/xi0ly3yT8H0dAC4r+
dz26xVgheVwOGgE6KGBcimedwjlXUvzXDOJFfSEqcJl8i6l0phj5blXwnVRUFjzA
0pfuS1Wn5poQZSBW3qSdRz0tBbVCbuX2rBrlOtdVM6Tj5WIY+xtmjeUjFbyH1hRs
FcIEpJxZGR5xy8rAzcegBWfhLJ0JPXIwbdrnZ9ZB6Ivbjp8C455RNBr2RTcs65L3
DBdVUP9IX0dI0qQPGD6EazswYMZ2+pInlD35rQkuM9Qxs9y1lHU2XLi2yvKH6CkV
y4zApXpHIImqttBFP7xH+XGYPUx8qz3CAe3GBI9G4AnAr9Sb4/thhT00DBNjmcTy
xgsKUJDMadAlOkrLuZbHJlNLg+CODTTTQEJmrdzN0V4/j6A/GMpL29dKjfPHq79F
7cCNZeP88FZgAeAc64MectPTdhYiZc6LAenzmEGLTqYwGAmFgusYbx5Bw3HHa8wG
7GEKLXf7Ehvhk0U3PMNVoAC6i41tgBtPGgoYMeDNTSoAHgug8Bi4rUktRKXd/8Q0
muxmSAIsdQgOQ1kN5ldpdBA9RjlzeMGD/uSnipNg79VpX8vQL/oJfxj9jxljFMVy
8U7ismmhM7j256J4+r+Vo0Lmc4wUKOcpWVdVMT9imsY0RsfE0Q7o9zPcMyXxzbO0
8Yeo5krZUv9SA+CtgoRom6IeQdNMbyTVg+LePIcflmWp8tlwGtaN4jaHTX6jl/mE
JoTPwoZzyVDNcuPsU5DOmx9n2iUB3DPgsx4zhtpyiES4MNCcdofyxzE+FzB3KS9x
ltaxVlsiGhtNRtwqse/6tfcU43RRZshmRDIhDbED8AAFl3tUqdhkw1xUp0mfN+WG
vODysACHWqVoaZoWjEfx/xuzXi/06jqTfKvev1Q5pp4xswLm/ZtECx9U6y6TOqdO
VJZDBu2tFoAnjtbAmJ4iHQxia7a+do+WqrwNiQZRhaEO0Jt8MhWaV7tQ2hWjpv6I
7UKfCxccsXu1GXYFMWS4vA+ytDmho7+4SeTU/dQa5DT4ST3NZSSENsGPYilnqnme
ufL272JrFSiAsppLxu9Mv44O5CWStdBrUq8rPD54VSvAai38Hn7N+taRMZg7Wmwg
QZBzYJ4E6hLb+Z3vScpNZGzB01oAm1nbShYPJ5lo/pvSyHBNAKDv3Nmq2u7b2fgG
/2zjs4M5OFAGFTosZTN7Rb7Wzeoxk7dWtL/eaWOOitsOw3W1K5M3XhD2zrSKEAUI
7kLKKj5OiWzzYGbiAFYvCulrMwecRUOnnSnBV64IDcZpcoUpfZZHRvTfMmQjicHK
zaTOfPb+20JWSlg760AMm/XwmogDclrI4QFL0oVio3FwCd6axhf12pb/DJXrH8jQ
x1H1KK3H/s+AZF9TYW3/DVcx8ifYyFvbf24H82EKhQIS4STs/l8ZpA7UmpTCYZmb
3rK+tIdyDY4eM7aH7r8ge1AhjpTtp63C1e9YlI0kan4+a2T8x4p6xt7dDgDW9gjG
sTWHHN4YkkmPj3Agv9X6ZpWdmPZp27MVFVOb8nBqjRdUjqg8STeOJOqJkZoDb6rb
3jKN0GInChCjF0nH0GxLx6L+Xf7QuSdamFb+wQzM5jAPtBbOErtIECZXRQaQ5CJ5
TknDdriQ+wuejIOc1h7lFuLLn8sTd07pWhp7yEEEvGwuHEUUNoawKQz55fC/C7wX
ke5cJYBN5k7b2TqPfH3kXowRSCt8dRlUE77i1Xkk1p13Yewc4e3UXwTuoq4JihzX
MTXHzKSmf0z7zM0MhYUWu+IGYHYuOl50sQOabqv/Uyp6O1uh3Suwxf87sSIIYsc7
ZCmHxoAGhZqrl9emlSws0V0RyZRsV6RCZL7EIatPE3HNWjfnJpaE6XqmUpU7vU3F
Ddorl2+VJhjnA5ukjh6bZe1rvFekCaW5r61h+E/gwcC1gV7NqmZ9KmO8U0Pu/vnh
lD1YqGLI8cHHDUlOGbTmZyvd6fkqTp3788pxxq8Nzuz2JKhWuu2YJwZM1vaoP3F/
I5TfMCFejGO9DS0/5DYJxvsYlbqpktGvDIHjtOcah7IBn/q3SuNHk0htMKMuiD+2
dvRrjtlGQXTpd01v3vfwDIKB+JLHCaA7FBk0DmdckdTwxAnhc4yRI7+wsi5gdL4k
mNDUvKSPv99cHyjZMQXTUt1xoN0QgWDw079v4WL18HqKTtoqwjjMXFJchpMtmkh/
/9ehE1BXr+UG5tvgvZN37obkL6TJuJi5E45DzVZBVmhxTCaN+zyRJmB7QWP8U0JG
e4WEz6rukTAn2YXh+6423tef+o3J1AUuM3ESKkHeWYjblHkTsL4lRMxDIF0De4WX
ANOM6q2nk0WaEDqfxiCpBT1daGIJqhfMS6hWxPqL1HUQtFWXv3YnELzcAeLA6zYG
RF/kaPSFjlfasdCKzuMufDEbDmUHh3v5NU7Veu0tIp6sTtXohShPH/1V4eq8boMT
LxfL6YymTuESlOmtJ6KaN3PWJdVwCfh+2C7uinEDgXwRMy9nvhmg59wa0FyqJtze
qklDKMnk1reCMCYX1rmByTxf8/rG7mpU/wGUO+PP4PUuV0A/XYHjMhEC3L7cZmmG
cwK/n70FtkcJf85xknWS1cREt+9yU5+iVXVsyeqX08434ue5EU4VJrTj7V3/TV6J
RYV1gotCVigh0P1g6/DhjYBg9yWoZkFIxmy1Ku/IwQ0vzxXetaVItEa8aGFBNJum
K+C2RWfX9Lr0zCAZTmibQLIYIAeZSyEer5VNOo6IhzjDQkmXuvY3PqtAEWb+8w/7
mph3sszcQCAFzaprSypkKNTqxMg4I6J8tb4h/tPYqUd1IJXlAeUjgsru6COogUcT
advuivrTv12TyMzuUwRnm8+TzkOYkj4N9VKD/9JdEDolSIfezasaYv6D2bgCg06x
CiHdH3pV21YGpcZUDWDcidpDAt5Pn3qQJ0RPAqvCrXZedXwVnX1m/hY5pUtpOIY6
81/pjh7nmFuNVZvMe/paJ4JOgdEparoEoUkUTvr2OttuXSQbptmlr1ptoRc0qV5L
PbJ+yXmdKsST8tPcwgpYDoVJYQP/B5M9HySKBViSz8xhgDNmep1agddh2cXmX1xP
6xhuR+zkUbNouYdraJztEBQ9BOaCQeWaEJzzhpb8A3cxYLNJtJNcckww82hwAuSH
AxS6+2OT50JCCIYg+yzL84bcPaPb68/UmTxpHdWMG49b3kJZBDslsUglh0Y7ewVn
fe2/C4Bhds/lccaHb2mTY2FRfw29XZqfAr84KSsi5oXtG+F3YTHswWRaPoi8XInM
E8sYit6H+u6SguhYbkrNohnD5gyQC3y0s79+ABpkuZGF17kYNft7EUFcMCngQMI/
g/bwovlRgR6QLoj8djgqbN1scFjEubsCuvsotBTfuE75edAysoWBQf+moGTPRFCw
uPcxuy1NOGnjYBBnhsbxTGue1yuAXyqfWa+ty3bfLdvmWJ2QXvLAINS+uVV/igfT
lm8cD2g5M06bZMoCRwOoC5hvBsRL27YtBAIOnJKMEmFQogxNjuy0iU0xNSS+sQFX
H7uZJRiS9JOe0PzStQzvFicyXA57Ms14v1n2O5vvIy6Zxf4Nc5OqiUt583VkUehj
dtflUNrDviyP31HyQGjqvWyGsRWRobiJI8tSIl7EzYAjSIiY8WG+9POqt79Bc/Pj
/LUP0H6AfjeNKbwBq+tlkwJR7MevYneiTwOSYZtmZazqp/qBbfgNnwSEQ+HuVdZ6
jK56GCOFu2a+41lEy9D7lOuJEmmI5AbAkl6jY/J283muVuc/E1iDthNmPdSLS+Ka
1S5Fl6qeJUWLX79EsMUsf3pXvb234dZWxJ2w4Nqa6xd42seepOAOaAu87a32XT9/
KeXYCq8wWSRW4w8jcuB/BIX/Kh7k+MKhMcv8wp3oAyGD+cUZNg3GKaJpIDXAlR8O
heUVsii0N6/eNKr6G4d2j1s+l5VgwG1vjBCW4lN0uTSLEA+YlqyfugU4wY6YzwDD
PztCBQL5tsOePkELQoG2+cBZ/4F6EFHri8+p8C9aSlyVkfBW09FT6XSoKmMxzgRK
ALUoqF4kxsK5PSV3CHq/TMCJ46gmf8RIncKPZOfoO7RX3OBiiOGTtSOarXShvA6p
DPJ0sK60Ew5Wr6vkUE19tiE2OGOk0qOU/xxNWyrzdP+M9v7qfbb3deeTGfaUK9lT
03RRShViAWP+t6oGKfTVyWnGXQGW1x13H9LF9LqjxlncZL9bI4lGQJLFeRUFEGmP
3bqgOEbk4m6Yb6Ao7AZTlIjTtXf3QtpVEv/ohj2/6FuVtF1+2kryqb48+rqXO3Bf
FbfhweQqqAFrAm6Itfq7pfiVUhvEgjlo845KOomfVlpTrJQ1vPT+Gqu/YtvkzGbe
MR5PMLvcHBwif/kTxU3WfSAr6JkKnNMgKERuD7aGJmY0L2a3FfkwgwRM3oVe4zaG
0KrYXXgxbRE3UY948VuvpQaw6GPbBePncWWovJeTyaY+DYxhMMfr9uzOUJLf8Bmu
cgaJ2unA3P0rGG5vZCWwYesgCITjaV0CBgP03PflO4yX84BiTSeOrQX3SflI51p5
bL3H/aNUiX40pp8q0pZyZ1yUV1P4Npqfv/mE+GMmELkbhK0lqRcCqzi6/iC2qhSE
65vKuUXSFE+kFnzHxCD8KLO0If+s35upzwCotrWrYWN4gBKO7IDgmI83VYUCubDM
zp4Y5J0Bjo5mzG+QPtmAuKSvyG5j/Z54Gp+ZtZ79u27e05JtuMG6EJX+iP70eXMl
NiCeiT+SG9xq75dQkNcMoOQ8V6qNNWW3fPkYmZZbWYCCAJZ+4JlBF+y3KaNXKRiw
xiR3Uk+xw/ayDRlEjj98DXfz4I5kIOZV6t51b4nYb6b7Ln+p7vERiTgM3K3t4DRQ
2Gg4zLOKxokGa//hf8j1kt5US0Q/EWsEgt1OixzMnSKIFiwcQ7K3JLdqtLS6oQSE
AnH+oqrf/GwNyn0VMDhxwKAIQ+HreuyzIIYt3lFPtqKm9qEYFSoJYDeGp/FgICx4
ICRT0HzlXNuAsRNgXHSkJ8+/nLiAKojFTsat5pFtvWHidaBoRfUTONNRjnuvazR3
WVgicTYZPrkJInBm6lE0fQgwl+YOHFYsqz0HgUn8DywNkApgjh/Z6cf/ldw0snSb
xpgtOrhjDekOFXZlhxx3PJos49bXxNRHr8LBvDef12XtDKcDqKAE8JNt7RTdN0gY
Q38g1QWcXeadl8Hd7OBj8NLKTTwDL1VPW3HuzcbUYneJR1du93FmMtPk//xE/QNW
RNJv6LIzC9HJVra63moOPZvNO/Uocg5WDraXgz2D+e3ULmnVdSo4+Gjl8+yAa1vk
5rByisnA3UTks6ibK4I1Q6YLuJTixZqovQVtbfHw7SpGH2/IgCQlqi1FSg4inlDf
5QPXefjFw7acDoKkSNRCAm8tmHZ2yv9l9hTj3zssJ5fOMZPNvW2TWfVREPHoShWW
M98HF/7zrJlGGM8WoaAU/GcbdK4jG7XI16cFtdjlGwCfLAqHolXPlEYF74D+reOG
hT+FyLMWu+WlSX8QvuBBs5eNefxHanxntJT9M1bBkThgiuZTNYDKMvH/tGUWCi7J
NkzpnMYQ9i6M429qUL4r0kI+ioZp//SSDeJdszaYIouGg2e0I5qpeWtqcNLkYVV+
nDmvpnP4gkmVGc/w0ESWod6SOcSwYyXz+mtFaMAAeZqzGFtzdWZndj2TlO6eiDbs
m0VDexqjmEOMV4pHgSfTej0A2BpBR6yoPq0gGd8LlUpDvsPMgYnUVDwarCve3BZ3
drJYGlnptwMToc95s7gt1d4NjNvwKkVa59OqQg/5IZJdMtmdEKasGdhiywznAQYc
Ng0oUYxmWhTg8fHjXhm5l69yMhqLUQZSEgr3tlXeht2a7jjX1SjtRFMvN7Qlm+Gw
3tMYsJuyiWQT9BwYKvWl1mJFirYLZ3elo0XZ+XupCCQ4PbwcT/fY4UrOaTZikE+H
xFu9wIVprdtqaw/IBS5HjNzCx4QCIEuKfALI6lpA58wk3mFcME2FX3GqYRrrUiXB
pR04MgOe+lI9q0HTS+1bO75xEzj7luPznhwGSzfUakk/AiUtKaBHOcbm2kUeLpov
hJdq8rXX01Ryw00rS8QVqAaqntrq+Yh5qEU5KmtTBJqx0Uv2E0sTyY7dIDzYvw/J
GXYEaRg9TJputYyruKCxw6saLEjhNmY90mj7SurBEiXxFwPr5bzO1u1R8S2qsup6
MC7aU0ISFvjRTiijsYU3peOch4oIKu2Hdqkh437xbjpow+LBQOYwaUQgBn3U/tvf
JJ0Bidu1AvxCFzpgl+ttKs5kgpvlDontwr5xIilF5diaxwfNeFk3QiaIUeoYhbon
uSz1Kkn8kIClaVD9G+eOCIojZvJFuzY49xFPKlfuIoSiSb4cVTA9CNnPqIUaugO7
NtdkGkD7E7yAQ4R8UOjSsXtKv5jf7MkiHti4Zwt0EiSuWXBC8xXCt0kaKWrzycfz
hnrKTtm/yWjtiMIBu7H7Mj6AvY2ojBRYZzI6OyjS0fC10amY9O0RqEVvLCu28gum
M19hU1zJFnBbQJjgXQHngwlut0fGQf2ODdB+QdnEbgX42ikgQ55ZSy6TwFkJnMc1
BawFELb68Ems7LOXnrw1+87w1ZYwLg7LXUhF98SxP9Pi7sdHAKYfMhbIiWuXUGPz
SSXgiIWbm3HuA/zqX+YrJIkJx6Cy1v+TPCBV0Mx+0Cz8QUMdSzAB/ddIQUmthyxH
CHFKf4TC8/EUdN+9+Q/2hKWG2/qrSBWaNCjewLO4i3cTe9YOl5skoEzYcJDCxj7z
3rMMJU0/mph8N6Yjuynal4gZOeEV6cB6TTJoqp7eLCiatPacAXf5DrOOl6dcV9D1
9YMF0oPNht2l0xJOQBLnfhEmBBi7X/CI0/jVBxpv8Axb2TsVBzKPypJ7RaU0VuzL
9ucCe8SzdZ246uZLAqD2hg+ZJoguxMa4/qEXQ+wv6SS/3pxyvEVbkJhj2ENG1SYt
t3FgxFz47n1mFho6LDFEpZGHTf+srGKFUjiuoUPKPl1sCX4UCa1KHipqzrwGMEb7
jXUDIOBYpLpHdcsEGJakVUJria5lwdtnPXaldtSOhvdcbuap7FEYwmGlzbbztt2E
FDfowJEkP52+d0CgmeFJ82nLqcKXLKtKdG9T9T171oUmnAPYpyVPIReIH1LxD2dd
sFypPhRata3zn+99/tazYdFkptbTZpuwnGyVvrPBd0abB1lbvlg5EG0IjFixIjLc
po3jUKVjw7fsZ0J95FUJnU1Ha4NVXUlL5/GinqsIsQcjGkbWQxgy3Z2vyIkZXKDi
iYakJCj5k8gQ9q9M+Nw06JKoh/v6ifiuppOqaLD0ZP+BgFV8u1otYxyfr/ORuXgC
bXM7MArNXUipqOTjhkYCPgdm5CW7rQEqmr55HfMZ6jDp1rKU3V71PUeqlPHKHON4
rCYZ0h+ygB3XPyaVoNinRQgkg0eREtB3XlxEH7brbAHMZSa+xuP252dcF4RtQ6mh
SOH92CHrOmPAcHPe1E34mpN3eleEcU25BHy/5zqhoWT0+VUzlbVhUYdNNHrc+72S
5jy3jkYD2PXJOOW2xfzt1fCrccoGJ8MBeol4NaOpO05Zv7v1U6r2+S4bFLBrbeqe
TxYD90T1Y2KXVKtYi/tN3QQAKwXWT0+JFMsTKtsgpgekP3WqbXudLpYV6nPiTP3W
D7wvY5VuCMrXfnmmDYOezUwH9EFEDJ9TtAqk3VhC0fdB0GnI85HuyEufuPPPQKDT
YQ6ruxR6s7N+TJCZEdOwJEN9xdDPc+J230YgoWEkivjcHgf3IvHlvxMDSFjq8beV
DAbYtxSBq+MRMfYSkvEMUPr/IKBo3FDFggprPRsOp60=
`pragma protect end_protected

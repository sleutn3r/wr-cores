// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VMvpgFfETj/JASidkbPZC4BDGoEwlthxvDy3CHCTOnlg0NGR2IxO2V9cR6Ucb0LJ
Cw9p/r8W7rJAkHWGHyNgpvXinkHS0iA1nqNXxm8QmovCv4iJhh2lqawV+3ZqnehQ
IoK+XZRXWWeWuV6r3W/X/CkwtnGiPoMWTxhtarIHNRU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 20480)
doOaFA2lOC4F+mT41xcEFTOvUK1tscRBcTzzgL70iwyUQWpCsAWXXncPvepfxo/O
t1SWcv4opVTseczS1zyfqX6SSjg1PLdy1ws6v/mJj77RIdlbvplItYvL8C3CaIIj
bCBAkzmIcHOVSQo1iW1zfgQ19VWTC+Hx/DPO//z6DHd5Xzt4XC890fpyOYuNJGoY
OCeIl/QLMsa5cOhJqX3n8gSOmDiA6q3IkE26AgfejDbhi8mHYrKEcyO7QYdUnNu/
gLZ1BkwaIZfYQfGqCKh56tpiU/tjddYfqJqYkeCxYYJ2+8bdcKmXgkqpiqH6INxS
fIbmtagr3IcKM4W4vTMz079cCFtFFIAZwJOJ/NbWlx8lfUD+evZ0aeFmYbileGjV
QoFdk8q/LpXRiUctizImXqRbWHDmdaTdsAoqs0TlTf5oUJhLsW0kFEcy8mDg5NoW
4TR8DVcUcTkfgGnNsCvMXzl1rQ3hPNKxhEsRVndXn7w8zP3aANA3kyLR2KjpqtJd
Jpia2xsVEHZjV8yb9QgHCOq2W/g/vQ1srNaMeWfbI8QL1MJuu0c7xCrDvxHHMjC8
JZcUtv8sqenDSH9BAAEBZtIM5YeSzozA2Sj1tOAEXGeN2Is1rEalN4whBX8OCcd/
DvPyMjzQTjTxrykfdNkriLUv3QBPftfsFCBd3ZmGyeMp7/tSRT9FdMq9xGdSHQDm
9g2V+LMxhGbnAezgtJwrWt4PElIc3g6l5nqjII1rw2K2EJhSZ9T/Oav7Evjr+Uk6
/4SldvmN/QyGhTiyLUMQxTYawoIxHHOtYTxISWCac+P5ynptny6DuHxpWkVbAmU9
UbbDzzpi/pRnIQlQXA3JYuttHtGGjb7Oor+Z6s/QwKWaEwlcvAumopn+DbM5hYtv
ubGSPwxaHXs2Ladu7hCFLGsuC52Ce5f7+VDQKgwZK+TM2GgiC27oUIN0R7Wa4w5J
vXVvocQ/u7gu6m2ErW+9JXgNdDIq5eCpER8rLYsK6657xSFzZ2dKyumPfg3tnBCq
dEjfXHbZdLYU2YMY8yfCtGFOUvtNXG0JbuFXSzKwSOJFXOJw0EWLlFNjCzwobuZr
fjt0tpsfifdn56uQYN3F22fBpo6r0sqM7aoManU9yL4GHRW4PUbN8DcxParVJAOW
fr/FWcV0611yYmAavLWbiIjjAlbnezVw25E2e4zSJxzHBWpASiRJEVBPCvMJUENI
AKtmoyXFowZSXynywzAhhBLl0yd1XnZ6G3A+eVb3EwMqB/AON5qlJJ+0v1WsDKhL
Pi5qp2VckZK1zaf/0l0pFaw5hBxPKS0xYlMbYRgKdXhXhTa3pD3SAu748Y9TEtga
ujdfGqZqLnJIhd8ghbIFb747Q9lLDONTr92XUDuZifw3RrYq/ZMT0n4JtvkgPrBv
UwQ5sh/Riv9HBr8vMHpdj8bUSBZ3wxG9JHH2JTtO2L2eMGPTT3LYvS5h0PuoWGpt
DASgszaPUYLk0fLgrHd5CVFq44BW4tkgatzAzoApXbksfexYmFgpWMWjzEbiLt0g
hB6gtldqm/INXF24KlOfrj8R1dq+ADhSnAuxP4mNpfkBxsjPsdmVmq8aW/GtFemJ
sTyM/kaILJRiKMDyMdyioY47J6T7TmwUWPcv48+TtHd49JydnH2izDDf1cT3TZ4b
L0bU83Mkn35256UwfPAGyNbxYAJqZ7fsK4hVAIezBLFinsqu9kzRxnxzbmjWGBvF
Hf7ZQ4DQ9OVDjDJX0nsFwZUntKyds0LxrfIpddA2oPM7ANVa02JCAA8w3E0f/2gJ
rzBzznT3bGRU0JyHPY+p5cm7ORnXcA7zIwSsBKVPGg4vq3lklWvjUfC4UhLxUmBi
FvCkWIt24JFMkgC5Taj2mcJOT58mwbSKnMhV8/3y6d5Kdv6VxasRVUhPtJtatOvL
mGQNq/V1F+c4UsZxpY15pzBIdZ6+sjzYsjDquZ5aK+DqmNpZRxIK0y23w/0c5ZTV
xeIvK336c73m5rWxUSRkok013IR7V2ldWmNgyBx8OfaeLuHLihHPusnPXKbet+/G
GB6NaY/dI2JmmNG5O6IMcD6I/axkmWXe/CDzEhojRlDrnIMMYKngJBx1CrFSBzbE
LMS6iVGiGewuKMUxseBypbbJzWPNCDGs6HB9FvGcvcm03eULqBnfIrDfOYwaJXpJ
s180BFB4EXSsWxLIYVKkKFzOcPjRPkBI7IZeXQ5xA1TDYJsHBWnugaYydam6XWWp
MptJywRhgLOa/QNDPfjxQdylmAWdM8lJnerkD5Gmcu/Y/15by2obQq4719MpeSTC
bqLWtorj6skffUTX9SVO2eGjGX0GTi9VHpeZzITSnbhFbCPmdaNCB4azndkF2x8a
eu2NKP3559oRQ7SKL/jQ6UGo97C3RCCJ1YnfnA3VKOPidhqJrhN6uuCiWn8tJDcF
cP+KfqOKXUJPAuAe7NShv9AJQ2py/Clyzh71CMK8ZopfppmIuxLY6HMJcpEJrk0K
3YnzkQEcmlpfbFy6gynNQDRkej+shB3ETla8dunDafFj6J07P/+QdeHZyqprM74U
RlYxXtkEQgVNMJpQIIlv7BNFHltDnQFgjyrKiQVgAHPUvyAjxtRsrq9EW+U5TImB
cpoRofGhxslMQtA6pEhJT5j15mTp+1iq5en1XYk/kh1+3rEbOS6ubhL/IiNrl9gl
7czqsOgamSjgacgeLWgE2j6vEQkUlTfZnQLJwu9cPjMUS6AaxqUe6V63ZJNlrQUw
DF4NScOfGwtTxf7j/ih3JQZ4IP7vWRzLpnrqX3XJUMFaCMM+EtiwBo2MEZWo+D40
5PdFRqfz7SrYrbOgXmlFVnLuUEkV1EeIX1fAbb+f5QMiyYhiPxheYadccZReFX85
ORhfZNeA0iuhNeQYrMsj71A89UxCY6o6X2Fi6CKgH61BtQ90yKFOwhhmc9XQa+bF
UcPUfgdbAPaPV4Ltfxj8kuVcivSRN3IjxbuL1rkn0KvlyFahC/oEuxyi+D++pNmY
jtuRFuChLrtdTjfJ8pZrTt46BZRJu8PSufgG/rvwPQZhF6ihi/tbyEcMXI48RZRj
naAQnhsTjRfd34FO3IfKbi8ZFtU88uCZAwG87Z6zXVYohaNH5XEl+L+3KRdssbEB
R2DQkvTjBwEV+X3EAMcR+CYchA7JcgjD1M1JEUG3+iAcXHvs4flJ3uaVTyLrQv3H
WxIfKaCrbJlpkYef8ZpDN7VWNpCAJyVspk1Z0Qr0dtOhZYS0ias3gX5R1MwdEdog
5JTpGaS6NQI5THS8rSpXGNMfOxnLVib0caLCVXZ9DSkjM0C7ENNFy+hJe13F6b+G
mRLO0QLv9Z/7m0DFuIjx3gzYFiuDbGfMwea0WnuxUgE9eDgbbyqj2ZHfM3vdZ5O5
iWcC1A0rgHpkTwH15OnNIBTWNLBMPhhWLO56Sgdw1nhOXGxtjfnt7bhseZJ4jZeg
+uCrd8XyktBzruABeS6bDcXx/gokTH6VoOxkXMNaGh0CCKr5jYz1ej+lvRNN9vpQ
ZiIgQu+dvgitz6Gpd3N5g706T+GWmN733QVYUWRldBNzXjxOQrdMeaBP60Gj3yrP
obR6YLW8pnr3yKS6M0PFuqKHjkUHxvARtGdlpPNMpFjbxOiyD07z8XrFDgllUxfd
diwDj0y7YSo8zE9XsCwDL7ThvoO7LadqKZrd7gjT0TyUsdT8lKsOEaHYB/Fn0xNL
MvLIxo1VVxgnk3jBxuhA/XbazE/zy2GOUCgwzeBADDAPdGBz3P7Cj20eVdVLHgnz
KWE5AWn+TuhAe7Oz6xdF3ZrF2I76ZuyUcNRZ5GGUHnEz+quBacI34FJt6u/WV2W2
PFOzsqMvll+sgrxDEKY6zr2tH7LxDkJhzmI1g2ExLdr7Zj3bhHpiTjEqzdQkY2k1
6A/Idu3p0PnHO08jhx6NAXy7cKMRXdk3nWNrwFIbc3f6qdPpstiPo/4LZ09xR/YF
z3jJdhkuBMpWnWXgCsLZmfiilLzCpTXfL+YZKoXp0ybVv+y/PwJzEN3sW3wJVHY+
c3S2wmNup3KW/OSYUZ/HRnaHWixAmMgmq7Z2L7TLPeUgeW8u2lWc/H5Or81VLI/A
yqz+oMq5eKDYrdDCLxH7Vrf31ASySCfxsDvALVqfT00RHFEcdrHatoASQ+Rl0pko
wpYcTp+/amjxj65TWQnb3VcRpo9wIDuLjwnvJ5STSi8ezGM+JQ10ZXKLBO0M065I
wpJPSlxVa91OnuOww+jVHcMNzUO/vX5UREL9VedbZB8pr8TYXqTWelpa/uCWq1wE
N+vT0yQBykct0PEQ7TA2XPz7ol+qHX/TCaPC9p+n4M0Ndi7UvaurQwCmLbu6fhFc
f7vcu9gk4mVJKBO85+wfTcsJ2AtznDEfzf1DmAkC2uJoiYvNJ4uJHwrZJD6ZLMAC
/t5pVb11OmWUC+NNn+3weAECX9TxoRwej0V64m79KmmsnkHED1eiN9LE/QqEEPwH
Us1tx2rQWSOpu51IkMz+ChjdnM92uXpXtjwQCB6cKKyM7zF7pJxNrtNGDGt/fL/y
5/Vl/RExPJSGi/cqlxHb1EmJjrebwC8wpN5WVIfV7r64wMiMCPn4EOimnb4gecIh
ln42D9zTF4DxvnbPDAODiG4pNZJt93vL/x/+eaQv/Fq44t0Tvhh4mhzX3frwpttw
LBXnFzGsn0YukfZQRj6+TqOiQiCVO4BBWOjwUERzb7OcPVXdtKTJz3l982O5Lxjf
u9IUo/LbAmDLNdla9vLN9dH7toVYp9evafF1JWTF7jekyRNgsc04qQaAcWQno6Kr
N8Nd/SKOc/P8HZvyHZ00NAhsoblzUdT6aPC2/gjYj/HwiKzRKU9e+kxj2vO2OtM3
nrAO70zRLafvdnucpH2gRuWNhUKqcl4PxTRrge9Wc+JowzvRneQlPGs4c/BURbj4
xSNkZLXM4rl5ggPYm+OGbij+08jPA6h/CMPrS7GwrR/oxC1zJIR6hStDDg5ei9Ls
P9bbdu981x7Vy3fhDAEx7eznnsZ1eJPFemS//c5C2FS75jmZhapd36vjlMnaXUgU
yakA+8bZy1lBSnfzEKxuHoTPeGMJX5osvu76eZsC9i2pd+QNqZphMtnbP/kzt+oU
s9mIzD8lzdHA42HvzADb0nnbot6pyNh4Ps1F+UcfYKGG01BD21sUkbnwRSuvaMFg
AKJJdm/Yr738iFcnDff+1UyY+xXALMtDmaiMsyyojl4880FQ7/3C6+ottGNg3Hdx
hpC2XfEyAFhDaGpHFJqo8fhSBlNhJxNSgpwqgy7CO1gFjRFmNe7kQX6t/+hOkPEB
r0k80kHYRe+koIh8v7NrqwQb6t4HIgcX5Dj+TCbAZBxeyGfyqathcOyxN8K8fwAE
BThOqMoxFYGwWjiyJeKjV4ELxvfiZy+FjX8hHbSzYXWiapdZZhBdIm65C/aNPd0m
/Z9Of3WMuRqnNwnSZnaA0uQz/YJZWWy06EAxJ8yIqvgPwwjyjBEuwvk8nSwFroe7
JUWHIDuVFsmQNGwivooxS3auIoohMj4RMIWsTpuHDXMcaazmT4YCjtrhUvTMB/6g
/RsTHN9OLW+MLfUbM1yqLZXaGHeFTvQdOMj0+gJzdftdqdtglVbnwr2a1H2eZ990
F9py2YhneCKM5/X48Y799/BGYa6TTiBKfaBBal8N7QZx+Wc2jMnpXvdjmsCWfY0U
48IOlUUdEk4dF9aa4PMekIr6ENKgsQBJrWVwjBYahymzmzzhr8tyVnWz3+PYVZmI
aZ4pYOVL72dJ6x5VAaAKXlgDpLKd14qHOBNTEHLsLEZkGcSnq12wB/ioleaQ6bQt
k29PUVzAcb99ZrC6MKCZXx8GBbIEiuWknWKrfih8h4JtQ/lul3IYOrOLobfOlkre
5m1nF9ktWW5OoVXdSCsuJA30osNWyAIhOP3i1/NYOlqCDXlrZs5FhIUMJbGWzvVM
aUcOk6EgbwcJ/9Ew6ZKP2EwcsBKXaxc4GvMQfVKD+msjaoVQ8SqWtwPcuG5DvH6+
iU7arTaJENPLqlGtI/L5Yvb+Jw43HshROukCnNJh9VlMP/7NuPe6A7mMsCSwq9mZ
dHTIVsRYH3bSgROda6JIWCiR4hHzx2EUKJsJ/lf4AGzt+Zu1P0kMuqMVBm0gt5Ui
PZhnTcUDakH+CTPgzcd9O1nib25LkUj3OM1bu1wR9VxoYzsnnfFAvXLLVsdgvpRS
MWe+Fbmucj8E8aw9iDYrztSp8hTSi/DeTY+E5mYnIWVELaBlZp3Oim3wapLJ2H41
sLX2fabT/PXYLBUkDgj7EdBZxNY9E7UeQ0+XtXwTA59xsxoT8oD2WsPNkihE4vBO
HzeDQHvl/RSO2TRL1+rF+On0jysPvEAuQbu4tnjY/VwA28vb+Yh1xsHoqXC0/qoP
wIrP0jaq6eHltQCrakOmTFlE85vI4LbSIe9sk3VdUFHr/ljhuHZ8AMkjRawX/CSC
H89o7dtLN5mYrRCtCRa6yv+I/Q+bfChwUEEkNWMGtQcAWxAKwxHZSV3nHH9gtA8b
vm95+z0nJ5I6lJm9fCo6dCNctkCicbj6Lm+x3uiLDjaAU8/6fAzpeEldHoGxJDWN
ZVb2yRqyJ4k2nre6+X3WVlR9nZWUMuOQPjC+rSQ0MloQH2XKWNDcJ5K41F0E+ZAE
4IWy6RgspWIm6Lk8rWeAkXg8GJvLzC9msexbH08pZKA/5H0XB9mu3sD78MrwzMrG
Fm1KGy5oWZ8WqpYolXc472zdQlJwqXcOrAWP8QN4R0n/5kULx8el7fkXyEuxMqgO
k7ZHb6XkGqDBL7e++HYEiD16FvhCA0g3FwNkie7fRnajagKhQpYqf74HqEjYarO8
l+v3AjSpyaufwapuqncgKlG0clIe7FSZii0EgWk5RXuuoUOvlSWblHKT2BD3i2Lu
ibmdVdnzDDcdlBdHpIGVuOaOGuJDMHuD5Yz5ciUNpnBFbhiGrbZ1licqS3g7fd/e
f4WZhVVPfZ4NSGBsGDux5Lt/0JmQaSPYmrIuER9JWM1I2LTm7rFgRlQngU3snjPo
P8N2ormQoVHegqlXQrdfgu3VcigaBXqGH+CTwfLZ2L6wfisrWmnSb/0QXks7LsqF
uOqHEabs3DY77s+dnT7dUaE5FvLwyhkj7DkFPWBptqBPSjeqMB6I1HC9dKXIasah
8Or3nDjfpNkmtwEcsolFY7QQmz2yH1gg9lhg89g/mJsy6gtwy4jBDMnp4iBWPc47
/xH2r9Xs9vTWzTKIGRr6jCDpbfHzEnVtnHhzon+qffcDHX9vLwDUtM/4lfDLIjTc
dFLvlskW6jpSQtO8SIeXXXhYmqCFDrq4orCB26QZRFf/N3qp0SzaFIMi2OVIpM+8
f4Jbgyf2CHPc/N9yX0ymmZejfo+VAMHVmnK0sqe4W8n22pIVxWFBq3t3J+au3FUs
KJ1CJN4yoAbYUJNyCIGkdhayHm/uEbY+H0K+dnF42CMM0+p6J8gQKBUsx3whS6dp
dssdHCuukGpvYxQyheGuZgKoq5akjeyr556H6laMgTccRsjE3m6W9JjFbtNGSpJI
DstFxEE6keCqItY7QXogw2HhRBK1UBMocuhCITNimNvwZmWdLkwKWINgKJHRm5XI
O/Zbp9JielzpXZvQNZd1m3GcJsw2An1fL0uOYyBIGjwKinRg3AFv1zRZEce1enJx
IFj9VXMFdj8CAuXUV0URv40QgDGJfx1hzca6fJu+bGYFp8FJmM5z3Y7e25HuGgI+
oGpKhb54ffziGXHGT1DFKofNF8dur1r7El1x/pbPopD4P/f4faAPTgBcDWDIvAtp
Cj75DxCLLfSWA8UiuwoQQ6pyDxXv7gGr68LTVylZivsZNAKNw6NmvLHGsgD4UBdJ
QbIQTiO3+5rWuWFaCKOKumquo4N36g845M3JfcbxBDir+CVFGd1kxSVJOGOJGwL9
bnz+AzqnxAVciaMQoJ2qUYTdGDXFyYQ2Oyjdu52P2vTpOEWTk55pmZgmYCWKvN46
2FpBeDCgvbZ8Fhk9Xk+iaI8OKwTrYlYTIJyG5Jz9NIihm5OIXO2kyPipbLj4gGcc
tkXbc5Aan/SQAvDszQPwo1LaHPVUwqmJuQ6Euq04LR+g38IHlTOvvjrSNySLZlRd
V1oobwQ/tzGQkygN/Q7bd8E3gvihY3ngRBY1hLqsu4pKSOjz4IzZHSu6AfQ/2Jy9
1SvPCPB9NnMiPVJ4UH4huC986KId1NnW47KYhk+7G6l17YmclPoEtr+ocBPRRxu0
RVGhi124fpQjoLMzVBPtGQV57BQ4hJt+ht70/j3dBUQmVkWp+9Ej2fLTCOV5eqCc
3jSCtJ4GJ8ix05dKWlRCCogJ/2EfeIyrnnMcebw5HQZuFGF8JzAeB+c9ETQcbonl
nXzbb7PuoJL3QFZFpg2BMEhhknJJe2/TygboA77NGG8+LyMFg4aLI4Bjxo+LAaaK
oKYH9lZIsXxVkWuYaE9APvxKqGXtGbAbdp2PZw8GsafWZ+GazVqcEy0DkxMQANbI
KEhAd5Lkd6jm4VY35TEM9y0jDNgB6q7cQeZbCvbkP1CvmTaoOfTpeeLtNKcV3eNd
d06i42gmysD0hntpT7TDbY48lMrCXzIyvRY71Lw9KUr72ucMIgfN5j/71gWTZaP6
PvKQZ1dJ/Dn6l5lktDIlhYUuQoYj0bP5ULqh9uwTRnQ3eVc/VCZvsYwXkud+8yRU
3mfMAYE5TTw48yenKjzqFFnGS5EXenaQVFrRsGUGqHKjfA8jOgBbCn/po6BEVQAy
eGMA5RjYrGNImOPsaLZjTTtOTuTzN4tu982qGQLHRhmLrw3wAJhU7zu7s1mFnnI2
FmF6rqpAvsNCM7wpnvP8XS+rCrY9iQJuux53o8jXI5C38bs2Mq1gGV27/2+HtQm5
1LkJkUewWksbdW2qPSvgq7bgf96QmKZrFWJjaHLhR4IBswwCH3+tZ4neNk7aa4ns
RWoGaiCuvtB3loGbsiOWe0ZYeB4mVX333AiSoexycrs5mlNFzHyDNwMsOtz/BArZ
FL+YjUNLRAb6W8344E2lGEnv95rs78rcC7VLmEtBUclASjDrkhdidXS6/43nnkwT
GP4HbkYAnGLNawg+xRZPNkx4TDEnylrGQAF22HF+HNk8BJ6pYi8UOdbtdtRyoYZ2
bCqgeUEjT3RIJgFbNPn3RgqTJ/ajV83yPOWi1WUOaEDVeNTBO9SwKRpRI52/glu8
KdMXAp7bhQ1KsaYTKe2BxaAz3WNk242X4zUxR1l7qX27eYMzyyNcneFIuO9JiQwI
v/XrgLopSAPyKGoqScrM49GqMlVFo5ynR1k5nKzrJae5iM5zXr2ioMy0/T0S4rEZ
dsl3sHducUvZ7S1XwC7VkB6LsXvoQEyDXEQdhF4oi2JfmRmpBd1g3eGFt/HIFGrz
ENZehqyllBvOHp00oPHscAgJHxYoXtL661nTg0ofaFue2Nu/hiDl2svGC6+kp7Sg
J9xqz13tMDGsAwlP/5rlW8ucZ7si9G896T7+4iXWB4Z3FbIHsFSvHGaYLM2mLx3u
sQbn9LaAwtII6Y5hG90Ojm4sgR9YI3IftPBxaaWhC8psmq6D1dKURm3Gew4zw0mt
Ur0p7TqR4va7jF6IuO+ul3y9EZ7QPtGFBdQNOYYT/14hnDo2BPHzipuQ4ROroivZ
zxlJv6KcYPxNeWHhN2PIkHwSyTMpFwo1TPxDzu21jUOVLjYnabYXBj0vV79r2K3x
99xDNORKjTQZAJQZDaecrYHF8QFo1vPAZdBADHX0jlIm4NiHvtORgnmoCoq4oOoZ
Lrwd19a7d4f7Ql+UIKxr0WNVJ4llrPniD/DL0AHc1dlqCZ06/3k/y+PakwID4BmU
Bj5o7uV6vllc8w9gZAzUhenZufNiY+F/iMf6iZl2D/bf8rpGi5XcP09zAlT6IY72
oCyCeo995U8Pw5kXefWVNQG7xEM657IJ/2hQZqZ3b+A1ARp6QQ/3uIoy3mPi2+wc
jEZYUrdjlFEd6h/bLv3ZPl/hJfMjH64os4YHQSLF+V76u+2TQsimBu/nTJmaJLAM
BNtdrbzNVv4Lak5wyXrkxOtRSChVRl0RAqVNCzDj4jGBC29fpMl4V9r/xU+QOxFV
DJkfAMm0uqRdr1TBDGs7vIagK885MnAIb/vl1+DF+jXsXh1uavaXIImcauvoGl9D
PIH7ZVcbik3v3aejTsnUsz7cDNjvKp0gmRRbfwDMk1hJ8YfJOct8hQVEMtZwHtAP
1ee2muDJoNL9UThCY8OsYEViw9emEj3sfAreO9Hh/m/nO6kkGX6p30b9TuspZbjW
t1MCuln4Uo6QXQAoA3x0CyWf9Ce09DLhEtaYbNkYcNWq2ks15buOu1g8Ekk3MC5v
fkm8dRoqG8TXDXjNQDDwkvedj8CIqG7QrBrGdFvLjHBTy4FcK5Uwi3jebnJioipD
vc9CovfbPdYjIXmAc8iU++FY/WKfucZyZO35ozIg/aeZePEJeZ1jdmBpdkeOTVTV
2ON57SEDI0PGRSm+PI8gMmpC981s7xSh2t0Bc+tOHyPlqckWjKtaMrObw6BRH/uw
oDALk+DObdunsKk537Tnz3yWhNQh7FRGyg/LHj1sXFpghg+kLxH5laiYLhGk/Dgw
PnWEMvp6kLspowDQXgzRcFs+M0qD/4dXvcGAJV9RG2KnxkOcIhEGC7LVTLQVjaQy
nc26p2Ngj4uHJkOHJdFeMjJyqMDsXA8FT3tksVQ1f3ddWCMJ7HwZNRXOZ8rodhO+
3+vE6c1VVftTXICONa2vqJAJkZX6G58+wEGt+RnFeRtQk4cxsRbjGv8fdEDIgZ5d
zIYmu4uiLG8Xms+W84UA3rBEDj9mZqhMjzpyLRiugUu2Wla/U+Aj8kZEJFKlHj8n
LFdLPpzDqE9xhRMmPT9vEU2FmmPtCn6M43bIZnksNUBTaIS8lIi2U2/n14HsKdlX
EhLFRCZZlhwq479mrQHI1q1zy/RiuNkdwkwqEksrWk+aa41Eo3I4PzlLs79IzyF0
1SOkRlqE0ADmyQQ9UHJ7PGkDK79l7WfuAsxrHouV1UPtDwPS+qc8ct0JC2W/E32S
9oCv5/Mgceaw6rZWBwPKShZW9SLQ7uZB6XZjoSz9H8iQLMo7mdWFLZvVvxbIOm/R
O+XIp/H0NYVfEnw5FT+6buQ/tQuqWojN1Aagtke9vJCmG8LzMu8zInbt2RJ4PH3O
MkhlEr5kk8+goZ/WqQGK7tr1y5edp/lPnUAzjeVmLiy86RUgMjXEsj6q0aIquxfK
NQHd8t1fxcJMvC2IxTEEhBpJ6FJsseOVEoka/cZWfdtAzAzWAzQQt9enpuClNAxv
eT0h7HPsSGzn0JyFlbgZuMYk6NEHrgppKtrdkTzG6NCndenmPRADgVJ23kUANT/j
1zr+/GrHQWYM3QzhpHXTXFf9mnC7QdrL+d2vfXB4XmjhS0harrpo1xSWko09Jp55
x3ArJugsbq/yAkVmuNXaPwTM7mMKvWqEx2NnVr3yzyQgOKQkE4TQ2bfagWMTnSWw
Znyrob8zOcyxtVstCyx0JNgkDVZs9poLgK8Qqt/hV9HQi0fbLx1IhCXAwcmQE1kc
pQxrOFNh3shk1AKLlys6Vo3CuBybEiUjEyyryFXWDSEAyXuJ4Ms7Ovd4f+9Eo67H
qvJBECu46IGMRulzEQAg5wKl3wOFNAnQFlSB4rAbvFem4MCNG3GqxhY8tulDxOaM
oRCNf89lFpD9+TrSsWDD+f0yehQHiyJgY0cLLGeMVzj5H3TgqOBG6o8U5LB/dBMZ
dV58j5Yf71zX1Jz38SRPCDMd6JH6p0sXzUkkd3pIqphtPAAgUczQmfljAcoDTMkd
NgrlK3dGN6Dmfl0yKe1hgQpoRSv8FS9FbklNfaoedjtSZXg17kQYjpbbuvzjwW3e
qo+0BcCssMNJyVjN1XJCD8HacaVy3zTlPusTddOKXjWfQBZnBgHBVHo1VuIMBiw2
GhlNbK69pMZIyGU5STVuV12Ijdykdo9M2GKgrRVK9vbypVSWLG3oGRFpEsnZpXo2
e4zete72qG0Q6PBa6Pw2uyZ+cEB+TyJBkLzeKiwxoF6EyadZAqBA3r5geJliXUKh
hLmwb2DCssJWTAfMqRxG+B/svZELOTGzhQbE/8obOA8W+3E1Vp9I2goJSWHFWs03
vSDN8qQLX4P2mnN1AsfdhlWKBQw91Cmf6homcnHE3sXkcDlwKmiBqIPPtDFL5mj6
NfHTmC8cLPt+yU7wO/odIv9s8dD8gVLPj/41wOVUeAFd6hZLbqfFeYvBUNwbJDyW
gyRXTIzpxx/VRkuxcJTxylvy8Q1Ucp2/qP/a06rTTceKuAabfD9z4O4mdWsM1MYw
iWf+SWcmFrYEg/nS23MBg7VQeuNu+7cZ97hQwBY0jgxpYhjZCtXcICV9wWDrNdqV
YC8qc8Ri7Ju+Nfv9u7I8nkSJ3SC5SaYVAmhdSwlW3Hgf+PVzG6RSC0eUDUMQ9wCJ
9NIgBouzYyJBeXi56dEgSbHoC7M1tl7XGHzBFiu1TzzmhUGkN+8f3lZJPWBg63kt
z6rpRYRhCdKAxaqWBsq6KLY+FbSJVe6M1emobGfkqpAYc/OSkTNHNIXGYRR0mkfY
m5GZ4YviBT4zroCb4wN5vEL1sjTM++lLbyBj4i3gkai3hfsISl2GT1A3/aC9OzQZ
pKnJ8bR+img1hkstSkI2bwC3XhzAG8mD/T0OVE+EwwUVRfWKMEwv8vyA6bmNa2Dm
LkSD3ayXQxjoqnSi7RU21RaBD5lvRuRc9ZV1zaqs9vllGeX88zXc+0UtcTUyq/HU
QYM40uQufmo9rfveFqEgcaM9R+BUXE8+CqNfMdoQwH+0e4Ssa77kKzOXjlZckSYI
9vwOMBsJm+JsYlBvBTkxXiCDeuFWiMfePW0KMXOMS8aR7J81M2r2Ewh7AglsBsCm
g85MHEIxZ6U+rUQDsFEIbToZ2dTNkOyTcXG1LdeKdx7qwkQof6da78tH9v4U2HLp
7Tj7+fcxqs8nAFX0HhqtDujH6UW0FKh20YmrrsoPsro9PH39PPYSIUU/X86gGb+l
Oq5Hdl/OSUxfeVpJEbnmpMABlTCeVtg6kuZMZjUHH60wIpuGIwyIlcMNvjqJPttj
SRG64WvbgWmtBV7DjOIYLNI2cJc5EBdcPg6dC9aw69h23N3j7dQ2sHLYJ0UPFRTU
MHYBPqZwGGJvzULpYjuUlMrExUUcW4ZT1WBB/JkXg2Yi8h2vvFrUuQ+g1KtlI0gE
OKUas4LpJAuMcbSeHmkIgaqpYQgejb6/l9pXTFK12MVJIvSXGT7qGYWYillrPypI
24wFjUWhZ1q1ZdOl5Zo9GFucncJxamiUEEUcZdYxiO0tLMX5ATVVtY6rUeHnHpKE
zJLbfSsRyLoKZ19GIjxHI1jXJhyDUDSllFsUDvALWMCPYooZ5CeouGcEu56dZu1B
4Ubnz0RzmQ9hmsjrOUiw1yKWk7bxl0BLCzh8gMcgkGnPmf8a8Cpsd+fjv/Cl0aFi
Enzcbt6IpW96uQX5S60XF6seoPvSdht4md7JVeFTNCk0G45uGxj/NKgu6gXANnHO
wvDh51YfkZmxHVnsrxk68cT8PPOOFiiOPIDodUmL9wJ77w8axVJUXGOP3W/i3qqx
Bx1mQlULs3/RVWBj33vL3h/R+aQ9knyCyKWl7H+PK5PLMsDERhxxGK5QAxFmWKpO
Ipl9PL2fC4C/tOHlWK4P51qLVxcYUPny/e1fFL9CMdpb/4IEkPHgiJs3VC+CVR40
YSjYFlpHkDKk0K30dnUM43YrWRKFGdo2WV0DLmATspdDt2EwuAP+vo2wssQVl2dU
Qxz8lZqNuMeHer+IluDXw00Ydx4I14jB46ouDibKag4UGTg7On3hZN6/RJBdaB9C
e2QhU3rvd27JXuYDusKf96p/3KrmiA3nRzpAKZ7g8Aw2BQ3sDArfQzqmRsbdUH/M
RJT8oXWtxz07o/d9pzhv0+9sAGoDqLENiJeANrCgzBOLWREGmNEvnssELvgaBnF7
2u9DR2pqj4mpmkHRxocAuM0sr9iJjjpZkpHu3ZgqrXgLkJCQlg3RczuNdK1gbD2G
AGj2wRhTFT+TjVtTnAqpmzvALq/xBODXdP6pEaMxoKhWFPdk2roRPGY6dp9avknV
DcbSR9Hc9nqEXKDUu/jeWno1d/s0+c6ZrDv00pUZIioaVR3YE3I3z4IiH2qBczaj
oHoWucZ3S7KPR/caqsurhs5cWH/Db82bSW7TKWkweyTdvLffTtxv4itI0u0zkr2E
aRiEC/Qe8+2R+4U/Bj5XVaHstg5NErwGCsokiO2VynNn3JN1RZOU0jbdVrFZ1l0I
t3u9vWLeHvQrByFDBMfiucUrX8wSdXRNp3DNttpsvLO2LUd90qwLnsIhEoPb/zuU
xeGQn+XpmD+LKwOIySF6JlyMSvM6GRnVJrmY+2corhnzVgBV00irXlvuFxf17Ijs
kzKQfSJStjY2Xddg2TlJD1v1ZXH1gHkLv03NRWrBeRR5Q8pymXAcb9zxrBYd4mkS
9gpKpXmsxtHAKyWe+K94OP0B7v89Tmk1pqsqabsP2RsJUX3yx9whWZ7EtPqVi7fl
myqTN5TOGDbVqo6v49ZuyCl5cNWEcFC0gT8KrtqhHhz9/clJm+a9OIQy7ar7y00G
HGlXaAMzhoPs4ideYhKA9q2cBW1X8x0Z21d5lrE3fF2dfU1YzK2w7MN9vtQnAvbW
AkYECIXrzjmScs1XzfXczib428Zu87x+7ZUtNxZjB9TxrMDAv0JVark2OoDdvyvl
gtcJ/lGF3VLHjByrzPUrbz3fuVpbgQ3LyPXRJ9rrzutSDdrM4pKd+DbmhOMibq6P
cTiox9wmhPsV5ccN3vFfFBCepPEsuzF7hzzxmDYosCy/gRiunzRndMH/zce/54TL
9qawLCi4kodPPrO8P/3w2SGmZ8QO5xIRy8vvBcQxRn+TiiYbLpZXcFdCdWwpOaax
R9b1h10pjpJ1zDyqn/eqhiHv4KUFKh8jEqiRrk04YWl2xO/gXk0WAV4n2AJW4Beu
UfqWHA4OSYdgALsIw2x4IOVRJ5dckCEWWB6LsB3t0wCjOjw9tseisl8bxEZ0HeGY
YHMY1mVwAqQk5Tk9Ca4ofzvf/aDxjMdoZwpEjNHI/jh/2lYqVm2RjeVifwRQ8E4W
IOzkcGKB7RBi26WNSptE+VUlbAxDYEt8dUOFOjfUJtvzAQ9Sj9PeH9tA/C/AM7te
cFK8DAXerhqaSsygBFCgyFZVZyNEfOufFWPPC8epc7SHiUSHx9iMSvR4G3jv41wR
OJi0wbaKGx7PvYQx8BCfsz58LY+njQZLLV3YBJbzw052HYSEKUmBFEjZPQYnr1Bb
j8MYJ7VBx1UFir+d9DMvJqLfCqnOTxDDmKv4fqqg8x5D1QCY3KfeKTqkWcHs4IYo
LTKq7LXD2fxiEB7GlNlBNDe7FAW5qhZ6qzSWnfPfVnUgW5ORg/oL7G0NuEH0cNDY
anC/rP4YSFp8qJ40Aql7wG5mXPkxSlNhIm2T4it9/jj8LCBAKvdfEOv3y5pkmSER
4KiYRABI1rxGY0Wuv6TYYBsTWFimgcKYLKVT/j88swi5TvgTeCBJW/iZIV3Vizqv
p1O1Ptg7kTL2YdlEOig6l8A/bt4koFXAjTR1BdoQzeX62oMmX6CNECVkZj7mB1Z8
gEcQTi034ooBdlsE+yyO7rVXFM+U5CVYToCoXJHXIdSLO6fjwi/rxCf5xTFMi6ax
1FBgFgRSjAKbWC7DAhfMtaeS88A1uuk8pfweAiWjStNo4+QllMOPskAmHOhZ/8CS
hsnmBh7iJ6R+kFalR0XMdyntwLD/JDMq5brHZU81j+dK2BXkCd4MsXcP9h0M/OwA
vgdXDmPo4UA0r2EzD0zqruviCRqmNGjZw2VVMC/qzzj3xffL+RPkGkhiK/RyY0d4
c/Yg36K6Fg5mtPq6p3Ujigh7/E2HtmqAJWP3okVjlGCIjCvr+mU3Za8BTGwfUOVV
/cExSdwPXJjx4pKCZ8VfaG2lva2PAEYSiVZidCcXAXe+KnXIX91Lkdw7mLpQQB5m
TJ0XgOU/7uaGXrb3obnM3wEmljX3UGVElp+UJs0lHQ0CPX9Jzj2guKJS+aNpl8uU
9hosHw3tU9p8DAV2vgx7bX2mpI9jDfRxE9yoGd4NJLVqVpBP/xH1YeZCFdoVPyk6
iWe3LMn2rW/LsAi+r7jhVti8PK6V1HJkpxJ37CJdFgXcSoGe2+R8I3mUokRqAImb
Ytf0/HC4jEi8y2RghsO13WYxqsk3cRYls+Wmwr7eN2Z/scHa8cjzZsQOTgpXNcYy
YsqZCRhgqo6rmn71vHu80N/u5mUMPSUE9lIazVRIC/CHb+hNIr1CvzovUJcvyEf9
mx/+vyMeodkvxvfSE6e0OOgkoM3Bx9cyK04BDxZlfMZ7/EqZ1nDTV5Fk1aC/mu8x
tRXCf34seFIG7E08TBBbjwyxXlQTRdYJ9m0oL8Wwi6069iUMXzgNP6KHnspFWBnS
kNeQ5qfbwbG7cy3Xaf8mowVDnYgl9J4nwsYeMXPDuueuV+hoi0Ej0+xvDKJ/OeaL
ODX+0D3Pk+jC3c237/eR9iQZ5ZI6qUpfzyfNYsiIf7XgNl9mIJaoR99W4ouU9tYq
B0hIpBrxbsWZwb36SuBDjapDzvk10oEriLDEjGojNE+zpcPhBSJpXwTvobHgwJZL
6YQCbcFc/DVHpOOMF9rppBn+90tA0AN+4d+4Z0vj16JpcSpIp7+rB5V7SfUcEpnn
1mK5brkpUCFcMfn7YOLW2Zvd+nGEpCglN64a3sYbJf0be17A6W8rWGh0IvqYwcUi
5GN5qWiffZdVNrsGzeRUSh37lkNIqPjU2tGz+i/QCkwmmlUPQXqDHFAYKQe4EC7p
mx+07eSJZCSRNKbi/UaT0K2okdTnw1DtLObGwCJYQT/SRGuaI+8sJ61Z2UIRHt80
3PTw/8vnkfDNBC2JmNJ8t41+NpWlU0ePH4Lmko7frPt4KPAMKylBeouX3xaArILL
PVAOY6576YfnxqU5HoGlFNe8/3eC7GP2Tz9l4nT6U/sv+Nqmyadfvg/a6G827JYL
NiHQO4Eav99q4zxjbwMKh7N0XIgF2b5yo1oSBoUYe/vUMakBFfP62SCivVnZRUjq
gzEpIuojnXJfmcOwxe+ov8E7Kih2VdgRNeY7zmPhdmmTxb0eht4IwHfJIuGSP4oF
bysC/q0aJT/F/gho3kKlJgxwZOrSH/cjeB7yMZkkJjLgHFJOuINY/3TpTcL4bNo/
7d7T4pyefeQu/oL0+nbwoCkNKhimf6LeYh/IntAW6nRCgejfaZ2bj26W7xatWvUH
yP4ZKXHfKTTrY3d/5lDZJTBNEilXBNcZI5Uh0Qqt7A3RUoaDlADD2Yot/jPiWeJV
EvglCo5D0TCyVtQ9jSs0DR71SSnSdHxfyc/Qhhsb8/UmQ4e+NbB5FBflGOlfKsTa
q9cD7bySWaBrdV8Y+1tKimRjbXPiZQOqIkgAo6SW72Jiu+cNw2Ek9ThdOEn7PWRv
BdtMG6DPjT32Hx1NhcsbzmGBfVQdqRf1+Wz7cpyAP01y1JWI6uc/fQZj0msINykC
hjQwTZoVP3frFqk8kQG2M/MuYJmoUtBqPTR7+0aFTvehsXNjAf7qz5d6tCFmFOXP
gbt++ZGS1PJnb9589KJV7YKq4qVFhC4xN9vkuHbiNKpAL5cUVBKnYk+8ld2zR1tp
MGDjEoulcj6bov5+04OMkOeoXjviGMHGC3hCeaSmZViuc+PMscQW3//haF0+xl6P
Vx587lkWAOUUuesoRYw5pTQzkozlZWnycxGjAJpdDmhVlMxdumiap3enGeFq5fot
1In/dXsm8sqDwIRGUyEVvviw678Hqdppfs75BQ7NB8NMeriOcw3K6ueqy9ortQdd
88NjXJ5KBnnKSxorsCZrlAlXKELoCf3kRlWE+eoUvmZHUq1gfax3rY8h49xZDyBY
MQLmCqv3Lu0QeEoie9DYjaI6EnsykV4NXFQhW1O2KshjIP5xP8cFyAP8i9DgadVA
gd+dXZcsrq6Jyo/cWvsfSF6/1LYIvaIudcr5qHl6hq0ewOuSzznoOrfpSggH3ksm
xy3UJC+9rmfRM0jFIXgghse6bDYyagUAEITF99HAhqOn032xgRKwoeF58Vm7qjST
EkpV4aRa3jokiKiTsrmY0FCpnfc47nuBWRyaE3V1QWuts7EjuEs60FZkon+La64D
P4JgaAPVAVQxD9RKQUDLw3QZRj0IGfPV/yjAiGe+XS3Q18R54AKR5dUbNrFvBtzC
Nvcnx9Y35/3JWJfTNe+7YZOKWDyjJ8IzrwtrmJoWAZBwvWMoKqp5pIN6b0xRuqfP
tu2IUeUVCfTxa0vC5Lp8VoS3IcBt5rblTu2U1zdcmcjILmJvaJkJQa1X9ah+UGsN
tIDbKTIcQNFm5GyjH2HdTlBBtWd6tape6/gN70voTcfSxL6Tpu1p/L6oOTvE9HhB
nXzQ0EraE7jvU627MtErJDObJglHv+r+Cgr4oQGNYLDXv0PxSCZlHAG/Ayn7qLJ+
GfUPP2L7IsRaFAKOagP1z5+GlZUwf8/ejWnt8VYh+4z5zMCdfN3QKGWEfM9uHOX5
RiQfWtpWx5+IoWhP0zuu6vo6gYt7kDY7Am8bph1Uk0mKQWudQHFr6/Fq9XF9Y/8G
q/EvKemxx5K2n4gDyFkUVDBHLKg3k0MrDBY292nTyUELtoJWBO3UkrPAQxXvsYVP
8xL/ua0FgxK5Mpq5vwA1Zm6J4l385QlaVs1dqiXSjqxEh0xpoV99TFdFjuGW4jQW
W+qe4hkXV1e3SntXuvtjYs4br9g7hBIw9MWlgb9e08l6jwcZZWvwETRjHlBv9t4b
7bORXS/eqqNHxKAiC6A04sHthbhJ3OPVSJNb16hnrKCrEhBYRxIIcxQc5eXgUjrf
0evWrINgKd0zXE0RNkRYO/mir8xUBE3EaMA7aqQaIU2kt7fWYx6AP0THE1Z3SSzK
NIMKoBCMPQgTaK1av2m6O9J/E/afwYDPS/PWD+PMiKSJ7XxTimBI2RGg71DPN3t7
k1GPBbKDAByssoQacTqbTWXyo+s/M8IgAzqsRcWssVzjSAOnK6JUhOzx+RrnyRw9
8XUEF76LHH9Ef5Nmh7INS3bnyJGO45TcYK8A7Gxl8nNHPOFIlty23yMoxLBRhDVa
zVEvhPQc3PEdcRe9JzwfbX/DO8zj2w2Qo7fVp5h5BHHC1bfEoGu40pwbPDOqUl5F
6pqVUfyfsSQa/c07lYlWGArll0w2aHNQe6Kbj7ey9MWLo63oAWzUCrtIYjR0b9Hz
oWVo30DO2OoHYnwA7EXyVVW/u+RHl683062MZ4OOoSs3s73tm/KAwc/j5V4ZxgvX
rzUacNpYJwir21aS3fFEbSrmQmIBgmyLx6yOiW85BK0AVElEzA+k3/MDGkYQSqKO
O3+YmX4zb3N1UqVfSR7ZQZVo1YOGJpv4nk2b4zMy9qmmR2aAukDbcl6m6zcqkgf9
5Mk4Tw1xHxweOBu6qic6by9LGuCPi1fBSJhykIzmp1YlT9KVAQF+4gLh9Ro/lIg5
drbLaFtzbJUI0WQ8aWKKgvqbiq7+hzhuqmV1Y5jgxntcjKO7/wrRUFyooxKLQIu1
TbQNhPGhyZpI4LVsnoOLFQXkBW4HhFc+YIvtjvh0qKBfCMZ14pE7T8Y6TNla5E27
TVDAzwQZTCx23uyv8EehrA+nLEVp0rOADn/Ue/myMdNlPm8rPFaDcq3Rv1m7bTlK
I85uKKZ5h090pIF2DIgO/5GEVaSslzXLTHh22URnMktzlDw7hrcFrGJo0TSUnHqR
9fFGRkia/AcelUjO0OZUwxEo+41FgfB5Jij5oJM0bleOCrAWFT0Wt+NKaIsk/iUQ
wUevZtF4KvTlXfQacG3cx566uj8kp7uSIbgTQoD0dJXGaGGVh035R75KjdHYGDed
nzFJTqjGahr3DMXElvN9SF/S1Y4xRjUFbLoZ9OlgrJxEfwqqgyMC/sJQ0tGo2FhW
sDnKhxy+wV53U8KKIs5Tv2255hLZK4tJJfcCMjAnykGJYJgSbQOQdZ/No8/lDfBQ
QhuJHmwfY64yRWk6DwVXgTAQjaO0P5lVsClTWBUvLFrhMkZJIo2KoEyqmvVG29o7
ecaJWBhAU3vrD55Q8vBSQ2acnFXoPHFglIyBG04r/0NT8NuqjtsF5HLZdVx3Pawx
lNhkTSjtbq+L36URpz9lSEtkw2WOmIRFld7X6X8lyDiq1DhM6+H3hmW/9fFPf8oe
qc2AGJaHl7jJCs0wSnl99IY8LwAS3Ijn6PVfJ8GJyInrCv1X5K8P4RKK/IPSE3Yw
scbFRff/5Cn/eRvHZ/rsR190sMSbDO0vSMZuKsK7ssX+CvbtpvWSNK3AYbLiDc85
YGfGeAaTzoockSTPGEPgFRnzWLm1LYJnTQKjKsczvVRm+7kP/q7U2cUQO1UbEmpC
SkxNnZiSK0Da6QAyn7ImBTZ/tkBtBJD5CEmCQvoEXK0PULrqalph8LtdalG/zrWg
WzwMnqjJPc8dmKOFv9SUj6+apO/Ddy1zO2BcLtzFOcrfaSPGQTuyjz5mk3bw0UPB
LOd7RvNX1/33ppQebMW4oXHa3S34gq9RYr16GD++UU22m1+6o+nPtVqNOlyH927b
yCqONd4xWaKL8bxk3RG8vxnYA4IJ0QTOa3MNsOJ5BJ4/WOafGNZSWisR/dfN1uUQ
wDf0DnonuqLdHrP2eXPHxduxsQY2k4Vi3wiJrQY5WNkWqclKUL7qBgew/bawtw0M
K3AajzLLxBDPww/BzNLyL7zyIcHgYEDjfw4z3TYnGniWDtMx77aYKb1uDN4SIJ92
y1c87Bt8pn3BZVfqrP4/PKJRrHI59kjQuFS6hrd+tKnHkp6Zldh3USRkqEWEmu2q
MqojYwqhvCCnguuaUm9s2ecKPOfLViiM/3Cp/R0ruwiITw87/NwrPm52Zd0e/yld
F08MFtkwjGLHxfFk0QjFbqUYBDn3te3/M1Fcj1BLR237NuZBrFIAqkV77g34dri7
RyNvxoF0M6fTmwbdWmIRQI+gKgbyQ6TdMlZ3osAF7yYZqXGown9x73PSj2P3k0bj
QOiInPf8no3L2mOl9vULLGXeqbNuOawQlyFWjAKplTZaJiuGbcSUKoaQ+6r/RVmN
l8KxTUG8OBG+A17e832YXfwW87Io713Wab8fGOgynW+h2d8t7c/x0ykU1/rLvnLZ
Jpo/bxChrNsqPiMv+8aG84RJxlLsNWZPwtGMqXM/UcNP0FBdtF39O7uUt/e6s3Vy
+Bv8Vz4OM9wx0S5OMgsIFNfjC0mivIJJi1vDJddknCpR8kWLEM0m7TVUaiJ9PPgN
SZKXu7wL5OEJXWUjIKTu/hskUYhFabrjNXRT6hGXdAm09pO+Y2cPKwKKGE0NqGVX
+IISi6dsVrVUuOisHuFMho04+/2/Yt11kSpZyB4GvdL2CudFqkSzJc+rhULK7m24
WyQgFfus6PFdtH41irg9fJ52Ya8mdwUqrznEkaqSl7fNaAtMpVl/Cl3OttuRu1Ow
FehSEe/lm6GfbM1YZfBoWTt2wCin1QgXKfbnX2041+7XyEiM3sNPwo5mCv9ko9q2
XjJ3WpyAL1+HI4OCm8GRFW6vLjTwzfCAu0LllRwFMil5OyurioVJcwwr3LtBoqZs
mJTuJXI4SIOj6ThbtJ4h1hI54yPvH7BjtmPNFs6IpUdSEAHjzQNoQ28QL+QvaiEN
gOUAUf5VUhub4Pet/yD5o6tcyoAz8QbhmEtfTA2kih0MyBt+C2fT+WhkDvCTQaNV
6MTZhNm/rz1mOoVwEIdmNUp83pDlpEZU4qoWMVzLwjEc8XH8jGUdoys1eL4r1Qe5
0kk3GanTEu2PZIm101mrI8oC2RdHokSTrjWDk9S7fDJsZnohrT7LpxLsley3dQ+L
c90/misTTX8DiGPOqwnOrojTmFj14wM/sjrDoTX+pNGu6MolvIB7rjTpcqj84GMx
CaAwsk64IUYbJYWCcZAPyfSNV4uumnwg9nIWVqejq7IXukKDmnIGQzbbZhACVdHS
MNWTy0KII1eDt7qYgsrWWX+efGhmba47CoFPP4Gb8XlFBrFbMavnmpPs3wHrJBr7
b+Pe7hme34jzO4bDxgGsGeWhq/Pug+ARC9aiy8L778jjc1YfGldbSOdANBRCB65D
UkTj1eNuqUq+fYy5Z8ojZ0WC4b5m39vgmrwiWrONNmZJ7yyvSjHKGAZiL+Awr8Xi
ZDSIaqWGP+QmNRDrh4QF9ysWIGGsDPYh3NcLy/wHF6dELbQG/t7VZSEm5ZHvpF5e
YxKWinHxA4Tyd+6ZR/ktT26jEyE2O/EcAGeVOg1Xsy3HMf019BcrDrC9YMUyici4
D3OUeatdCzPm0zcU7SB9nDd8VeOjbr6oMIfTQwW3Hx5QBr8rdJEi/NxR3xHXlBGj
fPnU0f4Lf/C0Bf6N0+9MXvCss6W4kBOX9Mu4ygrpA/v+ylcgHwQa+krCh5LVGhuP
c4DutkvZyXy39ZuG/QfB0hUtW6CTrB8Y8pFFpWDyv8qSlMXcyiKN9EdUnJ2UCoFY
t3aHh2457IZKDYTBLDuqlWHRjyxdZW9et1qvVNWzuwymdCEvmpYDxWGfTb59FqXg
HbyvyYgh8q513P8TNAqHn28yjTxQHX3qfVKKbAHDfeezHGmZZdlmMKsqq1CkBqgA
Z2xOGWoMzmqgrAjsTyG414KAJT6KoqZRVA6sp214qTv5r1t0Yp38Z5DiRuDTpfvm
hvQFHBro1glOeyjMFtaP8KA+Ea78hAlE0RBbt8vEwzQ/N4y5t+I5tgKnGJemevRh
4XUHRti28YsnDscsuQof4j4gYpp3qioFPtqivbkP7mfNNu96IEZmP64nsWasXARb
TRg3XaFTWL+n/gEmrhKEsLnoU1KtNBzg5mzxkLadoXfLZe8OZb756RAKu6iOYP50
UYvgqPImDh/DqiOLqD2BjGjJK/D+H07KtVGFuOszfWJm212AR+YqI6W8e7OIRMSV
pkLAVS5fcn9Uj0yxytl61x+tlCpvvbVxMuUgeweIHbdQmHEq1nTxVDd7qjGS6wLr
1PspFxElvikVLtYQWLDOPjzj4a1A8ysAhFR30Wn8GxASKfXDHJ2KnwYGwPHYLYRu
HZKR6qBcyYxxGTpeYxGFQtJkhHkjJInGXObmSFgWjlQOGGCgLF0yQMay4Z6QVpSC
gVlyCAjRuLq/e6mwzqs8pKa6OXSmUHxqwU4t1lsmf8eLZBaydoDYuz5FuL6Sm3gy
Z5E+/4ETxsSOwIwq7aHHdqa0vUapx1vM4ik6oLw3GiJghpFrVIxeAjsnlaOAI8Ek
LIz5WvxaJ205O8VLu3D7Jiy/nC8/WpPmIIvRBvfkfG3jp8f5rBMJg8F/6sSPlDzW
jzT9IXBOZybSXKifaf85vT+Vxv8qrtYorNWXxMZ4rcGET+GL+rU+Cr2aaPR1xbMR
KIvtNa2T1GHj2TtZgBjueNTLOWuT0QR3kuKW/oUyod5f3s1Y7x0ZHECXH9qh2XBi
Jn1HjhXPIjKxktD5aCsWCe7NXIdXeIGBTl67bHsHIi+h7WG3kOH3Ip3wV8X+cb6/
eL/o+3OfJHsdficCnwxaGOamhKn2Yp9KQLAth+ENUf4gBjxq0nftMvxWHiBHXGOA
AYqlq041XlOx2C0LxLpkxuvMdyKBYORKhv0mXWdyUfox0Ncls+ththdaeHQTC3Ae
H2nA5kTx+rISKAEGIipi8UWNDLIdMVCN6nePjkXVVtMjkBDL6iNUzlBqU9OMDQQo
/rwXujHqvH11X3bx6yWpldxCBZJnCTtEdQLigDBKWRlmZkjESnw2y3u8lpPNd7sx
I26iBHEJ918y68f0kg5kB8gPAX5HgXmp0z2HH2KvXWK+Zi0qSRs2wpka/rr+DfSv
OsbplJ6fe5R2gYcLwnzIgCyxi+XPTGM/ujEm7Z4RwlQz+q6TgziQXrw11OvsHS9f
YtEWYJ69kVzOZ1JDk4TEQkpHAdOlqAFys3/MLFG1hIc8p/wsSEGFtD9tFtzHqP9l
zFqa1nbEsB7uZ7+wHoLTFofaTSE5fBxOkGDWw1bXuURYSkv5p+qfVHsVqZJUepdg
RTOErt9HA5P8DW1dQJ48NMkb/f2pihXj3t3XXpgwqGglTzDP2rCepsFN3YYq5/iV
I1ZJyGRCnVnO1FdjWUgSWvpZ0LDvIGWijUKY7uiI8tiMs9U0VFUa0AYOJDt/TLmv
YYoycTAiho7sf/Q+dz29/X0Ci7sV4A3YLXVG1z7nF3rSSUEfi++bSK9zRSolFtjx
8pk2uUuob2faR2MzK5C4TK7NOCbPidOo4/pQQ1PjvrHa68E24WjuCYlxzHgY2DH2
D2xstSjgs+Tehz3OPFBBKQ5PDjs3TDrt6EucLWaExX5n+KXTtuQwRFgCbS0wGSUD
0UJIr3hkzdasP0FhZTXpe1DnM2q3u3BqojaYLhoCaRhSlDOnYJLzPuKi91/f16tQ
qM1x+gCsn1vVklHLlTy+TAP/EZwewTF9RiFpTolrIWIE/IsXAqBNk1u4NDCGdb7r
sO2Ogioq4WBQeianCRLg1tRgBXaQCNa1VmsG/6aYggqdhW3sgbPL+VxjADfIEWoY
pWuI3UmaUVyzqByn7kvqY9j5XHN1oiqDgKtarcqcKKV07tjstqF2i8zqtEgG0Sbt
RvQaowzbDCX2Tu7au4pc85qGv28+dgZphryK4K1CqOJ6TZzl9rS6bZGSXVVqXSZn
YpnR5yJW9vBMn5DsTr0H5HhqOc4yiV8r6U/1v58r1X8V+5OBXkyWHvJT/9972Heh
NZNCjfqYgSCn4lznKLVkgbFqf/WLByljNl7R/8EsR7o433hus5+99ChN9sg57Oky
kIqSTUdImpRdreh3sLWkaOxKPieAJAbInpn7wiz/PqZJCNLRSisT2n441AQRtSUQ
mC1d8xoc5IaTG7BI+39RDtuDu3eTpAsmmMhY9Gl6Dq2fpPUZVrEHA9Kyq1udCVDN
oBRNDqgKtkF9m/HvqIA95+bO5e63Fs8ltBV5wGO2ly0Vu9LQJXt8buNrQeF6LaI/
kvlsnvnQ2Ye0/Ot9QQxGlbpYx6HSNSUrUGn5csZVt8SCWVH7ncfMVx/Vj80u1vPU
qcHyi66GAIRp0t0FwcoWP3BvXf1DAtumOqS5zjE0hhWg852hJXAj2P6AexzuQltJ
vIY3KFTQGwo2CIVZkXqYmgF5FtSscaFymgiE8wlL9cJrw4xU+HBMp6ULGLjN4DBD
d44LVuI+TAnk18iAbB8S7/6SkO0zSa+9Xx+IZ8jFAufzWlZl8bvSaEoIcaRaLoTV
jd0T1pD73V5IN93Ony6hD0Twjej40L28PlFbNqkoV/WT9UlgUYe5hKvAUq3UDLwI
UbBL+J8XMVhGWDnZLdsAuUiVUWmqx0beKjcuUmRwmxtJGn+GdmKc6ufi6ETs9bI1
lSA2DycJa7+zsuspzPo4SQ4Qywb/0t9zijoUhKh3hGKQVN0WXYYfD41aB5tM4jo7
esP5aSYFz9MjU9J3MYe85tdg8fJOZFO1yUMSuLDchPFKlbiPETnBmLqBeJf/Xrz4
X3HvbshFP+G++orpQ7UGusM8n6jMjaw1WqwMvCxDdB9yRprbUpSIiIq9IHKjYEWh
27vaaZlfZIDsg9OfblSYWnsilARL+k3zqNGZ+WuhhIfnEiSsd6dhCvTVkgLwmTLd
q0dL8Vjo3K9bYqrUDVTSYtbzJq92j6pc35xJsHgGzDUtcXLzTqj8/ZAJTxjebjgm
1bQTFeiDuqLz5DMNHQJxq0AzuKQdfRnzI7JMibG+myW5zWbh6dI81ytTzkye899a
qFHzZrt2Fn48to8NaxWzwz3ZDDs4i/4heTEcAhePl1ANJ+8zFJDSl2XuqAtNYrgi
owc4v4n13y1oawVWJ0+Dq4YFMYpKPgFBWRCyt6EoNsvG7cRMNPbk+WqbrSbdEe/F
pd586XZJamJjGQia4ti9i/mDK6IaiSNs1JIKGqP0FxjtBojFJunrVsPjoaRcuqQR
ZzAFIm+THbFJ0gXIqcTyuV9Y7vLDgKwRFcM5OPvl5obWc11C7vp1oPfeszz3D8zN
ChNM2vcy4L+dwTBt6ECGnqZZ4mh/lGLXtFen6G0SV7HLDvlpmGKQjdg0tKspPunj
RJi6EsqBv5K8dRmBbAZNYqYW7AaZ218lvjB+G2/gC2mAJuclzTaIfP63EP/nBEvb
/I97BsoYRJGf6Pyw4SuqH4QfJuu5DYfUJnTZynA/Rgwfaa54O7xrSNMdYQL96NIw
fW1ZQxTNLcH1wVW3+03hyvtEsapQZFD0q0+mkY1ho566hoSXrW2bPDps6duMiQf5
XBF3l34HsptQHCL4d06Ec8tGBK82lS2A1E2JguzKsBpg2wkqkmU7oCI/l/uPjpP5
61IECbqeQRMpS4bU3xfG9s5UiMtSrqS7O1dPFspB6YSlg3ijVZKsooWGEbj6Mgx/
cQ5+NTa3mBNn+m9wtxtkVRmUUxgK/CD8Z3j/1tzgP5ewHjqZJYDg+zt0Nsc2et4p
XuYW4/O0TAyZHShefZk4eI//5VuJlqm1v+Vm7mcdelaDak8axwrKc63iw+uqY2T/
2KxMpAYgwqWae39nYbs4AvLA9cP9ZSSsjzJJau8wyvhukl5KDvipGojl8k+idW9x
x7hJWfe1TAtNPnunvtS/xsaR04JzkbtNzlKS7p0pb7tCwisncwZFgXFBHvVJc5Ig
cz3k3rR+UrPilqItXipCW30heHexlJlVU/5ChraJ2JQm+MJ02Jft3uiD3222wCxa
QTxB8G5SYtKlA/WOdKJ3PCGgdcBmCofO9EBFC33puxFll2jHEEctGyEniwWcRDEL
Jn1MtzeUcK6cb+eWoYBG84BsZE0hE2ig+AzCB/r04nF6nX5rqkvvyadTnJXIbcKB
/iiyssCZdQ4n3fM+xysVkWrt4J4L/8CiGCp6W1ME7YQmUCYC0owie3Ya76NH7qOH
rb/ZRBoVbQ05OM1k72ZNsCiIHmskxvD4KZh0TU1oE7qAw61my80yyv2xHQjUzgY5
gjlrmadI69BR3xTUV1BiZXVX4hAB6CbmQM4geJeY0UC99jfqARC8cV/lOjDTVEHc
5Iq9nM0BE9j1X53sM34/Q8Ehxgb15XST4KQNlpq6Z174tgFFoW+94cxwE56AUcOJ
5fNY5ybuu60UBs1PO7M+ziyplOMVLbEvxHG+Yx8wVHDLng/AKgx0Ls+9jutStLg5
3gjBB5i7h3yvZzD6EYSOXygRBeDMAtT1mwj8o4xhuZQ=
`pragma protect end_protected

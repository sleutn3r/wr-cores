// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qVzWBUPYuKrfEgFbB5fDLrqO8wbpEvkuZx2kRiLYDYUtVI6OgwcamTLWdcaj202S
n/LkKYziXbB0RYCoE7M4X6c6dnHoJntOloq2vl5NRtuLU/7d2y3U69lSnbKh/uIp
uAnSzok014/9uLgZWDPQABiWZjaFe01R+n+Gpvi7iTg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2304)
bYIigY7Vg/I6P0n2HXnhnzLmbUeY/FRUfbmOKKpSumcFjozh2KhnL663sZx++Srn
RAX77DKjA1xRTXt2Zh23jrJWTjE1OMEy/+NNVMXlIq66R9ZfAFgelG+4cEU/nhfY
9fUsmPNfVATFhPOZSGW6r+AT12wlFEOzmAQzuI4dJIf93WyTr/dUxuCddh2OcODn
0MhaRGdAOaT7Xr2vfG9b1cfBSavZPUr1mubW0WjckEoGW6nOror/cLRawpmIUaBZ
wpCWIK5LmN09jbf+TqoYz1sHExGirFNcsruKA3NAHDa7tRWxafXjlJ4LxJ0gDDzd
bZfemsiMR5nQa85NPQZdqwckDbLmLNzckz+NlyuWCwiQGier8whfvmBjRfe++kTB
aJuxfilz59u7yLsCJatWSWK+UK90y0Ygts4PS46MwgIRlVf7IQmZAJcM0khoWGC0
XDccaFjg1NhMpYLS2mtbSw6PvS7l6VFRcyolSD+YTfO8DZv+4tFTBybvp6jzkpvw
LyFVMoPBXZbsz+JQPVW7UwVDAT5OpHTyVHL1BZPSGw3ZPyGxAv2+gCyb/U06PvqO
TdR7bfcu7Lu0azLIy/MGjjxr8jsDX2KFCRM4z60sokaMbjCjq42OggeQspFAzy2g
4eq0oMRsJlc7etrLgHnExgQtW+lENt/5j5+nxOsfYa+5MC08AS5CBvmiuEeIL1fQ
gJ09oNj/bw/lduT8+EJN01zjIcz0gJU9cdHVKlDiQJPfS9XZwAGnHpE9P2vCcg7j
hBWvCRy05Moc7uaJVyhRufsTLZhin/L/VaoqcvL7KPel/0GV6zHUV32EMdWDz/n+
i8DOJXnF/6dxavm63bCvJo3Jt6NVJUNYRNgLnyQV0hXIE8JEQuNGXPR3AOfMTP5E
pAQV+WwC9KpW0ehJFwibYJ7BrMRlvPws3+UtEpJRxrWh3NiY6eVAagBkGe6KUoLv
wL2ZpvFkp/u4a7Ijnsvyy6cnxlo5dUYZlIMLFT3W5QiZn81B6WQGutKboMWMfb9M
Ex9TDiuYQwNRbwGQOQbiZLZspw1dUNTabj1v7ngYbLW8aU9lWthJIttCLFRnY4c3
NWkkBdhZyiCZ5lStZJSjmBZKJ80OSPCURXnYfTgHxZwP6yFq8+anomSrmwrJKIYa
ITZTWKJqJPTk/8OG1U9tbt5IyATx4EzhkzEQEPphgtyVLXoQoJP7Ko3YSKbn5pYK
1yVxfWbPX+M1FGLnzoEAE/yxN2mecPODlnmwSbJn7YZU6AbeZyjaUYE+daelOrtG
AFqeCPbBKe0wMYwuiuRCmdb72EMUQDYfAUMr7dw6aW0aA8Ww/zsNmtdF452mFUwc
67HAvRZlrdJnnSlfbi4sL4QB9qqMAx6AH6CCbXN0CEaB7DX51PVOwAXRCIRP28we
YlHGBSTTun9VrxtHntRDnDbH90XKCae3CfF5rdgrc23zEnAsyAg/1l/TumqXPmAL
nomKWY1gsqBzVRSlyV5vuvtblySFml853hoQgQtdPoMQoMuQtkdxtK+DKlDRimKX
h13MHEgoWyhhBPxOndqTfQ2JroUYyCFt90gxAwQ6ilZO993LAjMiiZwzGWoV2y7T
gBe4AgV+7jTZ9DhX+Es0mOe31lt6OwvQGhJvIJ2F6cmKxNSuPvz7oQ+mBLTEYmQM
8atEhsGssQ73QY5R95kQUyuVoun82n4Da3155cElSASb4nkU/oJsGUWwtYJ8kzUf
eFvp7F9LvqosyHiUFvyVssUy6toU91QZbfUUGCSgjy5DHggdRvnEEJ+T4WYxH0cF
NuWni/xUn9tErhYyGBKTUprgj6VMosflQuzh1i+8ucOapFvZcZIjPRSfRY3DaYq8
hNBmvZlnMORn4ASFVzN3e/0hPTjNSqz8g+WGKrnSSSi6npvN1D1q/CNS8lUZmGYo
jrFDa/O0qdu93ET8YSp5feJPpCdGCH1rriIYmH/YesMS1oSO4qSDeHbNVAK0otHZ
rZ0xoSnu/K02jovYbnMtyqErrW4V4RHDfqVZYp2QOEwBM9Tzp+Xnu56lmjfBCd0k
6bm1pUy4zbkgKWMa+gStHN3CsZzhgLrer6DJP/EOPwP5lyOMpSz1amaajp1gPui1
5sE1ErRTtAI6D06D182A3zOWqDepeX06tZQEX8kILHgsHtx9BNtcC6fm5D9kHUkj
jhg0ytsEkTXbxGtL7behisOq8JdSlfcKgFbspZh6zaJQEy3B6id0kn/M4rJwvZJN
LmX5W2wqb4TBIXJftbNu9vhOiglasTFOvnYSjl0XOhwcb1DPRWK+1sRe1Y2Ffmyc
dVP/U+bcXXXbHln1yinnp+WxjPV+cYU9vuE9C/b5idr1hbg3UBOG/7NLC2njTuXF
1FXoD3iD9iENEwYuDI+IbwelHgQpavqSkdehXiQpmmt61ePDx/8kSlIemx0ej+Z9
SiZFufG6b1KRnLe9XPLe4kcYyRaRYg1pXpMhCZ/1qTm3x/AUbLPUm46LuP7YQTup
6C/LLVqa9gK03qIdbN/ptqR5h7RE5omyjlZ8Z7FfVxSN7pvoU4WYBsFMEsywgu+r
7wN/ujgkxz6D69PtGKKpKXiNhCayfaYXSDOq3OAZPetE4PH6JAhxz6N8vv3uJGcO
w9PoLRfub+lqf/DmRrWDM1hGFAF+3E+RqZBCE56d/P8tiRKm2FygXqEXBDwQ0Vun
RNvde2EsnsFCfD3DV/5q8TRx+i1P9u7n3w4gaWDxDfaOmfTHXnXoOG4MIpDaNV++
ISSYkXzVICuILohqp6GWdRNy2S52ONbixxrgvBrmIsxc35mYvkyqC9caU6vrsJQ1
+5zqZj8ra3tz+bJVYgpYWt+mLpMP/1X+AJOqGOyi9KzG0w+Q0rlV5glQwwjbzSnu
hrvAM4tsda+VEZGeCw68MfKhicI28caFwfeckP6osBHdFr6gVGSa6VlRJaEkExib
s77V6nzOiEA/TCg4XsoRLc5cKd6kVVbV3agC9RA8pXgMXNstAmeqdIJe2i76meHu
hZda/thAl8x8kn6Q4yptQg5Br0yCBOXmxJkkn0Ofj0osaO6SBhF3p975/8S3DEuu
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eV2M8A4bQFwTTed3EPcBaINWXp+XHtnfH7jjST3k6pYA8N3GWpMooHqUE9PUpwar
8RLRuYwXyY7bsnLXbbySpQuiovhznH5C5u/ZX3g1QoQLZmhUVXQffQ43Gf6AfCic
SknwZpJaoCviw4vHYYhy3n+mQWoQ30+9IQ7jNMbX7uM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 123920)
xguECp3u5rWObdnu1JBGGuGfIjgEZoULILp/3wZvYvbLG0z6ANelLxpCfWVuMNle
S6e7NDMiPAZkuiLJShOn8xZeMntTSq3vnOwLFclC/NidSW0IEztYItR9bxUjEcuT
G9Wmj8eXx0BkgxYI3O/hpXHubkHczPT03YlpiUJl/UlEMkSKRZspudlBwG1FLrQB
TdlmveVT2+/qEz/MZkn3nCvJfECJbAmNZWKpz1j+ZCLg0Faa34+EW2EKG6LfpSaH
BIm9GqFwhb3kpL9fQ9npNqlRaEVXIm556/ZoD75NhTbX+IYPOBosmE0txbyzUp9L
bR10Wx+svYEKze/NklD1TLalPRvJGIJJTu7CqHGJL3PBiWGZmna3Kd8mqdMe+KTl
MWgANAISA5NyVuf7xbGPOJqUY400KqsCgvd3nOtjiUBC1U4pbtAGx5WeMWf7qQ7x
dSoCKwQXh46VzY/Dg1LaWMJw2B21QRxzvZN9dX0k1Iws7FMTv81YKppX64Uee0nG
QGxwaOACqqDzLK9GJkDFWsYyJbT3wXVru3OgQDQoZv8hzrI5Hlj9GG877Xy1siJL
palVGkXFHJge+geofk6fh/W1mh/EeVH/buiOC891NojXTmC3c36vInlAi1bPngQz
UKGg9G4lqcgryjgFV43Li6xOCLI/ok2Oq+3tS1bq0Giceh7AJ8dee91Bt9EOc25U
jNDVrmzgS8AVZV+E+3j21tymIhEL686n42gqAEBhGSrF3U5CISc3DUdfyJn9j3a1
aGuKotpUOfbiYwH9GiKwDY6SI741R0rO9h8LGXD175ET6H/zvFL9Rw1kEWVwBqEx
yXTYJ2+BVpd20+4mdC4VEZzrpp92iaWAGTJ/oI4maT4jyG0WK8p2v3Kcg5TKYjiz
Mk8jyCIU4xNCST/vhzSD6Tzd4TJdbQXGKy+QKpcYXcov6WdsrU6JSB3JxKxonEg1
ejm3/az8cHbh12rLfqki79PtPGgcwvYgd6IWrrtLh0tqSARpBA1zsltoq5QkEK5H
KoZFzNMLfIx7DOdgcAj3lyvvHyfEBV1FAUaVzCS/XhokGoP+QXB8kqUrjLT4Xhi/
is75Qux2WZh7Z0Z77cuKHxbrJNxONN+JJa4vls1BFqSHa8HHv07kmiNQNTxErRkP
xZjYV6Pu5gcwVaXKrBy2m7kkNTxiKbtN1lcU55ntz/z72tA98UrAB7kOIIR7mI7o
+RWn2ADtaka9vw7/+FsFrwnoCPuUO0fulj12QpafDDzI/YjetCiK/biPEpLbdvm2
8/M82oJerHG/katJ7CqIPEDDcQI0yNs+ntdNA3/7eIrNpqhHgmMrDFxS48z4Jz5O
MuEWkfXFF9SfxFKujxrmx5n04VyEuoJ/ce5Lhj1Xxr5UvZH6iElpvrlEtg+v+pZp
qv8vUyvZ8yi+wSbUT1rJUs20Pmf03ykrH6PG3d0c5ZWYk+uPr6v2pQOC65t/MXkT
kB8B7Hul7bM21CMYBlebwzj/fWi47m1y6k7j/BLY77Ftm5qVSQYsQHK/KWO5cc4p
JCrRl7dB4aIXBDeCOMIVTsgW9wFoQeL6wsbUPmHlHbrcyBWiwHDHj58xj5DByJNc
KsCqYujvH2bDCwcCiVhba4hf48b2OJNg+47CMa2unV5KT1eni8evWf1SxE5JtzuR
/dIB89Ia8qWgR3Q1yAT416NXkghQh8vCQ1Pzfx0Fb7PyFk9w5afFhwRH3iyWWmuQ
DG1tGgTIa+IYjicVB2yoB8wfIZQdEalvyDbEPMKdTfipdx7zvfQHR9vMQ5eJ2UUW
g+7w4vXW9HvDZ8xe4pFGWix9jREEG+VAkQScfOeb+/v/F8sRhWoY5mZDdrNV156p
VqkASWQi65mtCQNCNF06S6ls+ebQo6Q2wOsEAD4Z25z+uv8boWtPBYtIKmhBvKLA
PRhn8l1PPm9zJ1dEYC5VlnX6ulsE0fq5X/wCm8ja5rZhDCFSKhUwTZK+Ipv1Hx5h
ZdU2sI3IDtmiDI9HhYlqVaE2wDfPkTepAv4U9r22c1kacPP6UyP2PUFMV6ngyIA7
v8GmiWQyLEgx9TDlqGgU5pMY0d7RoP8WzEDNtrKNuJHO8hQG62XidwRIOz8NZ4LP
jWDfudCmnmH/iCX86f7NVeIQhGNM5zli4xyqLqKntcDzld7g35sKW19G9LZY6Dp8
6Hq5sqHSXSaH/l5gN+cDM6oOd5jqugeFL19D8lfmJK4W6lTAgv560cXbkRCSIPX4
aHn4OkRv2GOk1Pa7lsJVbq8AxE9+fQMo9+GaS7HS6M6FSKxoWStKWdFKrVLMkx41
6+6VKqyFNMKMbg/IXqyfJ5BQvogb+EYrF+XwnvEStnY1qjtYAXxi8cVjZS2OyFt3
QLUEx7GYe6up2tFgL600t6mt2XB4ohjTBw14GVE9yncWQt6O6Yb3krdzmOTkiju5
5l5witXrq1Vb1txEg4q22622gJavbs3rzGklAA55b9wO/ijUi8n1/eujgRd4UKHF
Fe1NJ+dLgjqbso0xijyxEsTXyachLMPiznwwU16z9jcvDis+adJN+j5HG+eyfoK5
nAkkzN1+tTA85JheCDtm4QGyaJ8NADh/nOoEwgKrKjFARPXbD+Rkj/VFUXQ9zDFn
JW+Xx7goeTOxGR0LtxzH8BJipbSU55qErDp1EvuygXRQ+WDJO4EaT9Sa90QbEHIZ
YQ+QaTPI0RIbZ/7sb93hT2hjF3gIzdR5fN8srSKly+uth4SVH1tTkOVTZO87n02M
RnZMrmnTp7ZAJacEt9lXs0A/yyUqDF94WiZ0N+ZYOvBXfiV4Zz2mwhH/6o6NbYq6
nj5vj6fygdKinZaLMRVj/ppKhSC+I3hg1pLtu16WOLxp3H+Zspvp8HeIA4qqRt05
llNuo2K7xptQAg6sSicKfpW4Z9ed5P2gXH+6jtR1xRvU3NKNmWGTRQ0OWMYMmssn
hBtB4NjkUUuMjg7VUtcvSXXQNFhOhkrJvRGl0kNSyFOAibze76m7nFl/tvCMafnY
JZT4N0mKtnBtcQ0Kse9fvuDV3xJ401pucXdQWg8K9aDq4sF8SDeMrfuNGRfVkpaM
u/o6LLkUTBohuB0DetpVwfjg9C8BMVZwDjpujtlr2BSz3q+27DDZG+Q4JDKYHYDI
+XjfOisn9Vnc/IXqiMZFZtWVVkZr0e8TG5l8dJ5UJTaHr+14R/QcPNxKs15A+8iE
/d9wZjib08mFIx0FMdDda5qQ62OKxboclE/T6s6MjhlOGfBbhrHQQZnKOkzWGNp1
CvAd4Fg0hO1t0dsodMyLJzGAr5RPRc3zmgTNjGPSBue4VVbPZRJ6LQM8dijO9BDj
hfU3qJF2M3SuaffQBcQzUO4mBTNoUYQe79Wq3L7cq11iIwAjmHX8BK2Av4WbebYt
gGqLedMb6VMYrppDYkIPqFUg5FdBNsi24XeD1hlkXEHCxJ0yf3XCbSWU2f6owAbe
Z9qtZtIPjrdtWD/in6pq7WEzzqgsc/U7w5TISNmKGMa9LleyDv3n9JJh/lVi9T7V
O15GtsQvDl9ophGk76rVqzlMAFhUoBTbfw+/fGn95yHGf7JNmN6fUKlr+ULjVm7+
oOuxmHJRJX/TzXredxIrkUUU7cAJxV36QbE94VrVjm9TDCyq2H8IKkw+GHLc/15/
7fimc39md7WEcj1AU9mOhoOaz9KVOVDDQADxoiBqXiUUsNItiAmxYQdMcXbOeaGi
vJB8OfMdc0ee+6FZOvyW5q428h2ETwDBiuzG/h0fgU9O5QCjDVS0fmfYt4zNfjx4
6/c/mUTJz7NO2jlOvf+x0ytAwomXC/itjAuNhEXXIhfORb7sBolyE7aop6rxe0HM
4fQ5A1TqCyUuSLyA96Yj9JUZeWzHur4+s18eRz1pwalfnS+MygISUzkEpfLiOW/z
82pW3h5WvzJ8AY8i1sI83Ggg+4qj3yh6ONkQJXFPYOAivsLq0f8vgeRXW61plrYI
bewe7Y2xbTRb6wIycB3e6/diVNM+jVlYWmg8uX/GFhzinhQujvjQo6IIGnHuixhc
ICQdj0oM8Qqoh2VdxH1P2h6hUe+O/aanC9LEZIW45l0XxmueLtNRw4j1FR1O4dUj
j9dDR8h9xv2SJ5VT2K+/vg2uKshYvq6Q+0RcsftPmpfn78ipkL0kBJYlJcYHIkSD
BFv7KQNG6KuBQ/ZJ3/9N/gtAJzH9XLy1qaUzE3a8d2S721/MniWUQuRb3AMDSr3u
6VzD2S4qEUn06Hs3eBIqRwRUk1Hl4qPiu4UE+siTqT9WPsnbxLooXkka+PEN0jH3
HnL60x66ElF9jey8K5sEm602K8dAP3sdP27JyUw3reXaytlegEnlopVheYFs5QdD
IYLCidEQHy/4AbdAA4UbuSNLCyHYpSEq87cHZbbvoHPegqWs4FWecatk/CLE8I+h
KBzXticlVb1cC+F4Vg9yc5kdqEbKInSWHK8gSL/Onhr6ZBpftj5ppTy64AMvYSqX
fzqItoQeG7u2Iv2UAgqAeC9ZB86t3Qvh86AEqpN7iBbinlm2hQOqCTAPef3DiVcr
xaCo1rkMLG4Oyd/+O9yeCzxcfG19yuOHHBa+sGlcRqZhlnojSa4kVS1rronnhker
HP8C/FfSMcvljpRJ8Bo1vK9DhW2fl3v6JKs942mbexQ/MO/mjIT5l5kAhO4j75SN
TEWzNXX7tQ9ohYJ78ou5lPFilLaX+o036DuQJtYMtIaHF7FMqxXhiVslgP4SQmap
NPD6nKMV2geNZrxYEO7TayMH59oTaJ4lvt1gZcCxGjawTXTcTaHimtQSP6uWjIvf
TJerllHvpF3gXx41iTABZoViQ+3abEjyB34zedkWSihDE1Aja+yRLDDLPGojdpnE
VyD3O7r7/5G+7vQVTmxt/aQs8xkk+W67p9gQgtVYZfQC84RArQ8wOtODD3zLAfsS
v9tKb+CfMRaViEq1pyUIuwUHauhIoQwmoRK2/hOaZpcWfNFE68aJxO5ExUmgrnoV
X/7+ESWKxs3gVaCRaTRmkUEdLc9bejo3ExJLad1LFx/cZKsebFJrLjQc8Sv+dFu4
vax5JSt77LU2I2tYqfVK4x/HUr3fBqV55Sz5p9a0YZlw+2x439GCEWPV+yNUr6CG
GuRXyDbN/jP/DuKuW9i+4ihgc7+vG4RFzaLsu+pOeRz0JzSjrhONKe95kwZ2Dshx
fg+GUOIFcQtEKsV3mhyPrRTHsGJw8HxvP1ZE0iDBQ1LnD5l+E2x3hUEvhFINql9j
fpQbqvtN6vvd1Liclwpe0NaxSz9FWs37tYQzXmUZoE8EXGsZ2KfctH+xJzbw8lfe
YJRgndjzOBe7DdgYwp4eLGMPZGIy7a30e61K74fgw7/dh9JAHu2+FL7LCyhkaDi3
vJgBbOnPIJm4o13dkbLvUPWbxZNqBNyWpmFRidzPI6BILGZQ/xKSxrB49NfUk+75
jsFaVC/FxaRCXphLuviMB87KLtX7/aR+2nDpHB7zMd81pwvW3/3seEB0uJLwjeAl
oBkT49wLzs3zDs0han1UaeK2Bk9ueBOFzDss6m3UzWZQklhrV28W19A2aO9isCBf
31ExgsTpHBy+SwZK6yP9/C0kqVGbV0XT1t35Z22Lt2gMwUCDMJA4ZzuFK/W+7Fb/
fpvLI8HLgyUsijdolPlbzTmR0dFOZ0Hzwdq6mkvtgs+l3eUIE452dEeBAY+Oe74X
Eqr9oIlCAPOdcUQNyiNTH5xok7lH+LQyfIJNgDXKRNrzqt6b9Ncl28I1uXzdKrY0
JVPbc4lMtGJkzy3Ne23f35z63V1Jpgb4HGU/wVZyJ78N0D2cp0L9aYOWjkGc0OtP
O7UTCmnNGj5+NzdfDWxlOic2m1EnbERHLAD91YkergFdKzcQh2kzZB0FxUHel3Pd
3WC/5ZANk5Bf28FxtMV/HWFGv3Odh1BozLvxY7C1u3Vinxp8aHhSmvdoUy69YBI5
0+Uo3UyFL2tfyqQZo64BuppK1e7010isnBnU3/o8BMcadM5vonbTr6Bg4L0S+5yH
lFa/wI0w8umWw5N+NZNYtaDhxH26lxt9qADtYQWzxnlg9nI/wJZresDq7J1WocAF
k9mK0wqsDlzIWWrTP+5FR/mD+vZ457pZNFcvyRR7YU00Hp/MudE9F+KgfiTVI+HW
MgvnKNzmcOQBjCyv+6Y/akDGe1lnvkJSc2UvCyl3jDXElTl3CnZpRXR/NEVJAp+x
X2jp95ixjjKHDbdj4FISlfiX1Ox8OiSf+ESSKlmfUmEAZ2bbIuWY8GXHY73tYFmJ
9X1a2V1WYSUqyJrg50xBydeCV9Egd/L2nCWbQxqM3/IIDHMipl0VAUXaKfaAq4QP
Et2a5j7MZ1JvurmmEAy4VITigZocp67HR1ixJm9R1S+5V+okvqyyqV8SjgQvxlHY
Fhng4/fluoto+Qs1RFZQOMZZcHtHhvpES4R8g4SDpGYnHPZwsrnQUzP5y3tseime
U/c5hFGgQZvO6BvGVzMuSULMJXiK1R9oJycBqcoovC6CbW1NZPUggoi8qHvw/Owe
vTSz7w4IrsDOlWN/2mHTAndVBOUKF64fjkrw7aAtQqhtYxgUYh6ZIOkokjbXa8ev
mNSVUrD0jRky5w3UzefTLRHQVR6xGDD8mlFnRoDlHIt3K8QZImVU0AezBpX8NEsW
GaVBKkwq7uQZ0V30ytJGCrPSb1vPUxz6KfVK6gxHR7/RTYKLKHaFsS4xMeIWmW5u
IcNc48UNiCBa9iuHLfu9RXX8Rt+p+acaaychB6Re18ZKuTtsRESAYk5dTGEFyg4D
5T5BlvT4MaUr4W65Lp03DJJysijkTV/KVNjqbXe5fOhQ25ODXyGT272ANM86rOLt
jpHVb1BxHIP9GvkaiTomgdwU1xLjEvrDbnXprKUxv/tcB88V9SeprHne+yzNyyVj
gENR4U+rpm8BIx7s3NKDb55Ja8pF2tx3oJ2tDxhsou7Gp3Fr/Ju1srA0L0zPwN2j
5AXeT430yLCI/ZNm/Cid+WYqtOpeE3G1AC3lI2avDqx2E5uXTyiSICfwO75gRyqv
Oa6S1JW+Eti+EzN6WV4zYdiNDWEZI3EkAXA+dJ97kut8ANQK1InmercJ8w+TDUOW
DvgyzKqTWMGu/5xHPLCdAn2nPtyTcxnOqr4Qz7k/AAp7LEfiQRgJrlTZBPRhXg9E
5JdXcSZXN64lCDvNwVgnScLqSQBJpEeENzJUoRheRZ3PtZ1evcbWtu0k2KbDRRYs
j6XQFMOt7enI/JZI9qNAwP80ppcIp4DPxwdo7WWVBgvTCiICVSySuWGjCPyh8nRC
0ank7j5Of4JR7a54LDxirgtLaiWWKHLnrh9IkuL7rv0RKUThqceLY5dWSS7h0Z0a
vKXtKcwOi9UlQK80IjDoIXRxfrkyvoovsMmyqix3icOHUftsmBhlH2kLlfvD2SwI
VzWfeuwACp7/tG594GyjEIg3ZvSDWQ37iQt9/Xyg/Qok8f4XZjtAlGiUGV5yRC6P
up6UOX1nzGwhJ+woe/TNC0KlOFk6yEihyoHms4hhiWjmSI2FPf+gtg85GEF74rNb
3JaqAXeRZypRk6DyZUReFkKOkXYQzJV0+qjfp8mCnRfCSBrUhUG0asMJJ/DXoAzl
egDZNrfBNbeo6cPvQ+48AjwBl9ThXf5TfWS0A89dpAutJHHszGcv56q47LmLhUjk
nQvh+4Hxz3pJBu8b3Vc3HFRiBOfXNMdVW1neIR749XZOGkN8hqAPGOPyVTbHZ6I+
5NSRiFVZp+tIBEVz/f4Dul6xi/E7E2ZhQduUANFaznwZs0K80+5mcZ54egdjVGNu
ABQa0zFhP6MO9T+qUSB2Vbf59H82jxP1K1CGtukNZX7fYp2acSy/lLCLprN/NOy9
GHdQaaSQOIUkXXYHveXrJqw1xwWOrOsRqsOM4WjG+B1LazGCqSfwupiVezPnigq7
aMecL+yF8NAqQ8jgC4dnHa1vnct/h51XicEfV12xFTjJyTcJ7WQ4/MYV3fIPGmC7
qvGMiMLPPQsKiDO7sygWnR6NJ1nNLAYTVchcsTMujqNIE+5vrNPLw2FWX64W+GTx
zJlZAMFqRZcSB+ut0w+mEhl+AP3prgRwxcJYXkxH+L1Cptz9yyr6ToOGRz1LtB2J
KOFHS//m6WPPlrtQIatWCJWZYqr2yhRLuLOdo/KMC3KTF+SNd6wwG8/vRtI9RyFj
qI9mKNW7qU9/fEfsdyeghCYrQt3DM4wqrODjsLE244uppJTv53WKXOwpI4bEBwNi
3Rtcwf5q50+eGlDAQUKkzIkCkJvNQ+fcUhQD7TgaNuQ1Yz6aupXCFjEz+CqolQ88
z8zjrvjRN63u+xDUKKLlvCVHY8Nx2QY27kU+TJZBsC7BDH2oRvFQRqQr853+vYAN
cJWr8SkE+1p8FSt+v+tLQBKq8/LJBwQOkuKI0RHWEujiqSEkHNLEgo0a/UVpdm7t
4ckpZEIWI/svyOCC2ronjgdVgifGZX6LM6hXcMZU0apPf34lcc7NZsD+X1CE+n0a
hzkfLYZhDEsY1iSldjL4fuTXeEvgqlDDEXzFYCFwTreTMknlpzM37qF58QQhxQBS
g8/HVnVn7Rl30w6uYxmIiUBGKbv3rQ4GBXxCjDgUfYhoEVaKy95TeY1sOZBMtIB6
psxA9+D3VWBO0HHNqKykuK7mBn2S4mSvyEXU1Ng/5msLydi7W1zyN+yr4/0+t4wU
1ra4mwgsJVylLWOveo7biifcJqegb0tPISIdXMJpoi/HtGnvSB4r7vp5Ta/uWWEP
9iruKSpREWQzNyzzoFUmVF894QjMaVM/Vs5HzpcHEoERz3GusdQtfVeOm0ldpSgE
G3X2dYbfEKPiliVScyXhfn6ClsupWw2f+VQ8go7lg8QVnq4tDK/OwhGZR4qNoMmn
UHSuWZwrUm+huaZaPYjhxtABuElj7S0htdWH2ZINhtWD4XGaJ8vq7IefcfTECGhF
gEUgijCWcVbl5q3HmHPftB14gBfy3Xx0enNY2ZR2yFJLLVSW+ispiC8t3lOVx71f
O5uP6g0sXCfZ8ZyDTeuvO0AyhPJ5r2PL2PVNEwi7ORSOCgM5N6os5VRKhV7B7Ymr
fa0B/PYHC2vOjigY1qnGnCMXnAPpXnIDayEq8tXRMcpCvpiKHzIiPQPZnDDdFyw0
FNt5Mifjnb6mlOO91I5RIvfWNg4uoRJOHyAQ5TDreO6uw2lLlW4dVT1xc1NLA6NY
O5coswzN6wdFuNzRIRqI4KC/ooMR7S/3G3K+gEy2xpviR11xGUh571T2xg5DR/cu
FwXJE2VjjF9T6sSKuPBmT2dnkTHKgJlNYJYtHXG0Wr1edZs9Xa6Ogsu1f/AKlJWS
CVoeO9TEkfc1wJcGGucwY0QhszdLgcnTYpiLWD2n6YZ9gXlPRUY1tgVZykn57li9
NGRdWPMsDoLE9Su0WGqm1CmzB6q2cTg8HvOGVN7hcZZDwrcR5Dj7/Asf0CEdYaDR
F0SFhLCjL0NTxJb653wfjyEjClLzhqsP0u+mMZOhrtfR/xqONgr8VWbi87bTxFhi
mSztAsQzkWwNwmmouLPo0CzqG4EkhJN3rVOKDizCoV8I3DKnptmqRhtMyf2A+XnP
1YIZdCQuAJEwme9iqMWtFaMbhIBlxTsP/+gIBdw37XSNxS2yOg7c8eP1MdKBP22h
zNiX3Xc7ZpxBLGxAHWfamtznMcRYtMHeuU7aCq1Gi7/MTO/nGY6DkBt6AaxVuUPt
in1tBFDa/BDpb9IBSeZMCWHvoPpt+FwleqBjqNzY78OaZBf1PhaJJoU5Avm4VEM0
28Eln8ZAsnLqrQZrEBCaIlT1WAXHCZ/rpoXDX7TJ+5K7KiDWpZE8iEeoen/1uwWA
k3JURaF0mL9QzPNvnbQf91e+OL0SGj9Rso1pHsP7KyhTpwBOMGUul7zjzm14+E2o
HFblpMvmiGnwinpUq2RTcGV25oMnHGZUKzSeRyiVFIJr6ocbx0bauSw9pXEFie+o
A+s7k5cjMPqw3eskIipJkzkQoGDppDI/sfD5ovjBRG4CoKJ/UwIysn5NHUDSlj1z
BbONmnlT2zMsX65y73Ds7tJ7vCmqI5YFIuW8wnHc9+ixKVGbPeNO6vz4WCAGYmzd
ByQ5Ax+b8Tn6lDMNYym8Shi2eM+zE2oOddPzMYE70NA2GY5STTktwhf9f2msGA38
uGUzCKmwTdr50PKL3vhFdQgc4Sgz/cvwp8njBKoqojS/wRBthr00TnPy0Dc8q4qx
RF4GNp8qZ4eHP+0y99cigS4R1xF/qTLNRAnebidBlQbOY6WKVy252QTHaV/loFLj
2GjiovddvzvG+DlyaahCsK+ROAYwdWvCmA/IJY+GXivgS6SdgJaj2lxiv9PPyTHi
57RaPDMUD9bgEiu63YulP8GMMEGafIR1TY8yBufjNq2o9ktz1Ogho+IVVyr9bFh0
JCbdJC1XFIOnFGUgTDEUz6w/VpcdCi+svz3/VTdLdFBzET1jPi6UO0cQWiD/NJp/
fiks2q7AsMtk9pn2REcP05YQtafoxCqG6+b62mq9Hxe5fSGmdLMSIh0ETo3wRatD
jVz/ER9+iz+95k9mSBQ90uPZ/Kdnd1ntpAfAdUOIFmV9msRBkSoKCIay39CkVYJM
mf23AaogkuPRQTYNVjvMh/XBmq4h5IlstKyK+Gg9hwfnchZ5z0tszndggvvXM8GH
C1kgn23k/eIFSdkL/pBO1YR55QkCesXdGSa6h+NuQuI0xhpxJyJ+EYexZvJxb/y/
uVUGkhKIB+ewc8wRhXvB2VSC3lhLEV60z1t4nalJNAhjV25wz3uDYJCKjDkomp0Q
kOdjCIOg4K9U29bEoL3v6oM+TG6JNz8GVwtHg9vZEpMD0ie5Orm0apYlMAK2AbXu
TXP1tBu1FvvXDmCyX7epwIDIprHSJOhGOI+5+1a9bJerwgiZJTigRIn/YAI7OgXc
cZSVae0xkQHri4gmNgiycX97+I43vvEhBkN5LtAeTjBAqaaxHrIsMb/zpE53G+iQ
Ks4UJq3JYB2PSSJAgqiyJFzY1d/l2g7+EBB3SwXLxxIDjxfC3DbAnE3TBf14OxEL
eu69XGa9xoIQDiHAKeICoOg/bfvTH4HtafUpPF1GqQOoQeuxGFg8hgiAG5iNuVS0
a/CT1ZXrE42CkHaNDgNqQvc/uyvnIGhzzXosgxGYIpzZms6NLWGn9j0YEQTyVsMC
ll3rrCOC2NKkTxtkXgHUwCz/ApqyFNPOzVqOonwcZX2mjjgJUyYwCPamvycZnxpO
hqZD0/dmXa4aLi0PBizMtbrmyI7Ce6cuyMIhVvOfbZKwOOp7wEmxqHDM0JA4eEPc
5ZWH4ym1LZsyw9PVBH9u9GcyYix7AZOA5GvsjvMlhj5xfCZbKBwEY99e8SJ3SWqc
hdWs5uc/7KeBt3u1+ds7Ev5gQw4IjaMwAdVjHdYYkPbaphogTCCBAcHCnWK7l2WC
Qz4OPxYRaAjNsj9tdbjOXTFD++yH+LayYFyftTv4HjmC+b3gxaWXOL8dVRpwF6xx
z3jy5D6PGdGZJb0LSJaY079by5QBlej1IvMxKjiCpxiBgLTlk4twLUKV940bDd5u
jJcw2bWIYZEgNWc/QKuarr4Y5SEqhTBeAQ2OTI655WZUNnDKgu7bPTUb1QR/0h6Z
AT1xbpEAMrxQCJ7+MihCuG9zErs45z4xbxafafsWZ9s2tbx4LxxyJFgWDHjyW/W6
X/vGoCDH/70mXd0+LUPAQkU7sqReB3T6ueZXoIzQYvqgOHy+WMxAAMwfwDnH+NQP
0EKbq1300ip0avsxwjadAX3/LgfPLNWS9N4M2WQytgQj1zZGkxRrJ6Tw2t/xmpfg
wtJacPt7ILSgNCVFPZiPqTT8/r493b5QBkIA5vJjOnt2He30gCGzwaFxHgmVPBSP
7PJniTY57nhPyCuQE3aElge8kjPEGGsYo+Df/XSStLKZKivOk2ryfIkWRe/RCbd+
hteZiP/LUcZoZgsoPkOmQBxkknxgg6Pr1vrQGguf2cp2l3vFkwDHU7g2m7TxFJgj
Z1MXxCDiDm35MOf5kRk2WcpIJcok21AbsDriFRsv1Ls5wV21C2jyvxUJ5I1GMDS2
hQ2opcFUQZ0MaSx5ahPvVE6AVpA8OrEno4jDOvHmCLFw8g6bFoulzfiqNRY46Xg7
GaN3tWTJP6tx8A3KTFxiwyTNi+iFxLtI6mEAzbMEXn4E4Wow/Rx1K47IC79+ckez
yxYssAdYcbvZVmOmBoA3QZdUWyOroF+egfJVcTrCYF2MenXehKMInxb4jPjo+NO9
nGkZoqsg8tnLvMXjjDXIyHuVl1skP8+4mWQEFBljuHvwmNHHcKU44fYlGEFMd87S
8qzegbqU4QrIKyb2ZT5NHn7QnzDdNhI1R7iPH/hYGcPIQuRwuzOZCR9wObl4gjd6
4143U5YZb2nIUFobBPqWrUqc2VuE1CaE/ZgkEvaXubAUgv4FYf0+LKR+aSNwF8C0
qVYmZOpJd5kykjhP2CeLkSPZBSng905wy+ysYlB4a7QGRgHDQ/3eXXcf5h1nUpm3
cHurqOWih7r/tMO3LCAcpYr7j0rQmPf5BMtz5CyVshhVtRKIcGqzqdlzh1Uz8Y3l
u6nCfT0Z2hpPCTGWrmkQGdMwH35u1MyhOrfslgufaZdkx1e9UBw9ibHzUySEWIJL
Om0sbRzm5JTzXRYASHsdQzSZeO6LveAEI1xsS4V1cg6BLvIOoysKi5K6MzUpMYjR
7Qw3snHX7Z6JFiUPWyoQEgOCVFQtxxpw8qG6IhPu9ud/NUWCugepwJIqHiWgpyUJ
JJmno3wrihsQeiPb+c38PfVQHlUHBgtDp9M76leohHT9gzY23R9yTMFx79f/tQMH
j+BYHjVcHcReyTV8NHjnoXV1yHFZroBIDjIjhgvn3mndWARSlr7EkJroCauVIwqF
GkTubcXsUNoIf6cV0VwBnJMmnUQ6cxHrUu3DJBj71daILjbwfMU2k+M5HpnVYBUq
V4QYmGoaXlA98a4JjqP7lXmp9EQ+XwtOVkP7YyZNbrsPGf6F3h09tIwHjUrLbqpP
zMlYlZyZe++Y088NR5X16ebuyM72Hp9v7Vpf2NKJpP86kRwtxZBG0RDHPmnrCuYJ
FU+nl4FNHarEe/eEG3BopQWs2rIUt/FCYXxIVRrnCBh2HPsBCAWKGcI4PqU9J1XZ
FHFAIm4FoaKzem0voAYs6XurRBmLQZJ2pjQJFAQveAtI+TYvoUG78X+nu+NM3dBI
KJ3Sloe8jPfte1x16BqjVf8SwQexwnzaVUTugsepBpmYkowIE/gf1WDc0GRjrFyi
Jh+yFZN9obDGu/lA6BLX+XH6N69Yx++Y+tUI1/l1cNxizOpQxqToEEhcKSC63xSM
o49LbrgRz3aO1tzry8XG5E1vFw5UeTq//N16P+2IRXQmzPcGV7VW6esVKWbjWs0a
w3LtTaWlwDmfscuns++a06Oambd2lsrm2Kk9w2ypZ/GjCmXa6pRet0xNeqTRV1uZ
tOC0JX7k6H2P1xHFraZVkkEUTrhpevMFeId52dCKZHbKqBxE3lXhiQShPSz5Ia0W
hiY/sG9F7ZoGXgUo5CM9X6X5EssVSx67UI+3P93lSnw6/yiM9EdxMMo+Frn6sPqU
Esg7LLnqzAEV2wVZkrGcBpQXQHEfGJGoqmYV47PDunIX/urTU4QSBs6mUkI0Lod9
5tXs6XVEYz8o6zaHwfPj618y2H5R7ikgMCCtQvo8buYBifS89lR45FzACQRP/CN7
+h7TRj1dz5iSdCBJd0/XbLmt7px7FvZlQuEEN5kJfkvN5VPac29UgkD3oVLc7erh
7cfYcnk4DCemg24Faa7axGcR1Lb5/LHPP6TNpPH11DBx7nDAFC7hpPB0EmTTiG5D
758rMoQFU6uAOOaWQQOdk+XGTZbfTT5okLuHi2+0Aky86Osrethtwg5DBjMR9iL5
vvEIpjz6X6RkZ4tgOB/1lpb9w1hngd4Q2yjVkfkc+MHkRuMYqpX+t4crOoTKrPhb
BZLY28zm6vlP34eyT2JEWQAIj0PacIc/A4UBGOCy/iYdUl50xFfTB5GIH7IErplZ
sTMb0Fs0v/Xo0Wiu1iRt499uCYShCmGvtpybdbKLeMFNwr6+tig8M0+CzJTKj9i/
ngTazFU9IOvaWoEMcU8cG6iCiR9Zakv0tTqbZcUg4Qe/rNlEYge+5QkmuUQ9FE0X
1bJPIKMctww3+yw+3rHpCpDAW3UG+XHvmo/w1ZrrHBBcXIHAJw1C46Yc6DvOJuY9
6oKLSEwmxOnZietLnZKTXsE0Z4xAg3CmDC+5ULZMXl8MDj/ofrmN+8HWvoDMvTZZ
RlpNQwJXFUKIIDP+sC6kjE+L5GVwgj+VfOS6PclVuv1iakf25E8ozzZXwXRKoKNT
RRzpCGo4E6jWxzS5yhfZgz9BPz+5UVMsgS3okpReQLm1l67zDIxmyz9450hY9s1M
NNIGukmPMuj8/uEi5Qqci/3KkJx5yXD+aht8HhMr8Yu28ExUhK5sCgwnroaegEzE
O0JNMEp3shRaAfkYPc6mjZSRAKpBho9AD1Cb8fbpK+ymp0tBzHLa8s19XtoF2eNp
L/0qLVEEXMCc0Aao6QLkg+qlIm0e5swzJZrW8lCO9wIhA8piJA7t4+ecTPKvuZ9i
DLVlDnUb5T9IT9ufjxu6ipZJ/I2/ijUS9MCWxZWFEd3rpQtIeZjahmxj7auejG9x
I21lZZinOAVWWF9AeN8qwwGhJ1GMbhwD3aQTfqbt4PBUjjqCGuhEvyn8KW1YWxzh
cKD0hJYjBhdZ3Lg9wvB3gjf8rRQEVenpr1HvCqwLPujN3343FV+OkvyfZM18qQmS
0nGsKZuck8jUZZTCVL9pItA4z1XzqzNw80uqb4gD0Wl+rKvzJpps88zhCJFz4W3b
jQ1QF6uDKsGJufCJMpcOcbvZgHyxTdlQwclpg0ZplcTPtcF7vIxhXei9MNe0zvFu
3R5hlY+lpgd95ho4NeqocnbrBpMtD2idwtC87SZiKXgLKZmOhe4CaZcRvrO19ttN
PiGSqVWc5NKSd1YBvh5NsOhzWaFc3x/IulDylXUQEBtARcONQxKqGLhby45cxqJX
UphV3waWMkmuUmJgtqvGbu58xpdxdUiTXwlcJJCXz4wLiJLV1OXTxxlyrMjljYi4
lKTSqa1P7DlFRIGSEhp/2ApYZ9Xf8wF1u2TGTyAbE9UAJ6F9bl8DAeDD7D1NHrO8
bGLnWt9lKL2w0pqeI3fVAp85N8o++4GQiEZbmb33+6mcOB+IrCm1emd43iJyGela
TCcMCPnBgoP9m+3NagnK4kj/mWzxoPjCJg3WEZDWpbehfwj9RFaUsqSXcfrJogSR
AsE9kHAk2gDoVibwTYRUUIimqLkK/lT30k29xDIHKU2xnDHM7pv0adhRikRV6YXl
J4PKTSIoLjNZ3nWkSevY2wp2uo2qJhR4NV+gbgSAMDTtB/FfRsjxdgRiF96EBcSQ
TcFA1LlRSSf28ieuxgmWYf1QOhX1jYq7lUm7QFlRHThbvdGejqbBvDSbBbkbJFKB
w0EDD/YcoYOn7PLB0CjyT/NPsaU9rf2v1iYBADPV17D5dvI0x5FVGymBTSEB244R
AvBAmZwsUbWOzE/iGuM9AZ6Id8LM6kyDgWcYVOq3H1Og3FouUH6OfAaUWb64LJ91
6q8TK/TEwwnncvbcYWGKxAzzV3RFO7111JgwC6a8l06pCdrvbPfU6C4RzTtflGip
MarxX/GlAEwEJjS0nk3mqhh498F21Rm+K+NSto51ynMjIcLXZ4f7eF0BVllegyU2
ag1ck+DF9c3G589ub9qlHovch/1EH0+rnOB3C5yDhcHpUEH4atdBUWLASYeNPUEj
qnvaOPKhXf98r7QLLvPOz2HT8F37JfhAbQDRWtbUelS/fRAWl5tzrisoyuv0yRKR
wOvzL4MBfRkq7XkWXJObD6OEEwm8Jlq/T2ld/1vsQwDkwuLPonuVeaYbb3lmYOan
hZbg9M1/P3hka6nK3iO2GwVI9Kp7ICOFmZ9RIBsOMxvVfM+fveNa5+MfcSFZiiKn
+6GjJGeLAO+RcLVoCTrnqzZG/4SGU0vp/8uFZ+SjV65u0zd4XvWU6WwnI6vnfQuF
KwBruBU553KObbBfl4aLyyRm8AtU5nMuBvBzKSNAtjv5q89aa4u/+cfRlwGojUf1
cyfxTnysGRWtf5tpMOm96F+BB5Aie3+IkWTmIXIqwaPy+vqMRw/iqzIZV7/+AE2F
XCIL5Xg2uQag1oO4l6229HRsRte/YJfuh7ypItcThyabyA+2XBkEbp5jNzloDSEF
KsllPJMVn1Ef+omG4WjN0Xik9OlARzataYcgdFoEW4mAPRKFRo+eK1CSpQ/ZaT+0
CTQnqQy1OH5z/alTtMwoWgh8w5EAGbUoZo2okwmSBb/KjoQKjkzYdh3sFY9bea+L
ZGmza39kZZ5N7tx5d6oKmoweSOoM4b6c7kqUQtkKUPY/mF7W6UhUBsfecsWWzB0+
Fx4KkSgQ/0rSQ4ViQ1kguR2sKRwZpO2eylmaa4dTwjQwO7MtfKhZW9UqPRSilXgY
3xLIP63OiiBA8f5ZOR0CvSaE+JTHGTuqWr4gRhLzqqsM/jptpfnYAz3uoaEG0Bne
IT41K3xvW1ylwozkQMVhhbfqU2KDa0TvotrX+R8DO6BnVbJn7nPhdqcnaPg5tXUa
OeTsUzGdM+yadR150QO8dxCPAX3gc5ih3kQSi+0y7ExriDBtfNjj0JN3hUX5JwVU
j2mM9foehjwf2EkknhHB8UKiNufNze/ORAG7/avfK5BNke8TeSJDoNJ9I5boElUp
eREVlb7C1hXgTGTSFsqJ6LolV7ErWtz2Dk69MnaArd5LTRliT6BBP0cfmCcXDZ2t
DV1FeH753ioQb7FJqG+5zhWzH35dlfVvreSYBxXjyIKG/wJ2E26MdyE/5Y1wN+l7
lglnGtYoVchmWW8pbbtvGJ65khMCBxq/t7qHhr01rTphnbR+Z1hAHsIOqzRu0Be5
qXWUZnu6rUO2pKBPUJInBNAl+JIRoXM/2X6bQt1/TuDNtbvlIzV363VSBMZ3oh7+
toS0AjqXHGUzmeFGOQ/+HK0PbSVOpf3eN+MuSttYbeJWrwd1J8m5zemyIzM7xI82
7i4RjtDMUPfP7EnFjbyT1mLMZnr5hkpyuoCEu4OZnz6xPcV72lIExCfi8EGsMATD
rSor5Nc9DfI0bD0n9C1Vzv1sSAHGZ8dlVyvDnu3agx6cWyknfGyKAvgRXCRATZnC
MNFIycR8Y09ieUR4Oc7VgArLcuy3AIV0Nu+hAqo1Urj+/xOPo0CJN7V9ELmjut2z
BuwjRpUEOVG0c3+6u2w8T1BKJTB9pKudADqgGLUi0Rxm3bsGx6bbiH7l3g2X2JAj
/nbiry3iSecfh0fcDtsr3nXxHcXezkv0j++f+wlH4A1aLOSelFmKZAWcvguW+GTh
0JS2X+JTQ+3tbbZDYkmEoFBPZEO8Ur3xGO0dcZiRGSfTWiySfE31fS/j78blskoZ
POoh+IX2gUqTlpsMHva/5OGVyn8NwAnJoU1bomX1dZVymCBXQWvyTOx7F6RYhs8H
JFb0d2UNzUav0puYPI1UzfIPansYSmKsX5/r3XGPrNtuG5ZcZ0o6hd8R8PUdG+Ak
+RHHD/U9yHzhz2b3LVY8aF0g4IhAlyTdUS23FJGz0aVjJXVhkHUopt1DKwKedymA
z5aVNLHeyp/nAwip8P6RO9wIuECG/L7iZXsW9K/p8p3Ltzqf80nMO0ieeBNSWleM
7hG1ufqj29xJ0ngwqidJLXsPjaimTN2QzweE0e4lRsgO+oK80MG6VsAt8m4K+Cyz
bo4QEOs9chD81co+pwu7OHh07AGQXJ6HlTgIxbOYxZtLx+BykHJK0P1rgVW1TGKe
VZf7F79b1ziC58uqVGiOnE26JpnOeoURsUbiAjRM3rD5rns6Oekg0CZCPCLN8l+n
8zyJpJJO2FFjJz3qu4r4M49rgpaEuJ/RREjjhbqU2+UbatRY5vafC7e+FrAoXVD0
wuQqej98xHRNIvDKkJTTncnV9NMEn47o82yYoiYegannGi5MTEUoPyGsWI2im6gn
f4o7Vq3lpYzy3pY/bNuQS6fNOtJQ1qg24jn/xFq9fm/QVnoIu/0TmrFWk1sDNIS0
JXOjklRHpntcEFys3UnnlaE3CWpP8CvajTcghoxTQ1/9NTsBDvfVsyPiTLrs+l1R
I0nG/3aqftoYOz0d8IxnIZyHW/kcFFzTMkTdfayiYRvnrwMowjEiyjY+KxTHAv8m
30i6BkwOT+T5Udtbf3CT+IIwQ5zqaU0TrFL6n4WD1LLL6+gCBqAPxRqDDp5dORuO
EyYbkposhkmlJutOizeVBWafJvXwBEayVJtTCuF8Pqbe0u7RYkLgYMXJjaC9A2Qk
+bto67DuulIILEhBmKkzHAXK2d/vdmL584TFSsVlpb4gbF8NY2E9oOvDzzvvYSqc
XNt2mkd9SmzzKMKGrdctnn93R8MHCjByfTP9GFMWn47bZb8dvd3ZGchiOJuPWREh
w0wGGZnvwXBVq/74zl3dWycqE91VnCFUzpADRKdh6tkBRejVV9RmkXjT+nGDzliZ
zkCnmPjjZX9BTs6gAPXXGIpSQZhG5I4oWW3AFePo2W3DK1byx6CsRX6kY8KEqs3w
k76EDX5qCHXaCLBwwjhraSCcgq4B12qCh3U+gDBLRVORdgYGdcureKeq4aBAgq/w
Tli8iSgOuKGHwCDC7BhS/5PKq/tOWJfTc14d5YA5yJrMKAavcdIKWil9+Ykzcp67
4ippSABc63YYBHWbuIoUswjSCO85utxrIH4aNkhleQKpZNwOzNdZ4sdsWnLthIMn
Zy6XTyPX9jHBiET5n9lmYCyijyH0pLz1znPQbSqVuuzg+BK9B4AGpawLVFiuejgh
sVogoofv78nW2O6lDg+na5+nvD4Z3av8Hh8aYrQfq2A35JpDxngu3d45m5f+vqQM
yDaGrZI1QXMdYIKOeNy6C19ONGWiMI7FV1pa4rTj/S5flgmvXJdvxj19RaH94Z/j
nMzcHjXhGmkYLBpTp6zZDKZnwc11eO9eB+GmgYYJsbWM0CxDMOXKogyMAcLi9XZz
F5F2PpWZe8eRNv2S2clZxIy65lXXXlDVtw7BtkshdLI2mzoXDd0oF9UibXrMV1Gx
bItR8S9Rznn/hkDGfeYqf3Mvmnr/Cp5/gpwaw9ibcJHp7ZUzOOqMH+5PI1QRiFIk
zaSHUVvzm7kxaG9pj3ztNUkPPb+DDlw7Ol3aTsoJc8zzJ4JzDpjaRch9lAgqLfis
M9vGq1tvWXJcqn2fEEh/CJzZMbm08XKUn+M+Gynd5HzFna9KgOoxPSHdWoER8XiX
ZZX8oALWz+q1vIEJbByRy/O+kx/UlNnG/hBddsUlSVRQz4ZfGP4wJhglddtQXK9G
iZlcrt7gzCLjoP36qCVvnSW/gulcRTuNyZL8aLlOJVu43+AVyqJb5N798fTvzE06
ItKT5yqsjH+YcVAku4I8KNAKvE7+gIGaY/4bPE6ILDPTm46cBP1Jqnv0od8HzUdG
bwtWc/+GKt5/iXl2onsTNYOVoBMz0swRVipFGIxTcRkhzvVjdErSxWlHBoMeSIuy
xDq+Wwj7t6p3n7sg0r1NHDd+VDeTIJGFoNAGm+N8F1WcL6CO4bq49i2PjvMoj33I
6aOs8NTaglUw7rgJM+xeUNWj4KqZuhpmrOUFlzIcr8xhW7vaL5rtslNg2WHQOhfL
oOwF7ylIxrhz/ovAfXqxkrBYRmATMVe+hRcLD9hfULuiDyqFCvSw9lNhZp80vjLM
8YMkW6bEmJ4Giyvmv8olHkuZNBAnU8V2e9rpzzDLt8jF8VBeNevRbRniZfzqzSdI
4mShrZzHr5QO78aOvNsisOdKiaUNHkm0qy9QrdmYWymFrnfgHzoiF+zmoGMZ8yMq
ZJ8gx+mR3cywEuMURyxtsvrskmlF9+DqnaypkmouXt+QzYSGqpiBikNyRlUe8BNx
ril/QqSnsMiEwWkU8LP1WgCOkQgJ9Lbbv85swage3tP5jWwznhYOlFF61niwy8x9
WOsnEsewuCEijHO6ceJb50G4E4QuKAlrvinShzN1idaheBfz4O85m7ssNJOh1lpq
sFp/wV80e5spEPfHTI3mYixVxURwRElcVIqqLNKmIxqmZ+nVgxKiaFeeCkyI3Ewo
fpBE0wOIKKExspFHbjQGlYBJfU00rXmfxs2F1Ysbkb25iMJXZGkpEMTeFEvb1QEu
edXz1XhvX+R8uyYHtIberlqKnyB1WeyWyv0/Nm7IctwkHcve/ow2/MMu5r6tfSA7
KoWddjemIaSG81UEHZ3qhFKDJzJaRONVW8ukK7rP3Dz58l+2s3sMyG8lI7U03iTA
kG67WUhQ+djil+VIOsZ2Jb9U/SJgNfM6Ydbc9MrQbU78rDUCpEdY1z7acKd4qr6F
DatQk5EwcH2I04pgVmJZRqTbHdomP4PMqHGE3iZ9spkjhTXqgDMRlhssQrrsTDXp
4J2Ig45N16v5T5ultS+iPv3SqS5NKbSh8vP5f/xxjVXRgjSOsgJ1cws/MDsd6mTp
Fg4qmNiBMF725GpXYCtfeHMw16MnvbTpZ21GtPo/yYeVKqzoTk+Tw+R3BzlL9F/F
0m1/7T0DNF+LJQ2nPIlb2larsVJxH6FeF1ESYgpus2FmnuNnZjD8h8A7w5U1ob0y
tNZUJporQMRnzcBLDYhGRR/zvsrO1sXaOn7hh7xaMPrjCN5LCtvVF+BtA2VRe+9Z
eqMzHhCTTXA0uhMQEm5MIwntPdFCDjU0eR13hDMrlks8XAyeoap4s+d0YXYK+Tm/
eep7eI4YATmEUR+xpWczmk2Oo773qs9RNNjnixp1TdHp3spQD7ifPIoygoGG7tGU
ALiMoo5+aUAmjiNLD5d+553q+V6UcIDT940CF+8BEEaFg7kZOdPPOfUggC2UD/bv
ZuIZqAlWuzczZrGr0qNMWZTfsd9xDJ+44/gSD6cN0eV9RJAg0NzW3Q0/v/E33gxh
3z9nhfkqKtFj56RmVStIsngOCorUiiwbR23NdJs8WPaJSdDU8DOzbcz5moHp6sEY
lke5cAoCTWeD+fI7vD3lfIyWQFguRGRYAQBXg1D+TcZte9Wdl2H7clQJMa0GJUKB
Yvke8RMLGghjfy/CcJMK5vJUTo8vbP7Whbl4UiSitZXrPBTQuhF9NNLcxwDG64xB
cMUhmgM1z5V+0WFmwcckzTTckYFp77JqoilgiLryyUvoxkBiYGlZphCPPzS/bKyu
rt1bZsVoFHLtLiqc4Mv1UNxaS8WpOwh2QSdj2G22Bn+KlRXFQ8BY+q5KjO2pVDfd
68wamiYoazZm8pwfh0IBLK26Cnu5aX12rqKCw3nW2NslJxR2Y0Pl/kNUJBcXr5cz
mYioM6VsCkc5i3Ahs4KuqA/7D9sSt4/SRnEXsBdBUv4XX7j1WpleBa/IiEsN0fJE
uj+cAobor5s/UkOoPD8/05YGQora7zfyF31Jo+akIOxrqhOqCzdGwJng4fYU9NNS
4zlTfE+LikVuaAtF44TSm2b8N4cVf39eNp2wbs5+7Be4wnEFVAN/fSX1bU66lScF
S9tor3k+0oUcPO+oEtJVp0gnr13pcwAEdONcDnXCdl5wkd6ASRNROtKFkxp2V1Ov
N7g1Ns8Wo1GCPKTtLeSLJ66r4BSF3wEQi6byB1924miXfvsliJPmeWL41QtXYewd
6QatEaXFhQPs+9Muv9l+uGyW0uZIXKwStqB9x79uc1bh1LCYK2X1aEaPw1kA81Tw
FLpdO/FWXhDMAuIcU4SNN6BipUKp8eRSCT/rmJnhiYTk3puuuaVyfB/36LUA9Urz
xP0CymwsH9RIIi2sn2v5YzwAxhB2tmNgMkJyrycOgwiLC0FdUkE3iSHfC3Y3Lsfj
jZQdO45AdkW1mZ77GYxml19zW94oAQXLJdO9/Ot0EeE+Yei22i1IW8prYI9ngKd4
f4dvgv7ndEgS60E8BcOu8IrvraUsxzLo2GeE9WxoiZL7z7OwP4aBhHwMgX5eXeVF
UVIG5H3xgeTJ1VIjy5XWdGS8Pu1c19ayBqfRp9h4bSabxDGLUcGqBOIqjfLqdFwx
p5prFMzTjDa7ZyDQjpiwWjXt0PVkUTya4oA/rcQN3HmqpJZyEcBZCUKVsxnNPz3K
MBmWPGShCZwl+XnMe/Ynq1Lf+tCAPPOE6mZw2r8qt256qXJ69D8zSLvBgXwUpTl6
6fgBtY3D3u90VC7xjgneRVZKab9KgGGLRh37OJk7Z6FOUdd/tRdacpVVLOm/GZYF
Gjcpi9pVDbmoU4XaALbTcQUmt5yUu/C441xEvcX8aot5MmUWfjY1a1AiI62Xz+8B
lqW3P7OmFQqgSYsrRFdifYw1JmlXle+Liw7oCfeEpO79lDVGtCiGFVN8caa7ZK0u
gZCm8YBSQODfz2peBw3ZJJZYq5lrTYWQGftJtfIbBNabGrNQEThrWlyYya75cCHg
cuSrUp9fxwcuWaLVP3BC49dEBEViISgeLIZJOQTAQAStjWtyL+yH3Iu8+Sa4YF41
NgWW80ey4dhBANtSyyGZ9/IqiMKuinxqhoPxuw4zj7fDMAkhVbtq/D6kSkbn7dQg
2R3KuvCCqFDGSlyNvWOzYqtXAVqgOdAkuCrLR73+iBRFFVLxom08Uta0++uinSPd
ZNhmAJoXuzYsTfbY35VpCuoBXL0EgXmwaK7O9gaCNkRpNvUDqShaJGeKp6vAI5TT
75YVUwqIKljyxYvtj8H9qxgcLWNhrEOYK87R665UlaXc+rIMpho9j8zs+5MflDQl
QsmDAJILhi42PSDuDcDtPLwu0G5Tpjm+ZNF5D+lDK/d3H42i/i7b9Zw3NN5Tm9HI
GJL9+SeSGZSa0fa/PER1GDtXRahk5v/k8z0sAqlqKM582iDjK8FCtWTot8gAn++W
pesfuk4q8k20OKlH2sBs7hJnlS9fwvyv9JGSLndARz95ZdwTD1GrTueEunXpFNWM
48AC537d15fsiuwIG+OMm0dIiSl3n8WdqKR6hzlxVxu9hqRwsQSV1tjmsOZ4c7Rf
VBvLqDcpY5ZgxNO4Ja/zxFIDaxfIlgjW2nQyDxZNp6+dKUuegQcQ2xpPIRvHkp5W
cKn6LFcLAYWUF94lJMScCZ/qQc1NmgsvyamAD3elw1l9hxJgMKKQi0ixsQ2pUkls
KowKTGuRW1SNS4YPfaTY0ovuudnD3mYOM3WOytgww48EaZxdI6Eqi/MKFv2T2BTZ
DBUO8XFoWYQ3uQvGiUlFoPAjgsOiJXokzfOugaV/Sm2xkShnsQ82pDZdPvCtqrzG
yo/XnYuGs0ooxTAWKpvr6X9K+zAf8/34mdWFMo1rQQo5me2kbtziGHrMrj+0hinU
tj/yOITaqvoY9x7jR+1hiFyuOOVh4OQ9Cka84S39PfbzSs2We9XPyEaT9TqVZ9Zo
Fn9SMrhIL1jihPdm+fyZANhRrKJAJpYnyH1wEJzXeZ4dTxJ3AhJaZ5qbTuR6hoeP
4KI96Z8Ruk62FK8zMrflrsQbeHO5KxV7FnXadNRy+Fk7auPGdocy3w3ovDyje2jt
2lPMcBpVyFyGbXOjl3QCbCGOL+LP6/2VQrZMGobQGUT0bgIUkuJM3OEnxIf+EkbR
E/A747JNPXG0QxKGPIIGEv9gjNg2YXkTn7s1xUoaVl+EdmSRzVx75K68WSkQO/2D
3O92vfxZRRZ4ldE49KNNiyG4NBpVqatmoIIHDIssPum9u2huacPvEpDhQDAV7e4x
ntaUoT1FBREJZn20yghLc2ljks7pP2u6GPtZa7dT7wc8GnhcyNSq93aCEDUdkXwy
2SUqx4l7WRkoBJwhtPHpn0RyeR2+Zl9jWoYPTzd0VLw7zUMg/9BGO337DlkirttK
BsrBmD+kRxVZW8L02Sj3B/CdanYnLOgqM6fZJPF9/dStDRPD65JCI76PUJcPkAsO
Qs388BTb5N46TTkWG278qJWUsqVPVswx834UcSS+ZN2wb7hD0/QfejZhRz4ZUm/p
POJF3+XCjXqJuYoe8j2+bheVu7da6gwyLgRT6QhYZXDE1bM0JAehpV7Jz7sciiPA
ne/QnFeGbYQevx2GM7ffGYwN6BKEehDTXWqnahirfhd8rDGxTYNpPCTunhjKoplj
YOA0iub+cv5Cm6iNkAnnuD6eK09S3ldei2Gef+GIv8DYp13IBVy6Eyr9cxMGB3oL
YKnS2mZWhighqdhWMrb0hHvqpEiDsGgDakygqTru+cyG+embQTP8eCYZ75wRVDqD
OfDnNnermauXtc2TGNB93reAZwC+8bO9jm9uoC8ETSnO+CX3AU6CQkxtDaYOHvNi
JnzbgKwiC3XaqWQgiM4AioKfbbgz8vudXGK09YRLnPzx/qJnK/g+c+Xqd+8eAVay
tIXo17pw8pyCG8+iWNuMiDYspMwVDwh3O/DaSvRuWcT+sZtQGuhqDzI4P4yI1ga7
JYRGhM8qexw2AM3IFkE3j+TC0rXwK8/PIBssK7pLeGjtZqRbvUNk1R+/UGUa+8pn
cNLVw2Bm/aBshu3tzMjbuyLvG3GlHrE5FgBTxq4JEBJT/0AQkaZl6UzcR8X4ZAJq
OMcjI9SiETI1s+VlvyMogjb/OabXkjzxOOGVMNvn68L4EYtEiOuTPVo6XU/V2LTJ
yRKpg0E8dONBl/NPb/TqiKdvaOfpxkzTzdBDNfy08xgdOgkgIokJQ0gLAa2FHbd7
xGSYXnrufTSeARtAtcDO/oW1VmiDmBEwJeoOA9avHMfXgiNRv5dLNoCacU5uIc8e
a452t96gnR+rrRod25nxliv5atXVYCfUk4Ow2U3E24mm77Q/o0BfJi5vaz9xk/py
t6H1XPoWYIvXqFsT6S8u78Ae9ptdyVBuQJ+adkyXvpDzM17/T8u+mI+EjLx+J4wq
RV8uolkriH7+Wg1VLTXMDHYoLom00Ixl7etUsJ9Zl+BOSpOBwLT+EWaoOMN7FBnT
84cZ/rdyu/UKy54fnVx6leeoYxP6BGwBUZ+qWxbSniO1FPA3SZvZvlRC6e2WgcO8
nzbRdm/H5DCVex+EOrLIor1Ds7Ht3BriQeXdnO0jcj1LJOG6PHs4j7RRrUhKGf71
Yxmt+RSz+jEGRoA16ME7ctPy4SY/t+IEAqZ4pxzfqhI3U3PCxS59aOLKkUZeRQlx
h/w/2I5O+3HKROPEIIAaROpdZEQln747hwSgaO9MZXa7pNah4n3bePdXUl/IVODL
jQOHrxMwj+Zxg3ky1Iuxigg93EanSmbcMSDNx+nAd+LZ0oJLW+cZbEldLoAfdUDG
LDvozL+qE+RC6TtGYp7D49DXRt6IfdCzXLwn5f72WjusTYjmaMWUylHIQX1NGDNP
uhP3EaJFj2vDYsighqLSd+9wRfZyBx1IEy9iuhUn91gQg24ZVHVJYRVS1U89mlGT
jI4R5Hqunb764GnEcbUom99t6FWdkwhX3ZGRVW83NifiHwaU1PCWtDbdmRN9FRt2
QvtbpCwifQoIHdIe7vat3mSzKlOdr2DHyU0nL38JQ8ZHxcFmuAAEQd7176BVUcF5
FUMb4//n9oejCw9myYJOG4rui77P/WPiVgaebE/hFbyTzw3leoVzRikdeqbUnUx2
X/EnHgO8vZvVWOiw0ka/b1bDWVGYqQCV39sO1tc38xWec9GWMAbnwudyGved3w8r
fW/5NqwZMc4gfYoM6a7e3bL4KPD0DLaWPmlblDnUiT36h0Dy6q4FYlV9pp38SVb6
3clTo9RN9AfZkJQ0FUU/TDMO7ErLvDFfmQrWJNiRmpMn1czPlh3cLqSG66AmgTS7
qESf9W6zlFsp/NnfwOsYEi39xJQmpNYBY6IcabD7QMGC9C3x3P1yyp3CZ2i1Oho0
3gbHtXM49cO6t4MgvMgHrnfe0mm6KZty/ynA0gZ+nLOt1qYEtNxvI9HgdRv12H/d
oAMmllZsFrfQB+v8tiANPjtYQKQFgZTpchQ4gci2R/3XivHjf0Aou6KQ1Ou9DD4k
K9Zqcff08duGpttfKoMru/6NpRjgfXvgi3kqHSMeuvm6hIQKrohuSaET2/pFx3ZV
ZR7vShvh1sJJLrWalzGjMLOi3zrAs5hO1s5TEhNY54P19zYe7z0UoMyX5uH+TAWX
efBSnyIo3ufSZGgdryjCD+gBdN/75cr6xwl0poHd2ZcBgLR0NzxOhPiSLGmTGB/8
MnucBZTtY1mW+abIJyO7cDOm08pdEoK1FLRHlQWrQW0CsYQHLrm6zaPlC8+g8QMs
chgO9ProTHRl2BD8+VMPux1dTUJ/ogYcDwLNEuV434KodbdmB4XwH6JTsU3R5Ety
eLYBMUuwZ6hRj3Tk2hf26p+3chexwsVJYHEBhW9z+czhquaVCHEa1BJbTbNuo93O
POs0QbK8slTH9MNxkW845XjfdmkI9I3f+YJDijNFQZ61t+yjYa77EF0/29xZz/gy
RLjutIpkJ9gyjt9L3/MpYKekoWjtmw/6iZeBo3rlDMy84bTgmw7ctRhj23AdA7Mp
hyIn3rROqSGN4jAmFtjHMpf1u4j4Gi/7CG8a14y2eqcrHFLlQauSHWPm09nQUDCD
HCBELMPGRQii7mVBgYwhsWKYyT6BlsM8TXQXxwCRA/r0GbiCwXPMR2w1Vs1gkoXN
h1KtDkarreikDkFMCTa0YIyIi3ZM2Y8o7Mnd9kMA2U6BlWm4KtAZM00xhgt2mZ4z
WUB19MDgrIMf3ZgsKbCdziakZpzHoQBY3DlGgnxWKZFHPKr4aX7Ap6MjZT3+Lrie
wqxNXAjha4416OO1lU4dJyYnz36KV8DyR/KnVYS3aPjJoYxDgp3JSTFKcjfrfs6V
k1O2BNgI1YZ/RVQQkUP1Hh36PwPcC9SLkmqpu3v55UMVGF2yV+uQtJ7ONBX21quN
AaRHdWVvz2t8DwQdt1NjVbJ5cCzTaNckM5XPeD/5Z5vQQhUPGWbjDI/jqq6vPlEM
R12HItqX51krPLWkG+ObZyUg7C3u3dFf7Yo0Fn6HaOcA3kBadQ1/vqVIMvRG292g
mpdZB3iEiwozJSlW19HY7Fw0PIGtXg8FfESQEqAkrSZkajmeGba+gc6UHgXGlySW
K9YaSfwrbZOprUv2V8pFtfRfgkWovOe9XZ6NNJnwRoczP8z97kyxKMbGeZNwCb1n
/sa5nXuESN5Q+1aahJ6yM5dhIiyagA9YrBOFbpShuaarONc56cWn1dIe5dVXyicb
oaPcXjxFecVqv2CwchZvLStOG4piX9I6c6EKVGIeM8WtSJ3N3uwUCdzLzZSk/RkA
XThufcV+wh0MU2rFBHG45SjC27TnNQDHjIUuhRFO+hK4iGcBOfdVOXRqMZpy3djt
SdAKZgf8mEBLqxy+UFPTDQKPBukS4R6U2J79qONoVUhNSUYvYuY4IhrIs5VVEAHH
wopy/vFb30/x2v31JUQrBCJ07n1ZL5jY61VfMdqLuQn6Zxix2grpAQ0OJR6ReRRt
xRpnYpnpQ/30A1LH7q3CP/Wsr13uxI01ZASHQG+JyFqUtfMzislJysT3PRMqyaH3
nLpC/P2VbSUFJo1s4D8aK6f4AqmqkAx4FakJL92MpzWBd33sXbqrX84DVeAYKfX3
N5eG4iIMDh/iNWGGryt3JI7AeLNOhssJVLuD8X/2TpgJOYNH3xIxLdyoTKX0CLTv
7xkOnuS44v+I/hvELnUpEjwg5HAecsZp+kJ0cFtftpsvgiE07v+F1mvOvRX7QVHS
Elql8a2W9oJktTpHvLwIUva3PPYW2F5bIQq0gJHD7DHI3SGatSMBq/ElCouPC3sr
4d8HsmADR8ZPj2L5v1Rl8pdezsFlHDVbUBYr+XafxBEipH8ndtxLE8nqGEk0Lo39
Ym9r7XS6EmUuAKVw2nHNburJQhX2oQR1V11TEPeU5Au+C0t5ExWgs3VVNF1+oeTV
x//wSyDMg7ym0Is0ceUgrUnscoK3zIT6n9anlgaibJYnc+Hyd7XGRUyy5lGO8+hD
hXwP+24hEKDy3xhnAhh5cZo4qGhjds9ooeQCino+nzfQ4ZwyfDpplT6XtDub6CRg
emS37SIBd6dmRRddOGBFvr+mdTGma4lRlg4GeVRUxNFaJn5IvnwFoeOmSFGeXGWf
MqqSYfbaCV1nj9ozDuFJ9dcSH3HikQIhAdM6mQxJDoYDQJ17vtI5Z5pC741oe89F
Eyj3gELq7AAkAws708FCiSzSGLI7KLd8DyEMhppQ7B+iixZOFbrLddoI3TN8bxvP
5X965MuBX5mBarckal4CLXjQfS8PI4M0yoEJdy1HHbfgXFlZdbt/Ha2s69cGSFWE
p0jz+cq++YiFCRYuKbZlI+DixMRPGiMSsprIeCHuqKP8BE8c9/FXTdilGE/tT8xf
2ouPDriUlNldRg1n71TpN3MTDDNXyJjGbJhbIroFNfl0FhV1L+C2SAGY3gNA3jwH
FpMOsMBN08DxWk8cx/RvWD4Og/pRwtObaedOMnCFTiTi4GgaM1h6P35Bqp5jSi6Q
J+CZHha9dsvmdbCNsYs3a6TUeUmI3locGIh4+0LVU9wT/pes5jQmbiPkHViibBNy
oCnf2oS3w+108I/i8m3XhoNKBeI+AcWtV2tpIkmTZB2JhbddCcdh9mBuzULugEar
4Zwpz1OjQuonQfcn4rpZVZZ4bsviAUsnTnkriz33vgn7RykgzfC4sj8/5R1JgAnu
JksrOV5c6EUnxdwRfoD9ljoHq3a23EuIKzgTnjMwV2rMW2HmnT3WvfdOugBknBG4
PU5ZWKv/5e7puYbowmnBeFZhMr6XO31omGTszyakq/IWK14OFvAp6k7gZT7RLvVt
9HAkE3jl8oRWm22Sj3IyT4RQ6pvZbVhUhz7DrpuZdBmAP8ph38OHVYS3uWOyI8/T
fyVgZ6MkXdhV0Dt2l916GkKdg73G2hEPx2CmjR02IWT+2C7+GuClwxJ7s+KnDPcg
M+tR/Rpce5J1x1PNwkuHl4vfXA9xhZyBlzx6XGJ+J4LRdt7Z2AlQXsmPZn+vHsJ6
I1KR8U9uOwo8X4+Pe+ljjbdtbXSP5T+9Ckch1N+3Mbt9HgEVvmS5UqjoLHqWNDqr
iSBh0NeBpjWctAql2YRCvcHejVGDUl/l0iCJaIvXdj0OpiYFBrWh5LRnuEG1nnmB
M1y6goVsGhCHTunLH4HAN2/XW1fhwRqtbqBbtuz3salaww4xBbu0iEtoehpjcUL9
JTBNY1Kj/htkMwDtA2aHDR/FsgKs7kkIlWsgI0nEwSd/HEq+LEPoF5ZM1UPO7u5K
Bbap9IqTcYR5iOP6mN/PRVziZlcWyRuSlG0/JwGmRr1NMWehLXFSX5qbcsjWSspn
nILjOdpBCKO+vKFG1yEtj5+G1dMXO8F/py3nFkZ0tVwWv/v2tppMXC2RKMYJqJA5
Yo38bsoT3BdBu3wfPEWuQB3ax6dzl+TBjNidyz4MggCfxPQZ4Yc7ssL5Ml+3o0+r
8WAM6mUh6FrzkP1z5DX05VuHAsFeojXlGtj6huUpjwhxUNz6EjKfVHtdUeox1/1U
BQXAK9oLQ2/E7Ltfa7zjwR2xeIGk7epwqzK0y8TfCsF5TlPZKo1pEsgdlctiLRQz
Ewa5GjWK9rITPX5BmqsAoEEyBYsqmLYs+Dh43kvxBBt1fpLDaHyofdYa8mR/Jirs
1Kx2n+EcWG1SsvNQVmJk/sX/IQwjk/OMx6lbAmecyuy5G5JXDp3l+GnMH92+oKm4
lwygS3pTnkOfcHD7lrefZbG4nHCltdLGZTX6Zxy4aRimvld+0rd2lUtb5wmaOQ81
wC1gYHPXrUJTakh5S2OUCP+EqBJhkxZs8DKbUtkX3YuvZCsllon9r4pJ52XaRfCg
BsQOgHEiVBO9suxOpBHG8hv7wIJncJrzwZk9p8IyQ2vJeImtWTIjjXhe44FVQ1Ui
1GA9GoHfR3yjm123pR6J3pOipEybxBZbVDyaWNe3V5fgwxKkg1SvKPEByM6KTcXl
yMS+o/METjcAfl/LE8avYj1IGicH4wuRQlp7SL8fV7zqP42vvI+BRr8LWxf9QpJw
pQ7S9V06NNm3FvWIvI/QqFN0vP7JYZVQ9MVmBE7+T8OCYtGD5/dC9kGA7i1ibAxp
3Mlm2XPp4iBxpdVNEyBRggXy+5vjk+f2vlLrXgm9eEJ6QBskeE2M32e8xDq2Vhex
0cvzqUqdt2EuAWDsETfvoddpah9c38C1jw9t2KBKVVB6GhrnId//EklvfvPjXuZi
FALRwvD4YlrWq53VYFWXEqsNAC7fZvMFQOjTCohi6GpndSfzRngJI4OsdzzcTQQT
xICNpDh7EvRkNE5aphuHOC7pL06QEkRrsrLfd61sna0fIx46SyuAkzKWZolxcKcP
fU47IrQUOCC1GhVoIqiOVTKx36LkzWxqL1EaMRHrd1hH4cl6fMzeuvtTbhCfSoIl
NpY9OCmOrs3vsgif48Kvvdz/Fei3ZCMeQzHD8zOAK57RMzPinDn7/k3U4orvfqUt
te9olD9KAAU9r0o8buKSwy+zw5fYyQPSaZJtT1vKZqMcAH9npox8wz8eI1DeslDc
jklov9RJgYZChKZ4TWXgujX6VrvZT9jDhbTpaPd/xbD/G4d4xlkOq/Ho8aEpNLjU
g3o6yf9ylbZgA38/M+bF1zq7ovNNT+5D6JkN33IS0Ty/T9k0jrEvX2e5CF5NbK26
7yx6yp1e9GAApGQ1fB/ORjFdgs0IKwBHs9oO47urRKjlssPp5VAgsFqyTxPIprlZ
MO9rsCmIyFISFYF82ot/zqD7NOCWvbZAYvvAYdD3dbb7Z1rTkcjm1zVcCICXZyoq
A5dK50hKzFNGk+G7KwjgSg0BT88JMKqMA4Nzf3LOvsAgOQYSJHRTNn7r05Fr+32E
67VwNjQfBSxuVoXQ/orekw6FhJNGQofxiTSb23x+OFr/mdKcvnKP+RjsOkvBGJjo
ZrBPVI9vx8xwoy1Ie1msAefDKJlwNKfcP84v+iyb2tr8dgauqcMedU2gg89vpKYw
8PI7iSlmGaoi01Bh5hRLvjP5+gY1jDqt8yWWlzeJskfu6X6J3bEpsUAngH60KIdh
2v0/cIxGUuJ8O5qAZjFEbv8cZA/1XJEMuV7Dw6+xtYlcTeKCHUqGMrqJMfY/kyup
geY6/YxC+sF/Gae7sdNgjw/QnPr+nzztHUiQku6WPMW5fJmPRzfwsRwKrN+/HdBn
XhFQyEpc1A1Eg5/57vCA1XM6mWCBbWhMBOBYbC5EXSh54cJFip41MPA5bbnrHwMG
4M7guncjdBy3B6FtuRdYXD3RZeufbQLj1CVx9uLvjeZjSzohR0Jx10asu/zh1OMq
WIfR5mFMHvMXD9bmOIxyyIbBoNxPrCmccRIvas+pTgHxnrA5MPe8Hj5L5rX+na8v
qtKPgV3uS94Tomln0BUbVNS9OgPxVjlsibe5nlSwfL2DDg8fOrLv+ZsuPCk1HBTi
IarGepe3B4syzlxacgTlwgU57EaCmmYJiEOl2yUy/aPmcZCyfZAAX76HJPmzNiox
RjVFgtbY1FlZ4ylwx4I+jrEwiP2VdPfsSw80CB4aDkG68bdk4CG2mZAvkp9ymc1y
d8KKTwdLzTHkjbwwf9vERaUtq2a55D9kKQYrmD8Tp4LmNbZNtAHrSQiv46a6qzIW
AxC5vh/9vOkkL9wKabYSnGHaj15k+XfwKlICjmsCfLk2dteH2pF2jC6x8xQgzJQy
60AERDxb6IMEnqsFNug/bGIbY7qJoeE5tGSEsiNkbwZpDcmJfx4bEgQHF0sxVvND
D1B3/sVA9LjMtXhSKQuy/y3buW6icjrQAeNeEkIjVYlQ753sbsK5leJ84ghpCFNx
vuVgL3wr6CHNJJFI4fFNmavO/I2FgM6Ovw2eu3mNk88/ensDUgNYstVb3Leq7leG
jGwdoKBE1ZL/xFtWYjgT5OQ8gRn340fEGJps0pT0fCCnpEclxDxWatYIiNRyg+TB
BaV7TW+w2lYQwJVEbSivHJE3gtdVtMQnuFhWHenEfr+FAeglTblwHmK+OrE7az4u
ODGMx42QT9hQuodB/lA+SF44t7ILxMuaMhqAWFQFZU9+mL9ycY3dg6RTCx8qJQmt
SdcCRlXCwD6dCeHrwrqWbhqjpkh/akBbdyz3OoxdZomJ26SIa7F59cCkElFEq37J
6Kh53Xc1z1TRwFvWKd9VLfiGWwC0SIAkp4uUCxf2EpMn4fYNs6TVSxriu8GCEB5h
FmYh0vqrcrnyxSDdauXJ1LpXlbsNFQ4Wh36LbrG3uyF1xWxUVgKDY9FsIHdCYTCB
QoksKzHXXrxXsStXV2j9L/KZblHRKj8ajgttUpBgatMBBH+Mo22Kir6z0rNgAz/Q
N0qrcjLu5xrjzBLZ3mxInYEAAnth7AgawDLQOoTU6DFK3f4vgWs0x/tvlz+Dva9P
qcxWXpBdexjsWNiO8CqSbE3FHFx0xmbi6i568EColI3RE2u0NQUtcRFW8IEQ5vOh
owzWDsAAGxf01erz6b3VI8YZx1GXLOjXuHa1DuuXb0vbY3Jaxd9GQ96ZMcDRjSJT
Kx1jn1PoIibfgIIDclZ97uxglDd9jqv6xr+BnT4AetElm9R8ifxe4j0LWMAvDOy9
4acfsMXx+MlnFoHrMZqD3amPqamsBSxxXhZjeGT0A2PNsYEA6JvHulhiII3qB0Oi
5PP1qERFyJQYklVWnmbLu6g+iRX/M7Bos+lvuMGAIK4n8+kXgsrKTURtT4MTRQQx
QqipLMn76bsMAnf+caec46ZrP/dlsM2eorAXa4KeAO2RTs6TdX9f/YodyVYNvWN4
OiRV7Yp99dCQ1wXRwm523vONCI4hPkf+xvc8Wye3niWgXGTxwZil6R4AMng2uOKV
nY9QVnC7MNAhnN6TFzRKiCQzutzQREBDlNB5zFbAju+Bn4whFxnl7BrqBUoxbEkz
BqKU+nIYDldhMsWkan1bfEPxfZWT7Szcqjbh/VM13m5R/gso0x7ltod873crb3eQ
i4K/VnopHqlpe1hJQueHIoy2KqIyyAn3Eer0zbbP9QHNkz83ZWdKrF/Do6giBJv9
urGGDL1gZlMrBDtlp3Jrxli9ha7FOBUUgFGs69BKI1cvQyz1YfQ4mRqn1l+rsGlC
HzBYsF69aOKR9YHzjaRQejQqGxqmTu6Kaohd0q9SN/9AeaPh1he9lhFd0Pk1Ow8L
ykftAO8/yGZRbF5AAlYcNmjHJfGKd8Ut+unwGPp6FTQQN9OXt7p+y4cYitUQLzVA
2rBzlUr8b0u3TE8nZ6e06NVHtaMQJnYeEJYzuFY+sXx5O/CoSO3wopJ2nPDibFW6
rODBfyhU3qeeGNwSZ9dHZSNcqBObSOfWLG4W6IWn79+5aBRPxiALyHMx6NInm15K
AA1eFslzvEIWkX5fQt3ndt8BEXElQeA4ntOPXX2wqmU5jcBFLKbgV3dUErsReP9O
ZQfYPjgmUUKuPfoiwi8U55WKb36QBza+m+ENvM0Ey4Le4p9C1R+w+MLPgQwQVkYj
fd+di7d+z7STHwtIYOs8knUV4oEQmuAe9HjZeCvisYx3nll6unBPFsx3s/l2SS+N
NVLH9vpfLlSdYbizpvZMGBKPQz+o+H3ykwz4+gS2qZColL/XYh6VAR+i7JCBZ5g6
AwFEiyY6fR8u/YkVyPNxA3XqJSpRueJqnJCn8Lhs0EzX1oKa50OY0eErO4KfFu0p
rjnjjGdqKvBQzEcQ2+cpRuSz2B3+YgZD541yE6n1ikvm9Res4kl2ExaYo6kFNYZ9
NJTDNTFsiHEOBPboMtmLAMSs8odO0S0qGzyIMIyV8CU/ozbWPL37Z4dliH/e7ABT
EJzYO+Q/gWcifSBlThf32kD5Lu5YrfOyFblwryAnKtgPgftnnN724tOtVzeddAqM
KRi4+xd0Pz9ZnBIF9sVeHee06Vx40lnr1l9PeXodKwJ03eDv66R4oRHrb7hPQXMc
UelvUdL6b7a5oTqqPWW8hB8pxHvz0496KN1iElYjSzBMWXsufqhYYN5jpj0VWEDH
QEa+N/T/1jNnMKteeKyb4LRQrwbUw8IIp4R0LrHTSX0m9sR8kxmSOZkiscac06NC
vgSvoC0ohdfNtXqkzST49ap22zMNYn+Y5f6iq5vWBqnCapyr2Lfu/dgbB46evGDA
1yMZdIy3KBowWYvxH6nrwaYXy8pMzi8ZKDdig+Kx9dnaasnpC+a10e1ELHidjYds
j6MVkHsonofw8qq+qANPNz4pDTdfVemt7n1AXUfpoBOIqKfVvNCeJMGXiduP7WFJ
lspIJQgnkgig2IspHGf0/TmmFewK2STI+kAE7ciwQyyI7pSkaLhgPLKZuKjJ/KHr
9chj85VoIzEr3D80ZabEXifBZH1tqVTcTcCecqmQPkDbhH2FguCVFimUGi9x17cE
xxQKUPrRzKmQzJ4kXR/gOK4hTcT8oPQ0bo+QNl6vgs2GCAb3kfaRqHZAL4eYtGas
Af7DwEKPbLp7X/Qgq2ZgzECUR2yNWj4NOyGAkP5KK/MiXtnKOY4tW/i3gwmIvF0U
+9gxWcfxfZlI8bU8dc6Q5SbxzWJv15TqqY/Uta9DVPmuZvQHZxQfZDBZweJLmBC2
lAPHa/PQe15kbE9p/yvEP8IXUwWH80M8ysT124Unb8x6NFsgZS1M/hxm1sHHO80r
pEN02EH9xmmWM7McPsB2IxXmHpDFb0W7HI7L418cuYRjivTMy6wuccA/ng8IF0lY
GeGuPPXpENV3bVbN+Cs6zUoCbD2y28yE3MF1Cnt5kMeJ7osN9LVmpDdRgnK2bACA
A32aT9IrPVjI4VegGkdQXpiiHOrmL7afK+uqJr1IWWU5VmwIRRBeUZ7uhpeKbSWg
I5oEiRSC2shuUqgDZFpS3jdCpeMRIx7rNKkARiyQ7tIt3cUQxS1Fts+XytieoDeL
orOqfQlp9WvJrd1DhAS+YSWtKNPeis7hzjROxIHQSRaMRdLduT8O5PvGrCZQOSf7
R86/QJZdO6Aw2dqiHMuC2DzwcJgz8Vey/+I/oWwf4joHOEKxMm5o/4V8luwogN6H
lJfKYfezJ276iKXFnkPoBQNCjKCWVQXpsOG/brOxoeUci34PJYqiTmLTfW04Mtfq
u+O6gNKOh8Y7PKSsXuTFv46sTiQn40bzc/Ww4Zd/YXbxtAs4lnpwUuksNjnj5lYJ
QgUDYHUMlqSW0NWfH3BAGKCUfXclPVF/aEi1AalJt/AzDmbxlJTxH9h9t4Q/rlLn
pOIFQnQqwnSk/0AWreY1rtYgBJdXXl6dr0kA1KVB1S6WuJegeCWJdoi3Mmkld1eM
2mCTKQfMBlxdNAUHX5LTldoGPYXbBs3LoCo+471SO7g8aRswuNDNAmcXyIzYaF2E
I6g56tI22HSVneuyInmq1xHmedfhM8JHCz4UWwEWxUZLrqRXlpksHi48pD2RLRqR
KCxX+SMpqyU3nKSYqu4umRmPokX/6CDxj47AcYbAAJg7dKDP2KeUAJ5dZw9WyU1p
aknUeoF0djgchUmDHISaFWinrYAQUIrtYCAb5LjTviPJ3qQu7b70YeiCBj9ciBFi
WPw57i0LvqS8Jq+DPVUQFbXXc8SPBuWW2habwoNDXx9sKMlqxM1mAsu7ipBnV9+n
dyv3VKTK2rQryUWVCCykPHOhUzKXmS7mXZlofRM7OrjZdFYseifaKFnOsy+Gaqz9
tgdeDD4gR6VaUFh7nxnbxF5IRwZYX0jAJUY+YdbWL1/IluwcId6fimJdB6A+d6ZZ
jiJzFUr36Q7a++e3PbGKSyFVKp2IEoeYooCLfVQ5kB1x1omj5DbRffsK0cjCcFrp
iaa5F/RVEvdxleo/kZ2ojmMEeudLFJyzxk0aUXg0lCl5M204sBgFg6ngah/r2GXx
0OX+zZXmxH/Ql7LGnhipljWFknfhsiwsgmYBal7F919BEnMhKLVaEY4nhSm/senk
7TGImFq0aVQ2QNQ5G6GUXfFP4MbDwvzgZw3ojK5O0fR6S3IkRNNjxfx5Nmroem2O
xUu2RdcxT2ls4B47gb2m+JxqnURhzPTbeLXWdUEYP2XS+ar7VYLOnlE5V2ACpd6T
sPAmxv94/rELcBkreZRiS1vhY46FpJ08QY8b0svbGPCC3m7Bt8iv3EARNzrOY2G5
x2d3NzQkhCcKCjvfXOqjVLxsJEgjnnTFglQkum2rgjyifyf+aobI6RrSymE1Kkne
qBnB2YXwcOhHYO0VgFB1+WG+IX4tugxO9rl2inZblogaW5Wg6I849n4+eFCScL7z
ZU1zE3HMMsYQxOOsVX1JGyjIFivk8tIj7s8r3V/lQqRippdRwbDAsz88nHt3oSHL
fiAjeC4W6ahwDcTj95WXjnD43ChxtNGtTxb7rJNftHXkCnS+n8IJsTEl7HZtuSy+
HkyLXDzJN6CJFApdG4jyj702eJXpRfaWMLEd5aisp9N/LE0FfGYD9i0bTIKvRFja
xqdbezqjAPEIIaPVDEtQnFkNMHcvr+COTHnrwR1Dgmsh+ST96KusnMUG51CJzf9b
iAKPK1pjVvV/PutyQsVFynsCY5WRNlMTVUwi2aIHSK+9Mjy6OLlSBkv8Y77USvMZ
p6PBpKZa7huJolYKJmWIUNCh5+0Mdz896bG3tMyF5cIuKK9dsOhro/FxipTzjEO7
pAoNDYObTq3sQ76K1NfcNRXP4Orecj08q4YRgNPcO4FgsCExAPFa6nBJD8n+9uwl
Mh2PW93Wvk/ildThJxa0ZloIpcuMwp1uc9arKw4nq7ksz6D5oqGBtwR9dM+vtS0h
K2VbCiVfSnIKzHtGxLFI+z1aTS5Miv4zS7enMEKMuDA4amGQH6V+j+zkGcwYMH6z
lb4cXV52MhYTG68nNrNBiKx41lF9lILgFpH2K9VdWV8sh2qaPXsuXM0bVw+Basah
2HhhKWkidZVGxVPxRUkBURyOF1tt/twWOZGs9fiShcHamxVCNcYJ/0Tt4eLL7u3W
ambo6XzMI0QqyzhhnvQ5oiIISY6dGEhPs5m75c3fQi1H+sfI8wagy1gkga/fXJws
FHCkpkyGLQsmDLX7sTjPLbqRXD2CrzDSbNSq8FNqZDXaDcn5zVfKGuhUQj2aFuaz
wLJ3cUEndlK+5yJbOl9osrp67m4dF6u43tW2ZuLepB/2RRLZmfJYfRtqSqPlrF6u
sC39FJobWdrNf0GnMAxLCKKwj+S5yT8ShhM8cEMcaqV4qZmQg8WyTr5HPmNTIGGn
iCmgLAPyJmfYhFncOWLLjHrc97QEF6POvsG56eOqNJwQC3jXYZC2j1rFgOXb82LN
UjtMs16my2ENvErHPIE4N5eGfD94GN8nSZbFLr3T4QBGc614OmPZUPP/2A0M00Ax
ie1Pb+QZhbUj17QRPY3DhY2DthetFtNhzrA0zug6ICoiTYfyGmxb1Pzl2v6INuQ0
ZK/sBL4V1VnO4fgZl1Rbwh7YF9lcVeTdVdfpPM98E/IHWDLwnpTeoLojzOB33rvk
hXeI5gbsXHHdtCSKvgAYQY+Vq7L3kZjgRM6zCFps1Zkv1ogNvoKxY5Riybtj28/6
HIGDj3/CT684Lh+ochcnTYoskS+Vn61l/caK80TBKZMTRHXgVaABrNNtRoKGK6/1
MGDeQaD9k6Ry7/++MeC3ds31/By/AEGYZaxnC6gJBd1kRDzNj/piSXyoIuHnpsuA
z3oXJ1WGijLtxUeZUhMvF1dEWYxQo5eT6tUPzJaD7wX8oEZTq75tEg1+izT5WbmD
707BOQPnBe5KWmQeSlFm6DfkWhZd+c8pXjCrO2D5ulOV8mR/Tte15ZbdHtVj2E5E
/U7QOV32LvKyxca9MCShf20vhI9O/Fbu3nessAywMtvKz3G382YrEwWtlrVDbndE
dpTGZ82hhwFIUmoJufh8rTN131XrawItDR2e7Ep2buAqtb5lYEQ1MN+9jGcT4dAx
Ju7DWw8vDAsg2H5jeEprjukY+iyJlFg2WbUlFHaQMHFSJu8NTIGCDnu/xPO63hCV
C7ayXpbpepoCQdO3rhecgPoNyMRp6T2Mcxb2WZ82IbzKSNgQfFIcfaWNKzEVmueJ
Q0rDy+p13ZYdsC8krFfcuoKQoVF/aqxYnEVoztInswVNkzp4RJjeFomi9o99d+CS
HSV13HEEHhHsdpqNwW3JCVtfX8WISr+uZbMZD6DHPZj0d05dqDwLhcjrGBtZ5oKU
LKCF0HAhzmBqqOROsgdnDGXfPwbCTszBWFNNdJ9clBFJOfIYTUoi+UjryYs242sn
R8emadG8VRYZl4A/lphSTytRcV3Z1sx4DXWgeOflZ3VURlWKVPLivaGMPFEXhQk5
jjUlwJDoG2Gx0UMILsHK334AXvfVbZFk7cwGVByBoR/YpFpRa+M3T91TB97DzbdK
45vbYP4OSEnqpCB1g8DP6AUb/zZAsVFUj84DlJaQdedmJn1ea0fyGDzFScBIrdVf
9bSS0rqpSYxIZYUp9dpwUgmbAuhbzRci7oOOqaEC7vH8myhYVQ/kLPnaUJnOhY9G
SkjgfEEfGg0lwxVTuT7sNwBjhs47/fmmnv/a/jDM10bc71gIVThkIlSOhJ888Bad
YMgx2H+YgxESM9Eri0UWPFvW29jnQ51EJ2FcTjpMVERAW9bFBGauVIZ88j7WBJXw
6TsFtTlVIiRDzWxfshjGlsNMPvTY5aGGnkNySRH7IfMimMnWD9S2cIAcHgj8F7zQ
91V872szsu9TNuemqpLZ27VRy4jcsVFidimzfPSw2pI4sk+PeOwPrOCosY7Wo0Va
VAXKK0GQeSaB/TpI2DEG6I1lgpz+7E44tJkiWI+jH1s042TWpzrjNkGPnMz/egpI
BRGGuEqSxIt861S88KmyTYwDkX1GpbZxrdshzbdFNM1ygNHVH95wDusFy0NK9B8p
DPbQgaq1+FAdzox+YPG75gz65pb87v8+ojoUWE7UPA04pwWBjH6KNDzc2KlkFj0Q
RB3U1eQSaiSenT1ZYMQ4fbBuBEWhmN3/ikUYQLR62CErcGz5jKlo3Sq6UuLKV5XO
XKGioeRQBAiCXXiajR9u+K43dsYukIUqfTbgIuzWRft7K0FbjFim0oSTt+ZAocto
RzEEIR58l0q0Qtot6ONw9BD6Yca/ViQo34rrmksv5hrdIIgf1NQ4o+ZqRNpe+fBC
nzU2w8WbC/Ngdzbab9jc+6aXWrzQO4P4PPRrUc/bFRgqM/c/VXoTNimLBZW0IuRr
TiWavIK7mf6kqi1CW3Rb7rAjBdqH0EfOUOmgKprsznIHn3TiWSLQr0kdFeLxjA4H
ujTv/jYU8n2e1Va2JprMuLzwhPsVNvd0ewFoMwzI4CDUV170cZRXqNf0WwWma+xi
B1BHhK1h2BdWQoDvEK0hi5j7mqkTm0B+gcnxYX3nbYGzHi/dbLtPoJJusP87xMil
/5CrUTL8CqoST3q7GjnRzA8LPmp07EmYOnnF7vAk099okVkfYHfcLmiKyFWXrawl
RK2NiWcpCUbXIpNGgCupQrGPA/nuoSTK7OaM1VFy0+UuM1A+4rmMydeK3e5WI2mq
WaJrmYDZ5ooYgNmVof0Tyx9T9qo6aJ3VYvNZTSu+8Xfl0jSKP0snKx5dSLaMIwv+
3vnCRfgTcVUiN3+Z1qaS0GPUU21+/b8sIqqfhkC4eQAiZx+Z5ErJd8Mx+KNSYSED
DO+5kwTsHOK791ePjqjJksjKEm7PfUBZl3kFMDwPm3ZodpZ9HvmAor9+PIkwVtQM
K9iqOCoOqAAm0rbk1WMeN5DsZh3GQ74P6jd5yzzA8m9Voju63o1McPjB+hd2o8ag
6JIaXG571qpU2yJuJdUJlEmXiwAQ+ysKDK8poURs1cnJTGM1bHnC3jyzFC7BDefD
q8G744jOJBo6XsvKjaQ7JuyuOLXSChUd+zDmZTfovUOd0v24obaVTbDIzIVHIvD8
sErmP2gfE3GZ26XSxroyBq6OVltki/YbE/glnG4sGBmwrZvxVauxB6f6rMoJPdxE
Nw8jjOu3dG74hVGhOIv5k0jp7fRjCGQQDDBbooCLCkDF9koVJRWoBX+e8y9HHks7
ODMW7nn3IW4r8ULJOnoCHYSGjocjFjHw3CXFrVQqLA27uv1nub5Uj1gbUPUr1IM/
9z14Nbas1SqCpI33rPLijeUVn8D0jgts99stZz3isokvSliJ1Hxe7CgTZ3+Fr0vV
t2MxLYWs0SaatZrhqxYz6QgS9907a5Y2pWFDhMnRDdGwx/Tb3CzANB/HT4Mtbb1U
TXO4lbDQH30X8oj6M7KdbNUyZCRRBsdHlv+wU4WdqWsy8czOQFkvsEyx3bKYs8pm
7DkJlAtFYOVQFEJ5Vs3sQWwSRNq3ZsbZ2gPj9+Llm/cX0aS+Pt+UK+vdeUMyX/b8
BewerKvUMOuxkFSnQMEEs90FP2BwypqNL59xMKe4BezrYaZnf7xweRKau/NVFc6I
Mru1hMGjjjgWWoRrTUrAkk8PzMdaZ0PD/WK8jK57RBhm4Yt2/o+qJFxQbPCTP9DV
kMwFMN3HPj33RhP7MzZJHE/IVQMscY3rZljOivK0uyMMWMJUVQGaaW4caK82LLDN
ohLn0V+MWTe4PrSw4ibWmmt98c87hC8UwV/vwjZgCWCbVY1g+vYxK6YCivsMYkHh
DjGBXtdeL1C8qDDhiGVhew7Oz/VqozG5D0zwPIHbVqzLxQ6gdOmWomdBkm2TZv2e
1tyCqnVwst+v/b8ZGJdgRz5jz5OiyDwoZ0fS27J+HOzyE8eN2I4nAVwO9QD5f5Hq
S//vbe/YtOf0JRgnEmgqKpHeSqkqqylqwvU5ReFD6RskEGk72kBzQFs410Siy6NZ
zSKtwLGdz8XwML3QC2Id7FeqZaAFYLtpcnewgTxGlRKVu+/Olm+dsn7xTqDIuqSf
TvD0jAjbC5C2ZFu2SqobvrqnTBD7dvG6WWZFbJ48Hl8Z2p1hnf2KXAf/Ql5OEJRY
K9duQyEt5Yi2f7EnUwDHAfvLaYBfyPTYa3XqN5tvZXW4tisbZS8DfNsbKShuHNwB
xW6RFbxGg6SOmdQOY/Ac9MzOJvswPaIgqHVkApuUn0pYY6+UfUjD11Fb3jOSwvJ9
XEyZe5Xv6oVOeTScxp6UCSIFe1k68SDAXTFHrMt1VByWqOgtLUO0kLklt2VN2g5b
mQX8k3J9kNfkyAMQROXgDoFhCdQ1TyVAxE/fDYNk8m+ksvd3MDBOYNQY4BK1frO9
szEdFR9Dqlyn3mU75oROBd02zcCdauwNe3gNyrszZPA5IeeDRgYD+utmaJIkWlZK
5M0bNJF8Z6xfloSLqATf2sdRTWL+KLfg5jLzrp1NhoKIp3HptLS7LU3kat3ktG92
QqPxXmjDgZqYtoWRUlu70dkIXwJzQYVM5c9nI74YuzVlQH4LqSp14PqQtPk/BduJ
lV7gwigK9DEm7L6nFIac+o+dzQb7iQ5eFE6bgePZ8d+uLLTWkY2sj5lRJz+93JCi
5XmbOfNdutjwmu5vd09NIl24FG7LdYJ0gyT5dYhp6WxrwwQiuQEF8eyAjQGMMapv
1RUW92echPYCk2TdLsRQW+K9JuAaxIs5k/3uQAE5/vlsTOD8ZL55UYdjgd0+2L41
0SMehMICMXdLSczTkZGHzCDSzSeAhEyi7q2aBGhpSym+hvFDxDvuXbo8OPvGwyRe
nHEScN4AyewenhK3Tyk33FF1WKficfqXF8raYBS+Q0eeUR/LW5hFN75i5a+lV7M6
k4S/tyaffRg4bjlK2hik8b8F8GCK+OFABpFj7wynZ6/sKMaKOp+5TeUvjdwD63jH
hE6TRN4S3EIwx80fEM8Y6URFD1v+NxYFqJPms/mSaqxAR81d59oJY6bjDUTUuWQx
NIYHsLuVqpz+Vb1QvL+bMUJJrTBj4HUO8SmItV13StcodgpFP+dIhhUctMsInH0u
zKE+VnClck0hwBAEnX3t/6VX41+0cRjrx8kaBZ1Ohqgc4bwpEU5bXEgeFIwtROuk
WUJVGVJCrcBFoc2wgsfEm3HfEPBuZofMw/UF8nksQnRSITXJDPuxKL+5ozS74gYA
l1mQ/z26RcfgreIohESBmNFM7BsV9D379dunB3VJ2zlRBb0UEYSuLg86R8nRp51W
GOBpwWJwk5TelorwZFUmMoFs6JO9WneYlvecrnm63ZzN6V+xDfYwhgLy2vTj/fcb
HaoNUGLW4YMAeq9lnVmVFZoK+10LL/T6fSyCyrznlcM6+eDNjE/hNu0JrAdCUJ9R
8IckEBCs8XrTrGYBKJqjcp2ZLtyXrtG8DI8z3Ssm5/y9FuI9kB2FDryhnZhIL4yX
UTdx7T4tjhf5AXRZ3xf/zNRfLXvh3iJ5Ao1oiQ3nCip/dc9doF2h1eGbH14+Tnfn
LsHPu4Cn6pXPf3iOjza9onPaugxP7qFz92XvfE0VNxe+hAOz/EtnLjbpvZ1qIqDc
CMaNH0ApkL0cAmbiRSPK3xxwZ6aBj8813UI/9XynN0xz5a2uvRBm9yhcVMfpOU/t
tHZk4ARIdcbpjmO4dotCpRuNsg3WJ6yjcAuYrJY9jg90RTRaiJPMO2srehINeRRY
mOwEcslpoBEhE389Pbt//pdVc6B6/6RZ26wHwPnlAQwH28kV48cGbG7P8ILp3xeP
3BUJNkDEfzdATp1csPDwDv69o8tOEdUjwsyh+Nijn5gITZ/JlrTk9Mku/s9kTEWz
KZ8kp9Uwo0obQWsXnxbs7BY+SVRLI6DfDxZAbkPE2cdE8F1fN08Jf/BTYPLh7xfO
7VCiGW8RjPvkHcd3ylDUvYryZTQTtfYRK5IyXCDtd4VT2g1PULj7xUyG0SWgzrB1
czdtj6GcHRwHnx55Pr8Hb5DaLxp8il7mL6TBuyB472Fqa3ElSLXUerlgRU3EiINt
t3S5CIuveESdDSeheZuPUqjSbVVEw1z5vPW/asV1pVau8IbUli77EQGngFZGUWqV
JUSn25TEErY/VxZJDXU6s7o28Ks17/RH1W+zp3OOqqGP4lMxE95Pt8hAy/Dn/3/w
pr83H88f7R09Ndgx38RlJ8cVv7JT/CZ4crx+pTyaQJjboR4rqbQRJNFT9kaeVh4J
XJJYijPqNKsCxIeNIsjn+irprcqePBbDckFB+8Rww7ycNZfZLNFv9VUL5pmKFs4H
K/DQ7Fh5+Wh29MNcz+fKf/ZQypqHJdXXiduTufg2oS+ldoY3gj1fYfnQ32m+Ey+b
zLspbbaVAfX+u9fOviSbZK8RSKYyFbirfPTetW749EHf1nROPPM7OVKqmKlvXGSQ
0iXTFxkkHA8ue/WkaCmjcI+XjmiIYHIT3UrinPeq+rssKAhRCpDCDSc6iTAez1Sp
v359vf9DoWDD+9ZrLgi4P4GuxWeP/a+pr2AfG2it4EhiCR0wZf2wLJ7VtCWYlqYF
xSZfbV1pyl8yS5d2Fd2sOdFIJgv7EkkMUNzpnZUHEixAQN9Kh6ZRnQ8NvW2PB484
+dO5uKPaogsCpUl2DUkLqWt8KEerIiGABluUvmJMhi4394bnqNpeZzib0+Zej16t
LiaqUihQ9Em0DZpHhGHrjlzsbX51ZOP+R/vbiZ0+Fk3PMyEBlJzvfgaVidbLm2tG
qBBvjedMgPlj0431dCD+jbJ+v3EfRVisHFuWX69Nl9Ih86OF1wyWnP/tEq71hn55
EIYOwimBLyOVBO5zJZQ/gW51BF4rNoowmHHyF1HcgT141b+RdnhW0aQwrbnF5Yr5
hn5O4LZcpP/HZlCo3OkBvhe1gwq907V+70MYW19YvhWCYO3nOVVJvZJYVrPaUudh
mFK/rcjfhE+HVa1SbfWBjoDcL8nhVr/Pa9iUgGqxNLOmDJVN3EDWkb+maCRiUufq
szSSv+PjonYgPvKfWKEzX8cUke+0Nd6eHUXg9VOpKDr0Xs/vGpmx/fxx5yXFbBT5
/p4NpvZsbkEBOpG9FqL6XhdNsbkIFd22zDdbjZbwDxhtrW477F27WwdrR29V9rCq
VdCzQIIqO6+sv+OQZ0BfwS5EUCqeZXN8QpOQ7M/+ig46+pfXeY9KnlYSMdnp7WE8
OGXKwu6hORoC4VfnOYmO+dU+mDFV7YbtBzDPsABvzm63oTYuhDDy6hEk7znEeWlQ
iDJexnnTwLAauJb2lGNs6EuBgVae5tga1vCj0W0knSNM/Ve05a6SD7a+xVXlHLza
8yyiN3ZauEJNHc9BKNYQ9SU8iYsetde2Bn+hKZHbZ2BVpl2TT/uQ1W7zlTtze6EI
Yfrl8orWeaU1WeKD4DEc7ruRj7cNLu9kSn645xmbNzVzciZqhIfQ3BdbwYCp4nWt
LZh7Wt/FWP14elPkAWxMTGAS74/gg9do/ky1AIRoLSAVecs2kH38eH07zeE1cj+1
kITOvLiN2MkUHk8SxJLtcFRIsJATWu0IJ5DgJQvtmdZvEoHujXgxzTstpGQK4JL4
gS+At96qcCNoFANrsBfHANvlFpjdtaAxIpOjR/WxXN1J1SlYMvlKqcjXYGM/Rs31
E0KFz3r4wvMkPJttMUnsq7WVFGwNXpKGkrJ3Rkx/ZU5nxoFBYQ8usjzDCvo4ddYo
AE6K+Ksx7nZO4uxizPCdE9zddVZF2iXK5lNZzX4X4T+Q5la68xEKg7qd5vEAoTso
J5yZ8UErWrW4u2sKwrlNLG0qBS6uLXsgqxyF6FXoh41M0iL3IA7lvak0Le0xE3uF
MBWaUJxaMtyqQXVx46OMHd14RsRH7FHaNTPSWaB+aQZcI1kyR+C9wLyIEEcD4QhK
IleRZY0Vugh5CoGsGCy75iy3QU2jOzJkCNkYzyLhqi4G2mSsv8yPttuIxZDewd27
MUUCJabQ4Dnvfet5nqE1zkmtSa2WFBHHstRSwMgQOU8UvLcY8I5rwHP/xgR0hu5j
J2vZESy6pZx/zr+CWO8KP5wBUzu+0jIx5pn/jRmbsDl6LiIAT0s/mjdZeSHDo6vJ
DI+eFTcxwFlxUmZx2vRyeN7fpkbDK+ECFYNLVdKMUzzpF5O/Ntq0X5hSbheQ8K32
bScjQCBbbuJV2C7YmnRBghTc+FiQJWtptuFt4TVXqDl09gTS/l+lsWlOdMaQGH0R
wC1A6MhygyNh9MSAzGkf7zoD9a/qz2mIknSKh7xH+P21H9bDfoKeWMgodCXL4zhk
j23LD+11FKhhyd1TDFSF3aKHjqRJ1yM4icM34uy9H52kIMCO/k8sDYO6/KnSrw+6
V2IOb2eWshSMGYci6w1RO5beJE8rwWAM+A0Bky54MgTwxHwFkFZK0GKWXpogFv5Q
IAwvMjFiLkFcrTdzD0Xz6FvENwX8YYmHY8l95L0Jd09DhyMz+iFpYIsheIskw0vZ
d5zlL7SGBBlIUeapUDLr7sci1rRVFC7TlkEkG4pE/lDpxZASHbNDqvYZHVxQCwIC
tPWD4BV/ijBo4qDn98kZb7yhadkAq9/jtpDcgA+1zF+wJK4Sfv5IAJhEc7hK4oxl
IDARwfDmAKipJ+5d3Yuq8xGuUwEzlPnHu2x/wUOw4CNUq5ghTr/HghKZiKKVjYgQ
tj0CPDdJYwLbfocEffIh4z5FrNH0ZSjZ1OnVQjrw1V/j4/HeaqmvDBGc0pbWdHvL
7zRVA3q1oN92ENGuSy4Nc3SHx9foim2oEbnCHXimK4iRXrI84rdjTdkrHV/TLQc8
3M8sfdUwcPACKQbmVdU8FY8oh3TE1Rtj4F8GNgB4qTFdrpeacWt31zObsRXo4+ag
41yB8E1gwRVSA/+JGejkqMoAKndjjouGRunYIDk6KwcupK/91IGN5QGMQs94q3Vc
ETgPEdjVYO2R/k0IzflvwzOc1z3kkB/c2Axmo9NXzVLihTB+inzUBa5MOAOCrabP
Qu1Yyzop9/XWCODFAWLUSFXqF3h1nAeukrOftWzW1B5CXEBKZr8sHSmAC6yktdyL
qDQPbHHgzsgSZjDLQqPUIM5Yl+WsPMWQsrwUaD1YckeQFE8klk4MlKwdY0uTswPw
g/nUeHw9v7ffCzrZIr8ADqYt2aZVOZbX96rJgyH2azU80cts5nxbAQej4NQTz/N1
OFRcKk4Hm7/a9r3tbzCovawjwNMFPIUU8zylQRlttwHRtlnMHKfDWjvhQI5BwF/g
1O/gT6XjkKRJ3ItHcHqQ67qKS2SSmo8q5rsTtfPI7JvHeUsSCKxrJZ2ZaVKADT0i
uCac+TxhqrAAksHYB/PAYOD/XXEeIdw+jgh2yGNPd9aWVHPrk6BR+vSsvQG8RYr3
ESEAwqSn0KqnXMZC1RvTP2y5+O9cFvIM/2U9PCpISTiVG4r07SreoHzeLcnG4mn/
RfqWJfwHGxb268IzEb4KYN9RcuR0h5B+JmZKh2/mDDUgP0AEydnPPP7UzxG8GYaO
XD3JbiUWatEeaxGSC0BQSBYogKVCvZNJuT6X7Wc3Rqwueh6tuTWlzmBUyOdMnbfm
IBXHZ5pq3FyOEjxEFcgH+PvlT2KRIJN7xwhVXQDDr+m9AL9THfDDEFf67Cn3SF1r
Hngycwz0oQix/HNfoukKzOiYNxQr/z0GId/o0mHwLw0AM2yoB8GlzLX1ViVlnkkQ
noVMTExRJbnjn7rNQXvVjjb4fmz3wMAJdrz1dtniVtQxjH75XvyysIhTHSkrbNnM
sKZ9zDRBY6Dn5DfU2ARcOsbQ3gJJP0n+ZRXJxpMvfA4HbexChUhz36TC3/X2QU4h
uuWh+54y8DSbc7otu2mPP+jTcwz6libBxyvDc+W72tGVfdFqfjuUKBv7DqsAmmxW
iU1mSfHtBlBk5GqVcW3XGXEYt19iiD6RvdUCj9/Soi9eD+mqNo0CEZiw47wKXB+U
QmqofzpMdfRWZbOuMoo2myx66HVK13QZlbHgegt+4VPx6tMIIuxXY/gPp02YwOha
BDacyy5Ws17NtalXcBOn7rTsiexNFjZs8qbE/yKibnQZ8ZvdMRKnFsDhhnTLi3fb
ZoPBAxtbnyoooo/32xLsoCfPheMX7uzDk+n6XNGaOSpuTvXPHC4RZ6BBkC6/5LCq
qEK0FOyHJCKihMVTwH9qieiIT2webZ4Mun95riAbBwj0cTZSgOcJTOJiXSkeT5Mo
m9VoEU2/NeiYbg3GB32kMJ4BNdztBmhAFKmeMa5BgErchrUKSeKYGqiaszKppE+v
bAJqDybqhZMVgWEMCJJ5JfBW1yarXITHoajLRAkCdurgy/8V3+BrRkNGkyXlYzZJ
PNfkeWHyrew0rNcOPzOVWDARI0JkI1rPxvJoI2sa3Sfc657gOh2txifYyfkBtyHk
SL8dyxHFUERC/8LAcbvXdALMQUqt/1e+VbCyuMh6s2e71qge5ewYqEtSIIDO/d7N
y02g7RYn32s8Z8IUCyyYAd3MU5vOvJacCznvEr7OWOee08ksITC0UCc7ZnLt3U48
u5pAb5wePsC0ax3nJ/WTNpIcUoPAufoYMkmEcSthoX+YxHubS7K2vpYZ93az3YKU
ck/NpG9dBiRExpnuUbpglLZM/c/TmgxO2p7zn5f8poHZH96YyG6a45uVukQLRi3x
3sSYoQ3Su8lcvT9czJdtjNBI6rLwogzhnmYWYdha8n71G/gpAhh9y2qXAC2EvqlZ
RN7+60Ty+25pyHsSpMcBJUTvs93TozOqHBveGAcaINsSzd4krioU646WA1lIJaCD
TOe7HEdMrfpxc4+z3AGwfa76L/D6/UEkdvLYirDZC4jQ8hg3VLiPH7ms9OrWFmYL
iX7BKH5ht8eArhVERoAF18dXU15gX4WGbsc1SGsmNMMSfI+uAK/jz3RTCfwKOVFM
jgnkAp92uCaO7E+jO8EEnBFOIf1REGeQ8iFaIBBO86eZ8e19A9ZrUXNBpm8h5V8D
ieGKASifqUxGfHSR+YFkjNdbC87ZJ+okPPb77N/BNfzeGeLtCKvKOiIsWtB33Pyo
nqS4HxQhdX6XS150bm1MSzLUGdm1b91haRb7nKXKCcgNa6+wk2hH9Y/HurkZEEcy
+6AntgNamGizgHiycxp7i3yPYNUQj+4LS9II9O4jlrwsAKofEh19UHInbDHxlxnn
QsUwL9ONa0W6KBBtTQNvg9LD2jF88l9RYGgLOTETc8EZ8OxRdNWYVRV39toon6z2
9EyjjG07gj4zbEcCH5M6cTIeFLhuQIFHq6p3vfKnHWtFAWYwaANN8McKQNp/u18W
jCLhcymwdOIYJ9IKjRaOJzuvfruPs4z4IynKycgSwteN4r9aYJfBTU3BS1gH8q2P
Z5pjuQE2ZUygeobL5Tw+pD+BLJ8gssnMTVIsGLkI1LqpCX2Av91N3WctJPbxQVCD
vVfCbnLG8GHLrGbtJrdj3q2PCg64vePuq79pJOedkEWYp8DsBZful/Cx+HaT5TZ0
k5V2q9Yo0Wue+2ZpzdmcxVVvSN+RUYu9uFT5HJK8R8bIPl8dWzj/XyMwZG5Xj9Ql
uUikeBbxCiSXd3VTl12Vi/JyW6yU/jzKHEg/GfivfLQW3DDAuITmSsEWNWIZRXGp
/6ourSAf2TcGYA7KL5JfESJETg6Rh7xQ3toRMSGWa7iIsGaWCELfLsuJ/zEX8mGl
DWx+H4Xq75D8ELxRzyYw0WwPFbrsebpDM+k+DkKlK7u2J+qyzVUwFIsnifbgsob1
kHhyUJcEhLCx8TqeKs1E4Yc2mOP+/JK0Yf4klwq9ccsNAvXEE49dZkHXUoNGPjvm
1BkIai6kGC4O8T9tL5LIRY5PMi/iu7c7I97tqxcb2CwSqgj9VzUxC/2LBGd7z0JR
e0VNKTmmEHoU0DVdHdQFwyg8474F7650z9vg5MckUohdSCyJqZDpQU9n6WeBeHIK
STez0dfvyXCHG5NW4r5nBQYsjtT7LIx1xmaPWHxR5qNqAjOIiv1X6AtYD5ZVc03N
SzM6vtwsCENbXnLC76uL8DwL2Yu+LaITkLKGdDV3hNsQNNFctgY4uHbd2/2c4dbk
G6XPZKLtgIhbHZsFhted3sTnKV2aoYgWr42LUobka34Os0eAgVS0oW5bBqzY253d
a5CdD4+xKK35wyUDe5zCIs926uxGhRoPhaD9AnH65Ucuw+61wtxbHWM1l3DfEnAG
pT5qt04ynGGwy2Q4F0FfAVf3aRTcfn4oCzHotNbUa3g2OZJJcldREvPNS816phkg
YPmG9iBSYaKXciQWL+yDkhx5nkzGYteySX+u78ZOO4SG0rYCKY0qaz6udIirBRUR
KsKi5D4q9J/NuUdBgmIRApjLJcTOVaXMinht58qmig/8XEQtR5MqHEI/9gvgz1+p
iBbTPJ7eV0tCLCm7SxJq6eBNrpfw8+x8YnVfXkSyl6Pr6N8YGwMFOg9ruGNPSBOh
1drlLwxr82ZeKDrymLlH7eZI8+QLv5BQmy5U5HaLyHQ+NJsejIXEAIM3AYPgQL1U
Uoiu0nFNFyCVO4U7vvWiPChpm4OC7ilq5waiqfw7smOPcxX9MwBGClzZhbg7VCUv
WeJoQ9c+zUWeKzjCQu7UeQiA7je6e0QMfW+fwOSjk8qxEyPw4gtiGPQPJ0Zw1d44
H9Ryls7S+1BmEh5Wapsi6mtZ/eb7FXXjCP8N/lyRDjKegZBGYq2E27CY1DNDqyVY
8fDagnvyFSVrYeEOXra6Pnuxp1HbX8vVyleKgPNMuTkoXtC3i9d3sACYPOMqjmgX
/7pYmNSpLwj///VBVzb16gq5xi8XTLRIq3z786Gm//5FfHhbVbQMOS3eoFui/X6b
Sda8eGVZTTSiPhOeRcflu9NtEE9VRBEvxGPkyK5rKdzbk1ZP1G0fpaNWVhQ0zOU7
6wnviJ0Bd+nF0RrDVFyXi7uCC5j/0Bfen4mMsGbkxLECpt3L78n6s6OoyIyXVSWd
YckqE2z15jz/24AaCGZyIkmJdWiyzQbIxFf910ofVgCZUcojNn2dohrTk7rHOQJc
fm6SwJQbgtK1CY8DRx0dqeF6hfWD662ehJjgDYE3IVMHpP9cuWOEI/JA5XkIFaL/
a9EyTAAKGFMsiEZ1zD6wxo+XNIyuvcamMN1Q1caJDyjxxYavDaHvzMFmqq9LcTYn
32gn2EUbOn8zg54S+HoTtddJYNSJDp+GKEQMP4CkeHkcCUuWyOSKYjz8R3YBIaNv
xhDE/vX5HRFqSvv84aOSutnNLhJAv8+VFVMGhe3oDfss53Nnt5/BU7mfneXKWyQQ
xuQbbuwwjk8E1Zk0CBtE38RzAvfgHFGVGoPDTsVAhvS7avP73P/DgVyA+fyVwyyW
+8+NVCeH7oiqPMkSDF5CM6SYAdeFRAI38qKoGPvWJIYUu78vjGnWmHeFnIE0CpVv
KcEdkx66AYKipRxYtVHA2mbzPf++QoC94MVW3D6L5fqFnbyDI5XaVcDyJfQ57Lnz
3vzplXBzjcfsc1D82ZxbyNOuLa0O2n1NPaDF5SC1EnKeT62EKgCVMts+EoDPIY+F
uZV6woRt9jm4FJcFmSuWHrTwA8ty+N0xeCVKMFfeIqHVtR7ohcQ/ryFCc3qoFiin
EO9VVOlKqb4gJHxcrQpfNtRxbkg4IQCGOPkl7quAwWxGm4bj1OhXF4OWMppcOYGY
e2r7p34pAi7/Ig6eHnor8FcgKoCW8LgTTTarLe/R/sUHHlGUQdBOqCwnX9UKTtw9
9r79nAZ0YISD6FhtpNu0S4VfpF03DNnQCxAr9X8T/QQQeZSMAzAHYJ8rAb/ahBAt
KIP6dWw1v9+GiVQ67hIV36Zkr1EH4dm16EnLlgT+iYjapU2JgtyKQp1Ea8CtvNnA
Up3q6rg8xH7F+LPHVTirzo9tUaS4bCcZ54rlGbKmAUuR4zY5AwKDeFCdBtMuGxAI
BXYawtN3qfBskSh6r2XHhznEUlmFF8QirMdBFoInm9H6f+XlAILN9D6FZdNNoO0R
xX61mmYs6pWOU8jFZZtTsHvipoKiFLtcoq2fzVtPBSJu0c432CVA4RKslINGojKb
DSTxslwpRNaEFtVR+69gT8endzkh2vnzM4BF520FQl85mohoN9ycY3DpOkCmflGF
hvEKZTk7SPxAt0fYNSNdqiGhjSuMa6oC21oPV10xHpY8tWbEs6ilpPDj342xgR/+
nijZHn6qyF1m5hU2JupSQfkh77QAO8VY2P3+lO1EX8tm/9yQ9BzzbE2SeOxMiyRG
Nhy7N2Hp5FBhP9VapC8MbMwimt6yaoDfzgd9NyjmTEeOUaZwL+4hMResq3xZi0gp
fQxP63aBs+x0gCDMss3GpmXQ1U4sY32TWvY+9IYJWC60vJArWp/7p00ONK0X4IU9
5N41MQsVtj1D3ZsiqYhG4TaksXO/DaLPWv1Mv4jrRsZOR4umObIcuJccDcwfXsHY
SXJNdW9ckFco33klQ1nwM1JUm/gg5ZnvcO8ln6ae/mk/0E9VZcG3SIDU+DdHYFiQ
CVinitcIyFYF/ZfuL8j4UCxdbis9nuFGy2rsTjQ2pYVt0BuCn2B2TJ6KRmrGo9J5
82itPsC0mdS2U2wsF7DBa5eDvxXj1E/j/oIcy164SgOOI0UFl5VcrTyrZobFt8i2
w2LqPQ+W97iHbrlVCySlhit4RprxyQF3KIZGMp0pKZFpI3nm4OoroqeIq8tC/c5Z
czmwcN6uT5c69F2bwctzIXWidN5IUWfUqc5jF275scGWtgL1qgaDBu+6DDJoS+vp
5N09hW9t2I1trmWBza07roC5FeBWdnXmak0xfEh9ccPqxk3Yvvf3MQL5454k7u10
lhVe7R6f9Ntko/T4AYPo5a2SgUtXZDFymWMSk/OXM0lb4stONBXIHoqXA5p27P3M
A/ftjAglS7PIoSmtPRseMHURB2zFEdXXx80WobO63MQ0p0/q3lr0x1NcItH4RM+X
8Qraq6CyhGWDf4kO1EKmTGfEXYil5+r86uYWa2FlbGwfp1y0ny2cBOXS/jCNv8E7
3mtHeyhcODE2BE28Vuy7teOmphCx8paK5V6fyaPk2csqZGE0e39vB/lxnQDJAG6N
8oNM1A7IGan3c5skNYFlNaXOwxj5n9Japk3P7uAazLtwYdqF65RGRyyuqxmmvhgO
VO3GWFkRKzHMVN8LFhLRDXMyOs3y2fSuD916Jzu5LJrinsa+cLf/jlItZYMjGaMK
lnpnbCIS7omZMkGfar1BUP+Y3QvVabg0Zbg5x136dp/pqnr8budqY5QdGcjm1KO1
n3zR9YVYP0Q6ISZlxxwfCsfY0ZVU7zCepZSLGUUlyDIP9XOc8zGZa7t9ubKEjA6p
8f2nLnfeOfPUdkKjkYrdPPgUgDhTCrHos+sBi/2dQ39JwrBM5//pMtokKUhZTZvd
cPvVb+JNR/wDOX2zteSYSP6B8MKSryvC6s1kphzs0HWGNSTb/qzzG+gSwsdfXxfV
yFtiziH0A4+Ipj/3hf3NAWuSRlt+2ZPMg6wHYW0glmLY2mYreb3pZXo3MqBgEoj/
2eM2Nzsfb799o4qNPNeEaCfPZ4Zgyg18Xsnt3Rp2DBLoTE+gIDjfa0G5MALaNjpP
eOWfWghq+DiVnqkZJX/Ciu0Ip/tNG8Q73QhornjX+PtzoaYPFCJNOHGRVLHoSwAN
OIFmWX26sLrDjo67LYBdRnlqInxyoMLy40rm8e+tvtoasYj/KG4KoYqn46qcTGvH
LWWp3xNQmlJkVtTaQD6jNw3cH21DeKmAv/v4kGB54CHN28ijjEL2enafMh9r6tqs
njOC1mJYAeWIyU2KB4LAW6yEmXq+WYEJF6xcusmj5Yg/yvk45fstGZ6gzO+/fbYJ
N0LoPi+BC7nJvR0zeQ/MfrsVbYUNeHpZWQwRpE8oA3Aw/SVQ3Oe5iy3ERaX9ceYq
Fyqk6q2CEs0UmflaQpIgmXrgQKhw9YVzh2YJH3DG/eDHzp2zkShv6g5yhMhJjGhp
kkIMh/ZOvoBjLsS3gKMzIJh36cRZZ4W/NOpZyhABRlGtenPlJIcPhQ85CU1gRbV3
4MzNjD96gNV7eqEmEuCv5SvTBsTiE5g6F5w+9JySpX/6BvrdlJRlqVlK0atve80V
NxkFpcj6Xtxkvc4wdCZ7v6J59Y1FAEYLj24MCAV0t/RoiDTCJyNWiEfy6gL+J7JN
ABRjlPcwH+KYvSkpZo142zFL+uTCwn9RwfjNhwZqRc9gueE3W5eS93FzG7+GaZkd
lCvq4bK2EGEnUCsp82JTUU82zXmZ1npRTSiK5ocYL8vcIOm7nS1LcKNmX3CLz1At
boG01Fzj4Pt8iyfpaI/GpJyj7+lUiUGSfHDidkw0shid9b30m78n1+9kYVe8CwZW
jXldrDGYsZJj54MvEapCEGLfhWqchJVptHKo0T29ujslrDNBzNG2NTd5tE826lgj
2/npRQVdrt2jh448rgJKN8hjXsdUhLcA1UfYSOmphuaqLwCLiQgOC5uG8iAND8fE
6eBLE8fINf6zkJSL3VkJN7jWYbnESNgCzaeVRyKskTbvdU/FQlcigKqrXs3/3U1i
XxP1tQRTTMXKcuLp83a/peXgV2NNnYhD7oA4sTgPBN0EOoxqvVbEem295xFIgpaP
2cGHQ0+5aCBEpiwHr7J9WHDDYdCRXz3LnNPS9ftrPZbFr5OFrOzhBdKLCkX8K6+Y
dLBIX/I/H3bn0iVJ5T0xyqlt+w1xFCotqkNHOZTDba9sgmbWoSd/Hf78Ngxja5p5
2ArpDalEDm2maOkSeB8QrtIn1dx250boVBcj1ne874CylUiSbsaxjzV+pNsrujVF
X/MpmI2U23CgdXOGWaD25BUc1W1XvCW6HJlA+MOLNliXqYM/X8mtYiqHotWl8tbW
LmM10S2lKRxvBACoBfbBqxwKHlPHf0XNSw5vjMRHnNYna1LpsnialLP5J8HDwH3U
SS1pNSV6oU+HTutcesMPsV103LyXFtbiRG+P61pGeRDXjCAPN1SedFls+5SQCoRU
GzTYETV/KU1WpPLnDJrO9VKvlYR9uZUB+3nhLJLyWdtR5ICnqJ1CTCaP+Tl1e4iZ
/YM3Fbqx4gijq4cOp30+n0cbi1HXLlzoAhkowAKaZK30NbV27fmGPtWqzZ7Hj3Pc
EedjzVtRIXvseEbfZzD0/8WWKClun9n56KcRaHny97+o9+jTC0ntruXKXF4V5feY
K9Gk6VbvsaAW75BNB3RDSeZkVRH03gDD2cxgwXOkVFOMHxk9+c11Dzg/k1CcEujv
ZxI5IdRM1FwTWwKW+E3qpT6pXf5nZCyJHCBGXoucBoYzqknFHeHKP0xJyL6iZYS/
hUHOClUgneD9oZ3FWeZIaaOLKk9nS30hUCs7AdVByexxg4DmzbXo784RrvnbYQPF
3EGB390ec8yR5ShD42NWu+cAo2QdNHxv6qy6IU4VT4HDmcVCQLQeYDh4MsxgHgrL
R7do8lpnKNa7CGajt4PKGyk1QcEFKO5KvebcwfumU9SRYQ7sonwtn5yorZojVKn5
OpiYPPue6o5jcERAoGkaZziXK7Gy7/Om0VgpoVNklBsH7rlYg8nSDw+3CXojWoSq
rGgGK4oykDhRxyilX+w7Q46WjQnJ12In8eXjMvIQ084ijkqWz7feDRtqRtUr86T6
z4Mhjjcskk13G1h77MYBImbLb7V2xwNOvErt//bfR/NzGFUGvPuEqcLYx/lK7ynS
zw4OytT63XGl7CtHrUGZLdgL3DX/iHmyQnWqaOFZ5jH5+xmmwTj6c0i53X4ienQc
y71oI3TEGmHmJYigK/Rw/YoEf+sdBC9gYF7IH50GuvUPGos6kezhhcQrxlH/45Qa
T/1pJh+5O1ZDzhWNdQCvj8TxkpexqHkXxe//obRcksHS5ukXqNWZRVvogQHM7JHJ
pXUD1pVjS6yj4I5ZPPuYSzpjQuYCpykHZhLa/aNCGNkNOptABE/spuccdvwic5YU
zxsgxFTfikjnlSbkVMn++oXDTDbhba+22Ybb9KlZSt937oh2vxToMEzXOtaPksy9
+6t55LY4pVrcrTRu9ecH57dJZPT4mmtd9b+5ZSXBNw41q7vsQw7kPC8W9x2wVi0i
kisAJLtIbv5xUNR+NBa3gcR7GPnfOtEW2MfBS53cezp34eJH13bHHXg4g6jlXTwB
365/fvq3yqvXgjs/su1JWQWya6ucVV/9QFoDI8S1Ore+LZzPW1x2uFrte66uOVrA
UQtEIjoSWIbvxvAqxcq981Bf8dkqjk9AQyMyTe96mSeZlOz4Zimak34IfamWi0HZ
/rHQCa3xMVKAJHiKMRFTNyTsnNthvP5BwdWf+i+Xpy/q+emAco0j2LYbUL3h3y3V
hIpPEYQyukLm0FkE3H9mH7NLu9RI8YnecB3gL5/kj4qOb/xO6EBO4Stpnt94ssfC
ktd/eGLGVDA1ze7gCnoS3IAjQv1h93upETHmV2N68SkkiPuEAU3mbM6idgf1RmTq
kwnrBVF3H1iwyBoJmcXW6k7BrMvbWXj0ChFMxp83+m4QOYgOAwf9pQXmLHUe8ROV
3q21elslCB3c8t3AzhhIKGYnO60SkjgzQwrhnr8YR134c/jGK1HpmoT6Omv0/Edw
CkyAMEM2wdV1RzG7R21qYjV5a5aHDYx1BfLyGxw5dWl/jQ4+nZp+E/2EKqNu9ylY
Ey2oSFgJMRVL6edQ+7aNGWnq6yteBCIIbDNDHINWh2wGebXpestP+IF9+I7D6YMH
XPaWW0W8Z/qZbck9zSHrZ2BimMsG5+jucarA7zqYOZUx/SNE1sH5c2atcArhY+Wk
C3p23v/PRER+ie2ZJpla6JdODkv/dgw+lgIWrwQ2mOv2ZcnxxizzoLAzwxoOMv3a
PbFm86XwKigc66M0YA/BdM/exQ9/8ak/rnex3GM7CAAH4jdXizyw1J/zAUUirxfB
YADuMj73GkWY+U4rU6JVoH70ci/74yNJwlXnO3NnIo2jIAOVs+ZIbRF8F5ong7DH
//rBikuuPAqQVYR6FeOrWwgpflgGJUOGkTgWHuKKYkUGCE4qnnViawQWZeCpB2AU
8irly4OgY+p9t6ZsQPqmJoaF1rKMBIcbQQ0BN++Fri9qv24ODlhjHqibHd8tA9hL
e2mwFlYbYMqq8Tn9gahC1MIlfmuO9XKoDHCzF6oWqRk5ynvy+8EDfHVEwziyMG1E
NnmNX7k2fAojl2sHDPzPfPSrmKHUeTWgJVaiGLVEUt7ZwOFXVHwOiCUL8gTDo0Dy
DSBHwoh3qe8txSLUjYQtBV225P3N9qC+lQ5DKrpMf9MZKaBdFH6zTn6YVfIXX//r
QanQH20Eo+mg/eZaSI5lDo+wLgMyiPQ4A31CjHnYsp0Wfk88SK2+mAmQno+1k4AW
n2sxBShUA/V0N8W4uXt+0Bc8XVLXPavUb0UcicG6HgpXfv1XlSL5JxuI63+XG+BY
LR32/sbzb+k4vNPy60WoTgqukeDPP2DRrlQzh4XhB86jTmzCP28yCdQaNSEw8N+C
dIGokDH98U49UCSoy0ZBoMLAdJs3qAMhn6zhXX2zF7LvbGyBYAaPgbpyscRk2PkS
9O8GWyugGQD50JlEbwKwWDztOcdTz81FuUWNlcj1Knz/QoKxNzcv2dPeylnVwAlo
havD49Q4HLp71iqdtHJd5J+ihL7j2VnkQHJO+r/+hEjccbohrB5LWMX+zWHVkeFn
uCIkn7OkJSRLDMMXexkGzNlg/7OxPya/9nvKjXIYwTfZbLDxIlxaUbrCzfv+PIYv
RRGZ98Q50udrlZbnY5CpwVHfvfEeNbJjImAzdwOGSN6Sl9qhLSX0qS52HRta/oKM
+IFZxjXQKXdFY1kcmkLn4158pn0qiDLPHjZcKXoIkT20SFCdttetozZ5MMI7CC7E
cEQPSDQ5F4DOEAijxm/HMjH8P0LDsTPW+8egoqitVYutneM9HlioXWmKcC1JE6/Y
bXUZT/r6e9r+C8NoWJrZzjXu9m88sNXgBdfBf/G2vMNC6EejyDw/l7iPalVKn0Jf
9SUXvLS+8ruai3nXcnfEHqEmg99LhcZe9rF3tKri8nzhP4l/iciiP/TgTIgjid3P
1m/DDLSP87jUtkjubjMPKsmjQiFOiFTFEVng6qWpHseGUgPbFRmtCPgeiDEhAn4q
zvBYmTRiO5wwD2R1PG/1GpDH0t1+Er9CfmPVntAEHJBw9fm17p76vi8ZA3jPiphy
d8pF9FQFSBA7j7hf+P1YmQH5ERE6DQCNihrNcx/S3t8cYeMrF0WaZee/jP8pCbf7
drrzqRkrTjqB/jLc4QN7PczEje/DjoDRb4Uh5CcGCMrezNwJmWw0V5H9pwNwGrcC
Byegy/AQuyFiDtw1HYoDeTfyF7eT/nIwziahxR4W8Ebp2N24TQlJovQ7m3D+bK9U
xycP+EOXcL4aTooYYsA64WccOySqni+lmXxCJNLWqBhYZXYRZtlcZ70dXBAciA6P
pFwcR2a8tYSoYTXmss92hcKIppiXdZLqf9u1YY+n8bmxIF7z5UBx2gV6hshPIzOu
SVEPWZQwwVsiss7MysMLEGeh7DXIAq55m4hjNPhWX21KjmeZIAr05bEcu2Jda+Ji
zKDEpKvHxBe0PHyWI4i5lsiH8f/Or0mR7itCrQT8KxftkA4geBUQSttOIx4VhAwD
R9o6rLWtUT1JXtbhaKVUpXKTv1rY/jIgYPMqW9SrLuVd51vvx1uOJ4DS9ESHSTu1
g3CAwowTUGSbBE+iY6AqJeM7lgvVa0EQZUJUJbF8TgPVdRWD3iHxqNWTLoQT/Hl0
mz4pSU0BzImPuflcDRCd5NP37qs8silmrZnHCWhz9mTjmy8KSF7Dg6oTtEwiQ2vk
lac61qPLrRUZ4g1PkUc5qjDMf7/DEJGBLCAn0db1qGUuwN8AwbtPLhP0CO/evPO2
kuUHBUtU9Rd2BRZDawxrlrkVbmVvQwyx+7Hy7QamyU1xPXiEMzTIaG/gHZ+u4Arm
9CjCpX7DpLSjhNEthG+2x+ZQ+5KvZIp1Haf2NwWuZhOXCQjo1Nc9sq+9lOsNKUYZ
jQhHPwiOKRJa5dFd4GuQ4o27Ovh/MGyvw5ikyQLICdBsc6f9akbh4lypXGFR8Lj7
gbHM0Gpi3l4ahMGJIE7hl83MlDRiwJoGuEfnvKUXJjBA5I2xkoS71vdbsqX4xjwz
CSUd67JoAB3JE0DeXjbmmOjt1Xf53ZdKXyLa1wBbgAIiRnQV03W08vr88PEB/Yc/
56EfZnpViGvPjg50YFL7GNYBsmdiYnP9vP0ycgsMwfV4yXogpnX1u4cFSUmhTI4e
898tIhYLEf3NpSWykus4GxTNalTYX74Rc31btkzmAsLIDZpr7IM8bPDaggAhhDka
9bEdiASclU3KV3uOYUXAa+NZkRRLalMBfA4IWY4k0FBXLqdf80ZlhEQPEA2pUiTe
BmGXXQqpXDs/BCNpaEE3Q7vtvT9PGGo6LFscmlOlqr09PWJSvd7mrAkAYJeO0/Dq
jwW32CiGG35NLsJtcp3OLH0VETFhkU3RbVU6TqMEevuxGQzQRna+EzLaA4YUROuW
HoS0oKq+rgzohDHq8QuLfaq+XIk/0rQ6EIftOTZONm8BGKZAuWowTOjGumvjkEkW
/NacqVbkZlCjWxnJ42g+cG0ZuvEKDBlOX/pI4BBHNRo8xIXwI4FAkBZWwrYQ800L
5Ba4vLBNIZsfn8aX96+qFCdt38Mlus0cgUbgHVqAYmZHdrnqZ0SA3gVM3eZeCzer
71cST0Dcz7WxG4HstJnTVimb4J5jG1O/YW8htK1XUSUkvnekj0vxPEr70nQ6WjWv
bSiQp1a9nw9sYmdCDRBSBODbw0RNf8UP0d9fjJpTs7Sw473QxMR2zhPvhM5Rm6ql
9E+0lVhvqOhvCJQmDq9RXWkDTzMK5kbssfcBCNkGtXoMuV7RyR3pJcLRAxqL5dKT
Ob4JOqcDPuCVbaSiRdkz4bT67JMivTmnV8ZzdFAiHcOnIev7tinvmvdmoabUWv9/
qYjKuMVnDsUhW0/+NzH9QV9nfqCwzOhEOwKEpuGSlPuneqv5X5742oX3GnWsfxFf
Wp1cnyHqgGg5C2+3UjDVoCrHQcCaPLflOi6qfEyHDgcgBcXWI8cAV2aqO9cLWJfp
wV7CQbpMQCR8DzRSFtCEzzQFdyYDN4BW5Cc5+U8JhWKAtNxR42Cy8LQz3l5N8CmC
QZkwZTvI7H1LbpKF5J+MRLXj/e+mJ6UbLgs3MSaWp4UWSamVoaYpB8u8bl21XwHU
lCBbXqROyG/OEyfy58sWTAN6y344SqZmIcaff116VQqjeK60Yq3m6iJiq2nzmfHY
2jqiGrrNo3xSZYQiFxM7Hq5qyhSXlNIyZQSAL9mKzcAsSI1SsoRx22n/OUzsCLmk
uKr/pFH4aNZ+dpbFBq1La01YDmjI2sah0JlYd+cfznpdnTsMUc6FbjIbysVIrP3P
RgT66OFvgADFRvo7XFv7qsr70VSaTW2fTYpBeVXZql15WByyPv/YTiwOGJLNjn7f
NsSZ9M1nQCx6u590C2uRdY/I0cFeICGEt2XDF7QW4LbuWBSo43pqP15o6oicQIOe
hDRi+gt3UVaiX8LShFlwLfZGNXkAHdQ2jJucn5OQ/IAhKiNfjU3XYPF19Aa0Q8Zk
1lBgySaihmXeG6xHcC/gX3iPupmCDZt8PU6dwk0yZUly7b5I22VCyXPIHSus3A1f
cytcTWeZYox1xSB65gAzZ8RJhkUH0EW99ZWRzx9RHnV+J6MxVWYtsIY1yKtLb+df
gMasTg43kPXIPoqwkFn9f/JyFtEjZ+43nZtN4pz6Uq2NyKfQBqGiQ26ICw+ngF/w
w1nK6ndAxEopTeyLjD46+oXV9mV3qpcDeeR3nQPu8NjQ35PvPO7+Lanuz4Lc+eTl
V8b/m3LrjdUJraaOR1bKBnuuZBhv3Wksfcmu2SQPanURWoXot0JaacnQp9VXBvuL
lc+bMWK1J6yV7QCkZazREhKFit5lU7FK++N8nQ9J9008f1uVXwoSJeARv/dRIx/l
VmsV2U+LwQ+npokSyZVlzUutUhIcZdcA7G2guTp/wvUwjVQKq/l6fGVhn4uar5y8
37KOlf/FiM0gwaPcoZmGr0/nPkpb7knLqLXgQYdz9Iai/vvrjxZ3y8RgOmI70rhS
dtCg4IkcETiZS//4a2XeQ/HY5JZkhZQunSe5/JR2KZtl5SQjK1IYaa1xcDp5GH3Y
vJLILngaGzff5d0U2j/GypuJGxvVXDGErPg6QcFEe7sneRJYneBBmDzWqoRLQXgG
WlNnp6GbvzsP9e/rZBj5YM/WaJ21AsJmX2JfYfbW3Ec9rgxpGNRbteNk6++9YbzB
CJUNhp9/6eeAgx9Pf0sGqe4QDSIgEnnOmTG7JqBKCqMg1np2eAbWblnorpNUgDYF
KOoFrhPO4kAVUGAoWpljLx4Fbpjh99lq8bogx8CIaEiliHupS47jpjLCh/YpeWiP
4q/ugsWXNboEIr1qCpjXSscRPAUNwY2bxlFO44FBaiq9ri/zFip0vvRPtEjnSaiJ
S1OSORa+HFxxZ+Svpp5F4RrIk47u/l8OzJjjc9+ibiIsNkAkaLjgLiAE2QcgTqG2
BJDwak7E3N8TwvCH10KiM8gj1RiVsdpUXmfsklasnSZuf16gmW7fQIEl/eAgxKJU
cjQy7fqUHQor3PE85Yi+OycSFNqg1+WjuvhtMh03VU0o5s5siy5gAmC2/HiOzvki
tgu4mgpLWafG17D7JcqxXvUBDX5VoZt05fXlu5/aLVXga+29N7bo2Mh7cjVaJ0Pg
IMJCx/+w/YmhXBQP82EfQP/n3X52/AevDsMPY3eihIuPxtdeWdtc3pOjXhUJXiMb
ommg+qwghT7d2LlUh38rL0tD0VZzqPfVhskDwDGmMXVAkW4ErrvNZ42X2i/LL8Ck
jgjs9OZK6y1yH9XibdE28DcAjRiS3H4OKFTifjUrn5Gf1L5nsjGwPxhioYG3DDaz
QXSKVx7aioSyTJqhzLBPNtkhU9lIP/Ta3YyJAeSaROkxn7JcVY2wfl1hnfu1Ln48
UOATCPOGtWQL/a+5Dvy0eJjIxLGTiaSswJTMdKk6NV3laZ0cXOdBEulfFvnll4NT
9IRkOgr+xnl9gNPCzjV0wqzKIP8L3T4tZk9NodeRpp4grdNsDJeadrXbnIZdL9gz
ivxGLxuJQiskAc8B1TKeYq8itZCgG2wv6asO6cD/C0vRC2QxICsmrbAkd2WyX0qf
zLQHwyId4z075UfE3gIiGEHnacSaudjzEyKW0ILj+NvmaY/71CcsKnt3I6Bda6MF
WhnRwBHkub/gVRxJbWj7WPVjpmu/YRyfmaLyuQtsejJ7X4BQL9bdj3oPouOb0oid
n+p/Tvd+88zKm9B/2fUEuN7qa2g8NjrEpsKx/9NmiiOBt1LwSS67GPQQLYqeQ4ql
3OuGyt88oiGdSqr9nLayV2x6dTUuQXDGQeQFapDzyfph3nvyw1pl/IS79gljMmpP
n2Zg+QgihvlcvlhjEmJfGhxOSX2Wgtu3TfBn2HY01YhG6naV9D3VqcbYCvNL5iUD
gMLbacnJhmWr9ajPYorMkZuQyWoj4t+gcmGMkPtOSbovcBkgrpWbeA4puNwPB7ah
eTkX1hEyBY47hWV7XoJEEF4OwO3hpWjKG1Wnz+oPDgUQiH1OwwQ/Gs9CTbNeIkHC
DIddJqfktSElzzKyDaABwRbegKUlXtZMlF44W8HO5vZlGoVBfYdl0P3MhObPlRPS
zenZctt4IWX6CIKN2DL9FLMiGf73GHUfw8iSM4smZ8jxnU4sfXTs39ufZC09cEED
cZHPbFxFiCNvjKFyAIKDOvGXi/Q6WvJVBHjt1TT2VQmVHhveDLuXvlRo8ReAtvlS
68YmhDRUk/mCtK0KSf0+5XHT4yCT+j8BBFODMW2DZgN/56ih2gfjTN3dGiftFQoA
y4pDcgnILq+pH/K49HWk21a5TWxo1RFdFa5UECkhn23zKSHymHBsrEMEXexbKGc6
pO4eQYTBs0Rhmli1WogA5nd6NRqC2whLWVIoa0Lzd7Eot5XKvjvpFM3ubt0G8uzT
B3Ez1tNbiHbmK9jt4+47Nf0i9D/YIjZsXp12o29c6cgVV8dnvWvH9xuMk/JMH5F/
88FBqpaMEQI2DimCOdvSGs5Wmnz8KcvtrkU4pH4ZHizX12lvNodAswyOfKlXbCYu
FC3AiIIJ36VrZy0xuHLZJQ2Jnb1EOeSD4QCm/r4RKvuW1ebHVxEkQuBT6wxGF5Uv
ez/k+0Ot4999Td91euJXUyFwavhbt+ypkmBhtKuA3tk/U7PNdP1wEHFAL5CqPH7w
mVPKmsCecyJTokthJo97MDve2QH3Nlaa1czDYnjiZ3CtWYZS/qG+mNmm23/j0UPL
OAf7gtDkwBi94yVeySAARQlpT63wW5Ba/eQB+2LAiI8yF4oug4Ko8vmuLcRV1j9X
EdUCUOFN1dHJqIWx7uMFa8gF0rAJAAX0jhL1zTO1+sPJbKaUSI1gGnvb6dMOSspw
/GVeychcS+nBw574BWPu6mz/qh3Tt9cS6NkAb2Qwb4Y4bZ2aBe2fdO96PIwu10Dw
hlhq8ps05xH351wfucqyE2QgtAGGHkPNivlqa80Zq1O97nrycy3DLR7Yrce4zMYw
MSA9kvXDQV3RXxX4A3RKTR4JGUIFPleF3mdVPFaRnUW+yedr/Ag4eVQ+WhxMCKO2
B3Zis/V2GbmzQTwnD4ePQiyDT5AuYF96d/ChOiWuaKl0OTRLAcy7OTx1+DAA/GUT
HpJFuR1lv261koDawcWTBCwYzJPj35FP7WJmiGb5Yp9iWdTf8CfVQ/w6pMKdRwFB
6QO4UmluHLCEyZUpSVjS3l8vQst6/XmatvxE0NcEO/ZT+EqE7L+MXW6dIotdPHYT
j3e5nM90x4bd67JmFSeAXkOY8mFZy5x4T8/VN3D0GgLOYqYTCb23zQiXTPkOlkLQ
eyAONUsjcFON6wediFP66YiBIvOVYviSI2w10X+YhqXAN4hjMFpLUvQ6UNFUviCE
qCDTLL7gprnT/dtEVjyHwSSlU58mXe3JoUCaSjFBN+CuJkwpAo8EwM2t0yRsWzCj
7lQjEVTYVWhrokWJvzFP/VVhhk80qvzcKYC9+5KLKt2QtpuZ8MfSyIp6JW3yjaws
njSff5UgPNhFmK842F9ZLf2uG7wVEf+Xl+5cDC/4JzqB1h//7bXlmkSZs1c2HSuX
tUG3CGZyZncMWhMQ7vWPaG53uCApMGWCnA0HZ3N8m4rZxHxMd+jeEEeGZrBlvdSW
cS50bBzcx9qUvblqh/24NnzHdeKL8OTkwJAy64Cj4SNY71lnwc5uFj25fUZnMMOd
ylj2iqgt99bmIhoyjZq5LkxIx2yA/aoqgEsfVcU+VuZe29htHkRBhGYviuV6XvpA
lYOCZV9j6j/KdFXyzfG1v9PNN0E/BxUQ2S+H2L5bXi3vo4lTeJa7Fb+veIu5jhsm
XJskRTEmnvc7lJ8e9XHkGZsBZIUsSOumg9LN1OTa+kwokbWISmV0SC2X43cSS64j
KCuFbrWuDLFcsC1sRAznPzzQaI2ssUNF0ZbaDbHXS1b0rAY1YgZvK3pWBxeE+Bfz
PzxysSH/bIwdRAomeAwVntmaHanbFWQZI/ElYaeffEqmiRNLrKVI9WERTCBV1Gb/
AR9DXIuzS2p6MXqTB2NIiw17zM0Zez68ZsPfN52m67nmqKn1WO5iyatPIcmO5XFx
mXGaWu2ikGLqneA1fkHTx+teS3zT7O4Zlz0+NjWsUuGEjF7JoRIbuvm4+3rP8+UR
a9GqfgmhdvtvMy3zz+v2mJjEfFcavTSKviJx841Jalc8YfyBCBrfhYMcoIQXOYCW
Q8sWHRrutqYYZkClQ+tFm/Kd/jmg4nheqNRWIZAqlNv5pLJmZPaJRVdLHRyjFfhK
Fd3Z52BfRPTBrdgMzUe44H/nmcQ3eFYwLGIya3CXmpQiuzXMyV1MhfxRIlfkxNDc
w1s2Tr/qzZIJbSnnuiy1b8mzIwblW5MycrSOyl6zFTp31odIB7Ww8M+02W1OSWMP
HYY2O86htQR/57+GVHoL96QM5hHpEqAtJroknKlEhj7xrSn5AlPgBhDQT2sN0R04
ePqVundPaLEQ0BmHqNXp0B4PEJdNqEexHnYjy02M2RXKIEyjTA9fBZ+d7QS2Xeri
psmUVDEtkfjOtB6VZYVyEcBZKIJ+qJWoSl96wNR79o7OTtM30IlTObx9OFJtfwH4
0kmDTc30t06oImPkCDq7HDDJENjQPZZLNZpKgAK7an/9Q93iUeY8bWYzGzxeibrG
HfeOGg2l0YWXz0aDt4IwFCuk7KVxJdDkamk0NTIMywZujVwaHHI1xzREWj7Qb2B7
W8p/PDE1A8Z2Yf8TSCiisiZEqWJJKQzmn+Bzb+EbcfJbLXpPzbRfo4OTA44AV3iC
jE0dSEBPxJH1G4UOmeTPzkCU6t6bXT4V6N3m34Kx5luYbY6gE/xBSeUXhKkQzYt2
/vPDa1yL2KnaJ00ppnTfoTTommqVQUS2AA2CqMKAp/0VzvpnKolIuWFIN+51cXp3
jWzrmEdHnl4n4XZHta+k0L0TCgU4PaN60CQbqgb6YKUbifHFDKza26pbNVxMoYO5
q6TE15q4D38+rvg6fLEzS+GmBhUuN5Bsxwpt8OXe19+eyh3wO4YYODZGcZ5D5J0U
3K63TL7tbWjDAcsUgMmOm7D3Zj0tSmF9HZbGtSpsb29/oM0aCItE3ncs47b9xtzD
84gLzJJZo5i8qxW8kTESE02ynPtyzIs82cVFUk/WnEqGabkgdDGRa8jiW2gfLrJO
VsITQBsnzVtu3Mo0eHVclxVa9y9Bghq+OH2Z/aH1vW3KphK4LVaMaEqKUyWKX9u6
vOCU6IKUfIPVddmz0ZaN5nIQ+fhGN5i1IE6wPJOQGLjbHqF/jQocPu/kNR0wDRhU
Ob4kyb966mRUgOuDP/YUmZDN16HFEYcqdMHQ8h/Ws12arYmI26ReJsy413YtIlHc
iIetp27WgoFCcE6noZDo4RCTeG0Y3ZYCnWqzpSR0v35swamr5gS9AfzngQiZDQDE
LiUuccAHwqd+4y2lunF1/jYiEaz0gmAD3UVsskWcrK903NqzWC2TPjD/FuczxU8x
HhKocuTaqeuXjofTviBjb+UtEC+BXSYxFMBYjdJUSQ29uogcXDMfvQDLGF4y+oy+
THIhaeho2Gou/4tWZ/l61fIAd2uqGUWvnFq0FCOZRFaxyEwon9TxkisshvJaGJwB
+2gCcDiw9SPVFlXJOZRdAwkYIoKQPT6DB/R7mjY2F6uTU6rftcfkNCR6MEudcIxd
y8VjXwuDDeDgpDG+j/9/OPVtwLLUl1ifkkz3+UFxX2/zUiE7kpdsUEnAUesieYOl
u59nBRCZpVwuH39bYeQcT64HzXUeXdLqu48ddr10CjjpqopSXXR0e70Hwc3RnFao
tAFBaxxcEHwUcexubH8xhNQczCTlRuXoJfZ7pKH1vUiLzXfBZ2YIlu9wOzQVHF3s
2yPI/C/hWF3tp/HiGh3U+kZ3T/Le6y94yXAX1smPQchLP6uZHOJk+UTb6GQp3C5R
wU3Pi5fYbP4rfp1/8Aue3LJrg2uU7/h0pA7Xn2CvCKZtl0ry+Vn5sLGZxF74yxiL
UowCADPmC6qT9+Tw1yAG4KKgFOUA4PZht5ApOOC10x6xKDjeMLjqDhDbAir5ryw4
/MJopbqkMlFfT0gMbnS/p10KkWCCxxEdyNxAgIUN/T1B4cXwKbCRC9qcTX3A255h
nsRnXJn3qfb3pDIEpOIKJgP8TKHD/BWxv3Xjrbhvwjm5RSn4Cjw5Mgnyvyi4vChp
U1r+GFu4pr6dPovfDVMtRbMdF30KMzXmc6ZfCR5Qe+qXbcDzhRDGHeW71NdyL1Ru
scppOfcfrKbZ7rTZg8mVfeiVh595+Wyiteq/PHyqbFp3nvb0ZOrWpUt8olLzEcIG
/qkH7FBWxGpgUUTa1R4WN6VXXjsHjNC9tO3H4d+zurnNA9DkW6bKGfh8yb9rPWsA
eBZS+OFBGu42aNot4u+NyTJUSlImyyC0lyTKlMPOZqABktgIGeMkbvNZ1V0/djfO
m2wnEpTU8XlvFeBuKCyeuUZbd95NFqylo+4fkG1B19Rs7gs1ahc/z6lX8Bm4btF2
knNZ3KicULVXIBKZbOnL0upak09YAnG7XwTeI2+fW9CkgDirSUrjw7k48/BrqpJq
UQRgkhkQ5t9McCj96XmDLRkmcsIGvcp6IiPxuANi7EVEKDLq+nEsapW3J7PpcMKZ
oLj2MscEZ+aQMnWseKG2l5hvj6Rot4+cZNIJ9D61GPZGxPWk03e1XFvKX8BoS2mQ
emflQzIGlg/SVMqHlhCQ9Hpa1y//W+AvABmy2U8UGGpQhnCtt5sCYTtsXhCtjgMl
q/EOivm/maiIEUQDzKBzzhkgmZy3P8A2n1h9Oq1ti4vud1PgPNQBPx1ZX5igGBQ7
oepqhi5tTdwR5ki3cqgE7WNTskBaK5PpPl/9QYa89H5nfdPUrmErIN9VoLXEaQES
ajXElrsrOIXIFpoXrHBDauVtI8SI6qAl56YOLOcJOsrnpuh5a5nkK6bgqOs2BG2s
M/R3MF5CyasI/73ok/5f4VR/0HuqhLjmQpdx+t5JpR7Um+7gtQmrZ0917bYScClN
GULQE9kxUoeMNvh4PxBHmRQn5fGADmYpakHrwWKorQUmktknYqYwBmdON0iujGk3
4bZyryEhIEK1h1wonR3BMKEyydQFvtnnkE5j3eRQ8QF5NaPTdwa5segmNaC/oPBt
qelVL8/bp7gxyr95NF8GrWpOp571vV5r4QhIuQikM3yN4Np68Ny+cD6c8trRfiLN
Wfne2WSwqRmTn7L3kKofOF6Kdr2ARklLBgPWknTo9I4zQSJJzijTuxprX1abPD0k
Cmz0UMm61XlltqhC9ceBa3YIErfRPTLzYoAsoTokX+nKxNIIl0+CWTaugb8n/p88
lzXj7JuMK59jkT0IwzNnEpmBogui+MrcRYEfEfzBahmu8M1Oywttvqx73cpPBZOR
ScowTANO8US6ITjv/IP082U0ks7fD9TZAruTCHSqKRvR+HwtebXL7TceJNQglPDB
OxyU2cTMOV/GTLUL58JPDM+i4oTsk012IV8coWURn400LBZ2qpTpTVHe3NkDtHYF
kaX9OfD8OHLzHK1jUqDVMriTGi8O3tVfQI7P2iVkfZwu6NMAH0Lo13/Zrf+d/TFO
13NUjwaEmNgWoYbvxdWtk8dKN4IV3lT6F031v8jxLgk5rQB87Jwe8Q3y64cMqYMt
UId4deW8M76FTEyC08uwbBeejiuOEPspjU4KtLNqNqBJvb3UjdHFIFXo/+2shTeF
npLqgsPG4aZH9jlxXRw/jHBftZ6O6M+2BZSPByOxBgSNmMrKq1VIqruip9WA2cdd
QlD0ZNJwnDbxsAcNa2qsoXvUwalgkdzUBMp6uOu2st9MZ1L05Yy4IqBwFw/eNjEZ
1q7KOcDjzrRNccbd0O9zuAiXDb7nSykJ9zvdMTXjkGOOV51OflsvPZTQTJNS76UX
0LWRAgFgBXHCfllm/XxNJVi5+XdJbfsL9G4udK3ItSdQOxrYpdWE/RG8U69x7PyP
xCRIoPYREDPw4sQhW0B4aJP/UnecHUV93wFTHGt8cw9+wihVUclIdJtbY/GxvUVH
h3LdmI4YSVon9M8CoZo6y9pAISCmb1Zsbs9r7nsvjykHQ04T3zXXu0gG0NAuSLb8
U17hR+c7+Sd5jgktPqXrA6sbRyyF3Fy98SebpNq4fUrYTFPCgE91cccHmqi3vDx+
9zNgeyA/EP/Gf5u5ozZorVQM0wgcIW80XL7j1vv7BDFT43pZtGtU1v8usGPSbbV5
1O+Q3YCpD7BrcvhimxaMXWI6R8dCbCsYm/xgCcgThdRwweEM8ociT8Fs16iQqhBs
I7IIBjDkwNqIzrvf1SkKoacH/lbaeuDK7IMT2Rpbh42LGoyeoQOZJ/YsQx/A5Lj1
3ZzwIdmkmp6AkV2DEEZ//WzuqH2U8m0rFCHxb6X/0GQVkH0MdlN60EjiMWYZTdtm
ocfyMba5hcSPlA1sKUudmu75TwWpY818cGPtbsTacBvl7m67To6Ch6clHfMed6gZ
DJQko0vZBuVBCKDxEQIe0PPp8HNJkvUb2TtB1CZaAvDkOkKXrzvYGFVFB4CDExmh
bgG+YcGcDaXpCtKufpPRPUHRsEkoXm/+U2EfgbezOCw5IjmqbDIx5oVwRxdNMvWM
u3k7ZLsl4SGFfmXPq8sGc0adix+YxKIsRnFNR+1BprTzDf/t25hNfxiS8Ho+r7i9
HiMb/W2iBgejVKAgF1LHVE3OdZCY13WZaej1+X8VNCMELoBCaJ0sA7JQwOXW3SFO
s7uBqvSf7sPosBpWJxLuyPqzU5NrNwSReQq2HSimBi4BwG+yvAtYzPuw6ELA1VBc
6XuUxwhypDIFmmG0WSAW/2BBN1WJe0iye+Aipt+1lukoecdF0HoN9zuhge7KCQBk
xU1JzWyR7y2A0Z5oaXbduYJss9/N4pafWuQnv284Ui4qDby2Sk5tcmaHAzsuaCxq
7D2kJlp9WfLC+nA7mhe4NVQ0gQOcRKA3cg8Ts54pjeve6715EHV+5WuKuha9+eHV
X/0o2EaoTYk4roJS7n50ZBkZJ4ChdBlN3R7zyAmm7rF1DlL/8khnkAMiO1HTt4/E
FCt4q6ZkGQYPqwZq5dkGsjztu0Apl1bNWaTz962iAs7cLSALP23ntznqSFO+QUY+
2F1ywcgMzjFaUQCLwTKQQ71ru0vRbZqsSizOEe0pjskgelcF3K/+4Kz9k6epowo2
1iAEb+HGMCNqWLsE6ljbFmGRde45VrtlaBmDaldVZpcYacLOtgB78ZE7wzF2wLNh
glnbBjlcR2EockqQ6crOO+Xvrk0AW7Fmv4nSXFwORUWteUhJsW2tLYYq9fo/HDE/
/MxqpTN/Ky/gxjE7E1jpSdFwrnwbXLW8m5FseuljnyXH83sf94fu4A8lT9BS7136
HdqSGTbhkwiEwnYvnIYhqDk7+XC2c04pLSOXP06IgCMHTwsSNyMiIqTFqcms8Wxl
+RV7eb2EtDDiNGosIRTXJuQb4vhkcP517f2Dp+7/f25p8Qd8CwdVlBh282s1HWl0
CGAxitHmroI6nhglMr/kT0v9NycnvvaTyGrpY/uVdveN4oRgex1S174zh6XOuGVF
5a4tGBoQj9Q3Ow1WS9ZKUJcJpG6d/EeLBzfAwZg8rsmLE80xtIawVJtkpfrC5U98
MwKit3w6N7uWBOadee27hOdry2g9rSuPgjNyp3MGcOSJ0EJfHqjJHVWjaGyqa6b2
VaAyfiIJV8u+MDHUXuGEz3my2WbmV08X0Jq7+7bNKiwkE4qtcu/zr37QPlU8sXVX
TaQ9DA+1upk6fLL7iKxnChMIXO0JtFvlhWCZmbs13kaplFjK/ZLcmC+rXNJfr0Ma
+wIpuedUbIaq1t+/NND6pZ8B3GzEdm8AFN13D7qT3AQefJ0um7bFhIbNNEk/Pog5
VF8tE3zBYxEN2GbLkcO8C02t5dplBfh2S1v2k3wkYhKz0BQhoZ/sbniOR2myRXch
+2Dvs4LBHsOwpA6U/+znOWNH0fcbRN7/lcThChx1k3Q/vd5qCItF2YbwsQ+OOLxd
J4HGQzHWo3LDXcGYEwuOULWOnbtpdP+A6ybLfnjzeLBvfsr+oEGsDIBh2kvsQIXW
3aDuRyVPPhHoe8/8oLlt29k8MYehUwybVhYatXn5Dg1VeFtCHfZ8aZWmP8j/uClp
lZVd1EP7GMiIpQgLzRlM4j1UHVJnvXRqUZ2TBG3sutgUjZQMTfLkQ0g17XzmKNG+
18anDzMVuvmc4aqknR8DRoKnD5PBDRn/hC9xMjIxpQLBDCVR0d3o3gbO5GdFji3W
8SZbhgvCNoYAJTTjD4kyWb6racF7A4J4vBcZhnd7pIDc9l9Ecs9/tofi09sX7qWK
SyGB8bzFp95vOvYM0wy1AyW8e0IFVTFBmrfnANOmZa4V08bbVB/nykJntWyK2Xvz
zYerf0i2yUDIJbZfb92fxYmSunu0K4Nvy1aunfnMsx0XOVbRavhTd3DaQZlqHMZC
RHYhhUHSeg7z4kqVCf2rVpmN9J3RyB9eK9ZE2dOwUwppoQQGTIFe5PcJ3V+Dqgnl
0WkmnBYtrHstrmlhxKtuQvDhpBPM3Aa0/INcS9+SlqLC31VH1OqKrgDWMcZQgvyU
PkW2l9UPH+G5J5+JOb8JhblrwabiOkJAZVLzIs2vhg7tTijXEyFe46DOeBheEJM2
63u+hwTKkAf/jjiImCtfSOj5E40Zk22yV/0pJ8UX03/6uaUl+HUKeMpvnx2DUaVN
PpaSl12pcs7uhWHr6oSoYzQW90VKFziIv6grZh5fJK+oTMdZ9IN9ehkz58IcUmEU
lvvzgn02JAs6217Men48u+7zygk32K876PUxf0jerbrs1cG/HZIjlPZKx8hUGMiR
cPP9wIVOS7KriyEgAfM8s3Tat42VcCR94w2TYUG4prpfDwDrFWNO5+nljf099Zlt
RtZ7dnQki6QRKF2GzdR2qxHEC47oLNG8pPuOOdZpe6NfAyabjuHWiGMsDQM18Ito
fVq3h/halOTRDzHesnCUHaZfA/DWmISunizX0NL5AwqmxmPL+A47tma20TDzxo8Y
OjbVn1Xcw0FuLjmYwv+cFsQiZGC7ifBwi199UzcfXC2Jv2guem/sYfXyAB32dqx0
IAVfVM1LQgi52/+eGInvwIGAt8Y1Xy083wfkWE0l/dnSgSWmhHhPTn0FDxAy9baX
TqLvycx9EPcSXReRv3MZysuNQ7exszutYGOrGbcf3fqiqsBAU0MP/xuf6MbybAi8
4cni/bxtUwaj1fgipLNNvSn0r+XLvmRR5i3YBoMASc/Nuo0tUDZMV7I5JZoPTOhE
0J4Y/0c9rJEJ7Qt1yOlQIEZ9Kc+InqXJtWGbsLReHQKyEBifjitH56jBaqVK2YSr
NdOXUWt0NMnF7pYG+vU/5hj1RbDjSwJGMBxHQfvSmyDRVbJWBJSNwswwFIt57kLZ
Ulu+YmBAhohDTFxR0E3jQJ6YMtP474d+if064EDB4S/AjF3U60ejZswSqpAqhv1N
4XYysek/28jCVhvgQqEGQaSLnQCVzUxrhc8QGUDnndr/JIZIPLE7YAKzNpWAze9q
kb7rM12lCeSUUeGCg3LdW1d5ASqyeJPBEU6saZ4h0R/ndjbX1zCLkoRnTqnxccPD
MzdDlMJ2cUOVRVwvsAfVfhpj6gIkf+01AX24eteme6dut1WnhYPtbTcnf62XVhtE
/w3iOLlph7+XDOYDTgbWt4+TSK+3hiJBWXStYHZ206P4/jsrsNizdiCzAPslvWsn
d1A0N6+8rrnuQgJzCrY3cRh+I+XpG4jolm2QUdnvknO0n/hlWubRrfV1++KgzeI3
qEDIGSc45BqUEDFuZgoZOrf35CEhuHG2mRsOdu2Zxv4Bq2XJGOKzWS51piHT1Ato
T92Wu3010ZfzOYru3fSV079soZ7aMEVQ/+8GeL6wN0vwIN+D/stEcXGoxof6Zhwt
vB27K1nt9huemt2ERhyLTr9noslQxiAU/BZe6zOwsU6uXVxY0lXM7wP/z77xIiaP
HCZ/AreADV8dGO0nCd6sHoK3RxxPgyZ89yQB7CNJjqAHgn0PJktUa1XVCHKvXv8y
qbXIcQXhsA1yAx+Eijr6yk+3uwM3hqysrwjJ4bRkGzt7fc2tIcJg3/bTz5meSNlZ
cOoat75QKD4UzfGj60rjeWFFflxVYl2Si1N8S+saISi3bvPt1NYJcNYHemnYnmyg
MUf5iJTMn0taYUVXH4ixRHvfRplwy4u0jYg4C1duA9Uly0zK6CisPs1pTDi/wvMA
JdHTXi1JcaDwn3lTcn56oFSiNYFatcRD3UtFRCnzoS8jXFEtEGUVA7zlmxMTpw0B
7bg70ey+YJHFaFBnzL3jlx+F++t86gznQifHTauS3983H03Ev02w4pup4SDjYhUw
6Rcj2DVIoqnuhz51K0Gxporuyp0B2vc7qUFTCwKDcezx7bilbU5qOcSVOZn9fPi0
ISnG2aKhrc0OqJXAMB7k96rO6bL/WXQh4vtlnEu+YiNgfKFSwFwzuZ3UiBrqf9E7
+s4lAhrdT2laG8fVW5LdYcqD9i8Yb53W23cO3MF1wqcPBr3ZDT59W3427vHCIyOz
/o+QWplUjzRnVPgZx2Qj8Qk/47Ce5kuKrKgRMX9WsT7OWuLq+/lhyt7/tCSzVWeG
miV9i4iyUsTbf0/syCWrlnWCxx7ctmRkuo3IZKTwYQOffeFLwwUOr8q460PkKNiO
S/1mQUcXONcobOsegipeFiMkB0fSMI8Z+4tLx6vmgPD+YCZrjeEoD753U88xUSee
RtkIczGud1Vfj3zvuM3u8P/IDMpidjdF7HNEvcbCnBKo3bEL+++N7hXKpWcO5+Qe
QJHyjgUAy3f7fP+LpMY6Y/+2IIuWLJ0MpNSaFjHAlJr2MVx2qOCxjbpFGWe+d5eI
bHLkt6wNOvX1eioszZ2UK8YAjf30LRBPj0/cN2XwinWh3UYnbOaJiu/9ZnnpwXuX
4TDPLKgsL+ik/dGpFIwbLtKEk0UcLNRM30VlriG5V0ZLJQOQRRzyMQai3q/mGkcq
gZ4Rms1UKkIaQ13bSuc6LxM6UKdm7Q660qdbEz+pfijA6RJ4CCWVJxhbDBVHyZVf
gnZRsL0YBrlRhYM4b9eWIIIJHIkcLjbOThS833nMbwYyuvLF5NXDJ881fo/3nSAL
ESzRQgCE9sxQyQJSDQtO3fhINx3acB/tKo5/MpHnCL/l0KYffXXxxG+Re2NDnN4Y
goI/8OUYjPS1EqF14coWb3blRp45HyZ2HVhpFVpFghpiYh78dA45G84xWuJg6PEq
EibhIshdZaTPEcSLtXD65Iz/Xz/Zon01boA3vq9/c3y3iQZQnARJ5zdLtUMAo9rA
ehzppCmJUFlWhbKuSp2XXDaJBgNXY9VLC2BBrPx9ujtdBNNkT0kQFw5JZx1nbguy
Vuq3bfOVHTFJQhT1M3+p6/51IAKBg2kW7NoRoEICfrz+Hsqui4QvRJXA+yddvoHF
NlNxYtE9lYwbrlIlYtgQdzZbuTz4xs9yMMC5VfJzR9PbhLM11Q15kjfid2AnJxKr
TQMfN41z66T4fJbWPtZnu+SNBykoDxGgaZG8Q8Ta3Qv6EjsJU3QrAPUknu/9mNhj
//QXzYuOCnhOVsIQqIDFrjWr5RcnsfVeZilxOLTxRXcJXsXfTa13in0Y8SDmfH5o
sXM7KGvsAkmhz9H/VqtV/LUpFlrh3J0nLDOIsoU8arP3n/x4NKFt/z/2U4tiP0JI
GyId6uU7mNboXcBEx+qqw8RL3BYupzXDDQ0q2kQRmGF1QZ4AGpXVQhd+IleR9hlc
6NM6rz4E7zgpB0fe17YQzwv0FOrLnEIM24Um8txiLIglykPdcpig5ujowWd83E/m
tEMArytxol1MG2mgnwZ5r7xUybcSKL/UI0yzzwYX9/5DL1Bp9YbnVWoZefuUZbtO
sYDGY47Eeg+ilPObRQz69UuMI7bwXK3OZu7ahZsxXdMjxsOaOrP+IO83vvBdJjf5
IxOKzmDU798C/VTcbfKXbP3tIlUEdsTedEg+z3Fi7ix7miijtIalp0npBD38lpqP
+Zq0dc2O7ccGRabMP8bc5BizCYfK/2/ahDE65zbKX+hDArhJ1pqbNoyvfUCzmWAt
fEzhGluhfA6U4cU9nEADjn0kIxHZG9/9DoSfLVx8vxjhzoLu5dyH4ueAaI+sMf8M
jZNb/x1XIfw2I+Fv08e5ibzKZwNZipebOV7Exe9xmEz2/+0+wkwKAmZt94YCLN2+
Wp9wXD8LM9I64MFldW3JaMFdvCIfKSBy8W+RN1tPQ3mAjfUkbfGcoV90V/J2os06
gQ0gwkyDrqCWWp6eBUruF4unVwXExtb3sSWY1iuj5GEkOACoxjZmt9b5srn3uvqY
EtqsN+SJo2a6pyjNi4VeKvtMhCrVZQBwA6y1rzTCU4WRZ0nt0EHRc3wnXfb8dxsY
XZklqoxSz7/yQ5HHNzuFoiibX7F0fyZROmfYaDs9x3B2h3kWa6IbGa3xFKq2JeZp
kQpte5WlwzFLW2VgqjoPAjUrvp5rqBluFBKpOi+E6a+zUN7e5pkZvmxLHSD0Wbuq
sTzviUpXM/nRjQFGUk9Pv6/XEvJTTtSMOtMJK5h251+SJtCzzBrMnzdQWLry5+Wt
VeYQvLwRysF6ZqFz3sZd/J2tHaYn2ghNwAL9R35DzyQDUMtJqRrO1RYLEE9KXoTY
FaRh8ea/B8MhtvKQObrdqCUDBbunHMEJ3pw7oyaX+NVjJeqWySLRAZX2jZxlDzZA
ZPJ0+jqVFjD8BxDdbhGsev9sObi/cpvqnVsixs3thVVwk2lhl5aAN3WFvMcf7s0q
W6dAdC6+z4wGK/vGLF2jqGcPqSrRpZoK6Q7Bf4aRVCiyKjpkGMQqGFNf8SkoKjX3
QGRKCr+APS4XjA9iLjMwpq8LuNkyGr2XoRcrzH9CJfesO1ugMIXKqFhMW/rtG6DU
v3bO4TPIK2t70ArzxJN6h36Jv2QzU2UuERCiuF34ltQrjyM9YGjV7RXpRgLys8Hq
pyU9HHtCRJaWf8tk3srFbzOLI+6izZwygy1wVYW1jz1Rsk8GXVZtwrnRqstGvx3A
bPUMi4D9B0iuv7SqZQevSdqKbgxTTlsz5gMQHb7awJlGOhzGu+nkF0wovy8SwxKm
4W71/dPueMX0sHtXZLD2U7Dm3Me6DyoaEKXPO3HNIIw+qk5pRjl6hrpp5FxtPBFt
M37Jnhd7521ZTrJDQFEvxK5Ic2fjTmwAKcp7bHyZoxnvQQ7EE+zHJLDTL71M3sgI
o4DVDqLWG1N8LkUl5BYIAdCSEWtmcCea78nSeHkwcM2OaE9If4LmK+ruw72eNTRm
A23yLEbm9rk/65gmMQzOAtTBc9Q7INcaGNdAuu6h/yI2V0b2Sb2kSinRdc2j+56F
YydSAFpEf/5MWKDxNLhnZgrjdzZD3RoeJsoUS9MkfrEUmjS5fz0QNtxeYTj9RbWK
Zxe4mIrx32wqvAn65lPBSj1wRKkT051F8ldBNmxJPi5p7csCeN7SJPi/xB73xFpr
dNq3MYreZrfSgvPyLQEEMBjKbyFOs3J/MnANA8iAnWpBViuD0KmCMBR9wa8QN22c
GK+ZTbw6HDLQcFEzA+8jwaQBjyUAuuSAn2rlWANsZ5MW9PIuTiua5rKUlYZYbLzr
lEKKmP4pti7YzdSOUQ49KILWOmWZDLdYgG6FeojsGmwqPDJ5SQMxRuJyyi0duQY4
3N4xnEjmtr82XGXHlwh3nF3OypPoEppmiep0GCR6Q2oJVPqM+4AWCyuYceuJ5TPc
7ZZDJIQAKKoOyj6SWnWLnO3fjszGAvuGx0Xftg920QYTIK1rysXmc10nbT0ITDP1
gCus4ynCoWAZ7q4IBOFQKTi2Yb89XbrOiBOOc3TfboVsBJRcR3imuk4jawUToAVh
gPm5nLiwdQ4+l3MQAtQeRCRXf8zrrmlxei6cTvUx3jK/V93Huk+Y0WvBBoXkxueC
zBAMKFPBAPvXfKkySRgxV9ph1PrxH1tXhvINKSnycMO0WUcxAQsqK+MUWoWPxHLp
SemJG78DDR0f1YTgKIsutXC5HYGfO+U4N+hTn6h6S752zmUAhZ3SUEW7Wq8uwWzr
8x8eg0M6SXwhmlSluK6JH8bQhjz5BC2pB+Ov27cDYXRRYE3EBjRRJhYp/zmnIRSw
Q2dpj/IPgt8ClvYbrZGb/V4LihfgxDLEgIvoD0uDXuBzlJj7G8ckIiskQosNnPRP
+L71L4CWwBHxNXnraxdR55e+pKVpK5oePG9/+jz2EPeTiBy+FXYgmC2p1FZ/7yt6
rAnDQ8HlZV3yPFMlr/pqdIhSY+0cVo7UQD8fRSx5Ttyu1AcXjAoi7CmI+Nis1S3c
Eb48Ta6vXEf+BSKIin2JgcoBV9Cmjl5tRkxOlRJBy7xJmmi5DQ8Qpb/Dg8PqUc3S
SdI9SbcYHZJg2ie1EuVaJTxDXsL87+gR3X9VZidBGlNYNHYQzkfy7Tv62mpkDh2n
CN66vUCsk/N4JUXx0a/yu0dANTTJppE0E9Z5yrFV8HcDCFkgJ8zv1o7LJY766z/m
DBYLXbgoDbKsRy8mdPbcDv5vJikSI1loGyyhpamros9/pcuTDE2+4H8U6ZyYg0MC
n50fnmYzY2FQGP2Wm2VhA/c7/6Er2f/Dd8r87wIeZOLvFHA70T1vID69egikI6TZ
Oy62iqDveV8Gh0Ngeh49afOHO8FEg5DgxOgEwVJlt1ccE5efWT5QY8zFJAhOZq1S
i91JpjbzvDKj4OzXRFS11WilrhsTIQ/NF/iu0Sm/koJsBm3hT06meIr4g7n55LS5
FvY59EX7WJWDnuz7LwxhDGpQnDRAVtzi8o9amZ5mflX6+46F5my3mmSeeSSh3qKy
RGJI4Mc9a4kagMgsn52r8UFgVl64F3MMYMx8lanXNNds9Qqgd781Fogl/7qXw5yU
nYbAuaIKGDmvlCFpp+zPjbJvH4UPgWck7FseqTC4QJCwltj6AkK+Lyq5VXZ6AeiD
JeO+XdVkh0STaOZyKBNVoF1o48NND3JWe5TEN617Y7LZLTROtKC+KL8NyzwLphdH
JqpoEJjKnQXnbZcKg5Ygwv5jmDPHhWnHYRAcqpDpg1+a4sZHisOb85Hdit1MZ8uF
Oa4iV3zrv67+ckqr8Ui+izqWT37djgLoZxNTTrJqIAEJsuVW3N2+n0jodEsA3Se5
qBodlFY8w9KA2tgNOA+4j5ogFN/hi+yllNproAI7WOYfb5KDaYrG8NY2Stji92/r
jbTcLAFcx+D1z02inlOg0vvBKRz75k5v4TPE7b3bTkZWa+K+KkNidCqcLybV+ozJ
xS2L8uScnsvLqyLsOs4M2fO+Pht4IqGkJGhC7ylEC/KFwju5w+5pqXswvbpXeT4f
HRFdrHR+xLFd/wD7cwvI78rN3GgOKtKbtwBtrNfr/q5sFFNnDCQ71Ae2fnoOp8ds
a4tsYkMwEjW5kzbxawAvPA7Vbaf1CYbNIiPT0MuSlOU4ek6NzQZBKBQDmWOc3Qsc
gAsR66mEuWGA8h5fHUxIRZyq1UsSDyovSvkmeTtfN1s3Dz7xvgP5UcgoTXCCi7Rd
rJDhwPm+XPeQIZvgWMPr9vVeeao8R6YEfi5NKComQg5Azh07liQPdoORSGsz1Kvr
1WCFXiKtaA4ti6uoCF2GdBWDdmJ7NLmOUX25DUfYvnu1VTWKabTgMiq3EUsPDumJ
6LFVyEMBgYtuWXjuCRQNJozkeyvrF+a5EX6SYJxX1w40hyZ/w+YsBBE0EqTjh72x
OzGSbBtUFqe0F8BkkL8A5s3408PAei4nUUOba3wINrriF1KjLu3ugyULp/8OoauK
2UmRv00x3ndgqOIGUGkcPb+egqe9uGizHBIQlgdeBRQkGWgwE5AZr/Ptx9dntq0+
qfOwn/XjDWdone+62J21z82zH+s4f+rhGKp+vwe7p38PqsTRdKGxpnYk18O/cP6W
HVPXqRxuGAr9rz582OjMOE1xd3ynY1K6NbICUOSdyVvqNd0GYJeBa0gktfDtxj2F
B9B0A5WqzfnmkF331z4p97H0cYSxTB60+F+Fk2OQZr0rqyRaXgIgLw3Cfkq2NjOz
v3gXh2JdBguI/bWtcEAJ+eExMf1zNMFrl0OYpH6zz0LqDJUCDpbNWaglFqBWFf1w
bOyK2qp8iywg+V5pzIS55d5Oyu6089GB0hjN6QJwrkmkA6C0IgxyhGuBXSbwI35y
pxkVQR/C+azBDZpAvgqBo5mS8noXgpbkBJIEsyiXwUNQ2tj6KbLBOQ3ZAV75UpyZ
41ZpU0wG3jQEjaKMFMwTzWCdXL4gYUbU2oYC1VIRdTGvewMp0BFH77PIykFWjik8
KvDQeVnBZM0Vv2KQTBvxzsxGPcmsJ47wpoL89T7iTFssYQNBTUv3FQ3b+btpB5qr
uXJfx6KwC1mETI3vcIr57aDU0aOP9GH/VsoAi/izQms0ylMWqgk4LWMTWrh2HR9B
JCmgRwWt5WeGRh/8eCF/0OtgpgO1dcRqciiwFj/gG42GjoxKoz48XX6cxnVdSShU
G6x3ecfgDw31MrMPyCQenpGHYc6M+X/SG1KAzCGJZN/jQ/xswLA/iDsNU2S5uqsc
OAiYpOXiifCtx96qtaaUnmgVVgBgbeMAExKCcresEpmArVDPGYNr4XE1rz5pclnN
GW0Cbfzf30ZvO8QxwsZq7coJUm6btsEvfO0TLb2THneGTSiS1i5nNeTV5wrQZRQ9
sMgPs++eTBZ1fsMvpiZQKxnT/C3wun4W9anJ9O9V7CYYmziYuGLIescACnBhnCPA
IpxVJkjDrGNJDCnRpEMvfVHUEA9i0yOlm/ZblVLZH/jdFEF0GeSkWoN1kh+1QHqU
NyI4In6Fyje8lNRBfhHf4n6BAI6iQ13lwnYChbVnrRhQh08YZ9xUY7sOH+4tyUdC
MIznIWpEAPBY18wJukpT1Vsoi6et3MMULXcjx5850hRuv1qDDdyk2uA7UtcwKD7o
ijgOpJjnAoxz7ZdPXSaPlARHEFjtEo07Bve18wl+aIEm9XudyIrV4fODhEdihplZ
Q3cEB08okvWtuIvtXjmSL02fCfArfJUglM2eXANkXRkWv6TzOeKTZC2tAZzwdfMy
bEdX8YuL2OdqZmohN+EpwGkNpK61lQDkXmh6EvcUqLrJLyPn2MUUcchGTbLTbvJx
qx9q+n9Uw8UM56LiW1XnFhCsdrwe/NKyGDXTIRZsjeFXXyz4Sjsl28E9xO7jWGzw
ZNhIjo/AOacABnGS+DmWI78fS5DqYkzs1QcV3vIOrFFGC43ztGiteRXSGAs/SU3A
HcasrYvpEa59UWDHjcDP73vmRHkHhzl1cnpLJ6jwEp84tuR1q3oYABtIxzy/kGB2
b6V4QvGbKOD+5F2x9Lkj3+eYfWrDjqJPg3y8EoQL/OQsX23iISFPy3HNyW/5DZjH
Exwa5bWwvQjkTgXBRYAnJZHoM90SfPc2l44QBDAlNkqA8Grn7B4rFEywWT7muMwI
qFPfTlXVtd359x5T+8V9UJdYBppKIcQ8hHv1cc60EoeLZZc2KxSMhYCrG/QLepue
cv7gjtgXggOwdOa5ekcu/CIIDVxHK35G6TDcW0zbfU7fU00GMeu3WpBVGmRTGMvM
UIWmjLcFGCrbMtfUhMcBRbGUFP2n/tuTpSs+O7mF1zSR/9kfIrVWCcomutiy99C7
O/brnUXPQbo+TisHTgdE8bh6O8AFTjRT2SUclmBluAIl80KPGwBQVJVVi54/t/oy
jZx6fhVpaNMChHprakkjxihHTHcj6O/0e9Hv3oruW8XXQOW+auPnbWtpn20tDWk7
nHu7ljf49HLxvHdpvJDUoqcg4JLkhw+ivimBbh/ooVHZ4hZi1Lx0fXPIeblmrzcu
rDcLr532QgVqXEPvC0SXc6c9UuBPBNfY9F3my4/ybhLjf9LYmJsGHERzpvzBDf6p
OVXu8pod0C/xL5nwrPjMXopocV5vvZq8i7gwM5rbowHYtTBf5Lh/y2kXrBa8Zryc
YPGKjpf1buvPhBLaJ9FDtwGJ2dcEn97Q61ZmStY8Aq7ZGa9Mbt9dqvf5ZuetsaNo
4w/So2i4fr7tDNAOVKogFmYYN00w1SWonuhBDliVRSMnPFCIltE6PFpzS471kItQ
TEhonf9KWgvyTi3zhLMVZ7+JVyrYBvBMS8wchR3ezJ+9R91Ktzl+/iwbeiELT+GS
UrIsoIw4XVYe/YpIatIH8nMyIdZ/3qiPHKXuLgCZbPoIxCmsMTth8nDCTWkCdess
hyAPd4El3wYCDLUqEreCubTV/XVELBtA2OP+4L/7oeSD3CZ/E1vIv6eIUZAtsxah
B29TlVWMo0KYHuMPPpAaZ2zk/9hUmSxkfx0SsEVEsh8KLzURmNjJuPL8smJf2Zgt
FL31HT9hX6QyzzBAvXecsxusk8vDglx8n+mCoFBXJhBE91IW4JQj2fYUBw6al9b7
YU0anAS6F1MsAvE7tWXayoZwc8kYCh1K+8N5JnWRMhkEgGeGQGJZH1zeRUyzYDrF
J615nEyeYpU2VxzR4OMgS4RK+G99B8uxSoHl51zwKZO5kb8CybRDd44N2qCO3++p
pETHxaJ/0AKHP5oRjjcpLVWJ03Zf9Gwv38xa/NfHE9bbupenjj5ylx4Lj3XTvlRr
20/nM28FOM2/Y+cypzjLQb5H/L+NG/4r0rz8fgb+I6LcxBk76R4XEmI4CJkPZMv/
5Fr28dWT5gHfdz+M6RnlwSuD927+sZiPvtTiUWTW3JOfcw8XX4gExjxZW2Zt0Aen
ajsdP+fgossRY1BY1M6RtthW39WBfjZOKW1v9LHMqzTo5BDL/B34XqJr+xaj1hGq
+wG2p/ErN6DhiMig/VTMX9B78c7QmxydTIDAI5uAHKuqdRdilyQlZLH9z/568Vnl
bxQBjpx9Ifg7Aynaiq8rnxyub4lEM6CPpi1NMA5jhQ5tjoetICnsPYieNBHZDW5W
jLVS+GJIpkPROcvimDRjcTMibnA1ly6JvdgLcdgLBzMQL/8r+cB6YfCDsRK/Dnof
3axZ6u0yNyqTqe3A4tIExg6g31XgQbzoFSn4yj58/42BELrHqmKMEeLwC74Ym1Wd
MnJQHUkqvO2w0iBWALCK7Jq6F6Ob1aDb1xRSFj5efblatYZDB+35Ny/O4HDA2l1e
I+ym/74kQZ31imOxp2il5dbMh99xC+Sl4RdSdI7BCSClw2Gp4aEwkNCWyAIEjt8c
8SzQvqsLW+v86PJ7ErpwWyGeFQ6NkrBjW0bm6+regyEuZ6xWdOFk54/cTkUic+yy
bDZ63Igop7ghzB87ZcyMu1vrzlBimvOIC+0iOriECnprO0kzEAJHthRFdv5RlSsB
uxFGDnoMhVbhqxnXVzl2zaFWbs7oocH3qqV2JEbCvwYDt66jgL8/cUbpIeeb2cB/
CLr5tUywjwMk7DdLdv79ys77nvvdrnv4a2UbFLltSLPKfic7Z77TTz2QZLXeRGwD
XWPVr/w8pTGUTnucZlmfeic5hFkznh5qTlF49u7PSGdjkdTHPrijNEHk9tFGjfUx
HNi9SEzZO6llNG96i9zkoxJ9x2ieticpZQZh8ffJ4jKCKyTMZ+mPfSCM0f/KnwIH
d1qEDcdLXBPaMT4c2YE0NhkfHdo3l/cKDhkYmXfvGhdgBrZME/KmgkD5XNg3kLwV
1t6dt4EnVW8HE8im6EOYbVZkAOlIFi+z6KTDOCZnCgjMLnPnWTubfL3Pkhf7RS1P
ufas51pXDJn9Xykvhg/Ib2XgSQUFQi24mxqCefTHAwLb/biooh08N6N1+BV4DdSS
MenNk/Kmj2DfJqz5drBNDnELjw9LJG5zcsEsFSSBtoM1lOkKJt7uHazcbAl6Sh8L
RdqOEfdTaG3Zw0TG7jWc/8ro7eLqP47Bdr8LS0nQdjc7xgM9X8stn+lq+H+CzmW4
fbQeLWxPI2m8xDstH9KP9RsJ9qWl4mzEMpX8qHn91BgnVFZmYPteLiQBK1yi3Q3y
V/0MYTl2+ZUVsJdEp8nu0605rEz1zzWd864dfKLPyAxDcIJpT3eQy5NFBZ8GYqWG
emORWr+l6qtBqnet9WOCzmI68O3+1z2ClUJyZwGroo6vEuMc2/dLigV/uwA2IKZ6
zAuvJvxxW+F+GzNQhZeg+uU9dkmZ+EQob1DlPrFfzaTGNn50HqnORNLr1sBluKZE
39cpueO36+tIV9Jy+9VDeghHAa2mIWHNTLK/d3HoR3bqfEcTaMZYJVIoX8FpTZDH
fuZS6ZD0N1ypB+2PIEP5Aurgm5wJSyaogBpLXmr/h0PmcJmsiHA2jDtDkkJOPb1v
xAJn3wf/4Q8CeHZc3+xXa9Ydgjaf2C2lfpaZejt8mg4KwnVi/XWp8BiU/lRQWkIM
WqQiqWklpbp+fW7oi0Bz8nVuWiMtPgXNtKnV+hOTjnr9N2XFWPa2maviDCAOiyN4
983nskXkbyHniUfIoeiktFoRAk6IQuM21h8E9bulzqG44ocWrnGfGbCG3DGmI6Df
+dYASI8JyRa8PLx88Td5YVuNH1DO6vsxDzFjB5ahwVxNfE7CrTq3rwqQwWo4wc8X
v+7s1wn/CtwTB81593KIx1nwAHheIIYW8XRa9MyLxRTtjtfkcZrW9XexlrcfNzXl
aNTROiQmnMpkBuWX0GCmJA0qGcGO5xpy0/grTHN2tt9FH6L09RRUQw13rrz6TnAD
VR1Ytvmhtm3HeDADszmi67bsX9y8GRQu588pBDBluI/SVfxawLEvPOwlud2+gBlk
8nbeQNwp+RYhlVhPKEsunmMD7msc4xMm24lrxIc34TkQpyHKOnI/UdNnkPZ1UcPM
kzaZMD24lDCnvGtSrm+bQhxQoyK48+xpviU/hSgbh6ySpsdReNlaqModFHoGRQPP
SgZhnmwIMO/T8m22W8kKOAPNZjqwhXrLvrfyQNegEm7L02YZ8+Qb0Z2Unu+qbFoF
mcqnEQ2u4VPqunla6pvIQyTcxSvrqbNBcY99bTTexVjmxxVbxL5fVj4w4fnRFn3X
klALlUjkFdK7dc/0JbH62SmOCHUD9qPMJm2DS4/2i0g7Nq7vLFu4/V6rnX6E7nmr
azt/xZeYWuMx4z5oVvRi/9LdjkL41ER9nCFTpUwWNL1gtxCLG1E3iPR37PZjCwGf
l4T5Gxos0LFq4XCdU9bqN3en5JYnhSywfDroF3l7reVb6UjeLdsbEpAgnb92o+OZ
IvxgJMQwDfLU55nv8YSK+vO7PFeZxbYpVfnkyy0lednsqpmVSluQ9i+BS4dypjVk
5XVAN2iyGXx6roubKOMNTX6luBW015wJEWZNC/wlLhGGwmbYc6LCbMOgxDCkt7cn
E4LDNRSbmBNxEHgvOlIHsCS/7mpuYv+qkbhMMzekDnFL+BMghgNIrer4RPLEFhgI
gCBX99491Jfc4+g2FrHBN2npe6I3I+bXcTZvsQC030RJtScD/ENaOj6i4tFgX5zU
ANSauGeAF4tA0ZdbnBmL4l9s21nKL6SiyYHzFvFesT2XDVnMJ0cYebuTEt1xP1kj
OqjB8d7QdPCtY7ev7aq29NT3py+ANW4gCgAcMUkKJOLQL3l7r7B6SUojiS/fXXJ2
d+NzMdrYP55TzlC5ZfecEFWXFX22qCpgCpqyfh8x2c3SYm/oSQNaIVjEb8Jraw30
3XgMeOzVpH2MM2Vk4We/E5W1y7XFn4Sj7pk9QWxR6eKH3zKuUx/lw+l5YPHBPrIg
YTp2lFwFhoR08snwGyg3Ig1vljngNUl1UEkAEVfM4WYU/JVrxt8x8gTyMis3hI9r
dC0bBvuVNfX+OyulMPSyOFE/Njo+0Mqgim/4J7r0I4z00Y7VLcoRTPvR2spSis30
b94CiBfLF5o9PeGA4CAsV5mLSHmwFa7XTjWLQqaUYO+d1atWqYavNxqJqsXouT2b
iXqq47RR7yztpClpw25j97+kFWwuptsbSH7juHwNQ5/IiYP4tG9TdWManFiqrFxW
Vn9H1Kzcpg2fBVWLwhb+tJK3CucIFPWveVE3CXie7qZm/ki9qRA59O9IhNOKmt7Y
edZLPhb+klftST2Kd8ityZEt2es0vSV+U5BaD6iXaG5G7114oLcIa/xu5c/AxFcq
jzoxRHLJKnkSd32PJQBlznYYz79LUTN4BkoJ5X1ghDWFwVKB6MKFZtiMDbcxWVVo
etUntfZA8k/YfgJ0UqSKfwmUezkgEDPY64BqzPvylyBbWCrSD9ALyP51NrYVp5us
veqWVMAJHB4jKbtMb2l3epRkElPWj2B1ZMIDlq79+Q5HoH90alUPIYl2OL3pqamU
vdTrNpZWU812HFYyJEOfllAQNOrERkEXKfGhRNC44Gtr78Irpy+K4dvbGnYBiWOY
rDqHL2dq/T3UfFg9fHalQ30ROcf+1iQ8e5x926xVjNPPweAk0TEadxFUHORxi4Ua
DcvD5G1yFAwEpx1lHKUnMVZ4XHhs8GSz/Rfg85k8OhHB5Pk82LOkV9308KK+6Y3I
3JTS9PlgEXlqpqiJRX6cQpMrFA5IO16hrS/beccnsBpsnLQCVfvCT1lY3o4kNert
tbl2JBAMogaHLuevQuu6s4Q7vDrBJM7rRohZ+Rn7SBvrBvwnKo94r8ppRQPjV0dy
I5svb2dFudcChsnKfF4I3AJCdUIqcTizj+Pp3ql5V+EZXNbEjphap1bSQlQFtwcy
IuIcmT1pkdBoLe6ornVGhHahNpplhkJ0UUez2Z33GiqRl8g6ZhIdl45ktJyV2WTW
YYxz5bS+TAhp/CyEUZ6KuCfnnDq7isfG/tLkc5BvwWnUKoj/+/ikWOEpX4aIZtoh
xSEY4h78QYZcs4f3+3Ir1Qn/6mCMIqb6r4S6Jx6Z9z9ZipqIVUimbCcQZvlykE50
TGXhxigfHyPkQnjThf8MWWbfLGvPoEKwZTC4pZTjoYhhFD2d7P6jsRFihue8/qdQ
+qhcjo45L3of7kmqMkuOmkWzZapGey837MSmuHiBKSJ1aUbuWFBnawkAICpp0PlE
Eyr3L0NIGCRlFzzFHSUlUjSL2PVdfJVYsIVlqlen85aF3k1SZv4tOlBlOm0GOqVr
srewRgSL9Lu3v5haCVUzlG5KRRpjdxCmckS7c2IeTJ3DEniaiyA8jCaWm3ZfRCv5
tpnOqvjN3LFto0o3jPZvk4fbjHP9vTf6knCJZ0XIXxd09mJbqpYdfiiVxaXVt2N3
3eGpeY86EvG/XC7yzRFToJELNIYGThFoZaMV0YPC6OlL58N4RafrZj6oYJDRGpdC
P8oUnfvYH80i3/FfVh8bW/hGu1+1RlULxo/wkew8RuuKSSZS+GuSTnZlpkb8YS8S
0/+fqXlesntX7qknrdw5/LHNrZc8rc5rFQgnMikjpkpmTsgzR5UYZJJA7LNdgOVo
0KNUUjNLkYBnQY6pBzlZIRRiHhYTGPdEuNwEJQ4jeaREr29f7mi1Q4fvi0rCSZAA
ssAF52MtMl6LdDPuqkEJ7dZ1Y9BNmBnxYFzxrNl6PAGjOXbzWT4UQE9J6plZ+k3f
RFj9q/Be1geIotu/ItuWRMun5QQr34Vum6ezqUKzypDb48NrJ/bpcxrlHPQUuiZz
AftOLzG5+S26P45cMvQ3CZqyo1upwiSXM0/8clomyspE31wnwCo89UpRmFdV+IBl
E/jFIRreT2TLegn/vXRHSpx5cgANeUWfzyd1tmD8/U9xiOwINg1kb8lpdW4c+Iih
/+Vu/9dLH6hcYq4/3TN9jyzGDAWW/y0pPMy27zjPv5S+YI8d0uKHX2LLsN85Rxxm
L9m78wsT7YTcaHUXh4wcqj1fBypdomQOxPTsHtEaqAALKc8bQR0+XG+S9zocbsJ2
H0eohFdKBv4N6f2D3BZiOGgMMsYAaDtiYMkQKjbtDMLzegrFEcX0BYUkBV7m3ZfV
wP72QqYCr/V4HiIVPNipRh5vS7haRUGvEpJYk0IXZKKT4aJSs8UxIbT6hiorjqEh
bOvuWizBkSKjR3hh0P0+DfDh/QLTDtzk9/mFydfbZAE+BWSUvNFCYYumkcq1mqNW
xAY+OXUItAa5bllR1NUuqi1ur0iyW7j4g2S9dAm3pc3T56OLMDG5tgzqtHwLVhPy
zgBuU6yu9y4Natq1Onupc+CB4zVxXtqGNA0uejkwju85ixjfymF14tKVlUnITnSn
PW8kycjpDFgUgMnVluAHcpwagTEvzAn4nXSq5sscp9oKpAE2Uobn2U39MmrsEZnO
qiA0VyPYQc9CMNXFOczZAps/fksDyk+j8qxxT8CtWpZVeIPoBqs7Bkjrprny4LU2
GergW0pRjZUrnffa8uXKElFQD6CHljCP6N7qcYlw1gAtAk6WD8/oFmmifEKrHzz6
ucVV8WIQCU4mtlEGwXBeVqVsogE2aSJNt0wIIpoD66dwAlj5fGBzB01H/+1pivvU
8qifroiCwF+S5Ozakt1fRn4ORWl/EbIgXQCS8GKmYomXa4BuIUiwpVapK1LVaj8W
brFP300Prq1v6ImDvmklgHX0hK8EaKNEPXfsALUVPMMo0tzQYEDiWVIODp7l0mFb
ZTdRLi8Zdjro06l9qn7mf4vkzkVvJb0Nb7E7Zel0zk9AUTloND1MMnu9X9C1d01I
ySHVXl4XmSZegxrcDHMB9aUQk0EbwrA9xyPYu5KaouVG8xZ50191hqAKHMIlWz0F
68Qe23gOe9V6qnsCsNn8hjmYjsDWeumo13VeKf2yfFWejgIgZ7XeO48TqBz983Ve
YMWDdveYNhFN9almOxtkSCoBbhgYm+TanOfjm46if106NZ+axsBscweRzpl3ftZ+
s5G94hAmwxvfzAqGVEukmxPww7Baj4CWD7TrIYl1UlSGRRvh/Sb+duuiK0S3RhxX
yZUbVBeYQ54lAwELK943k9LW7OtOI0tXF5jq3C1SjXPBUtTxldBxjpJn8eMwiMr7
KPKbY0zoJhpWV6V55dd7dGrDFVtWOkCtrtNTiEZf9OzKH8MgjekBTen+lNzTHc7P
6ctoNQEh+fvZhZc2HT70J6SqnEbMhJiF1vo4F3X+oe4aM8qqPKG7Q6kgJVsRdLvn
JE9SgMCVNSvFBoL2oSBmpeEMZSLuNYAMcQn7NKpNfpEKH3PUlE0wkjEZO+eejZ4Z
DuUw20MWW87sg5aHkw9IMdsU6V0jUvcOXi6+nj6udwZKqbpOcvsSbgQ2RmDnzajh
uH6TXn9vC9PfXVlg1gPwxKX3hFFGek3sDGcteA3wGHNQjuheJ8PabPC8yzzXdLmL
w3EUxzyExmY4FwQ35DsOCAifb2pvGHdg5hKSXf+LiZF5LcwhlcxAfKsf7sgisovN
7cJS/RlLkF2ZCOHqAQmnKVYJ/cX3M6SzVyhhmAieuX1dpcIOUqTO5UGCDIP9HquE
hns8acQpKYjCxO5YlzQk99vaQ0I9JJ2neG47E5CBoyhv4lw4FCvzpNvUjvZIAmzg
IC6mLwsAXdcHfq4MJzDKpgLbMml3ls/nBC4m1LlTsveVMavMEvTupI2QNUqP7JZ2
nh+oSiWn27YMAKLlJckn9PyRVMUsjar2CA5uB0SvXBXkgsFPNhf5fm/1G69u7tJ5
pXalRen+LsWZePW+MkqWyDGxn9dfHTV1V2QslV34pAMU9D9GTSLXpj6NeEmvmFCw
DfkFDGYqeKec45W1WJFgW/h/WzTJXyHnA9bFt4cpER9rEV01ZpEYySomZT+p8SYu
oOs1lEw7894XlABfWSMlQLMP2mBXtijE199fb3sjXn4jiwCB5qPHQfL1MOWajqRr
rxsNF8vHOBnolr2E6uVcY3LGk7D4UpiIDHTyTh6d9rqcEekntEf4oA7z2vQ8pRpJ
CVZASi/md9OvO0Uew9ghTPcjk+BRZfcLrozY5MuBNQg8yBUE9Kat+r2dr239yelz
sXj/pvz6kAuCEJsdC1jh+YIIK2yZWt8jvt19kchVHJhdOZP8iOqPK+bL0y53u/Fu
SGnkNRe8IHgkRXzrfzqR4487nB/4huhrmP+d6vhloKjBf2GpEB8P1Elte2fR6WSX
K2kwXeVk1AH6u4nG4GinGPiOn7bVi4EMb0zp21RRdgSi32gdq7RavgTsPX8Ikih3
n2eaCC4Zj2G+SWROOMXx0YA/IeaEbKnPXSj0iAHwAc+01EOQEa8S1ZhCqjoq1Jvh
ONsDjCk5Mu5/+FFj+Qv4XbiccuBr1X7PbLP359wvtbaE7/r9Drt4zTzvJvseKlCx
y6eH49mbplRVI2ZcYEzsU8aJnSCv68sT7IKxIWGkbjX7gAcoApFcxgMPbi+y+hCa
/fd2QuMrt3W2ywzxG7oUuXSHs/WADeyiCpSpsMs6DCPHyN07C/vyCyvhgFZnAUeT
VvDRihRj7hW35ekWfUzRYRcDdCxZG+S14T2AuB0LXGLj63CEOxr6k6pWvhoJmIJF
ESPRCiKINEzkO0J5ZCi7b6KcYDgYbOGokPRcNHCFB7vHBWGOZ8+Ctp5PiupTkg53
FYsSOrscjv4WipNKPXRpnvP3Ipr9JUHu4irfKazSCzZcfZtvvAG3i7a7qfcMJhob
OTCWi2qTFxM1Vzqdf4hXVIM4vRiR4LpCEPJxzppZOz0YSz95XYLwA7EiyRhB3wKq
PK6otZC/6LeWBXa005YZKyGIn/qLtdalQA6M5G/XMWu8rDt6VefoLjF6pEVzDf6c
Q/cPVB4N1vEEK1mL2n7kHJrvgsO2mkG+sXC+fDt0tHT2QUEmjaJz2OLJtgHyWHy1
YF9Dg7/MZZZoYNxz45Wd8bpvHOgFJuiI5JpkyxyQ/Tp9b3yM68XEK4Fxsy+MI2xt
vlSywN/PSXE5hdnv+fgnMsdlWkedey/vEu61lLgSJ/QwRgpMX9Q/wiG0fvyG3q/O
bkmn4/6ASLinNWeHd0o5TDHnWRQz92VguDG8UlwSjUoyuoACoK/nYJ8PQ5Y+IuCV
NDM8FnRxuWIuaaT9kPLFlGaCknUBpvmA/m6oirDaBojSqzJFTgUKWi7ItGtg4qHp
07jg4InFXiD47mWpNkOAjlFrsdw+Y2ie79KafLegniwigk9ihlw+rT/lfbTjHqoZ
egS5e+HSQvmQIovF7feRhrjmzzia/VChfwyUblpUgzBoOW8+I9vh6QJx3WVZieZD
CR5OdlZ4w+chZoifnxr5z2netFAwBwNFkCpv3YcJRpEhFof4xxiRCd9C9+2sxYsB
M0t0hv3LOwHBLS0/0Dfr14XkZnSbeiAOgWplZ9b9DOR1RIKb9tCkDQb2sN9ufkw0
fp/UEJ+fzqQEG3czjT7dRFTet12HjXdAgwKF3CKB1007ul9k2bLwS9T5Y7ujeUU+
2XQgH8o5O8geMOVMZ2C3OT0UlNeUQfbPO3QGAtdqEUxVrMYHXV0ypYe/eLjy6xHs
Q5cYgimWECIrRQDN0D601hmrkaFQm2NadO6gy4PcStA5m0tDCumXFTDtdUcoHvnZ
twuF5+A7zmVXYemmFjNF8vje2DBik+T7/caynCQpVxkWsphc98psqNdduX3jB/D1
uTVGJsyL2i5qmSmSqP3Y/+B95BS/FlCloQDQ4SUQX13XqEbQlLFMbXjHyKIj0DkA
MryosXlZIRyyahe8sTOjWnyg4ZH+5XNj4P+2UikNQeChq0eYKMu22kJhoD1ageor
l9L65eZFgzl5S3oGWAKYrlAgVr5xjoyXDwFwzP41WuNeXhAQR1QgwNAwkoiNozIA
1m5SsiHB9Ps3QoedF6C+uQ8UuXE/yQYG5eP1WlpsMg26faAxNawN+koY/0EeiTH5
G/f1YK2JiF0UQWcduUueqqS6vCFpsPsH96ifqEAVraNBKov/9tWK95pTMScWxW+i
+OGyiG3SRbK4ll+hmS3bhonf7zopdHQ98b7uLz8WAeLZrUx4lWTKlggffy/A/6Qs
81pvdue5sTcBhXpVW1I2M0w4Ag6bzI9IMcnMRICQUcCoJouPtIOAcxkqNAb5yXYM
fMco9hwkJc2Csl6IR21Fipbpp5/JuxgOon95Pv3UBJbmKbpOUe300qauQDZxl1lE
Xa6/Jbv5MXPqe1O33bb4ogvJ+PFywwq5VfPMhofvKzZ+3yeySsunv8AGx48RIZmC
Y8/DdE/Ogws5TqUwfMP021IQ1qXwbYNq6mPpN1GylH7CJrffuuQa1XAIe0YAn2tk
mH1QrZqgnmSU7Bhsda2o/1/mmWkAkgc5y13fBY6uLHcd815pSLSUa+wURKM//j2p
YlX1LJcl+7Wtz+nBJySW4RnCpxPSnoDalHSmTwd0TB5Ixc4zXhBn7gxIgdgAlpmC
rizNt+Fb2oTQl69wc8oIWVVIBDOITtq8iyjfMITTSdB2F+ZSf1eiLljLXs9DI44O
TiJhS7PH2918WyD9obFbC9v8UjxN06DOV07l9x6aD7XTV/6/vGzjO/JRLDh6p9Wv
zxSahFUqBl8YDSmYM0EOpmk4nFIG3sYjzEExZNs09R3wwQyKETHe6d00M9V9IBfD
KA9Q3vLLdlN6t9VH2Pkbr7sOrCdapAbUvz1/GUJrrl5hrKT6l7A5amdZpfk/Pstq
whVeoWJ6Ldv6DN74fK8eGSmoPW8tEJt1t69Cg17sA2GJh7g5YzHdcWfqEEQK6XUB
E9jwoAwPQ3/gX1GRy4cRlJlqZ7bZ9nynNPB1/+wHJWHRPg8eV5S6k7F+gXbyNWYC
X9YJcwuX/jNVRH3L/H2rJcmhtORYbL4NAZRawPSrjWgWLdUwJXbeOD2+/xYMvcWE
Ug+KYVVwdoyPcB3b7Egq/AWQIE52jR7XgsAon4BsU2qKOB2O3P24+Vt3OF2fUeGj
QND5JUC8dVNyVO2n6SFph2d4zGnTgF/BMNpllb6813BuANEqHNO5HRq78Inqc2+T
5tHD8f0HBoCgUhTXKoHz/8ksMnXtR3AJaZi3YMrJSO8b7UdpTrsBELVUO8sfLrC8
4KsnLfGkrz5BSia7qYrr5IbStBJ3cQazkCq3IlZY740O7vad7RVSgNMsjZ+sZ7VC
WxDVoVQuI0RvojhkkVkdGLEphZYUrI69fZDOxJvlzJLi/d4G/jUilzEJ72Jr82ph
ol6KecMxz4ae2hbTVCUiZgTz9NyttoI6p9et1qphbAnoZX1qsNHUKr/dRYVLUEfl
by5Kf+3/anWPBoGNLv8d+ixVwmb67IdkePdFKl7iorMXg5lG5RevmkGOW13eWmTE
oOOvkIWyYpD3gBJaVk4X3E37KQM6GkPS3e70K7LLT0NzaM5q20By0zCKBcGf9AFo
Uho21mjGofAArIMO9LYhzjWeue+w64yP7zr41SpCWBwOAfIb7ZnSzB9pUoz4s0Vr
EebcapYij4twIgj0zjQVgpVMt4xDrvlY0LGYPKA+gfmQ6qXhQsvGDqQy/ZjBIQKF
Fn+NIgFcnMJgpPU8AZpEkIGrxfRBJLLE5IQwhLDpnVwawLvscw8kuN7KATt0UOun
7YaCg3wInxqNtB/9PY5R82hb12JWp12+/jzQKC8RHzUEos5b8A7c4tu4rvqC/fOF
fSBnhp0639um+Miv7QZ19AExqejnE/s1wo9AKlihm8JkY94aVshrPzOq6F+NbP+H
ljddLKvDJCoY5CIR8V5XHAX5fn4cA+TVe8Yl4xKyZuwixkLyLt4BmZRKPuf6I6/t
bW7BoJXSy8KTDC0LGFp216IG2ORkr19y0KulyyRbAoiE7aheoc7/5OkgzIanMSKz
wDH8xP/bSYSZiNxrEpcGBUMUTOdp5cUXwKMKDcP10XotY/TJOW9sfxLeK65+MSZH
b/xjtyc+jEi7Ua9Q3bsjI1dW08uTOUIBIXH2ziHiTAV1aPr/2bdMo/Vm47FYOdBT
SYCbItcW6viRp9VQxbcF5F8TTs1ur+AETG3fVEyGodPqMGHlrYmj/9y+vfo8TBnS
A77Ens8Ygdt7QPSjT2o/dmtM4GJ+kpPhw+USdldfFuHhjm976pCpm99KazCVxeWs
JlpMz+U2JXSGmxothW570b5O9gbkOyb6SD8JXCNsiJqOwYeN7iVtAOQCXvc+TOfY
Vc6cVGDb7r8OOsX81TrrdjqZJ3Ulv0QDHDFhl6to51Enn39oVaJ3mAorVlrcP8Op
WJ4fsi0w5Dj1CyAlx1K/z+UtyzMkw6dKElV6FUObb9HcTSeq2czgL/PYPScn3mkt
h0j0TBXRPeXPqTUn3N56pZlQZ+etyRc1A/CpPsqsDxnTTSB9xrv8w+ciM38Qh8yL
04EluCzH5cPnXaTStcWFCFi1Y3dS6wRWV1nWrtOaVGBmlxD22EkM5rpyhtSKa1H0
VH2OGOMdz3yJv/Hk44+rC0owEikGY/NqFM8YGHhLmVIf1FZo/6fv1GJAwNyPkmh0
x7SYwN9pfmj00Yxw3NKV48hjFlqzPtM/Ma6L4OxrrTqUZrWUwmDRwZTjvhnubBZ/
QAVw3fPbnzZHe22dX1jNcfr9OwiBzySZBo4xWDp3ppZds5Wj/SuGxdKPz1JU1k07
NRvInV3xhiXB63O7JMa2MR5Fote7LNTzzMlTeHVmTu0QXoqKVUW9DRW19fnzIs2S
nd3UpTfEMuvsRm9Xh7lOqAzdYtM6zGGalPzj7C49SCOGN/qBAhgn3tXaJwRwhoLC
ycTSUYsOvpDaiTdH/zoVUysp9If+LESJATgJLVQlLR0PUjssTSh7suswKvUOqspk
xwT8vOsCE4GL9juPaYw20WoRGZqrqgRWSX+2eGXSHaSKMapWAi0OK4WavSRcSRmx
wHdoRGp6Z0gijQ8mHO+uhOAHtfS7FjImk23GsmqHLiMFP0NlBZPvThQgsWB8cNId
LbTLQ75CQpbIs/Cdkt0VEgCP+LXpCalNpdu3BM2CQ1rqj2gOpOrd2MhRju2FjWrw
i2JJmRjSDdNXx/FqH3eSxJQbJS1Gq4lygh0TxKSRxhTb6DnHnSZh8V+zubLUK83e
DMPVj1QrkCbC7dgROMV1+56XvggERUFOFihqRr+yUYoalPUI2qjAB9tBbiYIPPCd
9Ox33T//8twdfeN+YK/JIfD46VrDOVKU/CTkFj/pAzcZvfCZ262GZ8keaGWJzqh5
Xpb0OwZDG2fypJqFKyCuXJTlQZTzZos+6nr+781o1oROK04VCamY81mn44EpjVDe
2Ri/2siI6FkdEZPAHUH93G376DBddqwPYNcRpRSYIPS8KaO9wl1/GBTQrDEKJO9y
C2ZbVvtQRpn194H78TwY1FtbOQSRwOjFQa2x6+IXbSZ1WB/BJuHU+MUrsru7dMtk
iqKCCCbm8ExqN1XnnuTUEYJcnXOhmP/KBG6WTFdz20ZId/tyYH7Scfw4Op5st3R6
QuAzoUFDYTcClnb7d9k/HqhJDRWqW/evGvHq8SlxnjqytcT0v+vQZazagXNYA4C+
3TTjcu1vdbDcNL8dy2PtngD46ya/BqQ6BYadfO8IB3drFswdGbSPrEbq3Y3ScQvH
dQAi7YpG210j2UTYvA7xdaoYxyCJNS0PYKDLsxUBuwHlM4e0rN7B1lPVRA+zQMnz
H2iBXoJ0n+5ogVMvvZcdSDbBcKJ+3F8fWSmVS9Q8GXw4dr4uXURjbex8Jlr7/MbQ
X8wsJEv/TMQmmejwuwY8jZCTTOIooQtmWqZTvQdKQ7MOyjNS7yiaXI6lxlGqshOM
xynBhzM+N9pt2PiUhPS0Juoi36hIUCiTtenft+hJZ/+Zu1lQvPuhSuBtrIi2oAEK
c76JU+kXNfsXmuyJ2KE1K9UNGgBFeOTg0ZACsbXEFjpsAvHgKTIG1mCAxvzOwdz/
9rJU0a0AKw4HJ00KoQb/BYUTil6A5Di7m+qE0oRTNybuxScxUatKquO3kC2i2OR1
k8uGod7kJNFzE+xv3QlQciY/bcvngonRRESI91J6jUtAgHANoFcY2Uv1s75QcZAZ
SfvGJ1dJKyn1N73iwHGqXvPb+rWm5mb+qCLZLsgtF6oCj0XGMfUGYbuaoiz0WHaZ
3RaQzOPIACRT7ZSGUDxbucXyWREnCk7mELL4z20zHx8801/8hsBxTQGwkXyVPCVQ
/DOfNHBQEbqBuqqw/SxHfzFVDf2SsjdIgqkcBHUh78/IhDmOvstF/iZwqYhyvglU
QAcJIfrz8nVaTxTe99tpv+B4AFO7A3dvgKo9IoJpg3+uob5z3YeyMu3x3d4H1lDu
qLSbHbsVmWnXLNipuR+XHbSULbEXbHXC9OuM9wkw7P8im8nOL/viWk64ueG1s9Lt
zJ1GtgDf0ZrXT9mMSt2vVj9X44PdZMDijFxk8SXS9TtcgsroZ7RmEjA79M0AlOAC
QMQr7V3EPFwKsJPLdpVfV6C3sOWrDUrB9V8cYsCKy4fgi7agVkdxesZrARxLs6gI
EMs98OvTQyHMpYlHPlgCnFBrQuludQKgSm0NO+X2ciP04JNw9UK+nhwwFlgwVvkM
/X7gQOZ3n/LP7cOPm4oNt5EJCaPMLKGy+XaIz679FTF8j4oe3OtKwS+PchZvV4JL
ak7PT5CgwLJkVmjRlNzMeXfcKVIVZbhh0Te4Y/vvzLQ+s2xtx6uGbkOFysaFQ7t4
TuNNkFej7+ew5WK9dlgh/wvyTJRjeFCgaKvHofX31KQeOsqxe+gCIoSQJUShRwaG
hC6PwarpH0Cl9HRj/ogj0dF9BvkEHLA8mnRlHT6c8OkdTWocvfEL/qgAVp6JcmVS
J9F6JrI1F0yAE4HhWzeNsQdFzFKPFKhFOmNVvUKqOjRthvVYC1VhW78WxUoqbos8
NWuaBr5yRsJ9hJqkfsfR1R80s7YjTrHRbir1mgj0d/NOpbhY/+1tFKtNvr9N0ksm
g9fN7Tdrw2G0sH7mtIjx/UMYZhDn84J4T3W1ps895yzL//ty43pXPaMu4q7IgO0k
U7OXn+92fCBYydMVjHx1gkykeHs8uxr0EmYdaacN4upSqQ0fNx1zq0yC5drSf+y1
KAY8TnpS4dsbko8t0OAkfJAiR555na4+/7tECTLr9FXK+zuZlph6eTVNK6rq4hxP
laskZ20FCLI3QA0Zjp1vuCtxBfAxrt2JvjXZzPVaGJL5drJcsuqF4B/kWjJv3ARU
dPebWFGy5KmlevTDSEBvpVj3jKkbp/Tp3mAsKSmIjLHPcblrljmkybfPmWD67qNC
6x/2uB0tTx1nosyD6cvG8m/C9VADBzbz+T905rC4mm+LPSNsQdwRtOHT3JnuLDBl
f6QKu7AXwvgEnE6XDXug1bwa3FKmli8IYXBCkAIWLYJ/MQquoyNWpn2zAsJ3XpJd
xor4CBwec5q+V7O7pf6S4by+LggdnmRtwfItBet0aUQ6RzrtNnOSzHH3Q0D+dhRC
XmsSQABe4w9Llbw4IILEBJeG8Btfg1Tiq+++ZS65JLEDTjLMhrpyqhs6XASj4VCB
CT/xkFXMnCwKbODquORzKGo6wslF3H6zKwqooC99m/JfLxnOIFzz/gJTmm1x6PW3
h3xvtTZ66TLc5T4cAd0nOBtMe+VpyFOBWbNrlBRFE2RwltXCx0cNkdWWgp7POfxd
qe234NvLtjNDy9o8KUwDlJruNkkDmUr1xClEeVRJCJapYgN+eiwlhMEIAEs65opI
xjvhDMTuJOYa8oMOssuk81r5jBvAsOb3mf4GNyPX8NVl2mS/40TwEu47Z2yoIMDO
irzNA+y3YRgBBu27U2u+/uBl4k3EzbIST1WR+JCiko+HRdZwJi6uly7A74F+32EC
xm+KRR9q9up4yWr4emzk8tNasqxggTl+X/N8RM/HzBNHe8nAvN6iRW/ikfgYd9TV
D9ouriip3CDVR9dJGptD0/ZhAxurHJy15cAR8D+dWw8G+12Bj/qhrKQMOtv4BA+2
Xgcpaq/GEWjfYpUff8z7lh0TzOla58pvYCk/prTvHV3UHTCmQKdARf7rfT626fEB
mD3dUd8eKPNBxdjHBomz66zZ3EyAmD9MrDETX75R4a+HWHuBglwwTHhQInJ2sFe4
o22I3xdsSpq+Xua+vv4xY6eGjhKVGS3RLWuHqnNwgoQvs5Mf5VdxJz7qXkS4sG0j
tXf4oIUWIZ+G9SgWGIlJZBlc+RpfVzRnz0QbgAZHmoY+kqAg5QY0ehMoPRL+HQkp
3p1N57KTM0uRHg7bLnYbOp85KricdKdUvqj6vYfNUVzS5bl9FWf1+ky41oD0CoED
sHZz+EIp6GZzfcaU9xjoWGBrgM37OWauUvQ9zsui3+nDy75QOdxvnsmAOIeyqMZz
IkcIBL4LgcARblFEyIpY0NUXre/Z71d2qhcHe0U6Tv14SOchO6vcTl98vVpQRc24
X07pOS+dQhJ/npdMMD6ybsFvDCtZp/0IolFzADLfENgI2Wxxf52xzVc3MWFi0Y0U
G9B0cW/Pu4BLyWqr1W4IxPMlVRBAw0cYd1dQnqV1pexCvLpN8lnPgTIhSX7crjwG
y6+gKozg/R6F00ObHuAqPgga9AKJ6AeqOSwCy9TLm2bD61Q/WaDye9zLeXU0ong5
V0Te2cz3dpv1Fe+FQzssa1bN3ARBaxRaXlcgt4RBnP1UpQbp+6W/BwQwl2wu0mvO
bkwd2Qg5/JuFSXQh1CXSX81hTQpY3xtGMCygmexy8OA5vAPpQnTz87x5N044jycl
RZLkQfMUzJGL+gyTKESaQ0vbQck1AV5jhM1v++/TpBY3bpg6z3yJ7xCLrHgktt1P
fMDYpFxxyoBG2dxMi35CN5Dfpd6lW2gzRhcH35d0VOi8cnq2RZtbU4TXe1i27han
cJ9aG8Fcib0Xtcf9ajI6chBoIy6UkvJJMGxh6P/D3V9nH6lsz3+5MDYWg5kJkxNM
/WCQFLuw+icPiA1miIeXrw+7qSQFFh9SnxySHiwmtwuDKzZJf8hlHB0tTaKYlY3C
qcanOJmBdadyCHKMGcl+37A7ezJCimb9h08lLMn24e1Jk72SNsNETd0Z8R84m3fP
StfQs61JL+NBcgJxyWvlVEEYYJFsM00KC9I8HZw7WMoQL0THXiSJcrjD5QdZqiIN
aUaaEv+kyZCk0RpCVYT1Jj7GgHD64EpDHStIPle0Bud4k0DmW4HIo85Uhv9GxA/I
d74ftiSenxW68/Ebhvb6lO93u5iuTlIquik/F8zIr02MKNGmaewTvCr96TfmdgFK
ReiTp6owq3UOWeO1kSP0loFccR4FxPmdL1p+zh4yudkBp2s2V/NB4WUrDt+3Vfni
L5PHNh7Ojd9zalwTzdwofPRQfBEKcy2JMN4Sv/fVyv7UWEkAjqZudpibgnoD6H0F
SOZPz4zyEeQ8qshl6IhEH2aA/rBvCrKU9EneqJrsB8pQYQu+9o4gDzECff2PG6yV
fStkSbS43WxN9x0OLqcBtk1i8OAYclXCus/HDVDx+AP/0eh3YGJnEPjJoRyGwIk8
atW7v+wtJFVnLjFGvq6s+G17+ysX1V24q8CHeQbqs+LG3byt8e2B1bhpl1reb51W
V17D0CwgZO9pDl7YhUH6pGUfLvbN/EifsU4UsGXkmOzB3VCyE+0KiwNmZuAUSEly
LR/27cpx/+N5ZTVO8qkmXGZ+mrAs5UvAsbXEMr9aNFE0i5OEKovjy/lsrl6hamRA
6CMv5dBA+GeipvbvZceUYEmw5+8r9FA/NiwMNyqGgbZGeYcgeQS2DL35bHl/CW0b
GrV+KvFYZk2zRibqXfn8kIBHlUQCv8o+y5wPsROiZMkzS4r2NdKWK2T8Y0VpkCc1
1FKh/PzIjVcsRsh32afEsKz1FqVBQ3CrjPUQEIKqrz9/z/rGEMtcyf1J4JfDavp2
7o/Kq1uicg58pFRsxhi9aaIHRxdZtwE55X+KIsyj5hfFoId1INyoH34nSi7l10yT
jurmXUTqdmqBZfKojyG13TZSpb0H/s1yHdXtXuqUV2zgasvDnkQgJzK0aJsxP9ER
BRcRgili+O5ve5q/KyOKK2GXh3puIJaPS7NzRXs/uFdY9lxZbW7S1owTMQTTuwi2
On0I5Hcdi5a4PfwEP8fUEyIOPfs4693Yd9Q42EQLIzO+4gdhmgilZvd9NHUUkFtc
g0849wY3iCU4UzNh5MTFd+7bcAu0eDZ5APyatRxLbcauEyCGOkvUe37HM7hAkziI
cyPGJ6e4SQcPwnl+S6CV1pcz0JuMuVcJDRDDK67wmxKlFKljDSudHf9Ov//IhsSl
eRH6fQM9ojmkjBv9lXoNcbnqiF1Yt8TC5Fqb20RjO665toJUlLQRnRXAiIpMh/Ya
TxCDQFGlXcaN1l4H+yxTRjZf0nk67uM/bun4QtFNgceXiXmdj3MeJ69w22Bwak8X
Ari1AKV/BLUFZ3zE4ttJ4G2VjakK+OB4FRYfX3hMGEcPhnldgxcXzB8TpCpYusKR
Br2lyUieTEG4l3KfDU6/fjmDQICsm48wq4vQsOBy8NUnAR9b6OhPS9etH1icllUz
MQx00evcnxvPBowTtUjxl9Y5u80XcDThZsNZuBm6Ki7QkAQBt+9ZrZ80RYjnc5Wt
QiuwHm+vApCTOt+buHuBH5KhMf/UHvHnkugvlR9Rzww7piU43tyKBL4hhTxWAjhD
EXBfNZlZ6D9JrapyvQGuR7O1xgxqweZ8g4SDImSqRO55LdKyIWj58H5hbMcsez/W
9FPKe/VANIDBEBJXoWQ2H39rPcHN3hXoweUeBbGv/3BJyu5AT8OfXmSLdR6uee29
WuDpGzVlAU5God5Yz4o7/uzXwf8K4I/sAV//QhA673IoGxmPpGoY8P/Qf8Pd1mZj
3m6iY2SNQo8ezWebcT5u8MfJtxdmy4BMqgzcX3L7NCL3y+PtTkhKB5XKUGzQUlq3
6h9m7Crhqy8+mJRA4RRn4EI8lcIkeYfd0kqn75uOkwugIPTqI6zt+q8s3pkNTcxV
pkK/YK36DAx+dzbdwmuEO9Ltkid/YyMlUTH6B9ylCF+GV2DR6MCjqhjh5VN+84ws
XuGpCFMmnG1ZOuBGNfPfRRO8+fyxIGLpw+BR5l34qAwrFK9a4fKiW0GxIbgkOr4l
qrDDcI/YRt3yxYes3yo+WwXMZ0+JlVaz8rvThLEkg/HAhn4GhEAyQOrsiCvUx7V2
b811YW9dw390OGuHrX/GqsQCa+bbn8AMKWjzA2liKpfM+7FwRYIkqfgkPvceaB+i
+Jhyr5qVSEalW2b9RzZ5BvVXtqdDA/hGvv3EIu6KyIAvT2zjaPIWBGDqhTy4USW/
lHUw9sfjU+NhDMqTMayHj8omopFs/UwigolNEFvFgV2h/tr7cik1lfnFquGf6f9m
0Ik+6/daNTqXq3bRhUl2+J9nuKLp3bQ22rCxnZXoAWD9MfcozbZp9pVwcGE1BxzO
/f+J5dAIo81aGDWab/OaMIfEbjYoNm246IUioXSvPW6HRqOxUTjJPWVQTchAWBy2
KnBXzNJzO6TFzTJR3U7cWib+99C96q2SDl7RiuWbV2VnY9oDlNaY6WjHGdZOnxkW
08lPxQOgaitTX1tJcY5cf8qgJFNvwTV3RmKUYLZgTgNDYi1hYGxyQyhZRi0L5LGO
XpBIpbULxuhstSZ6fRbI+mjHE26EXTfeevu3EK+djCR5x/Dy0OjnzwGgE53VpbEU
cvpl24dSAD2rvz9rLzQkwo575ejW/1A/5oOVNvRHg3JVU2SGjP9KgkntToBtEfPv
BBTO5aK1PdnVWANBbom9loeKClITG6wJVqiCG56F8eVMVzWlHxOAAEEtc6GZ4fzk
7uNZPEAEoD0G7frtBA2KTRx9ANLbZxYyFwFmrlBRcrPHHiSWyuVINkgrGWqlxq2B
PW1AP9IBnmEv6lyPTq/O1ZXpqchgcXB2115J33QEKKbRj+r8Are4kXJxyXw1+sL/
VA7bkUJQD8y/MyF+LMJMDbfVMn7akDT5nMPMt0pPtddJ8yxie60M8RznIKwqee2x
5ZawwmgDoD2jDTEPL0DE2f3i8d0YUmHleWCXQ4Y17q1E217+RqRznkBjnyZA+X1I
XHVZK8GurEOUqep44Mn2kyV64sTbH0DxFcUZI0ADy9hlCCWtYgtlwuhGi8C4q9+s
vZLvrn1eKdEpJK2IQS+4kJ2ygRJniXyry5bbYDU3B5Bq17Xj4PCHumvStK+37Buj
vbwjQqThq9gmIBaKlaIzuADrsAOMZZY5kOu5GdUiVfDEnDyHD5B54hm3Zh6H4Nz1
HEPoU3/9ZpBS69rCIEelp3QvOYaho+9pK4bTkjMILuILErmpyHmldf1g0ZccgKOT
//1K1kNnCIwisc6DqHAn78/p5t2g10Z2r3rgwXmII+1zbDeohuTi2od6JySfjZ0C
qy34vUkJzyyC2VryzCaqt6p1uCpWGnikSb4MC2VtsaL6iWFiy2wCO55wFKCFYn1v
ojCu8r6T1O9ItecuX3EKwp8mhkwO4nqqdrIiZ2zhJP80EfIa0v1taZivoOAP9/FE
DbUwzjFtt/xT+3hXRH+cytEkXac8QJ8aWC8NaFA7+pLqoYdWmIOga1JTlC7bjhQg
SrUHeI19fGOAST4+cqJ0f6+G42usSew6MMNduNzoRF9e4jMgIpOXy///nPTWtfl2
cDb5Gtp9r5MqY77WrEKPCFnxCI5/llgRIwyUIIksL08AiYryHzzrt9OzPraJwvfj
qeDIA21vJ95FfLAz1f6EftrqAVyvM46OBYAmFaQm/yw6VOXz+++2Oyo9aYXTRNAa
Vce+ADLMFqROwAKUMw96cHqXip8fWbDoO28dWt+q63gdnjIlTyo3HERZyLkivFFW
IJqyEedhPOPw81WoDkqzHi5tF9aatGV68fGrbK2OnRST0c0Xp/nbrId5eLRGBnOu
78J6C0dqXo0R9VePWwh57D8A4pTqTFiTawWGkxqEcr0hC5nIPXC8tofw3Dxo/o8F
/6v1RVOXlwKKOCpDP2rYpE624pFoWj9ylT2JBk/NBUm7mpzNiERsjgM3DovKwlBt
p1YyreKOtfeWAxLBGRmyuCAHoxN7Xpk6anm3TDhOOaflnYFYuRMAvl56cag8XiuV
PK/wg7pDcutBvsGh6Y4OOdjkqCoYtaK1ppOh/P7avIqhWi/9JybUDWRF/OSCZb1t
UodOzsb4UOb4AqcxNJERTZmFMI4OzrJM380S3stEov598qqZ65iYWmWCVWqF2h4Z
Tv+6bl+B5GqmmGhlma5W0j0B/yRuElY3EK+2YDam8cfJyVntjy87S6x3nyLX6kGf
+N2fwSpgiUWfSMXMcExULKVrHu4UOBxu6S5Qrg2N74crZ45skIIGt3cH7GVeKEHz
EzJinfWZ6F9elYFrFVXDZaFM/DWo03ePCmxiFv2a1Y5CWzM8V4LBcdOzOB4ClIZI
/rtczi3HsRUm8bN4GVaEvwtOJh/PYNT+VZlZlHpC41iL513J8oSQHfLNIVjZ2HZS
qN5nB3F4KE6f2zZy87ylkDSRLilwCu0LNPDfmqvZrvAiVUAfrypRnehSqAxMa/OO
x3Ge9PzpVxg8ntyBrK5ofyFKPzWcUhZLZV7Vto29A3FUkh7o8xjb8frGfMaXJZE5
RQZu53LXBXSZeS+tkoNapXjVA5zprW3/91DqiBjxOs5R4mEhL8SzQWeY1PWnqEkm
yvqwNtUQmCGAolgyqZLIH3pzsNdfli22SnIwD5+bbehRBFKG6DFTHPzo5yI3MvY3
FEQo7D99Dxe3tRs4zO984TaxCRanWHzeoOQumqjdURl5wCr+jx8ta4zOJXXuyq2x
eZouhnQlXRzJ3AMQGmfBVpqw9L7+125cAyEfTkDwkDniupZO2nLtWvxm++nEEj8A
9YJoiBS/WXfl2hQlGcXxCWpKD7KWeFinf64O14kxyZJIf7oOTPzanriilvedvfki
PsyxC6UXMscqvhhbR4KCCreD/e93FkitTRPt0Ha4ZAHoLGvNP/F4q+B6N01+2dWB
sJvNUsDVHF0SrMMuaD3da/9874Om/lYcLIbEImhR1QI7GvL8ySQJBGdOb2ow3g7t
S6JUXrnmCBRp+jTrsE9yQj2/ESVvkqfKBwyRy15dxBIMQWumnswNA0ghWLXXnc8D
OS86CHNC982xt2FUXPuU9aBewmQAlsLma66cVIz1rMe65XWm4Qi7d74a/pzP0yMw
v5TpxWABJ025l89/e2dYB04HS4syuN5S2W/66xO443bMSSgYUf4cTI+x9AtF8jJX
lO5Vv3osZyRAQUOpIKWIoyLiHGlcdLClHYWkxlzFSnx9n7pgYh3xagp1lZgJSc0Y
cfDQxIoUirhD+VX/L/1ZKBIYFFVI+lJNoIsyWtjtTFLQp9lVKOrl8V2MV4tOem1h
qIx9epAUC258g0Q2nymRDLOLtDBFSxCIJLHbAvcTO05ULuby0K0V6/oSpQk0ci/h
XaXrktInx+vd4gXc4MjDOoqAlQW5OFKgBIhtCh6Yy9WQj4JSzn7MTqIt0mIqK0uE
Bq/GiSFXvbFJiiaRx59G0L7CaBeVKn6CqwFCPrvS4WnfL8yG5TWY9dm4X1ZHZk5S
97Y/qOETfrP9qPlU2DxxOVei3NHClu3P6XOmRLhLbMOQ3tn6icI4vMhCl40hC6GX
Ik8FC0fBcc6k0am7vN9bxPYt6gSVB3nQxMg3REv/U0IrUYnyc/19vp2UFubAZ519
47zIMcumkUoUOs8AKlGJpn+Frpwv8Ybqq7jBjbIuRyNw2+UywrwBSBACFCOmpE6D
tH9S0JT/RI0BraCK9lGnWiVBnufs8IBnHxHwRZQFwbEihNCzThwJ/uy/eNnrvzHS
sbKBE5gVRlW/Tu/65xlAjL+uHKsVt7ue+V3Q0RxjKJktse/YDSuAg5D4P+OD1e4v
+9VAe0c8luSbiNXHvp66F/0zBi8PrA2LtEmZbrq6DGKCCHChPGNMNHhXyk8OhAwW
ov2X0kGHsJbDuiOobciwJNbovET3VG6Dpq7QlKN/0ZhTno8VRPHUm4g2ZvuIhrwh
YEOA+qHim2nN8KqJ0RwdnMjXI1bSOi6HlSb22iN/HIRkUYBZuxc0kbM8xRUf4dt3
cfohJ0KMLH52o4CqTd/A7W7ppqwjZX0IT1QSpecHD7BEtsfLmgG3i9gd7N7yOoB6
YHLTYPvm6JWtSlNDpejfdmjCQeqdkKHbD9HM75khoxFJAxMinMdloHrJtBn+jkQS
ynUCcN377cdpgrx4NfMDYXaV1AU7bXx/CzQdG1Ax3fFsi0TYQQo0WWenAf30abdg
ZEZtrJc49ZN/bvQE7uaHIpfhk8cPPRmU6vey8sO6QyaqA0oljfWnbWBl+2aUVFZP
nKD+vKwTKujnIqR9MBVyYePnKIlg7cUrlpk1GrpYCkuDgzusdlCb7TJJuIUVNxrw
zbCUMYOvcsG3mfdW3AosoC38GWbtQjqQm7WO8RjJ+rMV3hFOD2nXqODRjdxSKXHc
WQqo/Ek0Y725rYAQib02c1ay0GKnG9W74F41xYxlde374fUVYfSKVaA9RHESgXxm
oxOqCNjKm5OPWdQ/o9QJRRchuXpcSKUjSwd7jfYGHIsHWmBM2aRIvVx90lIZLR4t
tJ9XH24WGCGAkthkNgtUxUqR9Sm3ZTXo3gpQsab4vUIfDkXRyjDRvoVIgMeQVym+
1tIuD+Jopg/S0CHZsf6pF78zEWz0TZtbl8W+NL1//EKS1rn9lY08+hS4N/HqCWpt
XQnDDUJqQo+alroDFgBnFsL7H6vxSvGKBtxqvP4wC9tpV4ipiQNVVWzd6cLdrftS
s4d2OUfZisDZ2YvYYvZz61zanLeKJDR8C0KDrE2tTBufybrPbBR9cnTicmRHSPeS
hmpu2xZ+g0db3/dwhj2bFsX+w0arIIZlsLw2RDpr41LJmP6W8SDzegUrY7zDg/IB
1KTy4jl2C9leHvN1HMbawbPy3oitqRwm5AyQLDBt2Hh3qeovqAHdJsKHHBfcFYrg
mHT2tc67dsmjE7BPsrakjciUIkbunwPD5HviIQkJup1wgsH8O6leozjlto0/hy9g
jC4ocMpFjS9efaQzobdGPV0MDG8PE3zEJEnztKkbsIrYqqSkv8otwzbaUF403O/O
LaqnqxN0j3wsNGc5+4gFWoi7BaxwZNwfVaxN+zM5BknxuoXz6+PC7rc5WOZe+zGe
/3k+k3qjAGCvxv3yf0Xkb89aKCROQLvGt3OaaaTZZGRYC1yBYVKIou5n+d/ol6oP
tQ828vgzCEkYaWMmD4nop5PIiUcAtC/11y+IGUVdfdF0Lluix9OAa+5cFpMvnBQS
Mgy8L35g4J71dmhlm78Iz12mLYVyQjIXt7gHzGYhOAj0X7xtqslsSTCZw86wZ5EJ
SI+Nr+T7dqSrXP59Hr/L548/Xg/qYpXOjqHeJeyRtRBS1rX/8VfBfQea5yBOiDDV
t1ryJH/pMZaKh+3SKGtFcW0MyDBIvHIEdUjXwiR8in+zQCc1qfA2IQlE4kmC0kK7
x83rXBPY3DOGVtbk9ZSdTBo2CFdLNugqI+bBM9FbvcBwx4NUTSqTSnPvswDYjBmb
njoKjSMh5CtUxvVYe3Frn1v6Xto5tMqKWnKmPXjqUu8tO7imNNV6I7teTH7qdv3g
hb4nVfk5BzWQ19S+4VnmGlpSw0VRL0w5Va8t+Ep38pf777eSf9T6qeJh+JlAlAKe
GJ5rkmtsmWN/S9EDPW6Rjg/LZBtO4nspP64vXRDrqOmIUauq0smd1bksQPxbhDhv
P7aQsdUBZ5urQWpxJG19KsWa2UHsp58p8euVUL08f+SqKfPoCSWQ/psQHEPmAq93
eu6vim8JeLJ4RVBAGRPDECqFA6mNPzCWl+P1YUgIRj2He7issulc2DMhqUnikQR+
qym2PjaWCdOYl7WPl69C232pwVuekeneC1z6SU8as6XGzPgVdpUdVW2Vby5RrivH
IhPvT8L3/2uMduw/skGy5gKoQOoiJItczE7KqRXgzHbvKIdrt7Lcfkgy90wVNhE3
GDRoRlFREfrdgHbr1enrgBH9MLrT1H/hXQu8V+UZ9AviGJXwfW4j9OUNFv1c0o+x
v/hwdsEjQWo+o/IiglUk7u9mA5dNE120oLi/0R8GBTFrJewcSdgMn/qupumrXeLx
78N13sBufx9Pp57xVPyTSPCpT85jzm12gA3PnMCXVpzzxq9K2DsfPfMgO/vnj+Mb
34+SD1PQRLUBOfc8TjpugyHsLSCofe4A3Xa4DkQOHA/RG9nMQxwMt5UDsvN2VOg0
UhDljlu5w8sr7bRiHa4lAlBPWtUOWubruCDUd1TW4bj9xB4tPeICHUBDqxNViDyL
k5G3wQgdwtpKExP865wsZcPEITYkqgA0VKkixuImddDsmuT2LwuyVWPOAhQQPIoy
Y2xgTuBxqQAdwW3ESxDwLrSGFyq3GIKRuXWueECoSeUyCrMfwz1Ze5bDzqWhR8Er
fsa15+UGgWjtjMzDx/3vJYnxK1ywEpTHKZE5dApaf+1l2eZcVYitR1cZ68c1x7xf
m5umyFRI5k0OKihOBXqcQiQjD7dcSo2R5hrSfnGVriZn/NZc/MajGeDU/ZWd9NY5
6DTjwHYrAGf9ujroMlNFrWpYGAV42VIF1UODJim12u/UHrt86ifhN6nEbyf6tiAU
JV1/V0JRlRf/t1KY53bqKcmHnl9IFYwt/lMam8qLRedjenG5d2zgV0kzh4pefgj+
sasXXYND1V9I5z4B5vY2gomq4FWIAn1UnD7zni0IgExO+khsx6dgHg63WGms29JC
RnUik0sSzN796uYYEvFbk4EnZqUuKWQzVkHWPj2Lw8jzWSPyQ8DmTL5J8y8cEv6q
THH5Vq9rmufiGhNt2Z1NyTiwRL9OacoNY3bkXo+h4Ktg3prsom9LaiyvfhPmhQ6i
zyQXe1iTBTR2C1hiLGILQlZdURrqsDNBEqlE00HsFcB6mXnhMiWD/DmJGdtt9lxZ
R9S6zCtY+IVZXxJSOOn6zpGCEUltln6g1E7TtgjnM0LPrMZuPL0H//u+dp7EYm2T
HsQOr3aavwNLxUdYtsHyP7D6cQhiTY23QrrWQDyEUd5AEu71AFAPWmYWg5rNajRR
xybXsJd071PRy1vC+iS3NOPjEOjGpk6qFSJHckZ76NIc6XihsqTtBGcMd+NjF0gl
v9P5Hp2t+aLFkYLTiA9Pz4rQprxwIyLxekEZ4l8JUEZxasq0Mk+sNPRUrpEJ2QEB
Au/dGGWJEgTUisxFyLhHR7hMfts6X+vkH5fy7749QTAV9Q8TnQXMnJe7qwAr3vyY
whyn8NmLBmx4rbLlivuze0BLCJpDGYGm5hxxewsYMUA9QsVJLtkjzeohmS3325WK
2rMXIyEMSmpJOZo0HtkThmReMDgIeaFVyzYYLZ4RO5vKLbQ2OxsNgomuhoRnJVkO
AwUTjCUw6ZRUWPb8SYfyjCXzP6fZIqRBM2wWEkGe6fIfgOpFvubxNcEruKDPzYZ6
Gx0hsMGN4ggLbFGicg1uOecD954kAYmqEtH/1rYYldviVxZDlnL5JgOBtYWKhgBX
ErnkUPSFGo6ZJ6Y/AgQkkmQESpVl0R1ZsDMHm5P6N5+k22HU1mLbzSiJx3xQLkYX
R3IvhNmcrW066ina28+907THhIGoBm6D8BQd0jxCWk0HRYEYTh6o6pZ1BubWnBRI
bEc8sturZEG0EJmucAKzFB8/c8HtWDZfQ3akyZC8zlHAz73l3x3L2HvdRvn6z8M9
+EwAFwPPjTmWfwQlzPKHL9b2wxJbDOz+07tWUMQOLc0y7uw/Xtm4dlZjap4t9hSi
rmVQPnq+d//YLQ3G+CwzRiTW/sOUn7sIN8NvZyr3wboHpMwrfgA+3YaziEfPv4C0
PjelbMolYvfqdDNr6jhc3+GXjnhtbKe0tq5NeXFmPwJMjjUOw+0EwS5vumyN8vva
Sm56SorLn1vkIOyPDE4kx1MaxWg+5rpolrmmH5y8CnWCTpDcGTFDcSPJe/MrbNQa
kcB8Sz7zLkbdtsQmGIivCYjo1roVjU3WQS8+VY8fpQS2LkWIzKpWdVVLN8stKl4s
KrpdoYg6Bx+r8amddc7F3lZxsktiyJApu99T0C6tCWtTgsOB1EoQxb0N500AqTr8
4OK6PiAt24uKYBWknVdh19T/0zLJIxfwiXwIhsImKqTgs3LwrgHt9HgKo1MiWzuA
VQ0UyDOB4dy6gL2Cc9wFNi8aY4gI0DZ2rEZ9rjO/QYzMvCLgY9dErij0Iz4GOAd9
OgLt6sj15zRWy22HzlBJ859j9JFwEixSdOzDxRdnO3KRAETUCoNC4PP50Wf+9MtS
qylkm2dkSMswmvHALESwnYfp4agSO8TFkwB3RE1RD+dgcky9KIiHLrpYRVdeyrV7
rBy0oo8JfN8ZyO5l6p8FXRB3nSL1hMXwrmFk8VkSUP1tUcQBk/Qwo1gEH/9RnTBc
njoOQOEbnGCCDgfymEz1SSoJlGUkFqCbIcun51ccp+mwnvUF1gSLGXz2dArCz8Fb
1rGTS/faYWflcd1oqoloZ8DTyz4TLGcsvTMhGN1ZzFz1sHUQqdedvZGQJUDKiM+m
4VWB/ieexC9+iE3G0QiGOe0qMAhxs5R4MYP7utDJXOEljqa+lcg/17i10jRB7gvR
8IosIJ2k/6Se3+MAEF9zXhpHkLjVI9KEx8E/tmH80/CpV9ha/ImbpCv6XcZIKUcD
estHOG04qmRUjuMqtMxRmoWtMljiiKvockX4IfEjMrzItwDtyoNmFlrQYJDswHqK
V2UFXCBW4HQBjydyGKhUeqqfiQGUFaQMBV/fiyxkVZJHGmj+cL23/UQpiHLT1NDa
6BCuXDP0sEJvSAtqqGDRGxhxoFOHOA/+iUnDFCOPYHTKy7Fku4ddzjIg8gosWLhc
nMVGA9xMlmReduJEZ+oZzfxu46EmHAJ9JpH1sV9AyVEWVeZUVJKB1/+JsqMUGENY
1F4KOgo4R3S58du7/ZOHiGrIrrdnKbqq/Pz8QltGPUtzRL6hp+k+XNECIV2Qcjk8
7lFIvD/vM1rbg64NIt0q1xurN/rqvilWVFyuGGq1Z3E6bSEovnwKUEGtJ5u/UKD6
e34ImKuVbdgaZAp65xA2qSx522XcYUEsmBtT/bOVr0ybYzfA0RsXEpk32kvAqSfE
PP+UyPQqtYt9Q0EpvrwqayhE104rug+/JTE2V4EHV8CxyzZ8HCab4tP7LD2xctHx
4uLpbjOZAJE2nZu7OXpbTsLJrCU/o0LacE086negvOlOfYeuUsNU2fulaq3HOSHL
ht2FPzjNNb2q7url+xHM/xVMwREm4yvAkAGvYX0ShBKNJzGrNYRWchU3rXuxSqFA
Y8Hb9aHxirkzPfZZrkZJmRldyfdkipz5WjsxwJsZrylRneGZOFhidrXNCNSC9shs
jZYsWpNeKtYxP52WuQcet0pWlTuCo3vV3ay8KB+rziHoJ/oJr/yMcxdtIdJqESIJ
Z8hoR22VSwxFZzNDvG5hdU66hxZe2Gzqzgkp/Xko+MjFT9Hme65I4P0ZVLhe4VH7
btXm+C2/lZLF1nuv9SbPevSmTOTi9853mHP56X4k8Xed1SrT5Ek/RJqvtmYekZ/i
FcM3AsaJV9XoFrghiyhZYfiP2CN0wrS6Ve7RfXzTRMeuDaXsBcYLGVPy4RJhCiGe
pchK5YDtCCf3Ew6WTLw+0IsAvymGP0ustbVCpCq0p3pnGm7w2rskSvLci5eAWmF1
oN53Ima8/b2jtmzV0z6YsXp/RmoewKaBX762WwlVf1MMQvDja8VKqwq0ZOiRiT/m
pbYZYTK17juwOQ39cNDhfSoK/Sug6cm3P0z37UmRdiEOEvYRumh2/eApnJCpC6/z
NGvvIYPy2Cg84u5kTtTlzEUOiQJUbQKp+u0Xp5o7BW7Us+REiKjviqhwdtiRTxkm
+bxQk+wrkT4r3wqBM/CE6AgDJxAZ6A8tIaspSa7dZfmMZ5GqquXZlI/Ib2pUeCJB
cYfvO28+yTQ1kOaKONoXoRoaClv+WtGGQu3rJzc+Hz54Om9ROejG0WIyNFTaPYBZ
6EnsXD2kEttOm0rW/2Zep1y4Gxirl2bwmc60hxW/5F06DmMBillX4QzLnNq+dOJd
PCvR5BoKESj1Pic8ZLH96Iakeej1nTo3tqXjzihSQajqVVkUPCeNeC/14NUV2i91
jgEAcS1VRC0Vbmj2v9WzZG/s6e+ak42CVg6CBzU5qZoLpP6kTGkWIux+rNQi+5Ke
b/b4Rk9HEH8hpBeCn93/udte0vNpOUyIiTleNUiJwGZN+DtKyFvJNVyRSnNXjbH5
+hBhICv5Jx0RUE3miyYScLx5E8AMbB4+peM3xuDvUePPSbyszytbJf26dD2rnZMJ
GxoBG2eGHBDvEETcBVOgXc8aF/w4Rdn1UY1h3Jeankf/bujJuctgByNw+PQYKV8B
Bpo3nL1lWYyDVEbnj5iewMoqbp0owk2sq4QLQPLQj123VCcYtwYVrh9wk7WlvrKe
ECVxLqW1oBoyBweNzyiwL52YhN0GsQwQyDkY1kY6N197FQ9qZOY6/QvdVtEae0Fr
B5ZSKp7SP3mYxlDlDIzSi73F59DzNTkJRh4b7LllPdq5neKrggpsEdHp9R3+FS9b
Z1MmHTcbiAP2ftffBcnDEStF4IjoX07aTQNQf5JgoWkRsu7dllvfJuo3WHNyvlLP
i/pRvaQ8pOpnHa9yB4lLhVT1CBihI9VrX7J5Pj4pb9d5HaIaaK+uA+YNrI3ZP3Ze
oTwxHsLXMfXyHn9HYJsPlrNYPfb5+ao234nUiFW7AKrSrMbxuZj8eih5yUqSNfDf
Zl2YqqnofV0hFjpedpsGjxuyx3Ao1dytXWuMExuLfgugef9X9HxKnqW4HxvcO1TH
Nw8GfLcALRT4k1+phGYT6N04SfKmaN7lHHxgZ8hwN9wsTcZJmTX/Rv6I65FplhVK
puQyBHlHlGZeyYlat8QNSsKe6c+XWyP9pSkT1nlyokf0QdM1wTqtirA3zeTFNjhE
ckNXbSpV2Z1kUGDKy+ue8e6TQ1zI3YQTqa+TL5ToKDNgukmRP8VA0c661LE9l5lh
7EfRKYN12HsRB68O4CiCWCiC6CPKp7tTHnErPTuGbiGgtq8fSwtOzgHEjGRGQQXG
W8MHAPgl1yS6HsgQekhkF0xjXd0cUIkuo9NzbR0MPQm0HujRoOjYlIXxUPS9kpIy
P2sre7gtoeqdIzOkFPf2jjRTKdSdhfF8AzUVwewvoVQjp8Ck3b+zfot5x8tzKM0M
N9wIUVvXlsSQOCBF35NsUk5Mvom7R06p2LopDvpsG5GIJCJm74oBC7mJCujw2pnL
bWaJoLkwvNm4eV8d8fPNtfialsv/UNfg5H0h9aVEntbOl8VeQEW3BkSyuHBd/QY6
TB0NUb2UGe0mRhueSsC9jWozCEyggdUhTjj+i72qjummthmTBVcMKYtHlGen2qC7
tD58JsheY3U/w1FVD9+PP21aw9u4R0BrHTstPqFgQgIy7isM8/FAKT5sDf3oaPSQ
tXT606PS6sbG4TvKcEGk7sFXf/5q/i3BrzkJZwlV+bbrdC/e9pV9LyNo65pLZOR7
0DPR8PKlu48d89TpBiGw2QJr1TIANgl2sf2Te10jcgCizOCB3Pg6lK42KeV0il/v
RXo6mn1qGp7ubQoiuSG5n1zPAASCNBDos9s2hJVyBODFzNsD1ZHH1inHiVMaOGnU
wr4k7espBaVqSqtyMgZiNQspbeqsq3ZjeyyGjRogIsyg44f4FW5uQ67rkxKMWWPL
cXvekvO0SW795NpKZd6hqnWyzQTWpyObrfuSdFV6YWXhXNwetZXbaHg4oAX5cc71
yGo/F+bvFdoYgaeC2vZw+gXWFkciAVmWA42I6zkACq6y4WKgD1M9aWycWNNwXMwj
5gasROAve0hdHBDi33iV5D0/lI1Oj6FC+04yxBV63QA7dVcfZ3+vueQsgluhcR9t
tl70AiyMIN8V9R2NCtxMzCQV0Qp7/0jL0UQEZMTJ8BmrzidVY1EWh3FqPGUHbRZQ
Qg4ooIz4DdMswoJm/bwMQcsXD7OcXYPE/X5wz9ew4yApva06fP9ephRwrF0rQV5v
AUyKH6P4En2iqtfL07tfdyV6BzXFmy99ZvfaKx5CId/pTgwvqBxF0ERJXJ9WNHt7
ffvkrKk22j/ci3bokEbVUGa9OjCZr3SYPfLCjpa6w9dV0aalheWDaMNES36Q503K
pvNaaJSgG8lASAhlukcmrdxn11qhL6WERRGvtCOJQGTwEWHjZV7Kst5fS4wuNJ0r
cmVmUy6X/rI0HTUnSZvrm6lxK9KHymBXTDTncSFBhhuqkEeQ599/VAkDO4FoxWsd
zr/BMS1hirhFudB+LngOgeIJJyVnqsIY/DExRptu3+i5x1dXiGOIRcbhgHvG6MK4
onfGR6976eThz6gGJkwQlkoQF95Jg5U8s4c6dHBGizWRrym1tHnSwnMjLST93mJD
+vPRd48ZqkbxgAE2kttAAgYHDR/6o90TKwiSys6FtoV57qf8tkZrIte+TKC69On5
ZEXd7dHrFJoOZxV1huq24AZz6E1BHh+VMP8EhsfwyibUFEjl16a9QbzBmm1Ij3fI
apb9hat8zPRm0Z+CxTLzt/yYKoKQDFKE+akwSXbJtX8I8EbqbFX3xMDZ1eW1q4Jf
y9PUSR/VXXNVCCmSVeFwLliG4FCOFvZz69K/+0MhqYhwqCNsRJFJ/tpXeLWJSx4G
lQYvPo7HMpbXk2k2OTOd/2Io8shc/S3zIzzCOqwyhu3P5YicGEXDX8zSQKBx0/fe
rmb0Nky6N7d4WBGL4TY0bF6VtpM+9sYzmkY8kBbbMZRJmRbuhlFvzrgfPTAwjEzz
qYb6QoobTlsYice36RatUGMy7NnxNxszo+xcqcz4pxfkZI67qiNuknhZ0adX833v
1m6xnTNqutcFom1KGx7asEGuDUgUmCGb3ZvH1hnJetFWiI9tE5aaeNuG9Em3Vke/
7cjNwG6mxCcIaKUfgDggT6IgovKhxD568wBtNi/y0oYGqgL/YYt2WAYgKqUARqDs
iyLIeKyItDG7KUHdKu+Ioe+NAaTFMjkSTNG4TzVJd/mNJOevR3o7cm1DLcLRrze4
hWONF786xPFcvKD4UxpbJw8G9Y4DixBhdVcpkNkaQWLyELuE62qCNoyBmVcAnj0d
PDqgroGqNGtgKjxiAcor6zQC0dK3Hmft19CjtJUrPmO5Xb6T4m5J1M9RpsRB6sx0
RDFRhyAFkjOp6CtseO7o0Xmdn4pYKV0N0sAdKk4fNiJRbsCnLMilzrcnTZW/v0wb
wF5BGQIqpToXao8Lh4bsiocddDqHRf2VQd6/P/CJiueNJPfRY305/ShLlmNGuLBJ
x3XmqbzjSQvmTSXejwZf+Ws/Rvg/Ev1pbnOHNZPpGwFr5GhisTwV95bSnu4VAuR5
sFQxhrEf1v3k1Oiy75Py5ExzL7tsfVNwBfXV2jIvN/haGEoZRO6ZCr2x6+za5IDI
wJjR7MeAxv+gc+SorujmK7EutiG5bNXMb+qmNN5ehLfwM16/8wkXO+7+tS78e/rL
GEWnM+IUTOcTzKNV9eSGPUiHAISvAd0+zGxTuzmh31oomSecvWC/mAfdPoY+VkUA
1lm0Wsj28XPprRcna6dgUzPJA4w+5LjaBj41Zj3ZFRI0ZCcHkgFjMMNxtZc9dMZi
CJCi49xEDVWOIs4bn+bhYuH3LD1sfJ5Odqg6O7YjZcSn8m/SSF/KJvuncethZHLb
EYVBZtTdwGL0AEhUIbLmcTvL6a4+EZlaLHj3C+DmXSLeRZ2Nlxy7mSO0tYQPANnU
nIRvzWu1QplLm7KJ+eeSBomC5KHaLf03A4Wq+26ez9YqJNejZU3SEeocPYG78tIH
SqkIdkszijfN2ZxCEpqxDuetbxe2I/kkbHn/bfywRRE0ANiczDfL6e2FVuzRE3Gx
JqgiHae2RoVedc39k7FpWtpTaQ26jgG/tkxYTbNtNJ5MUl8lmgwzBPvblZagRxRH
i0lvkODvAJ/u2BwQ37Z5w/ai2Z1oPXHMlIo7o+JgpMxLT+9/lxf0pSwE0CAICukU
1F1ClrJ4mf0tzo1MLu0YlQfYDO6G79LI4LED7NIo34b1V6dlzt28smEUUlttWG6i
YBMTW0MkT2Qy1AbVzf3dOtVW2geokwJIaq6pecEkpoatikl1nikuIjPpSBSmOHul
IEAgamqNmEtFsxXfm0aO0B4egx/wglPF1ZNwHkOosDQc+dUs4stoxKQ02kXX0Pjd
MCME0flvFT/XSosKkF6CMYqV+S2schtkO8jSduADHcpYSEyUk8yPk7wxJA/5DXc5
4v8xqnbNXuKmQcvMAiDMtGY6yCuA1/Isj6GqlQwFCd8h1JyZS6YmGOTLJqnwVnjR
AIkW+ODvEj9RT2m7uFB8Vf/sQg+zNGxtkM7XhElU3DnBgroXjbUi4qp8n9hj/WCY
8JLuUhXMPVF2v9Eert1vG2WTQCIFbpdmbvnllLcp87Wxj5QcWKj5OVDG18FkV7G8
hf8IisGXz7TGXjsd8Y8HoZ1OAqwFlw61ZrVUHC6nM1koYyfTt2pRp/4EWd5TcFSX
mGHjJbtFAJgzTxCbTs+Ji8XAmqVWjWZ3o89uIsfuG+yjcqIvnFhY7Zl9McPDXVdy
i+UhNbPX/BnWtl4Ut7Hh99C7rUBMhIYe0kcZf6aZOm1e5RDH3zsYRwttSePpvYYy
77N0YGB2o5Ror6685BJJppEHl6eA53z94RKKX3yyUQ+Leb9XHulEbw4Ql3dLTp6H
MPaRZMUkGwm874nyEXdA4hT17WxUbAfdRophhdvNn+LirPbHlIoS2L6qzH/PmiLe
ec2bYiZh7nidc9lnLTVgq1f5JXtAlhYqS3vJ/fl1LZ3cEmp9OGuEn7R/4GhiRUUi
RGCyLRsQp8WO7XiFkh+dYHfIkbbcU77w7/rZrcy6VkKWccx0d0sRyKq8Sj3JEqYB
+UMMi59I95ofHiBfD7haTsr97S/4Tgl6Jc33aJde3jrumhTuBWjNwpKk1KmN9Sol
onqkaZjOXVPQmLL6Zb0jZKDjHD0oLAApHyE7Ubnku+VunDwJKzVv+7Dj26OMlFpd
JBzv4JM4t7hF+t4nG/jxc8PkTKbQZ7QTwHhkn0Farz82YT7vINKKCuOVc0A+HkU7
a6R1H0inBEB9V+sAoryuMdkSk1XFnmO63Lx2NHt/27btP6nQ8IZZMimAvQOeGg9h
Ka90+Ujf4m46MdDq1MXHOQXq8DUBpvtSo6TNYaLpBlQiMEYnKilbhSnoRzB8Vq0N
JBFBfSUd8mxj5O58uEWpM0G7pWrR1WaBE+SESl8sz+9TfNE9FliFhnnljebnUet6
ms2ci08L9KXyITyJZUknpAtbAfcMZyo1EQzK2PjBZrdrSlfkBZUYQEfYD0pIsMOs
rCzyqOlFtmwxXth+nRgSs5/fRufRwchp/UBAP9FhLS95OaXTboUAqSkcpJ6hE+6o
CxnFKP9kkeKQijP/Z9Z6o4+NUxTByT29iqxa2IbOSDB5aL4Cxfzq+dy8SHLDQ5OS
21kZOTCOFJrSLz5BPJkSAujF0M3gj4LYPCl79CUnVBPhOjodsHloaJ3/8VjyI+mx
Q5ifRE6XP1nn9Scid/g3DPcive0vCJjWg2gckapkoUvCJ4tXQi2PHe4/4H+empuE
m4sdDYOg2eThoaWJVuF+jvwqe6F0v/9LBGWNQj4BnXLHAakTbRQlyWDft+TdPnR0
zpbZKskVLqSvCIvrPDrm/kik+uD28utaRXrYESkqN+fRtzBWMhPsJz0tCy2niaNF
YjootDV+ONybgTUSEDTN3LlgE3ds8CtG391PVqFSnIPe4F+Ld7uc7o+3VKndGSgl
KixL19hNIA4RQ1paNhsNJ+tGrzh3IC/uDJDs5U1htHwinZ3GqWGK75WB+dcd76g7
lWMoNCYU/VU3M3mzdLAfazomKEMtgKKt7Ju4iKrvw5X2odKup7ZU/mCnLK67FTF5
IMSrKMd0lwDNHLyGy/Ngl8CD5EkZrWoePvjaQ4pfI1J5CpUCfxTGL/YuenbkeAwn
oG1giJhqKYsglMgup2mqWBVwIqMb+6O1Am9QlvWfPFkC1kvEBBBQxNFMkhWH7pIz
/EnrHCTL3eH78IomCI1n0Z7NMqRIYPeYDJ4wTYLKDU2bVmne5ppgKvQ3iZwf6Pqo
ht8OvSVC2M+d0/sLmyQfnRC5f/9l3t//iBql95CDw0hwfJDsHxT7bqlHrwvMF4Vx
+zPy4hPpYcQ2BfEtHSBNOtENQN3jxRyOWRbTfymwO+umyZgCzU6uJz8UcMJDTXP8
a8cLfZE8a83O9k9i3iYZG7nqorwukREcQrWN2uhvVtgECxWaf9di0Gsu0aDJdV3X
0+AnImVHZ/5oYqfDgJaCLoZ1tDpY0rmVQ4061UbMCwEVULqsnr7bZcXevQG/Itpa
yk24NCJZx3OWID/O3h7ltAkKEhAwmIv17r+74mZmFcbrztv5STcAgMF/RuLFKp+9
efOFbn7Ompp2YIom5BlwxokbboTb4ja3ds5HhYUsDhkAJDgyQpcnwvBSTztuda8X
i7rj9CYKY3IYVxs+0mjzUYAWZgaRrl1+zdd4Mml4cD/lm+PK6/IRRdI0B0Heh52J
PM+kYUHMAJG/FtgNu6S1NxBqM7YYG+2rFeDp6tYy/je84slDh23V34vKVIB9Kxr6
d5TLvkuXjbgJYXDqKYziDSezoNFcqxdDU5YQ6x1GPmj2NauJRFwrnL2bRPKmGaWg
N9FJlVPXporvtGi0rv4R1A2ns/RnQVVbVMb/C5T1/2hocEqbw0WzqYRrdPANg/nq
FkIKRjBWPTIqSGw5/QNAVKoq8goSfF+7P9yhc0dEcGlDL3hppfWS6zSFyzFEOuke
EYonhxbb+Wxq/QMzrhV5J4YrZHbicHxKIgiMqArtsRN4WZ+H33hHbjepJf5bQ8AT
uS8xsQVozuFDR3Yu0zqH013t3DFxMWAvMeRM1t2lofdxXmDoQDHxfGlqFsX/SxIB
SW2r+vZ8lmQGfW4kFmaHHagqmtTGp4tkXaQxr0uJJG1OleK1tlxBT6D7rbPTNpwV
cVGgkhIEAsSKj4F9V9OMgnBI6OXUEb+czQYTlJZVDYt1JqsNPl+fqpyQc3ZKkFe6
ZpaLzNB5j5A1nRwIfZ+NqupsE+nxsh9Xv/UP9sm1npYN4BJ8cVRZVP3CfVvflL7W
oZwwqsT/C7WldR6OFDMlZm5pCMdnhn0NLeAGe97TVsaMKwCOO7R/Qmxm8q6FhRdw
g8TAWbu3se67vO06vqaLemeDlyBV1Q0rj6E334a4uxpHO1P6J8y680NYczt8HOEG
mn1Fx47ohOrz+XxlMDslXKYxyWKPu3wl/gbi1JA9MVSCUFZ6EDIAQWWDv0VMrGPm
xiRyjfXBbyGRiiIe84ymwetBtqH/m+OhGKGRocgqtn9EeY8GXKdECQt4GGtOWaEr
dc0Kp4mkEGpKvhs8oGoHZ/n5GkzUPtSzTvuAKv9OHOGUGrqOpiAEKo+dCxCIXGl+
tCoGs55sAN0gNwoG/CYmsRFPccRBt1XN7ExX9ZltVFPqhb6Fx/mPvs3XMTQN8Hnm
OGRiBMwGWjjFf6EykSGjc322/+83gR12c954Hc9z8RUEYM4Mie2C+euLAZgVjrMB
3+7TBX1WbxsUlLrJWQ5pqOTd04PNszOSu+KL5nYiOEE4gUO2K9T2KIXBv4YWW+2q
7ubiF9jGNvGJlszAfW7NelaVkrlf5m0d7xewbLCLqWJ6Qlw0iZ3HLqa/0kK2QXAM
ffOqzkdygNVhUK3mfVYmabgXljKG4QCjb/kMOrdU00fojOnQf7EdJy9kl/PaUFXJ
WEn6XnnEONgbyqX7ue/pZ5MgKI+bkoofdF6AsS5d9bB/7a5VxQQPy9jXkTz3X6x/
4nOPrtmr9n7EZ23CIQkpkYRpGs2Pvz+7N6mMtfF2/9d8R1POyczQu+JgjgUZfGPs
rcKf9+FRf6hzCgnsUtAqPAO8U3hb5Egzz+BzCm/uqiA2liwz27Nld6K0X0SYb0z5
BcttSSJg5fSb9dEh3VX6ydD8E8JcY+nFRTuJX327GLvhmlZLOr9Ty06uqKhn161n
SNM1AZlpAdmKUebOGrDl8B5HyxI3M2OIvjCYTCrPe1ivJYqifR/9/o24PEi/P4xH
ehjqadj2ttJnkx0eZZ0pwuyQEFQGHZWRVYkEsIhrGTz+xD528S5UmR5EY0Fac86a
9xPrP8knMidzUSQP/6qzWxqZtOlHpYsqdkIyni7sh3RvX04OqqNEUPgein1OKsCN
V6+yC6NomHKhZAXImxY9pDDMpHIckt11MakAtMNJMQqWsO0bcX+3SJ1cmdc16BUQ
BCqEhKI+DvLpS6QPyU0nmWueCtWXaAViqKALeeJimEN6BMV0sK0TGSJtTbQpjkeE
m3tYEqb0+M1lID5f1Vor3DdimtKEDqz326pV7AbOpk6fcXfJ1Lp7ISHgLJrXlIl4
D9FT2x8dh7bIb5X1oAr9x0ASt944dX+0yZ9eP6FJkmfd6YNEixjxbcJ/h5K2Ipr/
lShMiniKo9Es4nb7xI10K54Yzv2AmNIjEyAzeymm+o9KdlIH+cUsOLf6qGcQ3pWf
WQ9uIYL+ZHFrH5UqoIDdt5WwWTl0nNtnY027c0omuS9Tp+Fik4ipUjEz/zY1tUJz
GiTBHJyNyxEaq7ZVFzr5daH5vkagBO9Lza0HAPSoreNv1m2D+JZ8NqDyi2mOsjV2
0CJ15vkS0B/rpa7WbgmDhQ3+OIIQI7sfUe7N4zPqdU7U6qX/hfpZJwun2knkbjHu
KEObx8aB+EhyEGnslmKhWJeU6rZRuonT/OOYf+sXq7EOcGym4aY3lGNUD4aPwNAs
OGfidSc6lY7Aa3kmMmyPItIAAJkyD5B1M7kSClQIB+nzxMURJiwRrx2rE5qf4C6j
wdmqs1NihKTZOvCiO3tVfKGgq9KmVlSmRjssdN8cwiHU9zbPZH3FtfWE21fXhBt8
AozeI+NkCotqcanZ1RyTDU5xu/CELQeIfoHIr061FvuAhbR47VQP1K09T6lwTOLL
W/Tq+vBCWDa/h3EZJ9deMyFFibSbhooAkUjEiKC3jYJrKYUs8cdVdS534yYbbZpN
+yWgNJ/obu7cAh2RpLND7cRuU8JRc9LN4Ies44AGKnidLzWPXQMh8HF4QeVzOovi
zvSMnuivZqqSiyN6tzgYABF9bYqXsZbCfy3SlF+hJ/jRB0BGToAXjDGjCBHpgJTe
3FceU1V/NUv3Z/k9W7rlG+BICaz5/HzYsITJI2OpsHmzHmCPksFYyzfRSa1q4XrR
fcMoywQ3+X6+hNbipy4y98oeQzB3LhDquIZy2VVPlRMFNXwkqmPUYHhhQP9tUr1X
/Fi2l4Kbi7Nfe+cXj5gnI9Z4KaxBAkQiEbsZf7+taKd84QFnNa9uM9KyaQdHPyNB
XPQHu+PMZvVX2P1xmOlojyf/xNiTohz2aJ2wF0A7yzSforUozBmImnB+8HTI7+/4
J/DnHlDrs0hwR53OS1boGCbDhzOBq/sDkeYGDfHcMWEjcw4U3CjVe5AqtVGOEwUg
ZrCsCj5artP12Ks2OvkeZY5nuriPE2qqGO3oVN+FLpa4BM/n/9LAm+a+/t/XMu9T
zyACdY97gYBqmrpv8TLcAwyBPPg/DQtLfV74rDICgvr9BZIcTYjJPySUxTnBRmtD
Sbm0tWWqs9C9tic69Q8Lh/jm+ISvFBy8PDyy4BVs0+wIBZ/e8CyUslChzchmT25t
IRl34XX3AOmNeuEyKB9+6niNmfj3p0+a+jtl38BeDPzAzjgDF29msTSCQh2AHRLt
OSsQv9jgVt4JB1xXD9hWXmqIMVCIf4d3L28HBdMXPb/JAxwPxUuQnuQQD4X/Rw44
EwBoNMyOc3GqVdhJXqHBYsbmUurMx+rffxiSlHLcZd2C9Ax5p+9uSrKRMgG4ZnOu
TbjRLDJqq71ZlQ4RwRAWfb7MpVPf+wTpPl8RgW94jz6w5vNK04lAzOpiy/P21wyK
o5hR84LbcZFi/oXypYVcmFAOunJPhqcgAoM88ekYm+5EMyRUuplRqovg6ifm0pmK
zGZ46m8YxPwjaCbfyB00Fw95CtRUgzrnEVg11X5ddzh9gWsZArgrI5I22VUfxGjX
cFthp0OQ5wQeRMsRC+rPKaUYgNuqc4BZoja3MvF9INHvMeY3cq2jiJjEMlByfNbY
cEImBbM9+gtFLt/zbY3UWIM2Dq/7FeJb1Ba9IQxiPbVzEgmDQ6G6IjIoFC/CtU1e
17xtSV86qCjcE0BqPcNvgWWJ3HbWuPhFVb6+yzAo2M4QLfLUMSMenETZn/K/EFE9
NhAsQxHnO0I4kVYXo5IHGVpyzFqAwpOJj0DyFGC3KMiVAVEAktDJABDVa1vd3ywB
0qJv2Dn2WxcgkhujyGzhwzwS9U+Wa36KTSvn5RxVMkkzH+VJzmHjtYiKFeJw/p5W
aUNqZFezBXuVxgSWekcazon8RR8HBX+VvC70qotc8+7anHJ3cdCj4mU4GCKoOZEi
+Mb8jN/tDxyCEQF5rvnpGceiMXQjaflkuEqJarrR3V5O2UZXYl1nUvM6YcJXj4qZ
0gZ7r4NEFUjpWLvjUEqbBVivxCnH5+1QbQdiRKfN8WCxnqLy9Z/8PfM0JkWF65q8
3PI7ZHa52jFgF5cplfqRT6URRvaiBvVIlu76h48V3L6S/wtu2QnSxn8duPW5ID1d
WgLWImprP2gZdQd7P2tbDXYFaRgbvJWb9PtXi7OeP79A3p2beKwiaqmdOkA4dlvb
+2F7TAq9vLOEIvtX6R1xyMf1BsOHCLtq3jl4Jl85cZF/jOj/xulxwSYRMUDcvLbu
iBdjXQokaD5zGHsiwvd1VrI18stGEb53io0080NNDAUYdCZfdJkaprxIIaewg7PG
9+vf7zqOdzQ/uL24jzmLsK0rBDFEEhApErpelUbO4c8BVICNeP6e1M2/kDeB0/1e
p/LiQcyjA1gdBAYljCHNo3/IpA1jhjBykcblRhuULopPqDsqUluzjXpyKbpkWLme
LT5/Gmus5141ewACacZ7hcRQU1rgTNfVjcWx8EzDjgfZxFnoZGF5BPlBNBlZ2RSg
+F8f38zBr+KYs5d3kIrpkhCBmUwpRLVnNsM/A5T21a8idJDwMWHOZKALcMMzKbjM
TwBGEtrLVs1p1qHjOEUYysGcWfWPjWXthIA7nDK7eZlIGr57goByMc3mY3UCkW8G
DMxpAX3zvdJQsikdQ6PDP05GK7e4ZCdkvEsBcGc1NWHNlFhyJ9pDaiBZbICVhZZV
teFdWoNW4zh7tRTT+9xdr4uxuAiF5RxTMUzp26jfUapM1sJqT1dDqxX52HVYEyKs
841kaqPlu/HeyxSA7FP6MRvODPA4EXtgfz3016QvhpxVqa7gxGzobL//Xwhe4JJV
rnh8fex4xQVWz7YipAX/18SROOrPE0oxNq6RX3F4Peh3qiRyUx4XeGLILUDAGK31
L359tWgKOMZZYZOmfdi+Au6bm4GmZu9FtTcTphmi2aEIrVgsoJaBjwJDez0vg9ws
Oug5seO8qSmlHOZTS8fH8pxHEvKTF4FgrsdJdFTNb//tydt+BWnzfDhUFuP96GKb
8+N7KAlS1nzarWtwQUcy9yBdRHzGv9Q6fhlsXLjzWIQBCYEr2T/iw9ovAPtXNwxh
mglBigw+USwddNWIIApP/j5g6b5cVGrdCoFVEJj6SuEMylTocaXmUKhh05bsO0sH
rLjYbrLI66CRJwtw2gLnDMYfyjggPfkdbSSf2AcJyA/b70uMonGCeoS6t9awNfqh
6EHBR8nUZGzgr5RmDXbN9CrmMnaZaYjp7b74cNAJEBDRfn7I6fd9qOwgn0sT6nWt
j7myl/4/UFXky7k7/sfWhhPWlu4NUZf2XuDPhb0HyFP2kwzOE+wQ/jB8mkxSMv0h
6s9KfI2uwlzlgHjEjFbj5ueamuVRrd5X3IgwL3h4GqmyJM8sbK2YgcvzbZ83JNnT
zhSp0w1PtIJkGR77F1oW433TD8gNLOuTCwhbRao6DCJkjjvodsEvZXhNmxil6IuP
dtncyjU3mbLZ5MRkJ1EXmAFphH+3qG/wMinwkCpUxuYpUBQkxL/194TQDtmK+SHT
ZIlYJO64JIj8g4l49T+xymdsljMn7RAzFNcSRQhZS84GuV8YEED+zaTj5ggVisfO
iT4UKtV45ZJgjmIVFHu9x7RZBrJrNHuyWu16RzpZYcfbCqOjJg+qKCe/tVtFuL5k
+JfwXglHFMpqPEmxynJi+sxZpc4wG/c5DdKmA8SGKV5DVt2NE4WGIbQyuBJQJgPu
Y2DjVEpfYir7giTRv5AtOvsM1Vng3rkNrQYN6kTI0gb69Uw447wilM/ZBq45kavy
xk7zwrnPkZOwg72jbeYkZH0SaMfqMRHelUbh7lJDDLd3vQxfxH/jep5d0+50Al/x
kub0Sv/SI25K0rzPBAXULctVpdaiTu5o3VF7ejcBkW0eNPK+U2MVAj+sz8G0t2u1
Z4eRrIt17hoth9XkPaDDVefAexkgMqwTnqP5+H2KWFM6862WTYvVqyhJaxBdJYRu
o4EVWCZuiUnl8BWzDRJwdKi8g2epRZNw7HrVhEz6Vfyo0c15gIaJ7CzeNIr6gtYK
iObhb9PI5bqJaUqRI6l+zPPcU6ssugKA9AWR/0R86ONmGuAU9mub31F7gh9E9r9/
BmKUjKQjrh45k4p+X/onTWZdDy2cirx7cyn9apRTmOzTO0Y7y1nUfxalKgU98R+t
RtIr2aKxNYTUY5N5eccWvpCR1Tw0B+LBoF99gyQeqXFVH43HFuofBUNvYh3Bj/CL
b5RZ0rteBPXfZTvacOw507zr1QNYwtvNwSpWZ5nc/ZYBs+/cu2H2zu60AL7rsDeN
3l3u9KEQfy9BpqpK8kqVns8gCmLONmM/7ALDCcL2KCSqfqpWH7yLNdpPm9XKKVD8
Fc83vnZCLQ/jpbI+i7W80eKuPIAIPWRxThwNXq5caqvyz0bNsy2SshyWi2zVMAlR
/8zpY+zRTgCkWoeyoacNBBUIYCUoWKALUFaAWdHkfy9Sl4aM2uU+0O94JUnTwQXi
Xv9HMKjFqlW7sEuObh6Z0q35VzAlEFEW68h+dNkrFj4WbTocZW3RKKd5DeJTFM/I
IhiLZ5H/Uayyo9avKCJ98SvDEB4IMcpzRV8YzCOXj6W+6GdF3vjyQu0prWhbQ5/M
G6GCSlwxK0qDv/EnBXdDuwEwSXcKjG5WFgUUAArjlaSVna+F/obaYoAWjrII/b+Z
eumT2z7K60liosobjDeG40RMzjcgJfOkHgQilSoQ/2x0kFAien2MUxQ/40AaqiGO
UPa2OVtxi2GJRzWj/SueGjzd7MYcpTalHCM4J1lybAiwKlcO28tPtz7Auea0EsWi
vXUag+7HAyISgxcAz00GPNRK3toBCAPzJFk0toK32TID6SSqUglt+sLBA4G8bOvf
j9lmx/bQVKlErno94ru/2r3vfV7ejnlfAVJ9T3mcXlhBS5WHO3opP0DpHcfbUbC8
pp4DwybagCZvBXCnLlWW9u3KRxwHoc+mXoV/MkQaw885kLqDK9bGlrL9czpAiHpd
dc60p1kIjgFfK1ufMK8kSRlF7bruL0UR/QHU/os7gpS70ndG+EjiBKWfDuE7Eikn
kF5uiPDVafWHgV7nN2FC47e9eV/bYNPym8FSxmgIt0imrgaVjifccR4Xm3puEh5Y
LqT0cja0tQNC5zxcKL7GWUfSL9jxP7t4G3yU6WJp6z7wUxrL+jtas6O0MPQTYeKu
EGlZU7r/vgfPe4G180osyOz4uRkquQQrJLHtMzOipUx1upwgbdI+dQJTeliP0YH/
+MJJO01iO1E0+DvKemg/KG1ZI7B9qrfj2iqaifrTRu/288GWDYz/asWgxbf9EjEU
aCFMhu18JtXM2se/WxdU7/+F8J1FhZbOpPijtg0t4B6XGVzeCLnL0L0Ex3a2wtAc
F9ArPNjN+1zk2sfEWJKyp37NOpnpbFL6ZTaBfcRkticvh3rgl0Q8cDTDSn7YsYRV
tRBw+K6C0RqG3AmEVXxyQEzbrvIXWYCXDjFAwvveuNbLZcnyuNY9snTvqT2RxVFr
N6fynPu/W+zufCn+X+UjE3uKv09ZGc8C5do8VTtlKeLtJaY76zXpjXG1PmXEzorO
4A35qZoBn064atYDh/grtWzDNvfTl2wAbkJMFZW5KGRDvHfDw1DrpwbIaU/5rhd4
PBYGrzUAEAlfTG0p+B3I886zfcRRwwl0MmgSF80xbI9AQJoBVDSYELJO3f/0p2Ah
nIpjLa/uPgq0tMPv5Uuby6VYase+TIb4hHMpGJYc4SK4VAbClVFX7qKsZC9qZ4Ij
7wT6Emg0BXIwhiiTfoB+dIacJGN47vg7xhHBKMHzvZglZFycTmp+aJqzHGWnoalI
4UadE80zBpWEvFjRvswN1s2UQ2nvrCJDSAvLXmKMrkPxUamg4TmHVGdLwd8JUj5P
F7KwTyoIYK2ZSJ715tN5+wYMoTn2mBXqxl760Cr4ClVYwSTYROtjIbHxypB/Qbi1
mBmJq6prE2Y838LFgM4zSUXxtgwCvTETS+Wadi3U9cI2qsWoi0kqNWNuOy+UCDaa
uBpnB1x0PmQarbCQq29Q5g4U4prw8WaXyI/JNKUOOrAUskBezqaFT5X6aMl197nD
QYPnggVFVvO6em5zd5q99SQjYMNfyuUxZrKo4j2QHuvjzKfBauU5U7l4ryCbUXjg
jA/7VvVG7mleT+dI0HC6nOaZThUCtAnZpEj9Uub/YuPqGThUNu24E7xfO9RJJ1BS
fugn9c2AbJh2n7FmaBhj4wDqSREqrxJA0EIFkBrytHcHXRwSwwNr5q/1EW2TUgyS
CzWSHJR2ETJ+8clS516MIF0Rwh1dY6b4z5I3DSnqUQXBB4dS88tQ79LVwhHobH2K
ZQ8ZKgYF7n7Cr3rfmuPUMP3RgZpao+kPPpkQRfZRBLHaC1+boq1PePrcz7XPIL3H
Cz8tMI6T+UUgYadTtLVwKTMomygxg63sWkDbLKi3vOItSELAFxgpgMiNtPIl4GQz
3jl2F1U3hSACrMHWqkZjy2u8dv6riQoa5Y7kFAHMwEe+Ld3IXqcjaGpN5AY58ST4
VUce4yFkCXFQAVF2pL2KoPL8JxAyWxU8wrHLflxupCE8JpLKwSQH/nl5QjaQwqf+
KoGfm+7KbIauK2oVD2NzlAx1fBukyWtssOKoA8fJJzzpCTAHuxqL4PZ9ya0ZRy/N
cpxZfyZJXSYeZyWi06F+f41ioImFwtx8dmALuaTDqjpIrC0sYQJOAWol5esFTu55
vfFXPrXUKWneRfAat8IIdz/N3DrturznQu/F3FvQu84Fi8EW1w3MjyS4Qt1+Ovm2
0WR363SL7vhS0IVla/FNRSwWRhprrAjcqr0+2zf4zbI01kaU5AzUsZdYeYL5czJ3
xK0slRG7fUwP63vFlu0bXaYhx2IMgcpBH6c0HIGTmm3h4HHkNgvCRYhs22MwdAzJ
HQeEfXaVDGDlKH+QCUd3add9WWkQM2V+xoq3cUyUVhHPi2Fn+skhawahbPUVLr6s
IeX3AR0ikpC5UBulpgjxQCm2kUvlZ6wphigBtwAfIwUFjI/lgl6bRI/DQBWwwfhb
Zka+Llrd5MIs0U9BVFzz68H7PlRcI3Q/VeNEDDR7R7Hnn/l4xQdcbxTXv+XJuI8I
DbGccj5PPob0xT9aLwufRoyxtV/1S4luaa/eI8veNOd8nPLKxakEiTyWyf8uxUaX
ZInlwPuRLmPwllDtcdduRfv3jV0fV7bb6lRijzizJC9RxHN3/0ApytgAgD09JHOh
EFpWz5cbjjxcQTDkx9NGmH+d/s4Mi/hsR7M7TXwOfgLIkR7K0iFsFr0M6t/tPJtV
oIV3dNwwcBL9g1P+BmTqROVjFridK2dzITjMWqI9baGrEx+z9RPTfrvOVe2S1mNY
xRxrlSS2wkq/HyqQO0bE6/9K+Mj2Bok4QRzvWeZ48M+U/KgxrsrBabvcF4hCvFRt
53MkrGl8BzF312WhASwj8KG1MsywXTt5XSOjRY9yFHpkiYhh3s/cE5GGB5nrH1OE
CZE4/MH4Pt/seN3pCnl1EBc3TZQrYQklGPd37BTuq2andB4G30unCVND3GWnzPk2
0DSRxqTAyTtOGPwUzdSCe1AiH29kX4fC2CYFM/+gShZ8/rn0TXEbh3j0x8AppkXA
ocNdpUj6jwJ1SNMiK/7WpeZKxH9ldN3lMOxM6+Ol5O+IVD0uD/pY0e7rBRO928Iv
iPuzpHSINfOnedEvLKB8K5buPWJyA9pq7JU6wVggdrQ5b5bdvaqLlOUOIcLy3PFS
KWhFhJkB/zFNzWNHnhq+WF4CU6I1dTFbxTUagXUSCk52Wsh1EXrO+lFRK2N5PTpO
rfSfQrdTfDctAMlGIe50xxH1geuu3BMfGrMK6qfugtW/ZBBpavNmGEYjCJRMuJ5J
94u4ZK674iLjo4wuIrtbSmNmLza1u9Lm3ci3+JZAZ0zZ5J64GXgSmVLcviCE2Lb6
bx5BWQw/0SKKn+ZGfMVs2QPktRsY57fxl4oKQeAh1CZ/E7llu5NWZW4OU0UxI0fT
JYtTNihOBbQrszz+aIGD4MWiUJ6FiJRlJJuamnTf8JVJQYChPaeb5Lwn59I3dYeF
eoXwtuo7wQsH6O32CsnazLpLBvllW0O3zKe1BVd4LL2BWGC3Qzoonksp2FovUa/R
XAKRJha0IC/Q/UYA63CeDaPttFpvAikH3Wkt1q9eR60jI8bdDc7IHotaPX8/0Ms+
OF4y/aXWr4TQmNsMsQlvdXoY47FHJ1LnHTjY5FjOWVhz58GHY5TGqNvkFFn5L1YM
foVye+hmAa7523y5qQkds8eYLkPnJHS7GJnmMsSF8QqDk4iQwhDEIDajWeOv9LyB
UIyAbsm1ypr4h0thO4k5Gc22rSUtL2t3Cq9uGMctIzM2mOFQVa/uYiOR3crY7lHO
9QECf6aQsIfPIvMoHtEOH6hJK4NhKU5QBwCsUSpL5os3RT4Fh5PTg5EGTr0gI3aM
9U84ocaR9lI3GE1n9Mwr0W3YW/ygda5z60hN3+K/3IxtWfAKq0AfT5ekmWrvNTDR
vmrkQQd7SC0XOID7Z+Hr0uffx9YM76HyEPP099Y2GWrWAMGVn700qWw9LlB4E4o1
55GS98aU8w+6KZeFLwxCJYELvaKwBVejfyt9wSFCDyPsd4oxNtkJgbtiUtPPqi3P
nlo37MMoHyfeM5Lpvqm9Lh5uylxbo9LkVAPGq5z+McW1itE9T5VpGajhzPi/HNBV
4f4IurEVvbMw3nnp7EGEh8ju1Or5L1miEMTAo1r/lkQ+8vFIvQ4PeEaSv8DbU4w0
7NmzuT9NnpU/7aNZa2OYJPS9EK9+8xIVGnK6IQtJvViWUtyrGtn7E+hiElcy7Jxe
lQGqoeRmOvVVooGMtH9iJOyGdWpXvJvi1o1VSyhVnOlHN/Wj4Fo+xWdgXOxC98Ap
MY24lhJxSN4N+PKljcsqUGfJ5TEUe6Wgi9jia4qm3Z56KEsG9zXivWb1w71lhR9z
x3snSu1p9zsLp58C62+gkwFEiM9nMJVtN0I54gaRr3umuomsNvFH5clNA3EE2eDa
wAx/3KtZCikpugQ1pFPzPqdkgklWYd0stWcWYFF0HInNEaj5yWV3onxGAj3am1pN
qsEEk4EtPy88EO7yaho/3oM7rtvIs2NzhQwPjayW8uCrk13U6g8ba56qNmKWaxhz
Ps/RgMRnNKD4VuhdZRFF7EfQnNpQFFocHCLzowv2hEBKTE9pa1BgpUHd2LE3C2y/
ALr4JK/r4dKWIQ2U+eobCqVYMLkPdkwl3ZbxuHU66Fy2owlan0M8y9uCu5sJhlK4
5LcGAPKRyPcImMMjnsYgCd/3I3hPXaqyflKuukF29FZxBq/ffYDWVGQ8tKEAUO23
u6Q7NSVyKa7gAS5uCGiKsprFeDNixdSryCgme1wkHg8krZgwXSIoXDy9PUxw2Ef0
r7y12XUV63YJDPpS/vJKl9Ue98+1gIVAbQbpm7toaJWjxbKNISFPd1ofK89qaDnf
uxnhhnGflOtBp4zk13urryc/A1xDJgvZjyDKYGbqw7sjwrCktcdKpZMSrSMHPPHu
+KPlT0fjKl3RqDvfBYoGDbii/rhCgXvwKBbQYkKKIHOwsvtMjdq8gqTQj0sERvc9
2p4uG2DDvgu2+7zbrd7zwNJv/n8ia1H52+fCvUeckZCXgnfVN8ApKNGvvbpBZzTe
MH1mDbUfqkv2NKKaZc/JrcQbaeNvcM7owvSecyj9NB+5aXN4VckQD2JBoP1T/RSU
U/nZBIdPTUwB+e0iNq+MEaum2J3t5PuoY4+CXNhsFKzlLbK/JX2Q1mbdD6B+C9vh
soS0umxJ9DRtsS3uKlnrSdGlPpcWsdeSAmOlLBXS06gEzwiTy8YSSgDtt9hgulYf
h3+437G7UmyE6nJh5vBJpXNy2+AU/D7EGN4/Tcz1PiXcPUHCKgruQSF34Kt4uv8h
lBJtzHIacYI3WKSD/ES8yhaLvloH1crOlqtZlm/UmFAvJ95ba+vJ/s3y3I9rCZ00
xdJY6SACnXHy1UFqxu9PRuKxZRauhmnPV4TTZR0NdKgdGTYPFVbvR1Xo0fBq+V2Q
RFwD8A+Qxi9/XxelObXpK8e79F6fJpWsIIWF7uXVYY/6z5Z+gjRMlXJ8xnlGCnqi
InyL07cYi+zhQ3qqMfFm9rcoMbOnVWLCiR/wFDMwCpWKm3lulJii46o7b0FEFOuo
oW6z5h2JrS6Ej2KTfhfI8dc6L13AIfONyaMdfOmXXnP0JJx+tb9D1YJ1xZH2ywKu
NYJhePAlkzmahdW3sxRGLEe+ECmb12MqoCvultuDXF8jIt0WPvzXu0U6a6EE4Nr+
MTaKgZOR54jNWDPi83aMZgrCOLqIFHbIxkzx8OfIIJD2DaX1JOPrh6qyLNkVZ5qL
OmLtV+c4m75co9Bpi8f/5KOgrXh0fvTCYhg2V1p09kopFLGz5+db/357G0asOxJL
b6VLLgqe+zG687LN6Jx15kBAp4IW4nMYXyMbxPG2OAzUHe2LIXy7sIk+MSJe4jMP
sya2bstF15dOASCOMFbS+Mq+Y251NSrrj6p+hX9KPoZpBeHucZFRA2BR/fppyD1V
pdHdUV92Ujy1FnTJ142X5WYpVAUcYR9+/vl+dD/ZdQedZzDWPcHBPqNnz81NzmPk
2YQfHzREC/M7nAtd3s/BIq5jj4Sb+wvgx0Kl7v92iuA0CLiJ/libMoFWsOy/pjdX
PLHBJktoWDPgm1/QE7ZvzT+0RTrOf8N7j2cbb+BUE7lQLtUkzkfHMEa0s7ZftXEe
GMUdanmaXeatDKltdnAoulbubKRreMYdqCKAp7ufNXBWEQQWvNVBg7rJvgMOgdfG
6wDrt1qgqR0M5b/7ryrVTKco2T93zCxYJxGbxEWxh5rhLmKweOhP0IgdW7Posk8s
qeCyUHFssfDand9WcEM0kNkMX7yf6Qg/si8cO6MTmj/lHCql3P++rwJ4Ghn7dKeg
1ehdrS0J8/wJwm30eEoHoPLV0l5TH7eRmBO0bZhUbhM87R9Xp2BFO/6qUIrOItfZ
nwO251xYqEt3uooAXXvuchqru97SGjI21FYLpyjRwtC3GRn20izrmZoUt7RIe1eJ
CPpK4yc9EdvmaQEcIwCZUNj3XLVvvEAppOuxx8XgrYSF5kDLnNVxNARS0+z6NoQb
9PclwZobfW+wmTm2lGciMdAgB8vfXd2iFQShur9ANE6VetrgkiyT9zJi5aPI5+AA
6FDmJTvC0iFKQd9dvTB+1CUJZdgoWbG9n1OXQYunz0A+mrHV7gmxCy5gGLjQQPGF
Iq7uuW7Nrqa2xITcPIHdof97HBgAlpmtf2nUh5QfPD2ORuhT5n7P0EsUuAsx//RD
secyjHW4KSlnU6NOShjjPJT5rAf9QXEyd9m3mpjnuvPwu2KGXlC68p4V7givkc4D
S0J+XHgXd9ty7oczK4ZuM5wYZ5UjMF3Vwi7snpVVdKqR/pyYHIbpKFhdqWgpC1Rm
MPFUhRIZpinD/VMj7Jt8HrsqmGJncTevWzlMRtqApilwx9ZAFDSsFKjxH6TyrL9p
uNzM551oTLKs0hbnmiFEGg+l4YfD7vSQ4ZzXWgTt9iyHG9SXYkflR1wLffnAmBp8
LIP+SwxQPtGMyp0qCcvgHjHHfksEOns0VsGl6/cznAreqRy5aGv1oFRtt24/JXmE
Np4uMmRBkjQu3S8senA8cePxCdDoprfhNjqXbG3io7tWQ4G8l9JbT+RUOsqTxjdH
GwQIkCxtABtu1V0CStoyyanF7fBAZroD8btE/NMtxym79/+EL9CoGszfhK0BTTa0
zkw5PmdycByy/Ber0oOgA6M5whUnYjUFxWUfTVR2BLx4EcXErCVUYHU6x0x7trv8
mq+MYdc+JnzwYCQ/73w3caZPQx1FPucVKFUxK6eiPj/XcLt+/fweA106YXAJB2xY
zAKQLZHCzDuRWN6Bzd+nBCtgyO2TAg/MweDV523tU0VcVKwS9N9E92HoF4sUSnNY
yYPtVOowL5/Kjd1L0K5Aassd8jLiKClvgi2YYv+pQuRlgFvUaQ/6y0HGJbRHnzVf
pWfNW0PHtSmg0jbJhnu5r40BMnJoS26EO0CREIxIyUeL2ttjguPhonsvatFSAUEZ
hzy+6LdmiAWi3iUbn2JeEiiCXNP463zcSoSXUUKMQbfRMxotM/r2TM/dK67/iviA
SjbdI6RNlOoR4KKRDldpwLhSpEkpZAikOr2ySbxdB5skRwXoYzioq5Cd5/FREnlx
0D1443M62+NLD9jrEGcCHDH3LB+22v5/QLfsorv3yxrUJ3sU/cRxLjpQLfsLS7ae
rSFrCDOhi4n1vX9OEbWTzOrqg2hyQXhVRsw5P4olom1ls7ZNYp4aSx3+Qnil4k0k
Mhk0+IcU3kBFo5/a98MqhmNPnDCYijrPNDFNF8Y4miTwdVIcx+MSPXzox8AX4lb6
j+RrFWei2bsC9vHHuf+wVxY2psy97Am+wka/OaFISecO2wFDL0ZLiQFd3rloiUqY
vn6wUVzpkVZH1f+MKI+bofj2McazgGm/deKTgbVjM4Ga3cX2BI91kGiynJ5qyd9E
U8Xjx4YTmowuJ49/Zw3s9MX8FD0qRBxFs04g3ESfVwOP4i91g9SAyitktOEGcAQG
0JHi37UccZ4j9tWuaJ/sToBmWAO01qEqfHbBbsYiY6Pl48BlLlNMgieHHzW2VnQU
mYZWKt66DgIVOjbitUtaS+1/BvI1KnSH0uiOerltG+XX5KClLPsCIZE3BUMhKArX
5qoCmyTt+2progJeJhFxHWuGmhL4zIpSDobssovcYkF8YR0zOQBLyjkIsjDbeV7a
2TnqBeXD825GKURM9n+ZS9RsrxBjVDSioK+QXuIfsW8U+GuIYcT2911AyG7HsSO+
v/Qf+LxY09SfkrLh2JWE6OWFBkXtJpROY0uv/QkgjYBGp/g5sDpOltUbF7N4rrgR
155+BhhZgaw+6o3G41d9tsAVx0r46qb6/tfKYSs78/ZUQpr3rcS8I8SU25rHgPKM
f6uFOtlsD9laR0Ri6RqI8dn4Rlez7SDqEFPGvyrjw1Qzqu7vSfX6TZbU6NDsPeDr
zcCOlzWQEsyQf/I9dxWMqqnGhutFMfnRhkGrxcdn9swKjyTuQ/DpLF+IoBJ2MAwB
BeErgT1Z5+p4Vvdb8HtIKj3HKQN+sonN/kmQSgeOyDdBTC6tqPz8t+RtVsyNxEQ1
yYll8T3vo4C7fzIU3Lvf5O8j7UXqYba7nQs8XGHBQWdFbez5JrsLEdGhNKEGgqrE
IRaQAcN9iFkomVf6YK6BTdywOZu+0XA7Ey6EHjW1SYPd4ZNz+mHgxn8rBTQAaBjq
9095J1VRcdUZs1CKx9nvNOwjoEP7iwCmdwjW/upJRoaWMqYsd/Xh4oeSQxSubqQm
zj3T55TbKizQVfAfk+Uifzv7vGNf+RM5v1Sb06lGZGk+IqSzSXqTDcLX6BsN+9JT
ezSblvQ+DCKhdvFZzvwMwc1y4E7zzABGBUQpFCRzowmGznQPJ9IsCGK+Jg7Vdoxt
jGrfEAyCUnOhoFrvuMvlFnZvFQResb4aei5DpmTnxXFf4s++qjib7lPJcRW/bkpZ
NIsr5tkE/FQIms0m9eXSekh4My5j1z7Z7tTDk7W0RVu/LewZeFMzgUL1cpKXQMr2
vpXTTLJolzOkqkpr8ir4WCXKqH7SIrdBxQK4bThgHfABH9h2cW97jxYDjUVQAISG
6e6Jrb9mHzE8oZ/PbSL/DMw3NsTI68XH/LInPlur07adbfs75/px4YvGREvJfTfO
8Grj4QeS/VOg6Wk1fKfpd6g7gpC0d2AT4GGNSIZN8qpSieqyCirTuz9taVXJfo5Q
ThJkUmEzt+PHEqJW6BZ/uPD5277JBmx+6aWExlh5m1UugtttymMo9cdljYrEDwpt
N7Gsr4DO47BQ7WGIvihXJ55Dy0z4i81yoIGG//Hn9MASFSoiwIddgib+dKvy1Jkp
zhZIPJzq5+8acrXPPMBrwwjNO+/nXnd5F06v766XBEBMCSaeQ+Zm0uabIXj0hrvh
c/xBIXdAQpzRrJlZPKagr2XN77UbY2WFG/VcwTFVnfIHmKoB1y/TjaP6h9mcyD49
myYVw0mNyixOqEp3VLS3NyjZq2bm/oMPLE23bBhAUs4CIBuBTpIl4RSfXkg5dyfY
nVkmj/ezp1s12OigK/jQ1jJNi0fg5pCdc2JfWrS7KmHLh41oy7VgEcqsclM2LnzE
UDxIQDlTYHXhvtJftB959whNiL182E6/2WLLk7UfLFhMn64HqArGXl8axtJCFokb
GWfPxi9tBuo5fLvgGGqRFWC/5mMC93JRUvSeiyTAyOYNsmtj1xblh78qLFP2L4iM
4dZacD3IW244TeTQJ7KkE1T0LjPQIZc0bTwAde2TRCiSlQRslHkWTM+5DfbMrVdD
PZzaXy5aJsvWPOKErsbEr6CA10LgDXqQ4d5lhOq5M8YTLQM28eJJn0aN7Moc1/+n
U0bBVs3bPKPoABq4b81xMJFFf1zAKjg5uEo6F3NC8YMO99rBf6GPM5+54Ec4vPTl
vn9jER2K9T7IgNKpVrdIP/zNPaADurZonOwF6G/E7I4IRm44uUmMtas4089C/K7h
FkXwlNFz2ftlOQXEaODFVYpYy8Q3JKyc9c34guLonIAQgfy4vHE2KOPYtbZDQ7bc
N07UwCcWPQlvnDTGt7tTvquyblxZy3YI6fYVYsxutMtJILBUyUujV0OmespicJ4u
rhEcIYLliN0uaELCHGyRb0M0fiwGMN42HdpVKiwkf5qusfZVBOFw04o599GVTkc+
mEd/M75euHXRkXRYBFGEyIKFGlrVQSvGSRt2AZizsg7e9jIQgaq8IC8bcG7zWxTn
O8exYJdAA+iPb6aPi/rQrRqWwyS5vo7ohQjIMw9vYKjWXxWzt3thvlFPWXmGih25
7ee9LKBn7ho0qy4DsvCL1a968AToxBlTtgohFdA4mG7h5Ve9gMT3McwesC1ZZK8B
j5bSJODA71oMc4Q5HsFxeZmw0vaDAETtCC0bJHQ0cxRm5zG927AXIdbZ1Hq5Idx+
FNk66Av2KZDBn1a92DbtayWmN4KgNr/c9wCZD+RfixOgcmzhX6LSNbp4t8LhZZzd
NNeEHH5WX2BxOQF18cxV5xgdENiHpWU8zgs9ZpejEjureEQxhSP+OmhRTq1ggulB
pHKdL/gL0FtrdJnXvhiCpprjaOsQqqWcL8xuPUytBtaGaJTBJlls1QSDib8NbIaJ
alioghX47HHyl6aXGJrgGtpDtXK06RpSIKOMBg/bSq37pasFxacRcZz+hyWnYbdG
FdjfvdVytO2dBA6aE54yGGnJzCSpYKN4+ZkSGBP8mRguZmfhukv4+9+5IwBxenS/
95Nc0KMtJnvuCv00fHYpuJypdAw5V//8aAHkldJIr2pdGkgIg/qo8g4971pPGvYv
oo90qYQ3Y63O8Ni+x4p1WRNjAYI83/LGXoYq8JQ3PUq7p6+ZimSlrVkwx2yHkdB0
W3/0JuFcKe1iyB7I22MdjCY+PTefFExPE2I1M/hRIoj3xMFoUbHWJnM+AMm3dJAg
O01fbM2176OQS5zU9ctUm5Ws+upPlbD8jy2pcsbE9EFxIvBMO4ART+B4hI7Jtw45
Zs9CBNXTmhUm3b7zlriw3XZRMvbNcVOHqC2gUPjb/cfq4IzZqWJPVFFOvCIjXP30
mE3P++iQpUYrBN5mZ0Yb3HQO+FF6gXbAn7vAp0IcYgwAQag62tDPIVBYXal6mw5x
GBJj/TObV1nn4Q+85PIY+PFhOdLpw6eAwNYL550V2QuzpDKBP/WbXan60B/gLK+s
bQYp/JueGt9TrrLFenY8bFesQDmGoN5/wvWMaqgHU/aSsAWc+Gpwkttp+wlWlzno
uAW/qpuliUQC3YhtRdrXei4UyeHMAvkhSMpYvEdl+9VCl/UDXPVWVLPLu8Oc9t3o
BUg2UwdmO9ajGOdZS2Vx5BHn5vUT+QcquhKXwFvKM5J9QiV0yVkr3kLJl+B4aiDL
MSFPnBxVqp/a+qZwW4jCUGfxZtbF8bN1h0O7kAa8Bv9z3wpzR2gaDgQLBJvUydlQ
+5jC5jjx+rd63Xy9a54z9Ri2SOJHMQZy2qL+t3gI5GmziRAlIhI7R4d/cHRk8btl
lQnlxyerCufe9sIZ2DKTlWAB9hrJANyXBj0jDtln6vMp8S1yok5z/FUNb8nCMfIH
r8ghKOp3H7E7poS8h3pr80dh28aj9yoOpxmo8JUFUhPAoSvMtuZi3dapgQr61ke9
LeJbToNl8W/q30rjVv/o90zDgzchrNphZNgVp+ZDfERAjB7ijBFtKRvFGprfSCzu
7acaCsMSQIl7zH/Gw4KtH4GMa6SAoWlIodXk28BDuO4x3/ajy8Xmi+RAWUCBiCBI
uYkRbUifNqqR8DntOGeef1mr/ETyK6W1snNBxAnD4ivqxv7qrc6gt60jtV7wXhIi
hknQDKMWXrMZLCnZDuPwXw3xGpvLECJeTzovPwdv3V6bWQuHNc/E8vF3yrv1vd/S
+ckQJt6NrJiu5GQ6t9H+j8qqaLL5+nIB65ZsowhfZCrgLVfTJeGSXXiRCtNuTwp4
/foUdXs7SLlIPzhwDytmfdgPEL6o1D1YWHIcVh0PTJV9ptpRLSVqys36tKv+NNFq
vF639VrkbfeqE8P8ZcLTupXOZZTal4rJJw5io3JeH2V3sK2Zjs1hQc+5gzvlxZAK
fDTe+Q9ArBF5qHHVNxHlcy1i161khvgWjYFAESrr+1AQVhiOZmWUSmfSL/XIiDYV
V5+rQNMbtcKFrQOVaDkATj/kzyAacn02ghTG21UE3kLX69P4AXbJpiVW/JuvfLH5
EEFgHXIfzIIjx0CeM36Y2UK2HrnRvbsEoHvXUKpDhs1XUfPJb6wrTTx9vSdK6m2C
2u3Yi/zQ+ADuyR5EVVSqMIlWVOWc7OQj+2hT0odzV50QdpihU95i4T/RqjkZSZXD
pMJEBuWktoOSrIPpYtWqzw5OPhSWwvQgM7cEizk0TiM5UXClQabcThDyNE/BT1Oy
ph1Rh3mTYZB/e9KdbAkMhz1L8OoYZn6Sg18kSylyfwGUmkXftrLvgLzNuL6o4IDC
Inc4yxu9WvicMrQb7FOPeLSu2gqZ6NpCaMzZJ4TRTO2eNhzIrl6ewV2CEY0DUnx8
h9hgM/eqEyjQBp/z+n9oDCe7CLEOiOnnWwsVhG4rDzv6J6NIDBVr7Qgtp/Xv1aQ+
WBCSUTtTtDfDrOiUW+S0OUMTxrlZvG6+WizHtfwVqeAJueyCVE01mri9E8MUjaQS
Kjghw06HeapQrtZoPTX3TnU+eWB0UtQlgByXU0onWc30cTd32j6z+4wZ07rmgSMR
8Qw/5NnmTDqONfWtE4+Oyxk9giyuDUKnyG/GuETOVjoSnzv+DwYFaitSB5A+Wlxu
sDmJ82qv5uG6TOIdrRTVsRXVMDLv7QaT7+5w62m1WHBXjbGy/Ribmqp+7GvyLMdg
0fRVoD1u2d8zJ7w20t0nz7Xi6Qgqey1XW4JGlpVwaILYoqNmWrUu9mitXNCYXgCJ
7FbPN1E5FS7kJkAqCknBE92IqMoySlmozqDYRwLCpVhNi/4hljiRDf3abfFjVF8W
fjhjJ4dOZgT8ZxXlaqRH+5KeAKg8iZ4R0wUP8ald34lpEH4stCyI66VpYDd4LS02
7EZ5DCyR6EKd7pF5q+lFoer/viJqL2W6+TsytozUW+ecpVmeYvs8MsuQU/W+x9Qt
V568w1TtcSj6zv7jAXQXPkMO9EViSRmlqwaEkz2XNWFch86K4LRJ5NXERJxMdplC
Gy8Z0CowQ9ConqamhX+dgpnlzZt1K8tuJuBoxpYgTrNyYpNz288cSbvf0sJqLKab
DOO3wlTstIBRg7f43yjtpWgs3YQTqLVsjbxFu5h7a2FH+Mqx2f8fYvz7TkIo8eWp
1xKfmEPK22HSPI04H89szvEUwJYf4yLWX/3iZrNuX42P2qSsVRfYlRWlqTTVmvZJ
cfV+xD4hvicUVCsE1ErJ3jYWOCRg6rjL4I6pQZTUT4peOFiKaY5k341TuVim0iSI
fe3m3lASFl3XbcagBLT/bvwHebQKl5a9q40mKFOPMdGqM6NHtJUgGIpgjXyRptZ7
4o40J246pQxOHOaMrElOuIV666k2gedFtu2E093Hr63OXkq3VQzJolDM6P2yD8eD
9BlgUDKXnEyo0fKCgS3W3FCai1ApuZkFvIMDQCfnBawqWi+oq9dTOoA8MHOhKzwJ
/nc0AFUgbjsDCbqYZ2fR8vTXpzex8LDa/kuWRRZb+Fh/qHBsp1haxt+2Z3mO/AGT
wBsbRaIdABuGh3gw6s1NdQ4a0PO9uV/CIePT+ZWy0HV3pnJy4VubZuXgWDxdORwZ
GvBghLbG51JnU6YpC9NETrlSzigApLorITweZNrbN4Pw3DKm8qDIrqFHMtw1TAVE
qCzhnOokysUIOhe+s8wLaJgdPkwN+gHZnoHQTpaRYv5iqVLAGhTXUQKQUDbAU4We
dD6vjV5GFtHYSKnX31dey0upjy/BaQ+gaSIg/ywJaEgrWw4FBiFzvHidFjgjz4yd
y5LK1igtxUAoFdPKrK6+tvvEQ+U1NdTf/LsmGWsfsSPKjIsQTzF3qvFCjrumVYAC
2sZK+TkYuayJi47nJA+8tfp8uHUNuzJefi9yQMpmcJyqJii4BeTK0dV+IDhjjjpb
rpX9bVxFVA/NmoynXARIp7tboFSwDhtgb5nUGQyVdeWOX9Q+x/+DiA0MH9TbxHXA
Q69K7JkrTlvsMC9RRn4aBsKul4ePzPYktxMrxj3lz+jhwAK2ZCRh1pfbTL8S1q44
wF5bvbdnd86yddeVc6wf1N1CeV5p0DiRyAHZvO8x0K9J/Jw3h1JYsUb5aximLZlv
drvGjQ7GZfjtjteE39BWS7skO6y1uE8obe2XaUIsh2fL1alWt1uh8WKlDRgG0Af2
xLF9KyNOUUAUttPaojrppQC+Gr8tjWtBAbWyFfxGgaoAzSkddWeu2xgJ7yiAxTzw
iy7BndHfImosyHbqcst2BxifHymdTgV3f1IvZovxKQrAwsZTlqCot8S0mVZAh9SE
oUPCB7bELng9boxIJBK9MEFzPU9ChXg0YvUs49GlB5ZqQqc7AoqkSu2gv4jy5dol
K43xCikKVjbqlQThfV/szzpBnn/X2wBEVj3VqOlW+7d7bvujyN3UBWqhWtm/RKao
zP5+v31kMZ4hooraIpp/OywCodW2+E0Ldn5+xmKo5u4n2z3zrSVrMadRU0TG9puq
i3BvcJnvHKsAsm+TtmNVnoixCMjJW64HvdbTjXRh0RT61iD/ojcdfn46hCUQrkt6
YEwmQGh6HyfOmQEZxPygYyDbqr+a18TLaghogW+WU7W/CU+eu9DgwuHno6MwUIVl
oJnkCmdf7LK32VqtzC0Sdg/glwtWOMyJJTADWIXOOQtBA7gLyfwi2ekxJZY650Kt
dGVpBvp4xDr7a4KvKe1CgEvp8CLyBOW16ihyJ1kjoBXpnW8JsXuazz5q0rWfWrY5
/rJM2hiqK/GFqPZRiPgiHwM6KQ5WCEk3d26uCgKBAWgE1pUEpmWfO6JahyPsYDjn
fHKsqEklpXU5ebClBx0d7IY1e5bffW6cwiUUhVWQVd97zRdRTovDRxOhLNZsvgnI
dm+x8bH5TNWV1U2+38xG7p6UR/WLVkFBKFvk19SsJOfz1g35AmoqjzV5UktHVFoF
/uBB6rexR0bK9Sac1Jo+e5hRAtmDxY365Seejf/d/rb3ww9p+dB8aLaNgfwK5ItK
IGohH6FyHI5Fk88D8OU6L93QfexxiBU79X7lR6aLhApgRBMg0S9x3/wm+ZGa+rOg
Yhzy9sMXFVGDCjhOoshL1AKQP7tnfDaqGsURh3cca2ULQ9oaOGN0G9u9FTdoc+Yt
aZPYeZsMP5h/o2Jo8SyJUqqgjOqdMj/0xGOGLcEQNkto6GhkH2lYD6fQQ1KyThmR
s9XQ2WwMZVa1S5bTTyk2okg0C2l3Eln2+zjSh2P6w5cZDiqpoSjeIJHJ8APA0YYr
U1R58PeGZldwTYlcxweCjjsai3T4fVAIPZpJ2a06N/WaKsCP1Dn78e5Lgjf6DjpJ
GAMFTY1a2SgNWjzgooG1Vcziqr1rEIAFt/+gyOpE2bVIyzQXoVuCElnVOf7XWxVK
AOxayecpEpOh5S8gjb/qgQZm1joB+nnib13bCfsYddOh8ofdZpqgEl+FTUPNFTE1
xXsYia2tYPcvIUR5c6nx2E40diGfMWwPURz/1CoYVmaw2VM2aRj8KnVIrPMRPe63
/g2Zozbp+iocr6jziT6kQCU3nuO8GOuWGLvz7vRVusYItv2zEmK+ckEFrf+L4fvY
U6aamENS/F8Oo4ogpTpfTo8KiB+7XqoYnk10xn0MRu0TZrO9X2/g2FPlfvOr82bx
sAkqZh+Ki+Dh2XyLM2hzJy/5AHDryuXdLjBTGwjxalDbqfizKKZiOqu3sqCs2TWu
ApXNS/viZvlV5PvdFkyR7lbgIlSG5M0NmY7BfjghFsMl8wCuwee2XzSnjV5lXV0B
fLhoE9VyHsP4Tbs1dfuHZYxyp2d9PdFXBYy8YMKegdF51m6lnJbDgxnq0Fhh+T/u
WpMabPehOKARRsXwMoHvaKh+B0wHu8q0xMGOC/D0iDTaWZhEDSWcMUsngz0dBpHI
kZPqnT3IiWmNmFkxGwkL9E4XE+a4VEEwXlG1RMYzQZ+pZawkNdBYK2Enizrt0q1Z
f7QPevnRixRvIqKfW/cYeXoSXxxC4X01I072uz5LGO/uznncNKuysDetlEwhlI0I
NCxnOyvcTvt7l3MkLEBuwj/RsqNCflAqz+eaOgENKchkTvrTfx0QpdfFlowtAmVl
e6ru4Js5dFXfuPFtzP/TyU4OOuZQDVk3/6euBsAJ7AsL9STiFLzPA7MFy3zFzaAh
vqSrIS6cO/P7qKcsU5BdFKq+sAyDDfONHCjiScN/9R1abxHSDoQQ0nBPcEp+M2Bf
CaTuLi/MvRAwM0d3vCNpL0TtKV3LrKetw3RBGLDWoR5e3TFAtPQKN4kC0WexpdJb
z5Moa24TnMr/05Psnun1zlJMN1SlBJ7ezuTLDHlhIKAM4yjjzHUxSHzSKck9+Mwn
rjGd4TxgDgJYcOSIu3iwSGmdIwQqTmeYAFHFV/AHGQvPEVJKLGvCtjgkMkzZ7a6T
YW4x2zddfU9hC0nyeS1q7z23XP6ss63lJEZGVFGUFSj0XjqBl04TVNKGOtw9ORf5
05YhJ7A+pp+XpPPWEALbBmMxBzE/3MN2Rd2muL06GTowYcz+H00Nd22xQEEHmaL7
6YTaZ9B6NDeAARQyK3pjRb6BVkaKjFngeEd8snDiedaPb2IX9xOWgxFowqLuy/KY
oDkNmlyw5FsuDeVwHmXzEw6ahYAVTuApJOeve219wVBg912Wnwn9K/Sy9pgk53N1
aXYfunbG5od5IqeAay5xSfoWh08ZGn66DCOocvKpafyIo1qddkFDKyV3djgcNFl9
pXy9Hvqyum1UkWqfseUcIplmMxIuRvpYjBe0dUkj45eG0nAUO67UEMHJM6fj04Tc
Qpzmg5S3LG6IZ1sJigcOrkPw9zpavZTfVXiR7bpgNcc0ymL/6l0pisAkCgXcvSAC
h/LeNM3JES0Cs9oGxxqgAIOwzV4pu67pW+GA5yzc8X52JaLkpjEV0llh/He5w1Bw
7qlswIME7mLYEsv1PsewuvZjCa/mX3sNY/ySO81/qSacX+5gY054Kt6k4MjO+awx
azVh/kstoO3DiythNKFE4hwGYXyudqcWFcbaxYNotHDdze9VNBoQyh8Xl5SiXwzW
YElPTLJeBmQKpGZSxG7f5JsKK4TBbRkKmaZLHPW9+iUus4hXEJVpzwwYHxoLe560
f4GEo7MOCZVnNquaSdJE5oxbZaLRkC0099DCdjkJMXg+7rQuSbLknxupzZuOJrJJ
mwnnP/WZ49AX/ivvSMBqd5taalhdfqevDDLU3bSoyH/olcyv67fCGTADDo/CIYcG
aWwtQYVzPTGuZZIM9cumUkmVCKJy9ypNn6j8pohZcEdJfZQ7t9Tc0UuPmLwJEe/N
C3BE80cHgeoik4HRqqID+EnwWDUtFHoXA70qS8L60onUuh7V7Fxdw6y1JhxRyRMa
EkCa8A/8E7OVMVoWZNHrM0Glei6ct+nS8OotDPZfkSD8MQBEpQjIKy6dRDSHX/eX
y10c3LOCN0CEP3E/8CJ0IRE58rpBiFZ+OIDrNMH41Bd8ptNnZdkSZEm8sLzjwfhD
YtVQBJm7KQol+0ofF7/GBMtOsjuhE3v+R7u2gzPKNZrkJEsiOF75Ru/240/RLgDl
AanHn39P4B59PEEgHP0rEhCdPLwFaiCKMHxbyPytAGNDs1GLok57rlvoZN4nv1mD
mvmfltUk4XOIbOCsz56Zm56+VB/l93z3L2QZOipjkjng14P1tZrtQLk13WhDXlT2
Z4Zdu0ffbW+Kg6Ry4PtJnIWicJgi7ICvKj4Vul2ttG8JwMuYOFKQVAxUbKNF6AoJ
ZwXsqziaMBVnZZq+uvd9MG7SJjkrOs9GXA0tpg7CI/mZ1jvXuIHdMTCIiZd0CH+4
1nOepR2iB4DAzp86J8JRJK8u0TAwyhertl9aqvJUlfnAAuOPGpe0y0+X6M3sQqep
3KEXKn33v/rLhKMmO751dSC1iq7A9huvguV9d5AzE183uCezBMTFOWWDLNJCZNUG
cP1JyiHBEEq+xNBU71IGL9nGOZuOET8zpuYTwh8+1jf9uu8G65pHdQYZJe/OAwOr
4JpdpSxDnQadO16zR/UmVD7zW7T/XZN1lEfR13m+2UbNail+6Ez8ESlDzUPZjw/C
SFaEkQo0So0EcfheAwxY3V2MEKiYPv/FWiVhcP4hC5tLhJVqlBwUnLeXD2A33Jxm
EykDbqVLpknFKuNRuWJX2rhwfYbrjwXB+4FvFjy2eWsHbUGCmeisyAgljHwT7/N0
vKOJZUtVP0rsgxFwH9zXE5TG6eKi28m9tjgdVD5vJIp7zEUK5TEug/c+OnoswQ5a
Rh1PtP7LkHWEd1upYvDnNS0vttG0BdNsMM7yUlFswm3bbYfeVFq03ECTQvYUsAqx
7TwpxYqSnjFclP5BqZ6DZolft/WoI9BYeQRCE6+SS38/eZ5wOkW56IMFbr4bnfHT
KDPklJ8gm/iUj62HhzTwu6pXHLedh/zer8UbMI1F4GOCnW318YkIQT7q+PzQvS1i
hNH9McfIi+w49BEJQD2hzUTE0MlyqzWhuEw+M5ApmCWJHbUXgSBPI2icceGaDHGz
3rdVLTsT36DIpLX0Qp9pdXMcr34sbvc35XlySUY70ymDyAfZGXo5gjXNlWj1jkY4
QhTwLmgl4r/MNRZ23J/sHaUj9tyiNGBSeDQ66l6O9PGEpPfHjWN5+uvhuqdqMlgq
api5pciL/K/LnVKxps+ugSAomAzvSlZZChXJVFbbtfudGYX/cRmspbbgvA0cN1WJ
jp734H0NdkENfV9VZ2Svx63hST0dpQewyjpchRN29UWK1j0+0qflPndPsEwsMpb1
FuHI5tnycTSB5LsGpMxC7BnELfhkVcs2FIuu1spKqiCe/ZAX0bS4rf2OvoL4K9Rw
8kHyJrs1ZA4ct48p7qrMAhSMpnZqY7jWAURdP56InSrepAFnsokOghRixRi/HGRJ
/UdmtyxqX0Rlq2h/WfVfw9FN3VWdInIBkgT74kwzIH8fPm/EmSHh/5tG309Gs79x
vjBKM09ynJ+Dt3d3AuIPWv2XwanyISmF7fXRAMprlVDbChFhc3OPpkFcLOM6cl21
omu64/k4n1o9HCXb9k5oxmAokSNVHmaOzFl+gHdKO4Up5iFIuvLS+pdzq3Uh8WVg
ZlohuCem9XEoEckWf6KWrfzOVNkjOdddxpPMT/RK7hzEfHMTPxNxbs9orav6Wxoo
Ub6y6cmLzXEKw0ynqFo/eNPzD9JCUfok7TGccDpdO8xsuH6bO1vnTou6JRlfrLV0
dN+K6ngHCHHse1kVAk+eh5JQe3GCr927FrdPBgZu8J4ShnBM7ygRzvAf4K1iZJIu
k+qFWWq6jReXbq/u67A5LK6TcEsSSZokFHPWMkHZZO+8ZzgHGpM8JjnAbzMY7o6e
le/xPkDQLFj8/um9RT7wnVRYVB0QFMzzHmaM0LNo1ZjRtKct0eKRPXBNy5TJiSxC
+IJ7y27RyHVqIz0SJmOCgQA/e+Iak7QBvfDev/puCMc+RpSkZYymVm9nE4BlFMAW
UXhBwxYKf65Q7NnCJEuVz/ZlU9PECeQbu3QRgD7A+T/2KLmJ180E5C5KGX4XJRk3
w1Q6t5cbecPTDZZUS3cRIvKjksFIBvqDpsTFjB5Rsu5sYrFnC/sgVngieJ41Dn6s
CICUAVtHGyvcK+D2CHO19CbHn+eBARR8dcZWKuEZ6w3U8DuGRQl/MB2btLGj8U4Y
ZE/HWlw+yRGtuIGqH/0Azghz9BevVIT5ua9qNfzA4XO8U0jA6X58NDEz0b0FDO5a
pCWLaap7puOGN+njXfwvlF+weNjWguonLZSaExH/7Kh5Bg0twYuSfkM5VI2MbBBg
TjUH/L1TBKAaF5jeiDiNDK6nUurkRTSeN8IK2GR5HjFN67OgmZzjcNpYPRyY2gRj
N4NqcKtAzNVg7z/xV9AfwyrWjhcRfPdDHvGUYX4iHEje4Ed/DHUnfDwaguX/qNrx
KwbyA9xKmWxGAE8cV89q1NB6nu4yCn2KwKupDNfzhGJ/2udQt29n732dYEJKUarL
PvIG1FjNfQLuYgUA8iiycqJyfJki/otJ1z7e+JIsD3oRWAazLBXPqALlkPEwkbxV
fb090nokz4LIgxMMpoR/M5q/GMYOKYi00xJvthVGD6fpUEOx9COUBwEBslrraJXK
QnM5qEViXZIqLg6LVZdgMB+KEdQlhF9anKWMK9EedDXZQdb+FvOaEBdlvc+It5Gs
sLUkq5nJIXiruA36ECt9Vyx0V8C6Aa9MqlyH6QXUQz5+MIROtYPwEwZ1m5mjsNQu
KgkUfNa+nU6WRZUGaj8M86/ynf35RkVOa4Uub0HT6sMj4LtOOcEaPBR9La/VNfeK
fR7w/6XJm63s6EmHVYEWV2LFed3nteEr4sGgy8sqPuzWOZrYqgWNBsjthyGxxcli
wjabtYXX5QeTiRKNgUbT1GSlqfmtCYFzt4Q44lVZywmObOoPDmzCAMUm/i5JUr03
qcTTKPE5yp1YDKc3jMnE16doZxcpGypd8KsGkbwJpLd5xHJyFCtNGd90Y0RD0qCT
7+4ZovhxHUn36TM5G8oIM5C0jB2KioqDHMC78uNsHR49YihNoq1zjhEeyPfsDoaj
7jqebDTj4engWq1izJNABJ4D5T5iPSOT0oNiIA8bSaOmFXQc2fkyvcc/it92H0/r
sQ69Vrpd60SCG0aEu0AHXBeoH6dct6zKQLb/kDEfnozvPnt+AU6mMEnB10Um3bku
EFoS2BoDyRw9CLnjZEdC+VW3MUxtzQLdHkvDBau7jzvrSHWUIkfdvRpgHrDXcfgC
fLsIaTTDHzMnhst5Tigf+aqAq4J9FIcu9zjgImcZWnUKVWrpZZzYsBUh1Wv5Eyo5
/BbGlk9cPl5PBZf8kMg5iLpYH3BuluNdhl0rTpfLjjO47grr8DuLYkeYQFFSaP9e
89GOoUsAbNQBI0OZGBY9N/X84knPYoUtywhomHK8NdKFhegTfiGfRb5fEhB4Yi9W
gK9ntkyRon7dWLc3xkdbhNvopkel84Xp5Ia/+jru/aA8/hoKjgjLVG7A5tg/7Shv
ft02a2gmEaL3eoL/YM/vHlNrZh3bf0imjf4WdZ/rNAnkhweF1S06tNNSh1hRnyu7
eWsO+x4Tv2iMSbHat6/a05yAi8TDq5238gCgWDnjMpr3fKDJhUNprTSNJUNl5c2G
VEQMcOB9c3omOhu1qvyqNlihr9j3JI2of/RndMmSc+my7wwjtMwMq5R9TLeoaos8
eOlAaPGM2gBJUNix/omOAeRLI8h3LSEItv39O+CEzspkGfSCDCHLejLvb6U5nR8D
o+7yoYo6WbPWs8E2lyk5iqVTA5X8Dvwv0OeAbwYMTf8HLdcAxNWGlXG2HlwNgrbP
ylCx8XH7mtj97jPwDNim1w3xcpG2HWchdvKyfrLxboEfEJfQuEuwrbJV6vAV2VHY
hFqjkKLIovwQZuJ/Y/UqSGPgZqwqZPWkwky/1kg6N1QBpVyjMvKFiI/BhXpqMLQC
BGzDZAKLyQGT9cIC8eUNQ4rOYC/VfhHdwO+R/vEM5+u1QNbLeZwLzJ2eMUGRoywV
T9Rv8n4d08+S/gy2Y5ylJQ6WjOQq+kPUmy7t8LSbnQlgvWL1P6nRh+58/vYO6p7U
E8HefuuAXUWehkiZd+OqYy0S/s6+YflGzar5v2uJdoVo0pIic8suSkjHiu6kxPvC
NefokeSE16MJA1ximt/WdTPTSv2YvX/0Vfoht5BX5ldVLSGsDxypuC9B3CBlL8q4
Lfm/FiJ2/3lEQxlok5dw6TxGSD/EPC4VOlmw0OE6E5oZrgCCzisyn1SFySNMBlTY
e7/VYZej0GUJEAXKSxx2R1s+4qd/RzFh4PMXlyzsfNDfRYPDBlGVkvxI9DqCB2Rn
hzEjmDg4Jy8kyzdi4fozlfORnQ1xeqbcBWpexsDwYzPrwuLQ/thNWHqbzyjiM5ga
DI9BWl9eENjHJeoyvterfYxpgac9Zcn3tFo330h5efE4HhQBLq+D16bay+/7zfcQ
RDTFTB/bJg9IZn3dzHsDvhGQe8aFVyoYqpS31sqHI+pF/zNdUHlD/G/wQokwUN6U
uk/41dQYsWvw8XJFuFD/hVEIcewpInozE4LrhP2U/1Fw83dAgSj7ZxRC+lGZpatH
J2FQTAfIlK9oNuH08VE+AUVrnNXJNLOthnA3j0c8koEN+PIQB9gAWjz+j8ajCqws
SJA8rS6pxpZAb3bZhyr2CJYGEGNuTvFmjqoc2HAFFpI2O0rvny0CXK09MZAT8hCH
CylP8+TCUAi0+nPn345tJZ4XK2FwNDRGvv3mvTET7Q+5WqFw2RgHOjue5dFYhmqH
SXTkgedlPcM6exdyyIHQnOqlIQXf9o5F8Q4vg4bd6n3lwJk0CUrpm+dH5wTinMJN
Uy9TeLs3QnSnedfF61ZmH7oH3+lyhdnWvQWiCTUxiJubxBPEKYo0aqmLgoB1/qcp
zYaCCjza5t+n5CsUZHJR/nRzyhG8nBPDr4vm8x2mXWBqHv/9vbNmzXI5x5EweU1D
Yt/06eHn06rMkK32167cjhgdHvgMTDFcli9ZP4rp0qn6Ws3jxZ43GkQTn3i4tefL
SvhPhXJrAY+WdOwJn/GVZU2OLzn47z+ZsgDM2qgih2YdtEnkKyroisDBqDEMBGWX
Hc6GTXJQLvL2LimyA5D1ChoBCAao+Vlc3e2GaGJa1tPvKLYfJJ9ooGFrLpeogjS0
fEqX0xmD5Xkqv8v4foYYwQYlMO+l84z3uu8uR1NmGVMVSaL0LnlVlBppQapf41zK
bs8GiG5VWOfzfKflFAxTM7PZCuGVgdvdrFCw4JcSzh1ny+7VTn99vTLyC+InMGdQ
OfyRx20AKf5Vn7kAda4BozfvpzD6ioxiO7PIzxV2YYZLLZRhmacC1Hoa1yyMC5x2
6cS83aWlzKcL4iH7BfvVr/ejpJ1eQLOBIUYGsz6k0LBpwOCtbdyV8cR6O9x7yIKV
ZvyqEk+Lj+MwZBqkflE1n2nra9SNiZAZSZodCSUgaSKhRn37IMgfqH8th1QZqoqN
e++6fHV/V6uCoJqjBRVHn0eCgPOaDh2pMwufYOlhInUgRyU8qY5aweRClkYLgIt4
Bao4DvM4AawBz6xk9mEVaN3AsHbxwQ/javgzdksaN1y1VMMRsISk9C7rDSG/a81+
NzWo8ZxyNu9ftgYMc6mmtHl6+PI7rvs6amBstsTofOVxejQsJHdRG6ZJAoGX+Sng
+Bu97z7GzB1FcmXzSY5eoIvWxqdzwBAl/GpfHnLprNTIcVs8FrcY01nl9jNryuim
3Qz+KgK6zpJtLQIEy+R465E90HJBBnQrRZnp0w9trSp1z8A2E2NlX2x+31oDL7j+
7BZbjHv4ai5k9absqUT8FJXplVn4eofq1MAfy/GCmeBTjYq8dNNxg0wuwYt9HDcA
y8L/FM3PC0R5v8xqi6Z98mE2rDLvuXl7sGsy7ReowTRnEW1z/WqBdKegG+t8pzVI
SEuWlz2GaxppLvoxumKO3TUJprqOjjr07IM4Z+5z2T15ulOT6miHq33Ub/Z3x5wg
sRbK9JAOPJVtZ5gmfUq0acKimE6ZxrlzIdLdT565DfmBufBlKVcNEgB995xSC+/G
v7YszHahDBeTdagnyv4iUiS9pIcQrnUwGrPszJHeKlzAFId3H/dLWIg8KkDYWSVA
rAyfyMyKyNjP387KKowJ5TJTID1qK38KCIvvBw8ON2jXkD+8MYGPycNqe8gcdspo
QM1UolzIvb8n2vi5hlfV3c7YSopx154mtwQgmhlBTfrZDxg9BDkW9cIKc+5mkGcp
p8ibP2yiTHKs1HTq3ewhbbr2uCBGuR+3oIZ8MHdfVE3NDv6OaYPMmu4QFjM2jgzt
Jq9NBnJPK+B9crR9J+ET8yNrQ5ez0zEH5jOOHPwEhh+OHTyJnBjgOybObZbzjsmD
b/oLJiTvhtUTfxiVbsA+IVCNpxMIqH0GrqHlyFJdhqBn7s0+vNIi+2HgBbXABbZC
Cu2CZlrYGrQ+PETmpykESW6i363ZfdPQSxlT4MCIVOf+5TZKq9qdNR1aF89kjh0b
Mo0qNDMCf70HqzRikFtYgLOJwOafhCTtgxHYFHRVAB2F27uOW/8D8jw0lN6pMIJ7
F0sM9oS3V9LSp72kCRaZhzD7R/7/psRsBsUHILvtqgOT5LmNgLAeH5Z8IZ2chDab
dbLemEF9zQzUHfgakNC8sT9tDqAJsNZr5kAfPt3VQamj5NGmldu9fBanQ889dsmG
qI7KhXM6wzWuiwDAkR8+CsIfZe/7IJ/FI9a1+16+7J39FPQkDqpmu/c7LmLJlYzZ
ov894WCpyTkGUY5B/WcXad7a7GSAjYQJlgrbQ+DbgCrtw9VclhfNfgGLOLwJXBia
rKz7+9POKVAsS3rLkxv1+Z+2GtcW8i7CjwYMxpkvRPBWuYe1YGfkBp9Nnx6f7bFN
ek35RRK6/4TBRJcNyv/79wwJ1sMTMUNX2BgyLOHK5d+eb6LbNaPfkRG/c5tM/ubA
TxtXRfGOwGzStlcIkupUzNDp0faKm2GCBBs/EpkPaF2goXxaTj17sH4qI7IaQ2uz
rD5rtGGyL7fBusHikWlnoxQEjhoRhPD2YvFHPnB3Cf91hzruSX/Ge9QhSBerqvrn
AEqaLKBjCYnvrwV6Ln8UoodLlFOuiwwOnKQzL0Hf/N1BPNDxVBekKqR/EgkC4S3E
IF/ZbS4J6xlgG6yhIjsOuyB+3UZvIuOE9C8YlKBYLdtYNHfSk2+OC6tEm0XJkcQl
T4muiIiKaGDQBZp2mcVzESE6WH2m3oinFQmxyOmDfdm1zNoZHmj0lq1/XAcHYx3Y
jbyWQH+/f5SRbEYWj7JBj11bW/pp1V5+aXDMl5wlGoL75qp+f8gb8uv0NiuQaNNB
OgmtqdUMcq4er1yl1N+ZFGDY6JQalUsFVOV9hzK9LFRoEylshcoeKfG2dKofHyMl
5wfmW1NyMK58Nx7bEgj0M//dZYHGWzIX6razZ9WddgMM7GsOcIj+QbWNkNVwK1oH
Dhc7KYDvaY/otVN7ora7voNFC0x0EDvcHdb0wjWbCoCF9az1mHt3pHRvpfoMiG5o
AYZ93ojfGYXhW2rpao9b0yZlnMHntQoJNxsH9W2ZObfTGz3qpzj+qYnsGCr85XWV
dI7MaPKs/WnpLU10WlJvrdgvKgCL42LmzCHyV4uyC7GE6MTPZs2vAq4KDuwgpaR8
zb6N2iJIn6pcettw3X0GcXJnqqNzcIzCXMAY6Spaov977QdkkISVKeqwjkUYLq/k
MpVjN7qQ9BhqfRWr8U19E2/051Xoss/K7LHpEaRALaKugGJBhdpwxQpiuECLi0sx
Kb97gzXZYxa2bqgiD+4+QHBOc8jU/e8femWTuc3fbvlPspinr94fI2YN22KjHINj
97C9eL5vNQFir203Squ73MiQT4zRWdEgTue6CgDWlJX3WEIAGbDhDX+SBIR0gDod
r22L+eixmH4mMC/+Dj6eTAe4QejkfVlDepN1hzg9usRWMfyI+6zBJE7MZAELW0mm
HVUOFFa9+sqsU6PgTI9LAdh17i7tPFsc55Pyt44jgrfuPhrp840wa1xsl4LqlvIV
fFUOJDW+qsE+rR+yuO9RCpYC1SAfIqAoaPx4DwsOjTdwal3ruFRHNw1DK/QhtyvS
0DuHonDSSLCcZ0eFf3c2lfZjH/cB6AFM/Wglnj/fWTvhaDDGUMypcp1RH5b6Op9B
grGkHRFYy0m6W/nEVPT3LBWJAQO5NABKdbQWiu2Pj26Qw/ZM+a2LaOGr2cvlyAsX
5tVyVHgSka4uqoQpHJYwKD4XjfV3o3slX7tCbiqq3nwYwdxdQ5HWfbjZRUA7zY2O
NGN4aGTcqeZUGMTvUjT8iZnBNZOOZEAonPUu3bSi8tQbpasBT5scF/qomFKLZ1oZ
s8eETSUYvkHxXnTsQCWTljwMXYKevGq0e/MGTo3h0lCHztcAEbzYQtJtEREHxT91
ZNGpDg1hqRtjddFoTfdhg5jyUwjsXnh6j0nvwHhj6a4abkkCBxtIs6J5VHihh8Eu
lWDD1ItBTbJfL7pdSPIHbhVNTvZuP2vu0Z9EeAZqxc6qUjugqndrIky2G+krZa3b
Kf8JZibaMZx6mNUQ4rtXIoyFK2zm8w60Qi6ur0gSuicj9dPrM926vrha16uj7NHq
2Unz1ed27tkZKbIsu+3EqczwxSq5IgFAiZj670eaPfMP3tkGWrBjwViGJyM+rkp2
JaeL9aVW0GsEf07PqyuH18fQXlU0BwHKA4A+regjiyd7GxGuiW4+roKyvlBJ4QeF
lwSa/zPoqVuQIyY5gHHKgS4YaXE7OIv+KxLq+8pGjI1enswtFjWo8Xl5j0+52ZiJ
1JQ3NpfsQXurfv5jiEKoSvbhlhWHtBkNQcJMtlXTlY8oZRsBjSRt9umsZ5W/Rbh2
LL14PFD85OD0SGOpJ8SqeXkolJYg0tfrcfIEu8TL8Wph5QdLgCOZv+mund79QVee
wCtgARIfe+oyiGWQV0x0oVga3vhaSIpy8D7kjf5RlytJsLGYTk7GPVxp/SB5uAoX
BcNtV+QbJwwTv3pUtTUyb/Zva+YYqfgp9AaiCzxxqZw0w5N3OcBA6F7yR7o5qmL6
/SP65bWl83VkvMeQKNm1V7TON6IP1rV5oX3WnxzTAzsapUmEx5SSkSmL8NgLO/Su
rKcK9oKyxNbbEU3OLmQ6j87Cw6/rw9hkoM54ZWRlmuvIM0q5pGwpgtUalqEShZWW
Y7yjF779HN28cZK+07wxADNUVLer+9irRb24eJ9p7ZmQWGO2EW2pFq7czW+6UZUg
MHRl1sPEw9A2gURlM5fiMvMHzGQEWCK5c6ykv7iW3U0haCrn4EcreMp+EGhBajNG
/ylNyNjjSI80obcsbcWGiDQbUTZoYy8Eg1782owhcN0b33I8T6GpKa7UO/pF/UY0
MBqYkCUOQTeqwN50JE8V5Qn5hNZNWviDq7fozlWgUXR198qg9c5m1rNwrl7M80Z+
8IiOyKp8mNXlgeOxyCtASEJMiiLkQMnjLFOgSAjO+rhW/GuaWfbscjnQiuI075jP
5lxtiHjZAU6Pllzabb/v7bPJrk+SCrnUS+XvEaPaWZkaaPHdr2jL9iSasHZvlZ/i
ebyO1h/B1GBdY+WjLjyfN5MYXuLaTbwIMMzZUeQbEA/C3+HswvQP72sP9royEUCY
Z8pzNj7GJjSg7ifbgvY/r9RF3IgYFD2Z/ymmPDaCSS6PF9OW+T2FYmDJZX7Joij4
gGgMxY8r/+8E88CImtUvxoiu5MqSIBJY098XJjpnBMjTPy97KdxHJ6aXgpL0du6J
qPRQR9YEIwm0QVkHCU7H4lfvvX+7WbeWS57pEJhoxRNrJQlC1dsbtDNVBf1Je8ub
2cMUvYg9U89jjGdclqqjg+lz+EtPGqW58HsqGD/vZDixVZpbl2mEieuXt0ePNWCA
PIkf1lII5nmgg1ZRhGXxIaBJW4PkVye34jQMTqcFcqdIBYKPQqTsCA1YwD5uHuOX
yd+sh9Ir37e++6JvguTiyn6XLcNbp8KKvDlKUG9RdmpC6cs18uBuz1IgrGDDUPao
bfYC5v7T/23VgDI1QVr7JMhb1skXzMJlC9PUKneZ5WbRnrrV2+tO0yB4BVlykKJg
YQYf+f7CfsSD2aEMsUzR/4WYTy6bi3dXWJDLTXsHiADXxk2D0RRvx/xM0Ygrd7Tt
IXD6uVAF5a/7B5esorPpFLjqqlq5nlATvdQ+lJv7CyKoaugvSadNH0g3IyfK6U9p
bCchlUE4NINVufd0fV4eQjoXiYXSH9hLjpicBo0Ghkfn247QLEIY11P7uakh5Qg7
TuG/IVWjj5q7o0xua9Rxrzw2R4i+FS0lASR3QRaAYREy4468pWBcOIjT+5Kl4QaN
KC1JVVVzVeYm+xXwB/AZChe89p3IbGNFKdV4Nr7Bw4m2hZ1pBcdyWS/D83r6t1Rk
OllLWx2sZRRZ8nMatgS+5hA1SySKFTrANY9jnOVIxtin0tJmMbYyUm62XpXb4bvf
c6rGmHiooJdCnrC1Mu1+wK6k0LVO2VViYHxVbEs7BXmG/sDHizJ4mzkavmWvJQ0M
ZVBOIdGrfwHy+ItkhvS8T70tC/+vu3MFNfzsRRVmDFjwCRSQ1KYlpzFpQZJhjFQG
r4mL4JNPSc3gu5wUKi6t5estA3v0E9reoqDEcJaKrikwPTwIqpq5W3qFyBSNAZNM
Kn2i/Wx7ZViO7BNCrzTza5m8HvJIUx0K+pcQ476vrMikzB0a8ei7LEjlWHoMiygQ
pWMfp32LoJ7OFzAKjZ+WSHm9jZbFzsVcTpdzcGsPPUz0x/2ZGzUv/xcH/nDtAkEX
DaKOAn7i1T30KfXlZN2wB0/3CAqkWbcwgvYHk6NC/vsrEU5Tx11eq+fdPnZhIUNm
yZY8NebcSMDoB+EP9v4OQMRAeCCnAv4Phk8TLv/2QRDovPd6s8G+n9fPAtczGHF/
LCDCNF1jByM4RV4WeL8IRRqcYdJ9uCC2M8aaRoGRNZsQMKXt5F0JAJVlBcE65NGd
jzeblZI90BBxClq/kMXh6Q0DlrxxOgy01GCRg9FM5clRNRPbNDrZzT5ySf5kUiex
hkehkmqJJgoA7gGdtKCYRX34Z0cAQKC17AdS6T2KxRNiP5zhNZ7f9NCXGa1BYl7L
EkNn6evc2eXzgRODA9SaE0n7LwkJ4PF8d2TaO0OCDDHpXCxPC9HhkWW4vQEEUkxQ
JECD4wst/x7nHT1ldc95DVNf6KYmfpec1khLHXn8adTFDaikJXrlE+ykDjAb6njB
QOy3Hp9uj6bbgQXJErOvljU/W78WYBmaYl8MqIonT1wiDhA2l+liqdmSPtXZvl//
dEBuevbG+qpOUmcGlrnCjJHtXBiuUMCD5tvKwY7eTHn37qOWhZHSCBzLtpwiRQdL
u4nlbc8XPz7y68z1lj7vvVJ37c4oTVr9/N0y7m/W9GFBUMWrZxNftbBV9exAiVXv
5u38P77YmZqFwBB5RPBswqSGFmNITloIrD8jj7h+LLoEX3ty4gvWsxoAR5k1YUvq
iIbRPoSh33C5brmOU49eh/PhJzARIe4A2kMAk7acyGu4EtE7k4+rRAH+1ODSHYq0
zblMp514K68kQ7Gqd/5fG45jWS4BkS1hD+DoGbHlXO0ZUXGosUzGENE5tBlHvEFc
BuUwq8fgFwfTFT6XV6FOF8cEN8UUR8VUmMzMFevYlViqVYnbbUfsX7jm47ncKSMv
IeuRp/NHdP0jwu5TeT7l2bqPnGdNXqd7Q7bDO02WOSsl+f8n7xKPQCVbQYAkII1X
kaEcGripAjG3ZvhqQLiGIsx+bkYM0VxfGpms7o65Y43QLVyPh5x8f7D8YM601Szn
0SrPv3saPNGzSiWZ2j7LMbABVhvHf4qMLzYkgR45uJWQywXRfggdkbZ3lXoBZRUo
HyOjqsRELeUDdDWyCz9JA9FmkFkg1aYeayPjpLjjuoVzG3QAFaf4sPNQhY5dHnA6
p3+wN0HC2rAxT1xtt7FuyZjBBjT3+tqBsYM8AlT98PJEaGUnbkzBnPlOrqaw0F3p
WzgWVCCSbaitMw8411TYMB3nfs8zbMFSM1bX1hBVANvPGrPZkzZQdVeiPysB9CVQ
R9zv8WsKTydbQgcXPUZi7GC2/sJsq10kLsDu+yyf/+n5bCXJqwu7gqaSr4JANSAu
b87m68MkOwHvbZvoimJ/rGzuzI215rZYpQbhuxJwD7JC31Ps9ucTMgc8oJK8rjUm
JrnkTV1uZHfJAiNv+XZLt+7jj7Wi1erRoDw7MmAIRIC12JYsJHtFs6oZcK3paw3c
el3aDgUaYi0FHcGx/3WjKi4Bet8OtlYZ3CC7QBAhljYEfMOmJk93W6kceYt3eGSa
Qk1MjKpJRnmmtDAfTSVC4ml5aRJpGfKSchdA4Goml2VC+M6txIdpWtV8TwvW24QV
F2lZFssdVV6kNdPM25kbleqBXTMnso35UUXwGQQvxbhjNROYxTG8zXW4BmdGAbR6
Fn3eA3CFYbxMTjOih4Q+dATPCngpPHU69iahw1bIPlDcny5eH61J3Qj2w34LI9Pr
2kGzPyB5hCZOXEmWm9Zjn/3TAszlN7zntHPa2yznkPra3YPd1Cv+T2EhcvFnhL/J
rmFItktwyZT0GJNSYineJ+2taNf81a8blDQY7+sntUJX0OdDFV5cZrJanaQgpzXE
4omIN8mqOFzDmz57xexe89VbHIQYoSg99R2aXZqo2FQBuQq0sVpX9KhSXJ+wr1wV
dajc3cKncKU+S/aaxXBhNOpJ9Ff74JtIRJ3NwDt5fBc3GMoncMV/sTEx0Tj9/gaJ
ASCVHJVY8oNXSrCEq1lRP8vh6+CCADnItOKL5CEsI9Xw6+zxfztLHMZx/RM54l87
oCHl3PuQJMh5EwmSeule1idmcTSXdBjYr/gWV+Bg79GOihOm6CNb+uQ/21SC0958
UxyG/rwgRdgkM0XpGzpiMzC9fzlWuWupQkAGcqmnDNh9HhNwRirhLs60kxTtxNq2
2O5JwEEbB6/1O1apFZb5EPhmGuLYgoI0a0tAvhLj2w7ktdUXQGnrsyJjfG+y7QQi
jHaRZWBv2y7NNJFrqAyBo34rpP/sQgUU72FsnOHwF44Yy9pAvIWp7fPqGnmJSNwt
x0hfjNYrm1lM6djd1tjxWpL7yPEnnkzExCFW+udMvnIFhHM0kVxPA7GBTEfe2fIT
CbKn6U3MwkPFPwtEkTzyjLmeKaAFrDKkZ9K6+X4iYTtujOGZdsve9pw+mWXrDCKb
4lJ+rOjBpLO0eocnRZVTqgUTVNNp9gZ6C17GSEAb06Zu4J9q9EklL++WP+Zku1aj
4syWpEOVSU6gBOHGk6Paf8LuJ+a6XWKRwkb4V3H/0gcDTvFXlomsCEwi3ZDYEqvq
WZYB1VlQoNjsvM9kTVejpGX8dVQQaT+1Xswo/sKmDf+F2QpFRpUa7pmy4HVFVWZc
lVnV3kwkyPTk18ITLNmaWDsHNHscn6cVBOu5CAArzu3l8/bitK2L1gkdi/in0QJE
360Qwa9axohKR1yxc6wPDO3WC1TgNdPnNZ3TparHNUgiy4k1/6i6bflnfTbfsSw6
W3EgU4s96SHqTW1IFHlXnglDlqEWhoO7oaeP3KomYpMQ8Du7tN9rGHv2K4QQSy+F
E6T+mPKeLIJxm4Mhg5UaN5/JJfgnLEhznOI4O8PeTnZD0+AQKx0L4iPnirmJ8UKM
8wJB9sZlIeBPskNLTWDsyygKXKGanPRmfL3ZkBPkrRu2fqCuPYYw4nqDd3jpFD6Q
wSEtMZ5FgQ3VCvhdfbw1E507sMYUUmwl6Egrdu4ylZQKZKaKF5Kot9BTI5E/Fxtv
PkxN2p6BlDO6hquN+eBoAYIBG3TniymnUR422zOj/uUPkkW7RNn7MX4ZI0md1WWV
6+XM5VrFT253WQGJVNMSlEOGoqznJo+/wIO8Ro3QiLCn4AATZKexI3rLKPqoF8Po
rX38e4XwH3VtdCBueyZ+bgrezjVn+IjudFcIMoz05h3T7ueod6IYgqNrK2pf9XI3
vgDzD94FxuKy7DuKdP/u9pg48ybwzMuKSkgAyW1WfVLwdMIBnl6vWlhXi8YtcWo7
stw5xgihIw9oDt0kwW5z8M49m3L2NKnNuLyXZmkpEnEcW6XzYPREBb705oUOW8oA
OPjO7tKbcSYhajICk5CKyePOXZu9PvGN1jX5eaDnRE7v+f4cUF19/ZADpr4Rmyud
277Ux3VeEfyRhRv46A0KOUDXSvOgCt7eef7Pn+htVueRzCo4B/S9a7Jn92LovyBp
DNm1DZl/XLOPV80IoXsED0Uw6a9z8XByvUzWRyQotz6aqD5oxKWf+5k/uJW9vPpA
rCyNmUMpRd/9rpnfwDxus2+62+PeInP3yhaPvG/DzOhYhhGpa4PNTFxNhHwKosEn
pTfd11n7TNhpVlHI5PhiyKveUZ0T6tHCXSRcl/WJfOT6wAVwmOj9bXBCmb0BTBz5
Zg/SBGyVHlOE3atZeXMo6bbhhZi0g8QyL6W0CYvIWkxiy4nYHBALeHpuhc5l8bE8
5ZUX0NI7M726E3Zj6Jwswd/xn0JmB7NPMslpaMy5eslPWYW5neiFwZQ0+JQLjOBJ
JDYK7/g0TvJLg/WjjD5l24X+evXASK+H/HFzpJ2nGb00UgMrjOvvXj9/q/i4NePz
PbL+6jz/NGl+Fv40CCCZiLEKCXWMDLam8iADZPDI1t5rNHM9VW9X4EEUDNTFOH3W
j0us7cNj4spKRKXlxTY92SZd4tMd9/xfmjB0oUrQRwM3K37xYw9+6tbuQdTEBMz9
3wrVmYLaeAhTjUOH4uSzhoQZe9kcd/hxQL+R8/x85/REExjPxwRZUZqyTBKb3SoD
2+besyM8w+rU8UEoP5xcbrOYTnRz38yUvBMGUo30Lz/fxbYgOJL0zVwXdZJgbdme
GT0KkS+D+a7TQWsmxxrBRmlD6uUQWdcUXZR33ruUrK1mfB9IeGuDiK5gueOTQGMr
vKL3xlRtnO9ptVD5iGGzZ7il/VEhhNZje1bOk2EM3o3TKzJFzXaCRoLDrYuW7QPi
T6WVz13R+fkWkCjRhaprzH0eBOf4pmn9FnKmJAzo1iFMPCLxEWZIm0EA/ij9eAkl
urJlEiiwc8duBS8jP4nE6SSeDPtxdTtgVFOywPCWyo6x31B53sKfIWoh8FUTPWYR
jLAy/Sj6PdVPTy6MkCUDmiP6yzPyHYqe9edxgI5q9+66GK9t1Mr6ECnAv4jcTRpp
7Q8jKZ5woFcT2tlwepUFJzrGKwbpu+VELs08e9LdOWsFjKEV1J+cyfOzXp92oO3s
dE+SWDqZ8xHwpGsitixHmqfDFm6HRPAp1zOhNFzT3gRFvfW9bs8Pp3YpwbjXmxA+
CzwzPBStXL3G4TGHeWpmTwSZA3W/BE71drhLlNYIkYmGFy+bOsFdOmSMHjax5C0m
8ouZMWCmwqPaJjfRNY9KXka3HS4uBCHVHug5so1Ppmv/X34bU4ms+Nof4xEH9TRW
+AApNXBL0TkfyATfOVOMLmUqUKeyXVqhrOykvC+vnIM47cZhJlIZImv0L6fWI9EN
eq+/TaEnlqHZSBbXPbhTt+TRUCNRDsFMdu4G0hZMPImGi2Wt09MhXZyxdXlYs2Jg
r/DZ6+K4yGzy4wMcZMW5MRwx91BXNOMk5COdodZQQMKTXdfXDefv9Bk53pB6h0Rh
D7HZmnJzany0WGOXO4GNOS66Wz+50pBKLUVMmB/+Qh3EGtgl8c45kJNruci42TXU
YPFIDt9y+vCqcbiJ9IYiq1ngpytCKIkhbwZ/82soFV70IYfmbS60pB0Lkb3FAPK2
KNE+qieoQAS6SKGjMv9Hw3omSX7UokqW7sfO91BdRyZZpeyWgG8k1hsgWyPtTYRD
kz3yoTrKb/6xdb/0ynZDvlGTBs0heUz7cLmBHnfbNQXeyha9y423vOkVMwUnHBeW
/yunQGfQFRMGnC1zfi5LE1qXpSCa8691eXnoBRbjF1LyeNLvZf3Q03oTZyIWEhCU
DZkRa6KpJwLFRIjBY2UAsOezReEV0POuT4TEsDj0PK+QBa9dKBzDyfXLLZPptfsp
bZL4kczgvGIsKmVMz2egUzsBH9fazgvOj8HQT878WvwPGgSYXtR3x5ogD/inpRp/
/ovRqWubLT0jzPBLSTvvCzDSF8nYV25j7daYGlKqpMbWgs73b9t+psqt7rctgPzw
Vn+7Ez0FKaqOukkTwbZrjo56dbNTHQDFCF0Bj1MO5WejRM8GQq+nlviGHzR/Xr3+
Yzj7M5mIINd8jmR5/mYXaM9qIBlHzWV60NhqOyi8Ym0dc4rYSMW5ahqfw/OSjl39
V/PaUzDWdveNSczWAkAjLGtq6K/RwE+xLaY0w8HXOR0BY6Q/wJeclEaCV75mHwd+
GKz+wArN9jIOmZyZ2ZGI4ZAemZCL0UnuT3u02TgMphSAWcr/vcAJS7nu+qPW25jz
PeSkYDKJAyUZR/AGLt2e/W7X/PjQMomvP+i/lYwW1vm4e4WaoafrnBT61fNZa68Y
B9NASbOd2yGC+Yx7A808OoIfvjNcqHJA1O7mb3MOM7Yx4bGZ+UKDlxBKQSl4wqOv
vO89oDmNVyi93qw9WaPZeHEd3Fm3zGKjrGgF870ioSwNWk+xr6/I0FArRs/XMtSy
FMoqkKSWX1tZMT1p5ddE5RaeU+6M6P1VDyz8wymGz6+D+MW5dyfKAdxnCr5wlX8B
SkWBPkkX0X+2Q5ZIPN+2vLVyDjz1hso3flHIBHvO8xCQpV8KFE1r6O+gIu3ttqRb
93xmAnu5LQV4Wh44XqNMpw/TwkS7WOAX9oCvGODdiSy+stcFatKXYJe8qJ4eUypL
WzlDKDeorsNDV2C0Pq3yaYBHg+1Gxqj+zX7Y0w8lkgRwKWxpvf6Uy1HTNgv30tgI
RPDoWY8fXzxY2GtQDv6j+KaiYDNVJuN5KtPe4R6+8A0uwfA8mbSKavH2pbg4K1FS
vUrrZ3Ga+qZ0gvHt519h2qvPym7MEKgY3WcKIK9dRWQdDYAOYcUFiTfLGOHnQ2B1
gTAqfeLbkQcZ87Qf46qwx+CSa2iAHmgBT9ytZ7n3czQbMMnK7W6YCi+4grj9UbOW
JhzZgfk+LmpyYs0cLuBs+16T8Gng+I/jR3MeLaU2FYGyLWWg5u9UC3jDUg8IM1OJ
Ae4tPTqzRqASQh2Jn0Da+fa9GKq42LAaI0VhzMUnRVnpW5N7hs+LPDCK1JgvyoHE
LIWwS3+tn5Ah44iRAXcYEQUodnyCMqoClaT8YyTwnaADqWfE7T2optxdNTyk6BF9
sNP66dKGBiqak0K15XJCZV/TJ1QMaFX8vDe3cYmiwTYCKBhpu3RSTiUfLei2uMVB
8hxcKaXE8aoIO4w4FPD7L/4KuhNO9xesVhif4+1cGdxrohBFvbW9rscumGA/XW6g
n9ptQxktLMMHaKk5Ps1OcTY/Vuna9iFrS2TvjlfFl66ExusUsOdcELVHOVEJnCED
vk8ZkTTw71vrXS3YwdvM8ImRpEMjrjNGWzkiMSTwBejscyLgq4ZOEFmN10U7QXXC
tFnJt9TbPUqQwQi4GHD90TP4uBI68LMA16C41uIqRXEO5OrArzBKXfavtwiI+vo1
6ay9DF8w1umBj3Y5kW4m4/BH2y5hChFfBa04YCJcx2KhYXkQT2nqITXuUULOho9Q
SmW4F+Y2I6MZGudc0ojNpPBQsHewEZlgAIXm1UDBx+llnRwIrPUwLMnl+PmHd2ZA
533ClZVsPPEDEDlS6Sc8k9y8RxBy7bjbTI2mgMNBSntUfKWK423nnQ3px1sfQng4
8+IYtP2FJShWuxV4XH5kxJgkoijbc201P57AW++qJQJwsCwWi4N3n7JsDSlf3pUU
cQoDZDxl4y17cq9w1qRQjrsUuIDtxMMIHzNLSArP194qK+75P20LWMwaXUdaWbzr
zqJ20Qec2DR/WNAF5rt8xC0tu9AFou9KIsLIiacNAJbzb9InfKITfUbTj92S5z1d
Di4ldOl07FD+EnHR8W75qkrXfqcz/aOXSrZv3NAIeltEwx11Ka9bUxdBoAwzTAfP
s4xQEnd3QO58bVXLlUZGwGn73rQnrO8fUa1e1yfN9EaVJ57JH8XxtGJXsridPdCA
7XGKv2eCbQlL8Pac1dAoqq4wzVldmQGODKPCbxRnySa3o+HdRubI6NUZKhfeZlot
Q6eEtYWruuO5WfsgdtDwWlVpQBYw6cSdvJSLtOPny3Q1Jx2s7B8YQlBKsWWB/fJn
c2ICZwKos4TXL89xo4Okx/wn16ok36owLeg/lAbYJ3sCOSC7ppLd/42h0ap4Q3m6
q9UHa2X1L2JlpxKZf0U4PnZBmVbM/vNQTfq9x+eGvo6LyRrvI7/tKlhAjnKVI85U
8BGweBSqiRFhLWVRnW1RfNiDCaz8mJSHNAw343wv0UYDquc/mVgQd02+U3AhRsP3
wZVLDxpRmkaOp4zgQM/KNVPI/LUvGKTayLmO6ElbYuP00d3DZW5uaiIKfW1XViu7
o30dEjNg75HTK6FPxDRURqrRy4bLwo4t5NyMQZ73wd4oaSyRFK0zHz2jnIgA+GcL
ascpMJVVELzfh2z+Xfz1Q2As9xtNI7lI+huijH17mrDap24d4iiztQ/1bBbVmQ51
A2c4Ur5Zs4vMbMyQKOgAGH9zqQgl1cZLUubWQDvbqHdli+nY7KMz4fnIz7gPmKpJ
0Lw8uZ68JXm+jBogOQVUI2Pc2T7HY6QZijzgGd4MFUA3zmdUiWy81Qv/lZ+7GqoN
nVF/IDGLzhoN5dUKeSanItkt6qRoeSqk0bxj0US24uGD9oRo1G2qLYISv4z1eaHx
3vDVY81Z+RFERfxgfPSxAX+tlw+ycdmSCrVIli6Z16prI7LhSZJUXq9iZebNM1dd
6/HKq/MOQbjHrna785NzfS7FMIowFiHDn8eL4trAGNuI8DIkpiZaGY58rsZcA0uc
O8wazBgYO2BO3klFggHFzC7nkQQTPp0qOZGOp5LpMG33PttbWyjfZbjHYvVILfJu
uskCkNTNz0EdBYLNxrN4L945FKgUllIhozgjSahrypIOq2kSuzNqPYy1Cytk0+gk
pbmyRmuTiHqAAHod6SyCi+jybBnUBKkt4+geUp0hdA1i+AJKym8WsSUWjNaaUrw+
6lQxsHwF/7SCRqzmkEJpuQlb6FNh0oHwv6DOsHbxZFkhWkU65JpVTXELN77f+bm6
DIaR6Kkw0Qcn/gphVaxEoO38PTBOS6ErorqiTwCavE7O5gJhxNCWor6XdPH8Jx7m
c0P0zZ9ANhrPasYiX4WSCFyMSDd2OzdN3Ak4oqP6PaId49D+wRxV31o4634CCORv
q26pch8NWhQEL1Ut0uHWt8aq7cMhLMyWnd0zgI0cSSNKJRn2x+GftxJ+Uw+AOzoB
4KfBqbZEtBDheo/T6zKhUOSvwdAJ+bv3ntJvaTz6UeN5ODStXTxVPpPeJ9YVk23h
1W9n3ln44+Ag7ey0Guypxb9RkcXAAuiNTsAeuphY1f+keJbXdpq0zD36207+5bNw
4TCiaEs28zOwQdiFpXZS3iTY/PDlq4NDAGZfsmGYk7jWrQPqV7Vz56iarxZ6Fp8t
M27ydEU6sKf+qz6Asbwwct9mAyP34k6pCyVoE0V6VH6B4D/Jj/DvJBiCNMQnghAK
HGnkhiXvBXuh5M0k7F/oZDyAXqF6ZDFIo8NNx5NVLWnrtprkFVaRX0R1yCbgRAEk
XjmjxrWcz+X6/4M8erUlHYgH8QGA5lWoRVd9vpDLO3b+oOi0HIHf/TIFzz+llfSW
7dYydROwkXHwgBfBc/Qzw+lGsJRGHGRviINrX6KVy3MxaMtZG21Lu2eCiQdWeYJw
J594lPkiDwVPIf8E7/OriMF+bTVsFhvxrNqEZicKZ/2xFFdCufKvuBwMlw2jIJB7
4BTcTzHJIkXQ7XUnSB2DurKe2NRmGZDrsGoT7S74DQxe/JJjmeC8P0Zv4kDxxZ91
pd7DflIhiRa6JELme4AdW30mPSih8ESzHmropP7Ka8BcbOHY9lxOdX2sqE8mDfWn
kAeoSWUa70QqwL3wt46rT+bxlDNOH9l8jPD4l2zdJ3o2z0bPlGkSMr0SAArchAA0
8hQ9DRTyTinYJQr81MvwCEINvDG93IsI7Vf5iYk31H9xkDrK4HfEWMEDrLyyQZQp
0w8yMbjckahs3ymcn81e7kjPY/5fXpMJUleaYhFbNxFRojSAaXyw2RKkGqLFRuQr
OuASAj0suhOOzxRGEWxm/FIpw1LjXTiP1X/6yA/lYFEbfV0Pp4NcV7/gR3cMhk3h
qX2YCWyScgo60Qi+z4QRmfm3TV5QePc02p2tz/ivYRLeNtbFoYVOri/BQdWxPTT9
hZosRtX3PaLZwv6NEGeFZndFOkpElWBBMSODViNey21uTr3XrvDT1OGbTkA9NAKN
ELV5iiRqQL9Hy6tr3onbcJDnljVU9tunkB/1TU02yUxWJfOnQkAUrWkIhzvefODm
j9VUpY7BN89dORZf0LzBxQZ1uuamw4Oef8jFV9es9CgWwZIbaSCoEvU2N1u5mTgo
f6K32O+zO/GQE8j+mTKZffBvhxBQsuzLAnlqftBHBzUHg9XmjcTnu3a/iHd3NHla
rZeDVK+bKII62rq/D2kCzBugyRRVjezScuVR30AAseWkFibXX4mlDjOo3/VkCj0U
oAWGDicKuUbc/Mk2aH1zpB+Kwvmt+ndsBNXU+PNIkyVcJlhRgc54cksz7Ug+h9sF
arssQMdcV49TfKBKBnZ8FXxNpa8rktJ8AAW/o1MdJIVp3TkFc0unoL3wqHHGMr1Z
3Oqwiz0NI3n270gXt0hL48pscWBi+tt9Avaho2rrEljdUMzWcmlGTgkERqR+T8eM
X8AQkxDmSZ3CuVMJxGC9YFtTkkdRx+EYExK1E4i2/qQDlZI9d5GnhX/v4TGca0Gg
lNzQnbr7DTQQLm0z9F7kQ6Mj4uIfBcrZq8RQyNowbSgfIqne2u/j7QLcV5ANgGGC
Ak0NGi+xCkkkFZ09Drx/M+DqxtZuoRIjuy53Ob5Kw4FMbHPurJBvkuZLwbdVaoW3
aG6HNFn6zDwo5qVA2Ep7lHrbJG4MXwcur9oeW75T8ezwe/t2sd0Vli4gQe+cQL1H
7Z4lW7ierY/XnbTnW63ksx/gdj7MDgYADx1jamUlGLrBshH5U/cP/Ne3LALvyK51
WZMpZ+MxK45qlm/i1AD28LoCGVJV/W4Q2XEWcHEkGt33d0vPGX8+nHqmQUphxLhx
8ppB+PtghexSsiqxoFyqfmepK0gBz84VpSzsKMWmcHR/zEog0uDrqIvKYfDThF5N
PUHNSHXEf//pTWCfofF0FwJDyND7EoTSh+80iYMZMzfl9G8LQBXd5VuDEYlIcdVB
MIK5kvXJRqPA2597I/66/ABaLcEBWS0r4crVYVsKVMDh0cIzsWJOCsPXmqJFVVrx
PSeMdWivLi0AKcHmzBq9mk4xCXpr69thNOPWp9P/phgL1WAUt0BjLQbrA/qCPZUv
+AybzPHL/DgFZQlir+hqLTx3eFfwwZoCuCBe4RndzWOMoe4rEiFVCHLSB2KPiGja
JgcurjHYlMIQAKhT56vx3TnQXvTKSnyux0c/zjDmBUv+ncmtnZkmwNordyanrmIh
1rOYW+NHbqv66wScvzWKD9fQVExxF9H1q8pnZR+lNb2n0G7gnVrPtnpWAnGb6vP/
Q+ZSKYUS5hWjnJBFi/RxdDp0lv4zZV7C/sIu6cJcbpxEMbVQs4p+QfWl1ttglN9O
rupqfpM1/f69zIDIgmNsGQo3aZDF3myHXcLVuZgXn/jm+rE7M9zCS7XNK9nCw+4k
TNe2TdNoBHZ7TgFhEaZZYtjQqalvYDLEvYS51CLhmE1eu2AjEni6nCv3nxwOl+Cp
Xp4VaElF3xQjZW2onDdt7E473LgiqzymF0Y7hgowneXIcOjL8RJKlJGiLhOq+BeY
RNlvFaXVsWzeJyWIk5yM6HFI6KPPGXT1phDk+uKvHey28Q0jkopi8AoBFyCfOf22
PxLciogrveGJ+4sYTAxqWmB+0MY/GUaMaXyK4nsoaZVp/yHRlA7p5NgLBNQZFZaj
36eSOBuoS9U0457o7ZRXVL7PZEUAiZEhd3/y2kwmxFRCNKEwLe1dAmV6LYet113r
YqbwQtKqhoK5Qw9EKIEIyBW7Wm5iHwc7a9kpLTcncA0tjfjnqIm6xBXjOOPaaUEh
kBQhVhtyOKDjqOSK/OZp54NxKqWnC/IMcheIWQ0df/UiiQnf3WwZxTwxrvH8NUcH
VgugDRHkt+CkEny/BWegppLJ4Ir/EqUAYsyom7xi1e2bwzK3vmpTxZ7rIV4CbvRj
oIhaAWcJpfl6PAcZk+sGXvR/iZrn2nerNAn69qDM6d7+v9lfvwyBUzyUwZDbjb/S
AxpZCQtN9r/RpS+f1KXS/sjpepv4Q+s/bewqbfruBasTFdP0ApQXt2fOQ442+ova
txIwRiTQC0o6OgwBwW1Fi5Z/DXzKYXDevpK8Ui272FXsCwtzbOtuZd6pRw8cuiKq
E/ZL3/qZP1/weJMcCqo5MHXK9iqo3xK/DyDHAnAE5o/fjtfSVw6t887LPjfPU0QG
2ssUDDRW4Lu2xZrWUc7Cg7MfEUHKUw5mz9N74tM1pAtAyO5slzVpHhJ2U8g//5hh
kRKefzML6Uswf+yzqEWzXaeNDmdoo116guadgbxcRY2x/jLOzUBB1M/oP8fPvt8J
JaegId7/ppoQkooJhMiGJYk0zCGm9v+srNq+bqtMxoEs4OPitQ1PgfFCFjlNd+Pf
xv3SUD2nQ7cUnCd1D4u+6MtRzou2vPlhFeprNuTiYVGtEGvLDbyGMGg6gZcogVLW
qCCD2tMW/GSOqRJW3xs6gMg1CiRuombBxbJnbKJkoyWEwJKmAjWXSCowOHtT6Ygm
7QUxm/H3euV6l9sSnuVvpjpL0QPxYDr/7eOeKmI+hq5nj17bfwqfhk4YCK6z0nyK
ayX7F37387OPhug2zuglHsl7CSxgkhNyKAeXBanu/34AN+Df47GMoVEwPwwF0ccH
TQZ07FvTAb51n5HWArJCYXIr/ZlhCw6M/fUmX40RYpFdTlFLsHTsFsZl672w8W+c
6Z0MWm4MFvVuF7kklY0yAbeOS/g6QJc6sDGDJituQGpcSzV3RBKELXPClWarcliH
u3szlr32WnscbeBC5XkxB2g3oYDSt8zmToc4jP6R0d9JdpmA+3jeZgMjTCAsTrUV
kOvozAZZJTZ3eg91tlypp5MVIWu3M7RP2zu+qKHyl5nTVm1YmqmVMP1/p/GBqReK
tgT+a2Qxg1zdOCMRk6YTg31SDIwQY1miF+f9CTaC4lMiAeANQEaUVW4Hs/uJPzch
hOjEx9Teh9aCnWJHAMnJSMJHl8zUOvUz703MnCwXjXcXATJQuyk1DWmZqbKJIoM6
d9jrw4dG0vTaILieddVpyX1KXIimGq8Bh+b8Fhyt9ESsmo5omBpgIO2VaS0KXmSh
KyaZ/q+T+5aYk3lEa/vI36w+LkOHSjKI1nwxyNdbv0nB/WJu85Kk7OeAsP91ZI88
RNPOxh4hvAotr5+wzHv+uIsJVMIj7sRwecEPpPrvfv+hJbjj6r9bN7tIBy9u60Ti
/q3AKoxPtwde3YobNPzoYsAw+kVh0QbihjbB7V+c3cNI7r1pMbBY2M0AeXLFboxe
g6wN2KrBdA/iT7sbuC9grOf2YIQYPznEOIxNNjr0LCkUq0yONyszWwtqhGDmQ/Wa
hlnbUvoGmcATZgdL8PV1Kw97NyZ0ONpyg43TCJJRLS266sID8ZnUR7rQcl2mbX2G
vLT0vKvTn6YJw1BstJBw+hvL2rfNPsbDLeXaaZ/XDWy23fG4m9Jl4itiuNbwZv8k
x7o/BLX9xw6fbEY7WTJIpjrTySpTJf91hLDiXnbZWXzQ2rzna9hXeXUWGkknpFJW
kTII1bu24BCnJP3pTWzkoyLm2IFN2D2woy17tYZetV5C80/i22VAGn2SwvrhKpFS
bN8UZcRcadxhMiyp0sqtVrTWcnSBU/3AJYLgXtbAva2CGR3sPpbSdX7we01fOXCm
A04LFw+8K7hnn9QMbo41IIrlL2Hrm7dNyt/p+nH0hAzym5jegdfEInLfICPx4yhD
hs12n7fzSy2HcVJe+DOOOtUDgbuMHXSm0xYfuvcAL+3okOZ3RkQmWUN56Epa7B0M
UracRQ4TYRfpZ6i4zhPwCp3Q6YHRjeu/HTRN8hErJnrBq+vwziFWonfgb/E44fQH
sKGg8QBE0NU1ySn7C7vLq3iJ9atc3SbWE9UL4Q1Y5HWeFZ2aznEdsQr7SN/MFj0l
vDSig9i//JhBY2TXPHPakLl1mMVau4ngMAY6JgsahDqD75/dFzg/Qwbv+eLey5si
jFUhAa7ShQx0IcVTwXCzsOaMUX+WJ49FtdJx6fYuVNDLjvZKTmYI3DcGyqfBUVSg
r2d2GOw2zjKGM2b9wiwcLo5/G5CMIIksfVrbBFUXwb1vqAFbkLxR2tHkTugNjjd/
IhNrBuR/8pMkYleCk958Ti/V2U4UCTpK0/N/j+Zz9LBSX09IeiERtBRmyURK3mIW
OagP7O1Xc3cpf5YF1YlRr9O2YRS5S7cRrNLt+d+SLd/4jNoFruRUVjZ/Mb0mbxI+
RPTxtWxT/4syQ/+DkSWBGWz6dpiwU/ihbn9VDybbqxeD0kCtlPnhHCpqD24cOTpO
wDCfypgRHXAJ7QXTg8NYh2pinls+3hu9X7DxCPg/MJRGtROGthrsypM14cOxl3js
lyvhE7UOmt/x2yW4FN6DYbqrXIL7HwxKgkWfOh54mhu8noYNDzSZDmsdn24cKGss
2e+mwGDSs/qkw3h5iy5p2oQNAQmIIQ6hXT0UA+EIoazub2qtGIj6uzaIohrdJrk4
ehbLAmjCB4bsAOCeeUMydvQllQT5vTDGoplP4HewFhIMFtmdPmY2k8lG43HiN9+f
PL+BbAywllznQHA4lramV7AVEs/MXFnqqllErUnaKdu8DpXlADa5dtGO/7ObEiSx
9kmlPaVBO2NWd60sC9OHaYA2TwoXoklhmjWMAAJPhmUGjSzmebgpt6swa4jo8Mkj
wcvDjsEYcFuduBWgNy1zcDkcdnKleuHW5N4k1soXYX1ykb26NAQ+aeIqvvEZyHNQ
iCBpab+fU1IMOKyDm4VBsLQHaAyeUo9uJkVbqDordXqgn+AB69Ka/cVbZwVrsxnS
5s2OwrABMhDX7he7NvV3WOieWSrpnYV84yKNbhfN2m22ku+MfUBLOf2joYJmygsk
JVbYCHI2m/Pso35J+JndnL9109bBaGMQgO6r2L4IPG2QedC3+OfU3okaWf9KzEnI
rXDtTk1OVGVyKl0yhIxK/VAka864czYKcGx/vzRita5TcBb/VCCINKD5qz7hvJWN
zxjwf4h/GA+kqFSxkqmjIE1rF2VXhz2tmTeO0UG09gh5kllqs0z+5iNDWJEjzlhV
TvEY7IDRpRruUYqOEprDzhi0DDGL57zAfjGx6iJBwWBQXETlIlxEDvi5/aNV5lPK
4L5z9avU0BU0SrcXuaTKD9hHxGqfBBg7cKGJL1P6usUbRs5hBl7/TJsWnMriZzq4
jLRNN5kFENHpo1hcW5YWHfvkFh6Srt5fMLCjUSfV+8kKDqMtb5vmCaXINTrGOVTy
0lTSu8xT0+AkcQLinCxN91w9hCIjPDsJJgPpDzlwDyAUUWtsEkhMyodZ8BPbEIBp
8cSJtV0IvXh6ozwTHwH1uKsHyjTNc3A0vMNG+Rfgh0srkd4v6typ9lWHVTcJYxYa
ZE54Ek5m9DmzanuIHrlfICYjXbz0USBvd+Td41RtkgChRAaL3H+gYaZqQyAIWarV
DUVFPBO1jw+4F6gbnW3anvIwXEs5wrK2DXKJwhAXBfbr41xpiImpI2YPnxHrFrOA
20YfQ4pHoqVuat8f3vtErTvcWBwwg8vOrGfUyBCl1utXvsg4BAqtSiXx+1Acv8ex
hBrXGCiJQPBHmMl+M2V+wTtk2KX5331F/zMsZKYFzGqYowMnOrLG0Y+z5942LdKt
z+7ov1pbs43OgmNujAKIJ2bmPp0jXzbYZp1VWr6TKXM=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Mj6oZYzHIgb6VBKudKCpGVEJ8dX+7+6SdXfsyRRcC5aTlh/7rt5w62m1gVFwxdJ+
4xaUYLen00FZoBq3LVDOeD/WpkfykrOsWb/TcjxcBk1/fytncI3nl1oxQ/DnQM1I
Z4LadeAR6uZm5uv7vqN4kQRI20DPUOwgqJePTZhbWDY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13248)
oYMBEQWWewu9L847rbVwcSiFx0nWNS39Ca6g+kd7GtB0MuBLuO3PXeVnlku1pKOP
nRNfGo+tXA8n44kRzLTLxdLEJXpPFtTHzHr8Nd7SduksBiEierq0gQfUsgZsZBHt
rBHdemX0dH5cGbF3ArhY6apWIIhldZFv065WNw+dw8T/gsGCztMGa0Go4F7msNPn
rMG7Na2H04M0xFqkbjTIT5cQ1Nd0bXcnbFQIsNdG4g7NAAS/nYFBkVZk07EcVMQA
/diMYu/7/ZSkkzF31OHGf4yZXPfNhNVJctUkcxwZ0LynKlBZpFdadnp9ToADmqab
NNMKSLZ6eyuGDKk5SZa9/a5i69AzeWfqONqRpqGKdDMx+JQcJX6Bw5yQDucnhSS8
j15ZDXSUYbOM7VO8CWiW1wJ+8UhSpZo3IM3lSGnuQcFHav7zxMiaq4RFH1dXvI/i
tC6ibpfdXBtkKnP48niNUft4bEkcLO7ctmNncVWGSC1cILobLrultpXH/q04eQEg
Ww1LlTRXDYREI+vKCgphN7S+2vcq52WMro9Tn7QCCHT66YXnc7D2oXUB63hqkF9W
eMzuPrmhPpRX3cNq+eE2mO92dvHq7iEZS3NHGDZE5sGqK3eNUeeSJYVDwAjs8t6o
l1X9X0tu9gBnbHG7LlTypuooxGjfybsD3UWa9L0s/6DsxPBc2KlN4/uUkmINbEEm
mHY4FFwUmAxS1R90P2MwpcxAiBrbTdacutY9OALJdQXx0cp3KHSJvywV1gLsvAkS
OKmHxPjvZb6hWItrC2lJc5JHeiYcI2qm3kpW5TZ8q+yA3XpndXKX9DiLkBUq8GY8
bPzYT8eiOtiIl3K7mzFKgMs/omnwBrTYHh4oZvd9bqb0vUZrDv50jDRDvk9DIUsr
70AITuO9pPZJY1WxuIq56W1zOJVxCNwEL+qnecjFEcDgrO6uNT9/qH7eJtvFwgFk
XeVBKm2I15XjpbZnk87jt/diJK7LmJMNTE2UOEw17r6PkOfttV3o7DxUfy34pI9m
CuhWRoi/2plGn6BGbzIg6WeZeVfH6nsJruKW/3YExApNqiXkp87X74ptotfjfLj5
f1ZXg0vtNrXTG8F46qD7bqMQszraTzIYE4A8MVtId7BRTEkfU8imIWUaypyco3I9
Rlv/zQl4BGbDiGVp0UZFcfuD3XEfApaIyjRZdhCIDgUpcEfHge5sONXISufEFTc+
Ve/WgMcQAn9rLHv4uymbh5cqDFPD9wcvBHDeQslBOYHOC0zCKrRAkY8/QP292R4a
u9KvWbIdDkrP4zbO/Ewqc1l/eNF7zW2C3LHsSIBKdh2eGM6Sor1x9VQOonCLOLj1
Ifo9Dl2WS26QOCqUb5pnDSQ+/ccvFx1TC6eg38EEionWWv7aJvDqNmcd3Ygez/+v
jk3k0OAGDhtDtI8UJ4LkOZ2te9Xdj8rv1ciKGF990rjG4jOqS7MU3nipimAE6LH5
bWJaLu4iYZNCgoDz/ZPuwSBFiTGsexPWlByDVhAIqpYfOus+AW7k9L8Lpf14521W
STHW0dtIRA2iDYnA/QYskS2YBQGeDbcZPDhMlkC1mn9hn9YXpT1DBljdJ5TYop6N
0DLG0W8IlOnaypJR1mN9EXB/61eNgTj/iyDJJ4HATfWjQjT720QhlydZjFtpv9zY
h21ga5yNww1/C5rtvmCz5II6qFbGYp2P6mWUQIBCtGCQ5CLd+5oP7CkYtHyKST7E
NM7kq+bwYjBLlleiCSWjJpdtCsQq8fAPUYx8PqIfa+CLRMf4rD1voM2/9k7uYABk
Qi+doPT53378tG4N1C7adT6EzAg/JJ20XJ46rRWDwfdCCu5DDAerYvX14Ugr7MM+
91SgAE8ciJ5SXnHhes4ovG/oXHUp0P6W7z4jWDK3EpXu8UByBg4BK+BNt/O8cMXp
pJ+yukxV4IC10/sRrOX+eLN1p3RLlbSYvGDsJOEkmVWyaRoeAWU0q+jGoLBF4w3o
k/0TKmKAdpZ5KHvzX0OiDX9BjxLR71dZdQtq7dKnL3p51A6ubNwYIRv4Z9UL7/tT
AWbULcnGr1DxUsSNCctiAY80nR2/qCSQis+vlnpf09wds0Os4GJF80tBK+L9b8P9
VWljiGnQH4mq5L1v+DroNSH7UiZthXd9mqXd5sXbYN6aCH0O4y5whtAlv5F8R7R7
5ISVYRbdoP5+qL7UM0E5RSiSqvN2qZNX2le5kGi3ClGvvtsCJWOd/+FIYMJu8fyj
UMFsPi79hhaDf6batnh3dY2YY/YRnpUMuWXdBG0LzHahwdw662Kjs0EWXvoGIcc4
wgLiUmLyJFSkn+Xe/iMI8uGUnf7T2yf5RDuotv4pFsz707YqcGD0JSWPSU4FIITN
xAdHtOwt2NZ1D4S8j/FcYmqDv5yqFhYqIMfyO2a7wXnZTIe+RJ+TCJfDoocOhgFS
9yuwroW1OHHC1vh/3KPiKUkV+MGtYzXfKWXb6ILfwqY9x64bAk9MClevfefW2V6C
+PhnRuUOwv1P7jaKQEgHfEk+hDAZ1mL+IRWCy5bDIhmBmmgtwWqeK+NI8biLeCEy
aMhMelxFme/tlmkukChQUSQRdAPz+qCU64y6/mgB/yLXy5zJOauGD2Y5m89PsaXf
Tm9OmPYNQSPdDuFpLZmLnJX8Wjo4uSUyysbVNpoU5s+0j0inXUvoyJp8t7OHZG34
4yPUZgsy+tG7ziTvGh9hS99zvYAsj+YK48sfzJ4fgOSpsvuJ+i8uzSTHOyck0bSg
6/WrTmmDjOBQZm8n5r85/1z0ojXCIiA1toxVWMGWMUgsDDmYO/59dAnfdiHDiD2t
3ZxmPTnntBHZ8ln3YWF4bCcGCF0UrmiEwNxvECkUkqJ1loZLlF04p5igyd1whLwv
YjMcfpJWjz0i/Dgn5cumf8aO4HfxOSYT96d06wHfWZoeblwGSCMJD1OnTfx03uFD
YQ+iOGV9gn7y138ffXjBs+QnL+RoC2ohxMg+LvCOC0bKhA1PKo8W45h1ZoB++awt
4EW4wkI0hCjsLLmlfYGeuAmej4DOC9XtNRPvxoOudrs+ZlMu4mVo+F9GQujZAQGu
TY94IQsQZOIWCUELBGhAAI/q5mWAS8VnoBdlN2h1tV37KfAiKfapumOWnlEeMVyQ
I84gwXCsTmoxSPrfvdpc4Z1O5HaYhQwz9rGNBpbdZ9ho9uzAB3qoDMWYBgZpG0WB
TtDtv2ol1uZzeEInIzwwnPOhm78qdtg4H10zqnw0JvXUKR2aWPfSU+atJWKEcalQ
45Z9/sPMNbTSF3O7sSmQ0ePoUY4TMrYfG4D5OrRH/UKsBPRN6DfhgrCKuW2kmoXN
c4ySjTvYBGzu1ueh32pPL6Qj9io84tTgNhrrCC9HHtdMBLimNGu/dNXTTaE9BhH3
lm+upvxNxSxMW74hlpsqegd2/JUGXMbupuNtFmg/pKwuO9f/THHeOPXSBiaddSLR
fvakhhCXminyQQa9rTqHi+ypNhLalv8ldSTAdThmwmFS+yQIKaJXV4WisrFJg5kN
X7FA14HQtjEq5vUSZmTgcQMB8q9jV/3HhFIhH/sTC6JOAIVUy6IiUaYgcNMc3kK5
4xqoCLKQ3PtA2CWr56DgdKM3VHVczSz1feuVyym1i/Fykzu0nUAEqzhQSlkLYI9Z
74ABelQ/5+bz0fby7RoWtnNcBpTfjuLeT/p6mg1TaEJZpTXZ6ZzT23QyKVS3mmt4
p2h8TzOTkkblnUCFnQwO8aDqhNnu570iIXSZ5K7wFa4+lT3iRnRwnenvpvjjXCSU
DJy9KSSUKyWGzHiheWa9LaIhqlF9Iy49ru3gGvuHIoU9FyFGmm6cyoeMteEtg0aO
eLYjMLPrWhFGXn4O5FEvF0BYx6DmYke8n6raW01ubQr/qZFqTnkuqRjFzDN5mqYr
BcuZ16tIP8YIEIz5RGUVoGBYHFUYrbmO++TZPX2Yh4kUpn3VnJxT0bXxMvDfzrk2
eEflnWsgarJDk9Pt/2bbxr9VfYslY4pWT+6J8Y7O8Tuk+ohsUquo4FR7S1Y9KZSC
Uz+dXqr0WHwdjmLLDNJzo9SQCMY0Qh4EBLhpIchX6tcsYU8AIauoB2tdaBGmvS6T
HKndJ+t7ZE2ZojP5ptzRfiF3S7tySqUbOd/10MRpg763tWw0ksv9LH+PEFTIydZX
/B0n79aB7j5LLI12PobrO8Nzs3WD2m4wxyzSHwt5J8tGa1F/QuUcymJ4Z65eS9oh
mouQmEXIjSqZ3D7uSmJy49I/99pSGESjKgrvJs6lEqGmqQu/2J3pZJfKQ9jMx09e
3OeUdZKIcr9UgRGH7lENEBdmywNTS3cm+9YITM9T+INVx6dVslZ4ACKo01NzyD+K
PNL73gXFPClEGAR9HEUYOSEA6hbNmM2ZS9OWCAzFVWMrdaGg+O9lePc9StAv5OJ5
Bj/p/nRGSFGsZdBLBmtRQ4DkvEcGUzYMgsjPd2CkGo1UPlo5Wgjnx98aGwa+1/iY
Ezn8lg6/cVPJdNFpr+iB8CTz4I64UPDYWdqMiOkP8vzQY2WenwN9QM35XlFcVyxC
13iEyKQRrgHQ1s+CkuxrRkCMvQKMCoR5YfHB+sW3c32BWWisoWdzWu94NzI+0APK
ZGqxryuXrVS967jr2sTA5PX/REBGjAUpxiRRFq6NV0COc9mT+cr9x5Uoy8F+5OBj
bu7p6BZeb2ekj6EkeRZNCqpgxkjXWbcJ97X+Pt0QzIR5Wt3pDUArDDD/SEa5UrVE
fVHzaymcZmwySw3IevyCoHE58PeWYNWa8SnIT57Q3zP2WpfV5kodYLsut0noljSo
8EZtPSV4C38hL7x/WYOs5BP8hkeuAkIQonUdJg73Dk4EHFXOuTxbr0CDbk69GS7T
mwob27yKU07DNEkRZ3kkSOQAy+TYxsQGReXeNOilIX4PdcNBbFmoBSMkSXkR7QB2
X4zYLYWbPnlIHVGrXfYEYHTuQWDB6l/E0akIhJF/uhZvDImVS1rJBkDj9t16v5Jt
Ih88KlfJ4jIQKCZbRimcDcWxAKSTbUOLtGjX9blkyWN2nV7yzebqe2IJcr0cqUGn
xIKUrLN1EgjMWETFBrUgVzk6tE6eFl/IFeKvS5LzI4GRnDhSudw85od5+n2NsO+Y
R/LL7H7D7Tbqw19NmbbsIvJ3Ojlk/xnnVTabffyzJZpQAd+ILobcZFdn1qjJngQa
5FUk1QfFaX5Htt6TTWUJjy42whf9tVL10rN6GxIVVND1wpseKACc+WrNufdI5F/D
O25IinVU2EZinTuG4hqa74FBfIiRYiBwmuTJ7Nla25nDxD6ahAtOulP+lC0S9g8B
SbRmf4Un+fC0cgr2ezPL5UGkV3CN502a0Elwbz5XPEWEcRWDr8D7aPP+dk8fA8ib
oEzrYMsL5A68VHZkuMBT/El2d+bzqPfPgw5NOsCTtCRnFgR/+7K57fQy90OXM7wM
H/jtMS8oHhnVNDprnn2GDZWPqkYS+JxLfZz5Qz6mBqF0n+A9T2iBHPEmfVNlSdId
zZoeRM/qZjnIIcKhWzskC0ATjeEl+NSgjltUOewt5C0xYO0fXLxB46YzfCNv9gOu
zdqzqk2KBQforYyPB463WRtajLGY2p7Rlhxu/+PP4p2SB1Tes5welGtHebscopG1
fbIFzD8amKwKPK0J9YqD5qaHsAAuQW8Si9TNf5FT+jUIgPYcHBQO0T5EgGUzH4vh
DTHnCYt307usCX9q8ZnfAOsw7AHT/M/w8wqYBqJLzUdyr9rkTu8hGIiCMWN8u5C1
H67bx6NmI/PTYpSlK12e7nXyZ66bm0P3w38w2ujvb09P0lo9VRuLPp1dOjonJf0U
Woayh4y/lLxTQECCM3fepXTsTf4kSQFHrlsLGns91R9uR+hRJd+KqIJ2JX7r1V67
2MZsZB0t2Zl3vEdLTnowUljwPKDFpBOP1cJpOK2HUivJMyJx/SoMd7dpc6Ar5zjA
KG49kIJzIu3r/3IkiNg6cl5F2PAYh0PoFsy1DuIExLgNNIMJLEsFAm4R3BuiQUHw
8UzITNm/xXiRPEKBgqtqW3Wsq0lCRkId9QDoe/FbWLOeCSNudJyj16Vxxo3uKwK4
2SKRD0MNDtb82QW0kP6h7JY4tixynYfk1IcxBDMfnYNE30CLCmJf8cw/xB+OsjN+
yczurrKztZEqZZ3p/qmJEaPZpDKvUmz3szcrY/3gKc0ycdxn5mWRIq2nAUq0Y35l
a5oDv+Uf2Vg3o48LjoCb4b+6KhYuavZ7ffiZ5Dwiiy5pNDJqBCCeeezWPLsNJuR7
41YflAEmep2Meuo0s5oD7cOfbbmzqiS5nowzaOx7aMIOXpdjglyiYuzMtYoU3Ak3
qcO3LhWx3dhgIyZXrKWjfTovV3dXsB6LvDO21X8PHzbVGNi3dsD+TAAVu5BLAU5y
hh9WFchxKHGLm7NTSu2P59MypyMpx/QKfLWkKWPMWvLAHzCEACLApNcNXJxFV82/
9XHVnhF8CkZTIAtxsdzF8yZ3hpGghefuffsOKkJtFq9zDsV3WCeUGgd56Uh37ibr
D1izmm6tVSiuNwbKRu6HhoV+/C+jfqMw+uG7iKDNUCR3w2TQd/FaNe5RLT9c5PqC
/ftUEDv5wc96LCdcG6W6moSwJXhtncZ5lN/mkWS+ZEUqtzaEYVZITKvYpuVhy+o7
ULqwgIPcXcZKLo1As0H2V/HmTJFRVyKwkBpnX2mTsL3bYokEN97BtAm4rO8ihJrn
ZPvofaCutL/Up2SGD3BvrzhPuQjN6fsgEuRp4XIIh0J8d9KLdXhNyEPNIccmRJkX
aabXdLLerNW63PqzR+XUmmyqe3n6OiMTscH0+vEI14Bkc9WQzx3xMsyEL/yS69tj
FTr/GzNR7SNjasZU1loi4Wj8FrcX0PSUFetJpyoFq3T6cRJHFvwomAXvb0mqJ+VD
UuGOVl5HbQxYPHWKsby3VP8OJ96XHyK48o+nPc3eF8rg8cqfMAsdYQQ57D4Wwihh
T3GHaFVQyBVghhD3tvspAEJvGJxDI2ulZPXnGPAF79Ta8QxyG2yzOkkcBorH4XFt
I0CnqGlLZ6YETSzH9OPpIbVDZcaJp/6RvdF+3tegeTqmdvIZd/o64nJ6Ax5tvQvk
1u0+mhcvhJXgXAK7QebGIbevzDBtPh07Oc22XqvfLNMsLmTleMnpjsyL1so5EtH4
R//pM/WyzImRHs/kEK/DceNgY5zgoxOMXDpBt46uPvsBKHH731smM8xG+nUolaWl
XvEGlc6sps5nMA9WB6zwBBjrsfS6Tt3cVoLjyGqq+FnNSsxTRwABrgZmfL+03ZC1
f0NxVdY4U03G49JZT5lqZxzkFyLadM0rLnhqoBWzRQ4nx4BDCCdP5AqKzrUjL0S2
BXhBLmRZegGHhiLrj3fwFpCXOo6Udtn0DIXVGBGXjHkZLv2OuyLoT3II4G2OTWLs
PjuZTgLPBiEEyemOdyLHOffiqjC4ZFhAtOkoLLCFBaP14MK77f7C4/Wn3od/9UBb
Cy2Lw3r8IZvVJ50kCfZq0+tQ0d5jzTCN8gLYdzo3WuVrwHjzQjz4SKHjC0Qmc8Of
7Z+Mwz3v7r51TxMCEDp2oVS6WZKkisKcQen/UVPDpbhWF4cYJ6Px/4VCeMlL6CvY
bEe+2nwduEmYOFystxd9mED42VMu2088YGJrS7TcxtddIuV9KOLdgQqIUTJsHnwv
lnxTmceAaTurpJ/dYcWBAuKHvh1BPZYZvi3LHhFPrHnc6rSKQUYK7VXOZsWzyDSW
O5XsJNVAhbRTioUygqaJ/SgMIsM6UKtY/TfImORrMBV8o9ao8yEDwEYh+yvBxIM0
kl5TXOcqc/k4QaoUyFHdGXzsD0gghNrRdJP6kdLcXDKk9194d9ynEM2p91+VWgtF
TACXNjkc5dHirSr9tpz5SCw+B5/QDjSar2NsRoeteYRJHdQviFsDwXae1AX0PvZc
oXuja5MoAxSns/VZ9wTzi1R5ojfER6ELwbLIBnbZwn2KWtD9/Qr5C+GXIpVfMvr9
ssFkDW6Xw5zqQL3UyC/rHuhWbXyo58y6WORI1+pgukidTa6g3Q1tUq5D4IxBmAyL
NfF7u4UtMEwxyFgOO/fr2saODsBrQKibjcI71c6UhK2RrOU5f6RbiThxkuGfdlxG
cWZSS/UdVIsqUR3K6jZaTf0XnFz7JpFH9qq9ZNFIFWekPCi0qTxg/dD0HL1LGvOn
ZGU/fbbkXLN0QmHrY7DQnHS0Rc+Bs5mDxmCto/r0RRXJf/ieQMyx+cFCm4Q11h9j
JMgh6w+oeRvEoCjCL5yZKlGlm2VmoEPPbcujeyacDYKuo4w7AuFwPsAF4LBLPkJr
8oaFexhuOisogD098K6Z0wPTBRJkDsG7FSLQF881RpuSjGQoeRlvJvzBCQartzd+
cSF12FRx2VRzEtofwn1p7tDeEmHyb8iFbML/kw8nIu0YkI7S7CFaflCDbYQSZSoU
zuiOF3sNBsu+bHcG4CsyxhyChr5q2JAdn0q3S41g4H0gAIk33TY6IgL2PnpzvG+K
cxIv7PKGvOlqrBlH/8XMFPXJ8YIg15rcQDYCHzWS544F9wCdW1zEQpBspV4xKVif
WSpGIKln5FJmFE4x09agc3GYq54pqf0QiaJ3v0t/ubT42/GD7Z2vqu8thriT8SgD
pynLmNbbmV4cNZZEeFxTsvA8/d0nuPcPWwOFMB9Nl0uGjmQQL4pLluAnsNkcEOcb
R3co6sTJOuTuydyOF3H8fIjJEQy/EZqwlKCEQoRCmY6bxFOgjJ/986B+KQhEYVdk
wVx8nfHV4eS1tjDtPObusPRfTRIh9hzdlvToGbOkswHLkJK+gipYHQKy8hjjdpm6
2CYRu+50ddNzN+ZA85MzDPdUY/4xwnLFiQ1d6bfnRsK4JOFFAcmVM++Ici7K4DH4
+ybyV+WifBilxskh9MDAacji8IugnVSKalzNjKBnOBvxNHWLJPvqWqiTFdxKCxJb
ZVo1hzEgIqWCLztTX0n69kB6FIx7AnnO/eMqQkfQgR3nPCth1ScyuDWaNgNjTrdL
agc87wNQJxrJEz1dIkbZmzDi8QjxaKvMEjD7UyoWMWZvRw9O5m7ObrpTbGymMSJY
HJSDr0QgqT1V3K2uDkugEcKd718XMrBkMC5niAoTsB9o5mnpzJVTJsCYsAij/oqg
4Ols89ke1blwT3DAIgFH8nXSyLXvvC9t11ObB9FjgKbNyJ8D/RyOQFW4nOsIxzDn
pPp2aOv12ZCGmi800Sa3GX6rcXotvIxnRxiaBv8TKKUh4NOBJi9pZT9NrURu9SXm
KaDWOc9IILL6Srgx7nR6erK0lotvxERCZvAH09+unuRZTUpcRp/49ZwqjbTNcYyW
F2n4ULEl0N5/A9vIiN8I1gdvbQI1IrXOUHA0QZgWhgAzjsRvZgfmPzsBrUkHlW0x
NxAVDoEvkYLVTWsVR6jyExkV5aaURMts4Y0ifRzXEm6QSxZQ5mf8wttLB4VqM5yC
bROKg3g7xf4ttKahbr/3PQ+x6W+2QJWf95yHPlsmdX/r38OKYvsFtCSpsC67mtGs
Xxy2QwL5CiHIw4TihLP0UGBZHpPzC3FoMoueeX7Pev1am1UYSfuX297uYkz+nwGD
9Nw2h7mJrP5QgrNluO3M4PyNPW/SX8nFmPQ8nmbUb0YmWlXewz26WDP4VB4Gby21
o00p/SOpu7OzuAlp5VhVzXkKR/fwanQacUOloJxMeMPx2ZEcoEtMkA3b2A2iMA+4
JvUw48+n8xUzcbCR9BsvzrsAUyWd/sSKJ2CpdUsmMycD/AxYInbtvNOOUfuwNQOZ
XvStTYfGSe+flyYjcxDuVi1yy+YQxLgjvfvNOuTKYS3ANngZKk+fvVGTVuQSpBm7
vKOFm4fhYBCb/n/76LIwrorG5q4Vk0RAHLGTP2FwWXq0m2bspIfl9Fy97RWqn4Us
LYuh/5IdWjJ8lQ5O1EXegavTD5NA2O4Z7nBoF7+ZZZ8d4p9vUtYxptqBMs7+Tfd7
EU93G1nziTb9B3p2/0tOR4tJt1jyQ1HQSRIfXSLJHCWICotX00cDZgOC7NYwZ3Cj
OcepEvG7lEs10shOUo1rthfYJ7nwfp0ub8Se0DnCVBChTCNfg98NhwNVYzxohaQA
jssHwi2bUX0D9PTV3t1J9Btx0GFc3inS5BWDWhXlZGzOEA3DuzagDsdl0Nl+vagD
8ma7/Lw8btjh3DnINCgaS9PdpZ5dikGkw+RjqLAUAax95xLPXmXSnXVnY2r9w1hg
hRjx0ICFtTNudvWyVZ9OhWF85QcWIU0UcvrmXljHNyL5kzUzTRXRWP6115NtU4lj
B8AWZnfjY9RATafYUigEXWkirUVOP0uXnv9+Xf8bFoXgQPXN/qzPVID05AUIXc4X
Dy/2cvfgl4DiHbGg2/8RkmSpTFNU0AeLhxPZ6caQywznB3EVc9q6xskUpf1R78w8
Pdaa8PzRxG9FDjFANdKKPw0Mc73viR3jura6+DJvLJr8mhzdDVibvK/pwItDu4Ke
ekIhbVQ2xhsU7mIhQSO5q6/2OBaeazLxParkh9I2CgV1yyD4whdio7l7zXOXftuI
5zTeTx7pJvVBaTXeXM+g1A4JSjFj/AKu5Jvx8u9OibMy0XdkW93v1IXP2UF2dlAw
dKxHChQYkPKZhsrWzkuZO3UYxrcJRXNq3BIqM6Ti62gi5NzhQ12T5RtpxjrIqcC7
Z4XU+7WVVRRsmHeirZ9dsXW5hux7vXLdNw2zeQ4Q86Yz2+HHkaT9h1uwMKzGpG3g
ByxQjXw9f5wHJdh9NmwBAGwKbZbmvobx5uQhblrQeuiXKykPEg9gRHw0SkOxnikk
oE1fk5XQRL2zerPF2XXD+HVuphU4uakTRtVLb6/j50hsl1JUtoeda/8oY2DEB58E
IK+6YCG/CZBUq0GX21n+guj4no5V9T4wcg1wPSIMEBrDsfz2Y3WD0EyAH711TTJ4
FaTAWqiMlhHQe1rYJYuyNNZSY2t0qcDzB21qF6PvNO4EA5gkA235mLlPVptMIR5u
sKlN+cncFk9FlVwvP1p/M91hN+s7fAcnKP7xTh1JLqECGAPs2Skm7bp2rfkglRmo
RUCn9FfuMjgoX/VPChpQTgvPScCG+QzUamBNrrpCiue17wCWyDO8y39VAzSV4RPA
Hv3YkA5qbM8XalpDv0ioLPW/DuiNfNjfvAL5or4TM4ILW4BGvaYhn4Sqn0lHIzBo
wk13HhyUvyRTh+Y8FFAyPI8Co8e8mr/Pg9KgE1aSSRKorRispB6gknjnn/gkawTN
HdE1bfAuMwWLMnhi8YsyfvvU5IqFErQlGLv+qEsT54h1P+NIB43tCjHlXELoQYEc
Piy4j9F3A9JMXLix7GL7XHTuMLp4Qd63vYNbGvihC5wa4s4rvEBs2tg3Q25Cw+ge
gj8HLZ0d5FnJQDTHWyZpgLYSuT7S/8VCKeqL0piPe4mx+YN4/hoxarCGFfYn9gx7
vbkCEiEgyq6piN4uKM9/MPJHfVT5KwsQ71q4qp6+8lYU87OFsTcd6z0hQBLgD/su
XM2dg+sFZCbeXE+f6kT/lEb5hFFtNkONvO9IZCHkm6toPwXUf8jpWzPkJ8D1X0ko
ruGJ78zoTxD0+u+mnH+40Jbp0mm36x3kQoiMHWhTgKbiqKykbRmQmanASCLcOur2
wsC3Fvn4p0WlC0xZpmD+a2GpUSdRgLTjHIC1cpvfQrSje5+TxQvwzQC6WRdMMV0X
gtKo7SJ+hVMlxWtHalEU6bbBNFTbZ14DHr7+X7ks3glXFslWvhjABUpjiuGbqTW7
Q5wq04VJiezn3/L+vVDHKRS25BOxJYg05iYNJAM51DGDXITMxmTsvavFE2hqthh8
evUgmt0bqkisjkDMQGjzOwzDlQsFF8ijYKbnhsF3LsQwqfwmoS6PkqG2LhAEZYT7
EU0q1JGx0ak+tFAxFUJSfBbVpAz4JLkW7rp4rcRliE24beRlhaJWJ6o2fDq5fA0K
3mynx1C4Z5AIFAjAXzFMGSSEam2ZJbYTCr39KfUBxY+hpa47gWf7rbg9BqJMLC9A
Xlf+gOz868TkZoHZccWPZ6CiwLqmByC24gNFyft0SFICdtT4yuubWW9sGiWu3Wfy
dsE9JOMPm98l3DprzjgwGwpsuS2iItwgMSto7NxlBSVa1/VfoT44Z5abmJVcNPse
jfdpG0EcvbjFVDNgXmywd74DbsDEUM2q0v54vBiiQM20qzu5W4rzE1JOiEWKq3qE
2ESM3S34frykOGX0uiYhPVFS/iGMbRMCfrLB16Q5ZoKIu8D+5dmzieUx0m4KCpta
v9f34TqtK6f7L/Y4vfFqlCHB1sV++FyPJYiPrrSFHmaabPSF3nxj1Zbht3R9Edh0
iIUIOcEK6fj+RHCguY8F+7A6Lrpcpz2l8bxyHEePsII6eU/79ssLU9oc8iOoKJDV
FZZ3zJaBskzDGiIdKHO8Z7AJbKB5SyQHWhqWfA5dBhhaqSGpRxEXwUpFaByN/axD
JIjzgJ5hV5Ra1qOVeSVyvokcNOsKUI9lTm9YL5L2+10OvCXasArGT7xGK6f9hhog
BFyxVfh50V8goQRrGPLF7+8lYCi4sgDdJJlaa4FDyiNkpNm4gkBwjJUxcmtBfP0g
o/jzjTRh6TzISfZTn5OzGZLwT/SyeGIX9BOceps605eT+iWPPY7J9Rtc5iOPhIBG
8VfsJIyPXW9zIblkAmJTH2gdJgEmjnaAG874sQTlfvqytHT2TYqHMQsxFJ7pls5e
C9aCRILhtR+sSIz9Ndqo3jsEY4Ql5W1UV1a4q6nHVULOfiL6Tme/saQUOMuoCHyK
UCLKgdHl5GgIq/9rOlr4KOLFIstRNDi0D7PJl9ZyAot6Rkpe5tzPwY/m2Vu8JgDZ
h6iWibDkUB/sMKe+qIkqSiyuBthlPUgjpyzWs1TKX4qY6kt1Ty7xhhzlqP3SRXS2
w+nZvOoSZxk1l/XuGbnN/mc1qF4UAE4ZvTyKXoskVNYtWTj6PWmuuMg78ybCVgrp
SVOeY+0JiDeIqzm7E1WamaBVfupRTpuE61IbmawTsQbkkdjkpt0U1Ob0ftD4caBr
lE/Wdl/8Vku2U3GrZh+cdTmyiVS1EK2WnQvlzxcK4H/84mDHcTnwdkdpQy4+IiPj
OgPgP4Zlf4aT/0fPpQNmPSvPEjGC9bjCdEqFzI8JsYpV7fVGs4EWUSO2muCtF3EI
mDr65C979l0EFO9/Ftplz9E2vV5QRmFnx9LNf5mHxElPrKih0e9Upqr1E1SUxKTi
/v61IvrURgO2VVacRIvWRpfRcCOCjkP6bgCGU1/hXDx9hreeQg7lOcLN72k8MeFz
oJ/CLUn1yHnGl4BkpJAVQzcBnacYxUds46fxfd0Cw9E/VKl/7Oyx2Ml0azBNIIqQ
nQci1V65thFLPBYITNxYULVhXJMFxsUoe1Dkor5BSEiXpcc5ag5PGh2y0083OxD3
YGA+UjbIMKVRULDxjMCJN+BYrglU1VpRlzLRFP/UZff2cpjkBH7TljFPqdZXaehS
OQkPtz5ZrQy96rEO72cna7+9QKzNDCa4IG1PIOs+1KenD66F1eDoIWyy4Zwx3PS6
jnK33wYVqXSoccYd98XvCQ+BgNlmM5ge0aoRHiDCBelKe9J2JbeRPwDcsAPSqVXY
m+r8kapK/THH133Tip48JY3LtIMwgmHFjSu00tuy4SNsT89EWkOoYhlc+pBueC9w
sBoNkzDN4Dwiqw7Y67fpnRl1uTg5cRK3bJ3LfZ3Nfx8voTMFOUoBubEJYBrYxqx3
v43tofPVQJI10ptjZzBwMo7PxvURERnnK+Z1NSKLKiAHjIiXLGPu6Ztr8OpBuNW7
RMTd9kKZJnSA0mzsjuAa2FGpz44TBU69p/WixN0BjXLkbUiaRFrXciFa+yjmlwqJ
WnFbs4iJcgU5Hqwx9SKfLLwwReeDoxJICUVPR9gz01TXwkVNJKi712uki2/5Ynmo
VAIPeDN0huMMyuGDRa5gVrYjTsiu0BdeQ4yvCfTf7fe++mrjUpH4zE54cgZz2DmG
tt8FPM2cBuIr04sB8iki56fyW+7b5kI00E8NxMIO4TY/PjPALQbesObsbJJ9Gz3U
StMT7Fka+J/3rbSHp4aS0doUyA15zTi9sSumF5MXpkuClxquYBdvDO6xZ5SdVoq3
Flv/bJs7DwFIiJoX4uwrKV7XTao9e6nk7ugYL9n4KMP5MVBJuteKP4dLDbajYQuy
ExR8EBfQcGcSwFgd+cgv1+xxjoZIlcH3CjiBap/P7bbaTULT3M62PpDpGlvqaEA2
pRnXEmj+iOjLD2jiCHVIh5zq/sorru5dJtLUAOoYAXOp4XfI4N9V3mHvzdQ7LXd6
vAALWmN22SKPmuKg8Ck5bNDxpUOk3QyMv0oqoVipivBIN0VuwUYsQUu8jogT2nYj
reC7hAawXpyChMMlyDcl18w3vxeQSWImUdR4pKN3ux+wP7jKXZAUJIUQQb7ghS8x
LeoyhXOB8+XpVtoem1b5A7SI6FUKZ6MOaTLnlmKlkd+qm0mBN8YOJ8aYZryJd2Bv
ZFLDeFjtSUCFTmSv69YciL7+U6ON3bDMM7vJhSvbFE4azrMSIC3oy28RLT1EM31u
kiMebNU1ewojaLVaqQAJSZQDTwlEaPbYFZ7t5WsHid9pe6e6T7HXQkEEKPnkGJP4
+AHMtqdXeYHGqY58uGMTpogUJclylKMCA4Z6vInACOwtHn2Zo7/gMwx12N0SfEVx
m8y+74TvsjK1kgNSeOZCsQgOpB3tpnNcvZbOIqX8HI6X/4NzZLvEhvD5Pt0qmQdJ
vdsepmSixKQ22yvBl3Hs49dOJqR5ZdxD0IQ2NOd4V7vx/FHxUNDGlQPG6euk95LU
IGPeo2Pn3rW2b5N3Ri0gi4tk1bAmyrtJIOkNKjSVHQxW7Eo71Ui4YAc4aUEyxU/6
ypIfb65dfxvqwB68hOjeS82RTOIhUTQ3+1QjKjXSJ8QTEZhXYsx92X1lm1+wFLPy
b7n/Ql8WXR/PINQZa340EH3zQlHuFnQHJUffrcIXn4v537J0Q7+JasBd91QcLsLm
DuBL7dgga1bkpHCq/ANIiTE1O5QV5uA69NLjLML7mRqU4k2C71VX2XRgnW/yjMFW
GtELbLajKJsM0Du5rV1z7Ts7zWeg4v/kzxGPLVhVgAEhO3gMcyHcdJ+0kswTEEiN
n3vzyjsql0sntdmjt3rrm8lR4SEkJiJkhkZTAoUv1b9Hee6z2n+kZ3S4fIwXP0VP
u84ea9vdW/o8psqm9pn1GkSDJakWRqOMGyKVvxVjt3wpEk5OQTpNSWCcO/c8lw0O
mzigl+O2EtMY3RO2Kn9Maq9VTzd3zmPGeuPVAUB+2w9YY1Dq/y/SgDLzzwglZW21
EpMoVRJoBEJF0wyi2rHwdR9ChvjPzQ/H3giLW3Dc/+MxkVaovfbGSX6nIc+AqWpS
2gBkpPexumaCtOeqWrkW8PIgVQBmjc5abjJhWjFtERG/mqXaaX2Yy/DnmkUlO4s6
rw34NqlYJSoQyyi8gj2IWs+8lO2cPfYr1ofycVEeqx3E/PwoemjwG4XXMCbd/C8C
rC9YQ2RD4cnXSNPJ/j2+3egF92Sf5FWt8IK47MCS60AyfF0XlaQWLxMrdJWvHuCy
UwTUWE+AmWp722+ZlMCMX7GE5MAgu8r+WFCboGrn8bbkeqAoFghIdOrBx5mPTLh/
RQkge8Fly+AcPNkLB7JtixfuBX77Oe26s1TCGBoIzqU/SSkFiD0jrxXtDwhxSkk+
IuSQzk5tvKPqYY2WOU7IpTQapF24/mcgYez1LZbIPPFyI/i2kRP/HrSCBfJxsiBJ
i/HoxoPM6A+2WrIf0rNGEjiFiUV1a2CP7RkxrVJPlYBhbCscmQ5efxmA/14XuBv3
I5lqaEp0nCXQJaokFeqgX679XaZJdr7mg8tPqFRzLHdOtucb1k8CQkk+1Y+U+bJ7
RrcNCThHNiCwOI4I81r9kHLn+QzIgokV8hAhrqZlIh0VMxe19zSN2Eadju6U58oy
OiWq9a7w4AxidNB3GY5l31uaReH/RnriTUvr5njs+6cDUkx+hmkOSm6Hyvn4VaKN
TLVuhwm/OmePGvVVINdVFh79a0og9kad4ASBcdnTmYp+Hulv44Rat0TPCG6sAhVB
Q4IM6gIT1oyl0thooC7PC19UwL3MwZPJjvKAYtdOyMG3GMXu9SO9RVf29hajgdFq
3aQk7j90CELC/gUl15g6dXiwty8O53lL6SIKH7QL5N/5HWiCaYOf+/sSxcnVjOF/
7900Dsu2BxIRRzM0qgNnyNnpdEpQG1cbX63gpUfe8EqPFJsEFtAUAyk3ql4/q/As
a2OXGhYBc8Y3GiE26VZyF1aN5fGIXrtSxJxi7yDAnzYu8EM9mdVTxpscyEWxS5LI
IOi1TXlKAI4vWDJywRsh+HkhhDgMxldepLvA8R7UGWBMW8lVHQhQ8saHjSCSsxtC
Uyu5oc540dENDIvv1O2p8igOQ39OSAvP4hTCAHbj6sDFAtbMCEU4o+67usM5GN0A
DUFTP+cfbRUZY99j+8oK66VRpp/JnLwZBvLWX9ZWWUfx7y5XiLvDhDoHE9qnORKA
OqgeCjw3BSy9/0ljF+jq1PmXa4KBjfGmJBbIaa01f0wLyF49g+j/9wm8GYOtiptd
NstdvxWaxBJEFBECmt99WqXVoPPSYDxOQtbvtH+exhjKmtLAZI5mQ4EUE0CC+ha5
dUKvepr7CkHXdU/VwMcqOcflGQGQSw4s6cgKbJGqa5DN5ERoM/DDo92CdfpwT1Hl
0cmZAkaNOlMoBrgUFhfSrq/HocSIs9IerXCQiIW721LTgIcvw/jYO3u24+T9HAMQ
qEtfqtfajzo17KzyNfyKZMNFWW6KjVcxLKtpJs1STdkS4+HaVrfrXgtJLnN5O2lt
KPR5D/oPmaF8n7K8NGDEQ1dv/HlIgSs3POQyOw+iSQTsWzqYYr7pIqOKQ300xk39
FlFKA9JLEpvm9pW2Vd9r8AL9dn+rrTkaXt/JaSOgBctup+NM/lHcRk8Qy8B1x3ii
wNdQtAE2tctAtB0H3khUj8ASrCKT3USlFq+bwvAey8ObsRaGLSwaiTkc7JDdXwX9
tc0ufOrERdxcQrtsxA/xAZAns3LSBVcDFXcL6OAa+L1LfJNTsHPUSURDXJ2yaL65
9SIppzFIN/PW1Tz8gD1HXiFZGiFSUCrTxJT5EVqKIahvYVFXnS7DgjuBmlQxf3B3
SiDBG5L3mQT4a0plyl+lRYKRHuJS3dTt8Lmvyb5FA6joqyM/Hg9lGSM81MtAHH5a
s9CgDkSjZ1+LuiMHY3Lys7+N1WVDij+u2rjhpRUE5dbYOCjv+wNrDgfVPGb9Q9lU
SgDme6UV8P/dSov5C1+RV7t6LeEL4N9MJRQ4tPc9nTdoQz3tQeAtSMnTYQABjtpU
4Op+gis1WldQPYaZRAXu2WPZs8M+CfSB6+DzesGqjbVHlCVF5ljvq4qJmNNQZezQ
VFLp5ihOzi++bpikkxZN/mJ9Fg920JTYReDJwWgl15NYoU38DU9Ye0wrWuFWUUC9
UzhPQJz4vToSNje0L7sjq9uQf38Wa+1rdiZ/VVu0LhdvLV12VyDUbwXXomacC/7n
y6v6jtsYVSYjilnmJA+s+ctXHRbYmkMl/U51H3o4kHNpLen+jk65BKD4Reif+ght
`pragma protect end_protected

-- WRPC LM32 RAM initialization: --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.memory_loader_pkg.all;
use work.genram_pkg.all;

package wrc_bin_pkg is
  constant c_wrc_bin_init : t_ram_fast_load ( 0 to 32767 ) := (
        0 => x"98000000",     1 => x"d0000000",     2 => x"d0200000",
        3 => x"78010000",     4 => x"38210000",     5 => x"d0e10000",
        6 => x"f800003a",     7 => x"34000000",     8 => x"00000000",
        9 => x"00000000",    10 => x"00000000",    11 => x"00000000",
       12 => x"00000000",    13 => x"00000000",    14 => x"00000000",
       15 => x"00000000",    16 => x"00000000",    17 => x"00000000",
       18 => x"00000000",    19 => x"00000000",    20 => x"00000000",
       21 => x"00000000",    22 => x"00000000",    23 => x"00000000",
       24 => x"00000000",    25 => x"00000000",    26 => x"00000000",
       27 => x"00000000",    28 => x"00000000",    29 => x"00000000",
       30 => x"00000000",    31 => x"00000000",    32 => x"00000000",
       33 => x"00000000",    34 => x"00000000",    35 => x"00000000",
       36 => x"00000000",    37 => x"00000000",    38 => x"00000000",
       39 => x"00000000",    40 => x"00000000",    41 => x"00000000",
       42 => x"00000000",    43 => x"00000000",    44 => x"00000000",
       45 => x"00000000",    46 => x"00000000",    47 => x"00000000",
       48 => x"5b9d0000",    49 => x"f800001e",    50 => x"34010002",
       51 => x"f8003e61",    52 => x"e000002e",    53 => x"34000000",
       54 => x"34000000",    55 => x"34000000",    56 => x"00000000",
       57 => x"00000000",    58 => x"00000000",    59 => x"00000000",
       60 => x"00000000",    61 => x"00000000",    62 => x"00000000",
       63 => x"00000000",    64 => x"98000000",    65 => x"781c0001",
       66 => x"3b9cfffc",    67 => x"78010001",    68 => x"38214e68",
       69 => x"34020000",    70 => x"78030001",    71 => x"38636dd8",
       72 => x"c8611800",    73 => x"f8004487",    74 => x"34010000",
       75 => x"34020000",    76 => x"34030000",    77 => x"f800004d",
       78 => x"e0000000",    79 => x"379cffc4",    80 => x"5b810004",
       81 => x"5b820008",    82 => x"5b83000c",    83 => x"5b840010",
       84 => x"5b850014",    85 => x"5b860018",    86 => x"5b87001c",
       87 => x"5b880020",    88 => x"5b890024",    89 => x"5b8a0028",
       90 => x"5b9e0034",    91 => x"5b9f0038",    92 => x"2b81003c",
       93 => x"5b810030",    94 => x"bb800800",    95 => x"3421003c",
       96 => x"5b81002c",    97 => x"c3a00000",    98 => x"2b810004",
       99 => x"2b820008",   100 => x"2b83000c",   101 => x"2b840010",
      102 => x"2b850014",   103 => x"2b860018",   104 => x"2b87001c",
      105 => x"2b880020",   106 => x"2b890024",   107 => x"2b8a0028",
      108 => x"2b9d0030",   109 => x"2b9e0034",   110 => x"2b9f0038",
      111 => x"2b9c002c",   112 => x"34000000",   113 => x"c3c00000",
      114 => x"90001000",   115 => x"3401fffe",   116 => x"a0410800",
      117 => x"d0010000",   118 => x"90201000",   119 => x"3401fffe",
      120 => x"a0410800",   121 => x"d0210000",   122 => x"c3a00000",
      123 => x"90001000",   124 => x"3401fffe",   125 => x"a0410800",
      126 => x"d0010000",   127 => x"90201000",   128 => x"38420001",
      129 => x"d0220000",   130 => x"38210001",   131 => x"d0010000",
      132 => x"c3a00000",   133 => x"379cffe0",   134 => x"5b9d0004",
      135 => x"5b83000c",   136 => x"78030001",   137 => x"5b820008",
      138 => x"5b840010",   139 => x"5b850014",   140 => x"5b860018",
      141 => x"5b87001c",   142 => x"5b880020",   143 => x"38634e68",
      144 => x"28630000",   145 => x"5c600006",   146 => x"20210020",
      147 => x"44230004",   148 => x"b8400800",   149 => x"3782000c",
      150 => x"f8002ab9",   151 => x"2b9d0004",   152 => x"379c0020",
      153 => x"c3a00000",   154 => x"379cffbc",   155 => x"5b8b003c",
      156 => x"5b8c0038",   157 => x"5b8d0034",   158 => x"5b8e0030",
      159 => x"5b8f002c",   160 => x"5b900028",   161 => x"5b910024",
      162 => x"5b920020",   163 => x"5b93001c",   164 => x"5b940018",
      165 => x"5b950014",   166 => x"5b960010",   167 => x"5b97000c",
      168 => x"5b980008",   169 => x"5b9d0004",   170 => x"f80041c7",
      171 => x"78030001",   172 => x"38633cd8",   173 => x"78010001",
      174 => x"28620000",   175 => x"38214e68",   176 => x"58200000",
      177 => x"78010001",   178 => x"3821f800",   179 => x"58220000",
      180 => x"f800317c",   181 => x"f8003932",   182 => x"f8003928",
      183 => x"78010001",   184 => x"38211814",   185 => x"f8002ab8",
      186 => x"34010001",   187 => x"f80030d6",   188 => x"f800370f",
      189 => x"78010001",   190 => x"38216d18",   191 => x"58200000",
      192 => x"f8003635",   193 => x"f80032bb",   194 => x"34010000",
      195 => x"f8002dfa",   196 => x"34010000",   197 => x"34020050",
      198 => x"f8003382",   199 => x"37820040",   200 => x"34010000",
      201 => x"f80035c6",   202 => x"3402ffff",   203 => x"5c220010",
      204 => x"78010001",   205 => x"38211830",   206 => x"f8002aa3",
      207 => x"34010022",   208 => x"33810040",   209 => x"34010033",
      210 => x"33810041",   211 => x"34010044",   212 => x"33810042",
      213 => x"34010055",   214 => x"33810043",   215 => x"34010066",
      216 => x"33810044",   217 => x"34010077",   218 => x"33810045",
      219 => x"43830041",   220 => x"43840042",   221 => x"43850043",
      222 => x"43860044",   223 => x"43870045",   224 => x"43820040",
      225 => x"78010001",   226 => x"38211854",   227 => x"f8002a8e",
      228 => x"378b0040",   229 => x"b9600800",   230 => x"f8002c5a",
      231 => x"b9600800",   232 => x"f80032a2",   233 => x"34020001",
      234 => x"34010001",   235 => x"f8002ba7",   236 => x"f8002e70",
      237 => x"f8002ff6",   238 => x"f8000550",   239 => x"78020001",
      240 => x"384243f0",   241 => x"34010002",   242 => x"f8003259",
      243 => x"f8003e65",   244 => x"f80028ea",   245 => x"f80027fe",
      246 => x"f80025d5",   247 => x"f8001fa8",   248 => x"34010003",
      249 => x"f800059b",   250 => x"f8000556",   251 => x"780f0001",
      252 => x"78130001",   253 => x"780b0001",   254 => x"78110001",
      255 => x"78100001",   256 => x"780c0001",   257 => x"780e0001",
      258 => x"780d0001",   259 => x"f800207f",   260 => x"39ef43f4",
      261 => x"34180004",   262 => x"3a731894",   263 => x"396b6db8",
      264 => x"34120002",   265 => x"3a311888",   266 => x"34160001",
      267 => x"34150003",   268 => x"3a105d6c",   269 => x"398c4e68",
      270 => x"3417001b",   271 => x"39ce43e4",   272 => x"39ad6dac",
      273 => x"34010000",   274 => x"f8002bb2",   275 => x"29e40000",
      276 => x"7c230000",   277 => x"b820a000",   278 => x"64810000",
      279 => x"a0610800",   280 => x"44200008",   281 => x"34010000",
      282 => x"ba201000",   283 => x"fbffff6a",   284 => x"29610000",
      285 => x"34030001",   286 => x"58320004",   287 => x"e000000d",
      288 => x"66820000",   289 => x"7c840000",   290 => x"a0441000",
      291 => x"fc621800",   292 => x"cb031800",   293 => x"44410007",
      294 => x"34010000",   295 => x"ba601000",   296 => x"fbffff5d",
      297 => x"29610000",   298 => x"34030002",   299 => x"58320008",
      300 => x"59f40000",   301 => x"44720009",   302 => x"44750004",
      303 => x"5c76000f",   304 => x"5a000000",   305 => x"e000000d",
      306 => x"f8002738",   307 => x"f80028c5",   308 => x"f80027d8",
      309 => x"e0000009",   310 => x"f8000516",   311 => x"5c350007",
      312 => x"34010002",   313 => x"34020000",   314 => x"34030001",
      315 => x"f8003e28",   316 => x"34010000",   317 => x"f8003048",
      318 => x"29810000",   319 => x"5c360009",   320 => x"f8000066",
      321 => x"f80038cc",   322 => x"44370003",   323 => x"29c10000",
      324 => x"5c200005",   325 => x"f8001f5a",   326 => x"59800000",
      327 => x"e0000002",   328 => x"f8001f61",   329 => x"29a10000",
      330 => x"44200002",   331 => x"f8000213",   332 => x"f80005c3",
      333 => x"f8004027",   334 => x"f800410a",   335 => x"e3ffffc2",
      336 => x"78010001",   337 => x"382143f8",   338 => x"28220000",
      339 => x"78010001",   340 => x"382148a4",   341 => x"e0000004",
      342 => x"28440000",   343 => x"44640004",   344 => x"3421000c",
      345 => x"28230000",   346 => x"5c60fffc",   347 => x"28210004",
      348 => x"c3a00000",   349 => x"379cfff4",   350 => x"5b9d0004",
      351 => x"5b810008",   352 => x"5b82000c",   353 => x"b8401800",
      354 => x"5c20000b",   355 => x"78020001",   356 => x"38423cdc",
      357 => x"28410000",   358 => x"54610007",   359 => x"78010001",
      360 => x"78020001",   361 => x"384218a0",   362 => x"38214e7c",
      363 => x"f80029f8",   364 => x"e000000d",   365 => x"78030001",
      366 => x"38633ce0",   367 => x"28620000",   368 => x"37810008",
      369 => x"f80007f7",   370 => x"2b83000c",   371 => x"b8202000",
      372 => x"78020001",   373 => x"78010001",   374 => x"38214e7c",
      375 => x"384218a4",   376 => x"f80029eb",   377 => x"78010001",
      378 => x"38214e7c",   379 => x"2b9d0004",   380 => x"379c000c",
      381 => x"c3a00000",   382 => x"379cfff4",   383 => x"5b8b000c",
      384 => x"5b8c0008",   385 => x"5b9d0004",   386 => x"780b0001",
      387 => x"396b43f8",   388 => x"29610000",   389 => x"78020001",
      390 => x"384218ac",   391 => x"282c0014",   392 => x"34010004",
      393 => x"f80024ce",   394 => x"fbffffc6",   395 => x"78020001",
      396 => x"b8201800",   397 => x"384218bc",   398 => x"34010007",
      399 => x"f80024c8",   400 => x"29810010",   401 => x"44200005",
      402 => x"29610000",   403 => x"28220000",   404 => x"34010009",
      405 => x"44410007",   406 => x"78020001",   407 => x"34010001",
      408 => x"384218c0",   409 => x"f80024be",   410 => x"34010000",
      411 => x"e0000006",   412 => x"78020001",   413 => x"34010004",
      414 => x"384218d8",   415 => x"f80024b8",   416 => x"34010001",
      417 => x"2b9d0004",   418 => x"2b8b000c",   419 => x"2b8c0008",
      420 => x"379c000c",   421 => x"c3a00000",   422 => x"379cff08",
      423 => x"5b8b0018",   424 => x"5b8c0014",   425 => x"5b8d0010",
      426 => x"5b8e000c",   427 => x"5b8f0008",   428 => x"5b9d0004",
      429 => x"78010001",   430 => x"382143f8",   431 => x"28210000",
      432 => x"780c0001",   433 => x"398c4e98",   434 => x"282b0014",
      435 => x"29810000",   436 => x"5c200008",   437 => x"f8002fee",
      438 => x"78020001",   439 => x"384243e4",   440 => x"28420000",
      441 => x"a4401000",   442 => x"b4410800",   443 => x"59810000",
      444 => x"f8002fe7",   445 => x"78030001",   446 => x"78020001",
      447 => x"386343e4",   448 => x"38424e98",   449 => x"28630000",
      450 => x"28420000",   451 => x"b4621000",   452 => x"c8220800",
      453 => x"4c200006",   454 => x"78010001",   455 => x"38214e94",
      456 => x"28210000",   457 => x"296200b8",   458 => x"4422018c",
      459 => x"f8002fd8",   460 => x"78020001",   461 => x"38424e98",
      462 => x"58410000",   463 => x"296200b8",   464 => x"78010001",
      465 => x"38214e94",   466 => x"58220000",   467 => x"f80024ca",
      468 => x"78040001",   469 => x"34010001",   470 => x"34020001",
      471 => x"34030004",   472 => x"388418f4",   473 => x"f800249d",
      474 => x"78040001",   475 => x"38841914",   476 => x"34030087",
      477 => x"34010002",   478 => x"34020001",   479 => x"f8002497",
      480 => x"378100e4",   481 => x"378200f0",   482 => x"f8002f73",
      483 => x"78020001",   484 => x"34010004",   485 => x"38421920",
      486 => x"f8002471",   487 => x"2b8200e8",   488 => x"2b8100e4",
      489 => x"f80023e3",   490 => x"78020001",   491 => x"b8201800",
      492 => x"384218bc",   493 => x"34010007",   494 => x"f8002469",
      495 => x"34020000",   496 => x"3781001c",   497 => x"f800024a",
      498 => x"78040001",   499 => x"34010004",   500 => x"34020001",
      501 => x"34030004",   502 => x"38841940",   503 => x"f800247f",
      504 => x"78040001",   505 => x"78050001",   506 => x"34010006",
      507 => x"34020001",   508 => x"34030007",   509 => x"38841950",
      510 => x"38a51958",   511 => x"f8002477",   512 => x"2b810048",
      513 => x"44200005",   514 => x"78020001",   515 => x"34010002",
      516 => x"38421960",   517 => x"e0000004",   518 => x"78020001",
      519 => x"34010001",   520 => x"3842196c",   521 => x"f800244e",
      522 => x"2b810048",   523 => x"44200148",   524 => x"378100f8",
      525 => x"378200f4",   526 => x"f8002ec7",   527 => x"2b8300f4",
      528 => x"2b8400f8",   529 => x"78020001",   530 => x"34010087",
      531 => x"38421978",   532 => x"780c0001",   533 => x"f8002442",
      534 => x"398c43f8",   535 => x"29810000",   536 => x"282102c8",
      537 => x"28210010",   538 => x"282d0008",   539 => x"5da00038",
      540 => x"78020001",   541 => x"34010001",   542 => x"38421994",
      543 => x"f8002438",   544 => x"fbffff5e",   545 => x"442d0135",
      546 => x"78020001",   547 => x"34010087",   548 => x"3842199c",
      549 => x"f8002432",   550 => x"29810000",   551 => x"28210020",
      552 => x"28240010",   553 => x"28830004",   554 => x"4460000b",
      555 => x"78020001",   556 => x"384219bc",   557 => x"28840008",
      558 => x"4c030003",   559 => x"34010007",   560 => x"e0000003",
      561 => x"34010007",   562 => x"c8042000",   563 => x"f8002424",
      564 => x"e0000122",   565 => x"28830008",   566 => x"780b0001",
      567 => x"396b19c8",   568 => x"b9601000",   569 => x"34010007",
      570 => x"f800241d",   571 => x"78020001",   572 => x"34010087",
      573 => x"384219d0",   574 => x"f8002419",   575 => x"29810000",
      576 => x"b9601000",   577 => x"28210020",   578 => x"28230010",
      579 => x"34010007",   580 => x"2863001c",   581 => x"f8002412",
      582 => x"78020001",   583 => x"34010087",   584 => x"384219f0",
      585 => x"f800240e",   586 => x"29810000",   587 => x"b9601000",
      588 => x"28210020",   589 => x"28240004",   590 => x"34010007",
      591 => x"28830028",   592 => x"2884002c",   593 => x"f8002406",
      594 => x"e0000104",   595 => x"78010001",   596 => x"38214f24",
      597 => x"28210000",   598 => x"34020001",   599 => x"4841000e",
      600 => x"34020002",   601 => x"4c410004",   602 => x"34020003",
      603 => x"5c22000a",   604 => x"e0000005",   605 => x"78020001",
      606 => x"34010007",   607 => x"38421a10",   608 => x"e0000008",
      609 => x"78020001",   610 => x"34010007",   611 => x"38421a1c",
      612 => x"e0000004",   613 => x"78020001",   614 => x"34010001",
      615 => x"38421a28",   616 => x"f80023ef",   617 => x"2b810050",
      618 => x"44200005",   619 => x"78020001",   620 => x"34010002",
      621 => x"38421a38",   622 => x"e0000004",   623 => x"78020001",
      624 => x"34010001",   625 => x"38421a44",   626 => x"f80023e5",
      627 => x"2b81006c",   628 => x"44200007",   629 => x"2b810070",
      630 => x"44200005",   631 => x"78020001",   632 => x"34010002",
      633 => x"38421a50",   634 => x"e0000004",   635 => x"78020001",
      636 => x"34010001",   637 => x"38421a60",   638 => x"f80023d9",
      639 => x"78020001",   640 => x"34010007",   641 => x"38421a70",
      642 => x"f80023d5",   643 => x"378100ec",   644 => x"f80027d0",
      645 => x"78010001",   646 => x"38215d6c",   647 => x"28210000",
      648 => x"44200006",   649 => x"78020001",   650 => x"34010001",
      651 => x"38421a78",   652 => x"f80023cb",   653 => x"e0000009",
      654 => x"438300ec",   655 => x"438400ed",   656 => x"438500ee",
      657 => x"438600ef",   658 => x"78020001",   659 => x"34010002",
      660 => x"38421a88",   661 => x"f80023c2",   662 => x"fbfffee8",
      663 => x"442000bf",   664 => x"78020001",   665 => x"34010087",
      666 => x"38421a94",   667 => x"f80023bc",   668 => x"78020001",
      669 => x"34010007",   670 => x"38422e70",   671 => x"356300c0",
      672 => x"f80023b7",   673 => x"78020001",   674 => x"34010087",
      675 => x"38421ab0",   676 => x"f80023b3",   677 => x"296100bc",
      678 => x"44200005",   679 => x"78020001",   680 => x"34010002",
      681 => x"38421acc",   682 => x"e0000004",   683 => x"78020001",
      684 => x"34010001",   685 => x"38421ad0",   686 => x"f80023a9",
      687 => x"78020001",   688 => x"34010087",   689 => x"38421ad8",
      690 => x"f80023a5",   691 => x"34010000",   692 => x"f8003e8d",
      693 => x"b8206000",   694 => x"20210001",   695 => x"44200005",
      696 => x"78020001",   697 => x"34010002",   698 => x"38421af4",
      699 => x"f800239c",   700 => x"218c0002",   701 => x"45800005",
      702 => x"78020001",   703 => x"34010002",   704 => x"38421afc",
      705 => x"f8002396",   706 => x"78010001",   707 => x"38211b1c",
      708 => x"f80028ad",   709 => x"78020001",   710 => x"34010004",
      711 => x"38421b08",   712 => x"f800238f",   713 => x"78020001",
      714 => x"34010087",   715 => x"38421b20",   716 => x"f800238b",
      717 => x"296200a4",   718 => x"296100a0",   719 => x"780d0001",
      720 => x"39ad1b3c",   721 => x"fbfffe8c",   722 => x"b8201800",
      723 => x"b9a01000",   724 => x"34010007",   725 => x"f8002382",
      726 => x"78020001",   727 => x"34010087",   728 => x"38421b44",
      729 => x"f800237e",   730 => x"296200b4",   731 => x"296100b0",
      732 => x"780c0001",   733 => x"398c1b7c",   734 => x"fbfffe7f",
      735 => x"b8201800",   736 => x"b9a01000",   737 => x"34010007",
      738 => x"f8002375",   739 => x"78020001",   740 => x"34010087",
      741 => x"38421b60",   742 => x"f8002371",   743 => x"29630018",
      744 => x"2964001c",   745 => x"b9801000",   746 => x"34010007",
      747 => x"f800236c",   748 => x"78020001",   749 => x"34010087",
      750 => x"38421b94",   751 => x"f8002368",   752 => x"29640024",
      753 => x"29630020",   754 => x"b9801000",   755 => x"34010007",
      756 => x"f8002363",   757 => x"296e00b4",   758 => x"296100a4",
      759 => x"78020001",   760 => x"3dce0001",   761 => x"38421bb0",
      762 => x"c82e7000",   763 => x"780c0001",   764 => x"34010087",
      765 => x"398c1bcc",   766 => x"f8002359",   767 => x"b9c01800",
      768 => x"34010007",   769 => x"b9801000",   770 => x"f8002355",
      771 => x"29610018",   772 => x"296200a4",   773 => x"296f00a0",
      774 => x"1423001f",   775 => x"c8410800",   776 => x"f4221000",
      777 => x"c9e37800",   778 => x"c9e27800",   779 => x"2962001c",
      780 => x"296e0024",   781 => x"1443001f",   782 => x"c8221000",
      783 => x"f4410800",   784 => x"c9e37800",   785 => x"c9e17800",
      786 => x"29610020",   787 => x"1423001f",   788 => x"c8410800",
      789 => x"f4221000",   790 => x"c9e37800",   791 => x"15c3001f",
      792 => x"c82e7000",   793 => x"c9e27800",   794 => x"f5c10800",
      795 => x"c9e37800",   796 => x"78020001",   797 => x"c9e17800",
      798 => x"38421bd4",   799 => x"34010087",   800 => x"f8002337",
      801 => x"b9c01000",   802 => x"b9e00800",   803 => x"fbfffe3a",
      804 => x"b8201800",   805 => x"b9a01000",   806 => x"34010007",
      807 => x"f8002330",   808 => x"78020001",   809 => x"34010087",
      810 => x"38421bf0",   811 => x"f800232c",   812 => x"296300ec",
      813 => x"34010007",   814 => x"b9801000",   815 => x"f8002328",
      816 => x"78020001",   817 => x"34010087",   818 => x"38421c0c",
      819 => x"f8002324",   820 => x"296300a8",   821 => x"34010007",
      822 => x"b9801000",   823 => x"f8002320",   824 => x"78020001",
      825 => x"34010087",   826 => x"38421c28",   827 => x"f800231c",
      828 => x"296300e4",   829 => x"34010007",   830 => x"b9801000",
      831 => x"f8002318",   832 => x"78020001",   833 => x"34010087",
      834 => x"38421c44",   835 => x"f8002314",   836 => x"78030001",
      837 => x"38634e74",   838 => x"28630000",   839 => x"34010007",
      840 => x"b9801000",   841 => x"f800230e",   842 => x"78020001",
      843 => x"34010087",   844 => x"38421c60",   845 => x"f800230a",
      846 => x"296300b8",   847 => x"78020001",   848 => x"34010007",
      849 => x"38421c7c",   850 => x"f8002305",   851 => x"78010001",
      852 => x"38211c84",   853 => x"f800281c",   854 => x"2b9d0004",
      855 => x"2b8b0018",   856 => x"2b8c0014",   857 => x"2b8d0010",
      858 => x"2b8e000c",   859 => x"2b8f0008",   860 => x"379c00f8",
      861 => x"c3a00000",   862 => x"379cff18",   863 => x"5b8b000c",
      864 => x"5b8c0008",   865 => x"5b9d0004",   866 => x"78010001",
      867 => x"382143f8",   868 => x"28210000",   869 => x"780c0001",
      870 => x"398c4e78",   871 => x"282b0014",   872 => x"29810000",
      873 => x"5c200008",   874 => x"f8002e39",   875 => x"78020001",
      876 => x"384243e4",   877 => x"28420000",   878 => x"a4401000",
      879 => x"b4410800",   880 => x"59810000",   881 => x"78010001",
      882 => x"38216d04",   883 => x"28210000",   884 => x"296200b8",
      885 => x"5c220006",   886 => x"78010001",   887 => x"38214f24",
      888 => x"28220000",   889 => x"34010003",   890 => x"444100bb",
      891 => x"f8002e28",   892 => x"78030001",   893 => x"78020001",
      894 => x"386343e4",   895 => x"38424e78",   896 => x"28630000",
      897 => x"28420000",   898 => x"b4621000",   899 => x"c8220800",
      900 => x"4c200006",   901 => x"78010001",   902 => x"38214f24",
      903 => x"28220000",   904 => x"34010003",   905 => x"5c4100ac",
      906 => x"f8002e19",   907 => x"78020001",   908 => x"38424e78",
      909 => x"58410000",   910 => x"296200b8",   911 => x"78010001",
      912 => x"38216d04",   913 => x"58220000",   914 => x"378100d8",
      915 => x"378200e0",   916 => x"f8002dc1",   917 => x"34020000",
      918 => x"37810010",   919 => x"f80000a4",   920 => x"378100e8",
      921 => x"378200e4",   922 => x"f8002d3b",   923 => x"2b8300e4",
      924 => x"2b8400e8",   925 => x"2b82003c",   926 => x"78010001",
      927 => x"38211c88",   928 => x"f80027d1",   929 => x"2b820044",
      930 => x"78010001",   931 => x"38211c9c",   932 => x"7c420000",
      933 => x"f80027cc",   934 => x"fbfffdaa",   935 => x"b8201000",
      936 => x"78010001",   937 => x"38211ca8",   938 => x"f80027c7",
      939 => x"78010001",   940 => x"38214f24",   941 => x"28220000",
      942 => x"34010003",   943 => x"5c41000a",   944 => x"29620010",
      945 => x"78010001",   946 => x"38211cb0",   947 => x"20420001",
      948 => x"f80027bd",   949 => x"78010001",   950 => x"38211cb8",
      951 => x"356200c0",   952 => x"f80027b9",   953 => x"34010000",
      954 => x"f8003d87",   955 => x"b8201000",   956 => x"78010001",
      957 => x"38211cc4",   958 => x"f80027b3",   959 => x"2b8200dc",
      960 => x"2b8300e0",   961 => x"78010001",   962 => x"38211ccc",
      963 => x"f80027ae",   964 => x"78010001",   965 => x"38214f24",
      966 => x"28220000",   967 => x"34010003",   968 => x"5c41004b",
      969 => x"296200a4",   970 => x"296100a0",   971 => x"fbfffd92",
      972 => x"b8201000",   973 => x"78010001",   974 => x"38211cdc",
      975 => x"f80027a2",   976 => x"296200b4",   977 => x"296100b0",
      978 => x"fbfffd8b",   979 => x"b8201000",   980 => x"78010001",
      981 => x"38211ce4",   982 => x"f800279b",   983 => x"29620018",
      984 => x"2963001c",   985 => x"78010001",   986 => x"38211cec",
      987 => x"f8002796",   988 => x"29620020",   989 => x"29630024",
      990 => x"78010001",   991 => x"38211d00",   992 => x"f8002791",
      993 => x"296200b4",   994 => x"296300a4",   995 => x"78010001",
      996 => x"3c420001",   997 => x"38211d14",   998 => x"c8621000",
      999 => x"f800278a",  1000 => x"29620018",  1001 => x"296100a4",
     1002 => x"296300a0",  1003 => x"1444001f",  1004 => x"c8221000",
     1005 => x"f4410800",  1006 => x"c8641800",  1007 => x"c8611800",
     1008 => x"2961001c",  1009 => x"1424001f",  1010 => x"c8410800",
     1011 => x"f4221000",  1012 => x"c8641800",  1013 => x"c8621000",
     1014 => x"29630020",  1015 => x"1464001f",  1016 => x"c8231800",
     1017 => x"f4610800",  1018 => x"c8441000",  1019 => x"c8410800",
     1020 => x"29620024",  1021 => x"1444001f",  1022 => x"c8621000",
     1023 => x"f4431800",  1024 => x"c8240800",  1025 => x"c8230800",
     1026 => x"fbfffd5b",  1027 => x"b8201000",  1028 => x"78010001",
     1029 => x"38211d20",  1030 => x"f800276b",  1031 => x"296200ec",
     1032 => x"78010001",  1033 => x"38211d2c",  1034 => x"f8002767",
     1035 => x"296200a8",  1036 => x"78010001",  1037 => x"38211d34",
     1038 => x"f8002763",  1039 => x"296200b8",  1040 => x"78010001",
     1041 => x"38211d40",  1042 => x"f800275f",  1043 => x"3401ffff",
     1044 => x"f8003d38",  1045 => x"b8206000",  1046 => x"34010000",
     1047 => x"f8003d35",  1048 => x"b8205800",  1049 => x"34010001",
     1050 => x"f8003d32",  1051 => x"78050001",  1052 => x"b8202000",
     1053 => x"b8a00800",  1054 => x"b9601800",  1055 => x"b9801000",
     1056 => x"38211d4c",  1057 => x"780b0001",  1058 => x"f800274f",
     1059 => x"396b6d18",  1060 => x"34020002",  1061 => x"b9600800",
     1062 => x"f80034ab",  1063 => x"b8206000",  1064 => x"34020001",
     1065 => x"b9600800",  1066 => x"f80034a7",  1067 => x"2183ffff",
     1068 => x"08632710",  1069 => x"78010001",  1070 => x"15820010",
     1071 => x"14630010",  1072 => x"38211d60",  1073 => x"f8002740",
     1074 => x"78010001",  1075 => x"38211b1c",  1076 => x"f800273d",
     1077 => x"34010000",  1078 => x"2b9d0004",  1079 => x"2b8b000c",
     1080 => x"2b8c0008",  1081 => x"379c00e8",  1082 => x"c3a00000",
     1083 => x"379cfff4",  1084 => x"5b8b0008",  1085 => x"5b9d0004",
     1086 => x"b8205800",  1087 => x"f800020d",  1088 => x"34020003",
     1089 => x"5c220003",  1090 => x"34010002",  1091 => x"e0000002",
     1092 => x"34010001",  1093 => x"59610028",  1094 => x"3562004c",
     1095 => x"35610048",  1096 => x"f80028a4",  1097 => x"34010000",
     1098 => x"59600040",  1099 => x"59600044",  1100 => x"59600088",
     1101 => x"5960008c",  1102 => x"3782000c",  1103 => x"34030000",
     1104 => x"f8003c5d",  1105 => x"44200006",  1106 => x"2b81000c",
     1107 => x"596100a0",  1108 => x"34010001",  1109 => x"596100a4",
     1110 => x"e0000003",  1111 => x"596000a0",  1112 => x"596000a4",
     1113 => x"34010000",  1114 => x"f800286a",  1115 => x"5961002c",
     1116 => x"34010001",  1117 => x"59610054",  1118 => x"59610050",
     1119 => x"34010000",  1120 => x"f8003be8",  1121 => x"59610034",
     1122 => x"34011f40",  1123 => x"596100b4",  1124 => x"78010001",
     1125 => x"382143f0",  1126 => x"28210000",  1127 => x"596100b8",
     1128 => x"596100bc",  1129 => x"35610014",  1130 => x"f800280f",
     1131 => x"34010000",  1132 => x"5960001c",  1133 => x"2b9d0004",
     1134 => x"2b8b0008",  1135 => x"379c000c",  1136 => x"c3a00000",
     1137 => x"c3a00000",  1138 => x"379cffbc",  1139 => x"5b8b0014",
     1140 => x"5b8c0010",  1141 => x"5b8d000c",  1142 => x"5b8e0008",
     1143 => x"5b9d0004",  1144 => x"5b830030",  1145 => x"78030001",
     1146 => x"38634e9c",  1147 => x"5b82002c",  1148 => x"5b840034",
     1149 => x"5b850038",  1150 => x"5b86003c",  1151 => x"5b870040",
     1152 => x"5b880044",  1153 => x"286d0000",  1154 => x"b8205800",
     1155 => x"b8407000",  1156 => x"34030000",  1157 => x"44200002",
     1158 => x"28230018",  1159 => x"b86d1800",  1160 => x"0063001c",
     1161 => x"4460001b",  1162 => x"780c0001",  1163 => x"398c4e9c",
     1164 => x"39a10001",  1165 => x"59810000",  1166 => x"29610028",
     1167 => x"37820018",  1168 => x"28230000",  1169 => x"b9600800",
     1170 => x"d8600000",  1171 => x"78030001",  1172 => x"38633ce4",
     1173 => x"28620000",  1174 => x"2b81001c",  1175 => x"598d0000",
     1176 => x"296b0334",  1177 => x"f8003f0b",  1178 => x"780c0001",
     1179 => x"2b830018",  1180 => x"398c1d78",  1181 => x"b8202000",
     1182 => x"b9601000",  1183 => x"b9800800",  1184 => x"f80026d1",
     1185 => x"b9c00800",  1186 => x"37820030",  1187 => x"f80026ac",
     1188 => x"2b9d0004",  1189 => x"2b8b0014",  1190 => x"2b8c0010",
     1191 => x"2b8d000c",  1192 => x"2b8e0008",  1193 => x"379c0044",
     1194 => x"c3a00000",  1195 => x"379cfffc",  1196 => x"5b9d0004",
     1197 => x"b8402800",  1198 => x"5c600005",  1199 => x"78020001",
     1200 => x"38421d94",  1201 => x"b8a01800",  1202 => x"e000000c",
     1203 => x"34020001",  1204 => x"5c620006",  1205 => x"78020001",
     1206 => x"38421db0",  1207 => x"b8a01800",  1208 => x"28240008",
     1209 => x"e0000005",  1210 => x"28240004",  1211 => x"78020001",
     1212 => x"38421dc8",  1213 => x"b8a01800",  1214 => x"fbffffb4",
     1215 => x"2b9d0004",  1216 => x"379c0004",  1217 => x"c3a00000",
     1218 => x"379cffe8",  1219 => x"5b8b0018",  1220 => x"5b8c0014",
     1221 => x"5b8d0010",  1222 => x"5b8e000c",  1223 => x"5b9d0008",
     1224 => x"b8205800",  1225 => x"b8407000",  1226 => x"b8606800",
     1227 => x"4460001a",  1228 => x"40480000",  1229 => x"78020001",
     1230 => x"38424a14",  1231 => x"2108000f",  1232 => x"3d030002",
     1233 => x"282600e4",  1234 => x"b4431000",  1235 => x"28420000",
     1236 => x"282700e8",  1237 => x"78040001",  1238 => x"5b820004",
     1239 => x"34030001",  1240 => x"34020005",  1241 => x"38841de0",
     1242 => x"b9a02800",  1243 => x"f8000048",  1244 => x"34010021",
     1245 => x"4c2d0006",  1246 => x"b9600800",  1247 => x"b9c01000",
     1248 => x"b9a01800",  1249 => x"f80015f5",  1250 => x"44200003",
     1251 => x"340d0000",  1252 => x"340e0000",  1253 => x"780c0001",
     1254 => x"29610000",  1255 => x"398c48a4",  1256 => x"e000002d",
     1257 => x"44410003",  1258 => x"358c000c",  1259 => x"e000002a",
     1260 => x"59610004",  1261 => x"2961000c",  1262 => x"59600008",
     1263 => x"44200006",  1264 => x"29820004",  1265 => x"b9600800",
     1266 => x"34030000",  1267 => x"b9a02000",  1268 => x"fbffffb7",
     1269 => x"29840008",  1270 => x"b9a01800",  1271 => x"b9600800",
     1272 => x"b9c01000",  1273 => x"d8800000",  1274 => x"b8201800",
     1275 => x"44200006",  1276 => x"29620334",  1277 => x"29840004",
     1278 => x"78010001",  1279 => x"38211e0c",  1280 => x"f8002671",
     1281 => x"29610004",  1282 => x"29630000",  1283 => x"29820004",
     1284 => x"4461000a",  1285 => x"59610000",  1286 => x"34010001",
     1287 => x"5961000c",  1288 => x"34030002",  1289 => x"b9600800",
     1290 => x"34040000",  1291 => x"fbffffa0",  1292 => x"34010000",
     1293 => x"e000000f",  1294 => x"b9600800",  1295 => x"5960000c",
     1296 => x"34030001",  1297 => x"34040000",  1298 => x"fbffff99",
     1299 => x"29610008",  1300 => x"e0000008",  1301 => x"29820000",
     1302 => x"5c40ffd3",  1303 => x"29620334",  1304 => x"78010001",
     1305 => x"38211e28",  1306 => x"f8002657",  1307 => x"34012710",
     1308 => x"2b9d0008",  1309 => x"2b8b0018",  1310 => x"2b8c0014",
     1311 => x"2b8d0010",  1312 => x"2b8e000c",  1313 => x"379c0018",
     1314 => x"c3a00000",  1315 => x"379cffe0",  1316 => x"5b8b000c",
     1317 => x"5b8c0008",  1318 => x"5b9d0004",  1319 => x"5b850014",
     1320 => x"5b840010",  1321 => x"78050001",  1322 => x"5b860018",
     1323 => x"5b87001c",  1324 => x"5b880020",  1325 => x"b8604800",
     1326 => x"b8806000",  1327 => x"38a51e48",  1328 => x"34030000",
     1329 => x"44200003",  1330 => x"28250334",  1331 => x"28230018",
     1332 => x"78060001",  1333 => x"38c64e9c",  1334 => x"28c10000",
     1335 => x"b8610800",  1336 => x"3c430002",  1337 => x"80230800",
     1338 => x"2021000f",  1339 => x"55210015",  1340 => x"78010001",
     1341 => x"38213da0",  1342 => x"b4231800",  1343 => x"78060001",
     1344 => x"28630000",  1345 => x"780b0001",  1346 => x"396b4ea0",
     1347 => x"b8c01000",  1348 => x"38421e50",  1349 => x"b9202000",
     1350 => x"b9600800",  1351 => x"f800261c",  1352 => x"b9600800",
     1353 => x"f80034b2",  1354 => x"b9600800",  1355 => x"b9801000",
     1356 => x"37830014",  1357 => x"f8002633",  1358 => x"b9600800",
     1359 => x"f80034ac",  1360 => x"2b9d0004",  1361 => x"2b8b000c",
     1362 => x"2b8c0008",  1363 => x"379c0020",  1364 => x"c3a00000",
     1365 => x"379cfff8",  1366 => x"5b8b0008",  1367 => x"5b9d0004",
     1368 => x"3402001c",  1369 => x"b8201800",  1370 => x"340b0000",
     1371 => x"3405fffc",  1372 => x"34040003",  1373 => x"e0000009",
     1374 => x"3421ffd0",  1375 => x"202600ff",  1376 => x"50860002",
     1377 => x"e0000008",  1378 => x"bc220800",  1379 => x"34630001",
     1380 => x"b9615800",  1381 => x"3442fffc",  1382 => x"40610000",
     1383 => x"44200007",  1384 => x"5c45fff6",  1385 => x"78010001",
     1386 => x"78020001",  1387 => x"38211e5c",  1388 => x"38423d90",
     1389 => x"f8002604",  1390 => x"b9600800",  1391 => x"2b9d0004",
     1392 => x"2b8b0008",  1393 => x"379c0008",  1394 => x"c3a00000",
     1395 => x"379cfffc",  1396 => x"5b9d0004",  1397 => x"34030001",
     1398 => x"34010003",  1399 => x"34020000",  1400 => x"f80039eb",
     1401 => x"34010000",  1402 => x"34020001",  1403 => x"f8003b98",
     1404 => x"34010000",  1405 => x"2b9d0004",  1406 => x"379c0004",
     1407 => x"c3a00000",  1408 => x"379cfff4",  1409 => x"5b8b000c",
     1410 => x"5b8c0008",  1411 => x"5b9d0004",  1412 => x"34010000",
     1413 => x"b8406000",  1414 => x"f8003ac2",  1415 => x"45800005",
     1416 => x"642c0000",  1417 => x"c80c6000",  1418 => x"398c0001",
     1419 => x"e000000f",  1420 => x"780b0001",  1421 => x"396b4f20",
     1422 => x"5c2c0004",  1423 => x"59600000",  1424 => x"340cffff",
     1425 => x"e0000009",  1426 => x"29610000",  1427 => x"340c0001",
     1428 => x"5c200006",  1429 => x"78020001",  1430 => x"34010003",
     1431 => x"384243f0",  1432 => x"f8002db3",  1433 => x"596c0000",
     1434 => x"b9800800",  1435 => x"2b9d0004",  1436 => x"2b8b000c",
     1437 => x"2b8c0008",  1438 => x"379c000c",  1439 => x"c3a00000",
     1440 => x"34010000",  1441 => x"c3a00000",  1442 => x"379cfffc",
     1443 => x"5b9d0004",  1444 => x"34010000",  1445 => x"34020001",
     1446 => x"f8003b6d",  1447 => x"34010000",  1448 => x"2b9d0004",
     1449 => x"379c0004",  1450 => x"c3a00000",  1451 => x"379cfffc",
     1452 => x"5b9d0004",  1453 => x"282102c8",  1454 => x"28210010",
     1455 => x"2823000c",  1456 => x"44430004",  1457 => x"5822000c",
     1458 => x"b8400800",  1459 => x"f8002bd2",  1460 => x"34010000",
     1461 => x"2b9d0004",  1462 => x"379c0004",  1463 => x"c3a00000",
     1464 => x"379cfffc",  1465 => x"5b9d0004",  1466 => x"f8002bc4",
     1467 => x"34020001",  1468 => x"5c200003",  1469 => x"f8003b46",
     1470 => x"7c220000",  1471 => x"b8400800",  1472 => x"2b9d0004",
     1473 => x"379c0004",  1474 => x"c3a00000",  1475 => x"379cfff8",
     1476 => x"5b8b0008",  1477 => x"5b9d0004",  1478 => x"b8202800",
     1479 => x"b8220800",  1480 => x"b8402000",  1481 => x"b8605800",
     1482 => x"44200005",  1483 => x"34010001",  1484 => x"b8a01000",
     1485 => x"b8801800",  1486 => x"f8002b26",  1487 => x"45600005",
     1488 => x"1562001f",  1489 => x"34010002",  1490 => x"b9601800",
     1491 => x"f8002b21",  1492 => x"34010000",  1493 => x"2b9d0004",
     1494 => x"2b8b0008",  1495 => x"379c0008",  1496 => x"c3a00000",
     1497 => x"379cfffc",  1498 => x"5b9d0004",  1499 => x"b8201000",
     1500 => x"3401ffff",  1501 => x"f8003a7c",  1502 => x"34010000",
     1503 => x"2b9d0004",  1504 => x"379c0004",  1505 => x"c3a00000",
     1506 => x"379cff24",  1507 => x"5b8b0014",  1508 => x"5b8c0010",
     1509 => x"5b8d000c",  1510 => x"5b8e0008",  1511 => x"5b9d0004",
     1512 => x"b8406000",  1513 => x"28220330",  1514 => x"b8807000",
     1515 => x"37810018",  1516 => x"b8605800",  1517 => x"b8a06800",
     1518 => x"fbfffe4d",  1519 => x"45c00005",  1520 => x"78010001",
     1521 => x"382143ec",  1522 => x"28210000",  1523 => x"59c10000",
     1524 => x"45a00003",  1525 => x"2b8100cc",  1526 => x"59a10000",
     1527 => x"2b82006c",  1528 => x"3401fffd",  1529 => x"44400013",
     1530 => x"45800007",  1531 => x"2b820060",  1532 => x"2b810058",
     1533 => x"b4410800",  1534 => x"2b8200a0",  1535 => x"b4220800",
     1536 => x"59810000",  1537 => x"2b820068",  1538 => x"3401fffd",
     1539 => x"44400009",  1540 => x"34010000",  1541 => x"45600007",
     1542 => x"2b830064",  1543 => x"2b82005c",  1544 => x"b4621000",
     1545 => x"2b8300a4",  1546 => x"b4431000",  1547 => x"59620000",
     1548 => x"2b9d0004",  1549 => x"2b8b0014",  1550 => x"2b8c0010",
     1551 => x"2b8d000c",  1552 => x"2b8e0008",  1553 => x"379c00dc",
     1554 => x"c3a00000",  1555 => x"34010000",  1556 => x"c3a00000",
     1557 => x"34010000",  1558 => x"c3a00000",  1559 => x"379cffec",
     1560 => x"5b8b000c",  1561 => x"5b8c0008",  1562 => x"5b9d0004",
     1563 => x"34040000",  1564 => x"b8406000",  1565 => x"b8605800",
     1566 => x"37820010",  1567 => x"37830014",  1568 => x"34050000",
     1569 => x"5b800014",  1570 => x"5b800010",  1571 => x"fbffffbf",
     1572 => x"34010001",  1573 => x"5d810003",  1574 => x"2b810010",
     1575 => x"e0000002",  1576 => x"2b810014",  1577 => x"59610000",
     1578 => x"34010001",  1579 => x"2b9d0004",  1580 => x"2b8b000c",
     1581 => x"2b8c0008",  1582 => x"379c0014",  1583 => x"c3a00000",
     1584 => x"379cfffc",  1585 => x"5b9d0004",  1586 => x"f80026d3",
     1587 => x"34010000",  1588 => x"2b9d0004",  1589 => x"379c0004",
     1590 => x"c3a00000",  1591 => x"379cfffc",  1592 => x"5b9d0004",
     1593 => x"f80026d7",  1594 => x"34010000",  1595 => x"2b9d0004",
     1596 => x"379c0004",  1597 => x"c3a00000",  1598 => x"379cfffc",
     1599 => x"5b9d0004",  1600 => x"f8002bf0",  1601 => x"f800339d",
     1602 => x"f80033a5",  1603 => x"78010001",  1604 => x"78020001",
     1605 => x"38421efc",  1606 => x"38211ecc",  1607 => x"f800252a",
     1608 => x"34010000",  1609 => x"2b9d0004",  1610 => x"379c0004",
     1611 => x"c3a00000",  1612 => x"78010001",  1613 => x"38214f24",
     1614 => x"28210000",  1615 => x"c3a00000",  1616 => x"379cfff8",
     1617 => x"5b8b0008",  1618 => x"5b9d0004",  1619 => x"78010001",
     1620 => x"78020001",  1621 => x"38424a74",  1622 => x"38214770",
     1623 => x"780b0001",  1624 => x"f8001981",  1625 => x"396b43fc",
     1626 => x"34030000",  1627 => x"b9600800",  1628 => x"34020000",
     1629 => x"fbfffe65",  1630 => x"78020001",  1631 => x"384247b4",
     1632 => x"58410000",  1633 => x"f8002b42",  1634 => x"78020001",
     1635 => x"38424f30",  1636 => x"58410000",  1637 => x"296102c8",
     1638 => x"28210010",  1639 => x"58200068",  1640 => x"f8000ae8",
     1641 => x"78010001",  1642 => x"38214f2c",  1643 => x"34020001",
     1644 => x"58220000",  1645 => x"34010000",  1646 => x"2b9d0004",
     1647 => x"2b8b0008",  1648 => x"379c0008",  1649 => x"c3a00000",
     1650 => x"379cfff4",  1651 => x"5b8b000c",  1652 => x"5b8c0008",
     1653 => x"5b9d0004",  1654 => x"780b0001",  1655 => x"396b43fc",
     1656 => x"296102c8",  1657 => x"34020000",  1658 => x"282c0010",
     1659 => x"29810000",  1660 => x"28230034",  1661 => x"b9600800",
     1662 => x"d8600000",  1663 => x"78010001",  1664 => x"34020000",
     1665 => x"340301b8",  1666 => x"59800040",  1667 => x"31800035",
     1668 => x"3821450c",  1669 => x"f8003e4b",  1670 => x"78010001",
     1671 => x"38214f2c",  1672 => x"58200000",  1673 => x"0d60010c",
     1674 => x"f8000ac6",  1675 => x"78010001",  1676 => x"38214770",
     1677 => x"f8001995",  1678 => x"34010000",  1679 => x"2b9d0004",
     1680 => x"2b8b000c",  1681 => x"2b8c0008",  1682 => x"379c000c",
     1683 => x"c3a00000",  1684 => x"379cffec",  1685 => x"5b8b0014",
     1686 => x"5b8c0010",  1687 => x"5b8d000c",  1688 => x"5b8e0008",
     1689 => x"5b9d0004",  1690 => x"780b0001",  1691 => x"396b43fc",
     1692 => x"b8206000",  1693 => x"296102c8",  1694 => x"282d0010",
     1695 => x"78010001",  1696 => x"38214f24",  1697 => x"58200000",
     1698 => x"fbffffd0",  1699 => x"34010002",  1700 => x"45810016",
     1701 => x"34020003",  1702 => x"45820026",  1703 => x"34010001",
     1704 => x"5d81002e",  1705 => x"78010001",  1706 => x"31ac0004",
     1707 => x"38214a74",  1708 => x"340e0006",  1709 => x"316c001d",
     1710 => x"302e0000",  1711 => x"34020000",  1712 => x"34010001",
     1713 => x"34030001",  1714 => x"f80038b1",  1715 => x"29610020",
     1716 => x"2821000c",  1717 => x"302e000e",  1718 => x"b9600800",
     1719 => x"f8001295",  1720 => x"380bea60",  1721 => x"e000001e",
     1722 => x"34010001",  1723 => x"31a10004",  1724 => x"3161001d",
     1725 => x"78010001",  1726 => x"38214a74",  1727 => x"340effbb",
     1728 => x"302e0000",  1729 => x"34020000",  1730 => x"34010002",
     1731 => x"34030001",  1732 => x"f800389f",  1733 => x"29610020",
     1734 => x"2821000c",  1735 => x"302e000e",  1736 => x"b9600800",
     1737 => x"f8001283",  1738 => x"340b0fa0",  1739 => x"e000000c",
     1740 => x"31a10004",  1741 => x"3161001d",  1742 => x"78010001",
     1743 => x"38214a74",  1744 => x"3402ffff",  1745 => x"30220000",
     1746 => x"34030001",  1747 => x"34010003",  1748 => x"34020000",
     1749 => x"f800388e",  1750 => x"340b0000",  1751 => x"f8002acc",
     1752 => x"78020001",  1753 => x"b8207000",  1754 => x"b8400800",
     1755 => x"38211f18",  1756 => x"f8002495",  1757 => x"29a20000",
     1758 => x"780d0001",  1759 => x"39ad1f34",  1760 => x"28430034",
     1761 => x"78020001",  1762 => x"b8400800",  1763 => x"382143fc",
     1764 => x"34020000",  1765 => x"d8600000",  1766 => x"e000000e",
     1767 => x"f8003a8d",  1768 => x"340103e8",  1769 => x"f8002abf",
     1770 => x"f8002ab9",  1771 => x"c82e1000",  1772 => x"51620006",
     1773 => x"78010001",  1774 => x"38211f24",  1775 => x"f8002482",
     1776 => x"340bff8c",  1777 => x"e0000008",  1778 => x"b9a00800",
     1779 => x"f800247e",  1780 => x"34010000",  1781 => x"f8003953",
     1782 => x"5c200002",  1783 => x"5d61fff0",  1784 => x"340b0000",
     1785 => x"78010001",  1786 => x"38211b1c",  1787 => x"f8002476",
     1788 => x"7d620000",  1789 => x"65810001",  1790 => x"a0410800",
     1791 => x"44200005",  1792 => x"78010001",  1793 => x"38214a74",
     1794 => x"34020034",  1795 => x"30220000",  1796 => x"78010001",
     1797 => x"38214f24",  1798 => x"582c0000",  1799 => x"b9600800",
     1800 => x"2b9d0004",  1801 => x"2b8b0014",  1802 => x"2b8c0010",
     1803 => x"2b8d000c",  1804 => x"2b8e0008",  1805 => x"379c0014",
     1806 => x"c3a00000",  1807 => x"379cfff0",  1808 => x"5b8b0010",
     1809 => x"5b8c000c",  1810 => x"5b8d0008",  1811 => x"5b9d0004",
     1812 => x"34010000",  1813 => x"f80025af",  1814 => x"78020001",
     1815 => x"38424f28",  1816 => x"b8205800",  1817 => x"28410000",
     1818 => x"442b0018",  1819 => x"78010001",  1820 => x"38214f2c",
     1821 => x"28210000",  1822 => x"584b0000",  1823 => x"65620000",
     1824 => x"7c210000",  1825 => x"a0410800",  1826 => x"44200005",
     1827 => x"fbffff4f",  1828 => x"78010001",  1829 => x"38211f38",
     1830 => x"f800244b",  1831 => x"78010001",  1832 => x"38214f2c",
     1833 => x"28210000",  1834 => x"7d6b0000",  1835 => x"64210000",
     1836 => x"a1615800",  1837 => x"45600005",  1838 => x"78010001",
     1839 => x"38211f50",  1840 => x"f8002441",  1841 => x"fbffff1f",
     1842 => x"78010001",  1843 => x"38214f2c",  1844 => x"28210000",
     1845 => x"44200022",  1846 => x"780b0001",  1847 => x"396b43fc",
     1848 => x"29610024",  1849 => x"29620038",  1850 => x"78040001",
     1851 => x"28250008",  1852 => x"3403007c",  1853 => x"b9600800",
     1854 => x"388444e0",  1855 => x"d8a00000",  1856 => x"b8201800",
     1857 => x"4801000f",  1858 => x"29610370",  1859 => x"34210001",
     1860 => x"59610370",  1861 => x"5c60000b",  1862 => x"780d0001",
     1863 => x"f8002a5c",  1864 => x"39ad4f30",  1865 => x"29a20000",
     1866 => x"780c0001",  1867 => x"398c47b4",  1868 => x"c8220800",
     1869 => x"29820000",  1870 => x"54410009",  1871 => x"e000000f",
     1872 => x"78010001",  1873 => x"382143fc",  1874 => x"28220040",
     1875 => x"fbfffd6f",  1876 => x"78020001",  1877 => x"384247b4",
     1878 => x"58410000",  1879 => x"34010000",  1880 => x"2b9d0004",
     1881 => x"2b8b0010",  1882 => x"2b8c000c",  1883 => x"2b8d0008",
     1884 => x"379c0010",  1885 => x"c3a00000",  1886 => x"f8002a45",
     1887 => x"59a10000",  1888 => x"34020000",  1889 => x"b9600800",
     1890 => x"34030000",  1891 => x"fbfffd5f",  1892 => x"59810000",
     1893 => x"e3fffff2",  1894 => x"379cffe8",  1895 => x"5b9d0018",
     1896 => x"b8205000",  1897 => x"40610005",  1898 => x"40640000",
     1899 => x"40650001",  1900 => x"40660002",  1901 => x"40670003",
     1902 => x"40680004",  1903 => x"5b810004",  1904 => x"40610006",
     1905 => x"b8404800",  1906 => x"b9401000",  1907 => x"5b810008",
     1908 => x"40610007",  1909 => x"5b81000c",  1910 => x"40610008",
     1911 => x"5b810010",  1912 => x"40610009",  1913 => x"b9201800",
     1914 => x"5b810014",  1915 => x"78010001",  1916 => x"38211f68",
     1917 => x"f80023f4",  1918 => x"2b9d0018",  1919 => x"379c0018",
     1920 => x"c3a00000",  1921 => x"379cffd0",  1922 => x"5b8b0030",
     1923 => x"5b8c002c",  1924 => x"5b8d0028",  1925 => x"5b8e0024",
     1926 => x"5b8f0020",  1927 => x"5b90001c",  1928 => x"5b910018",
     1929 => x"5b920014",  1930 => x"5b930010",  1931 => x"5b94000c",
     1932 => x"5b950008",  1933 => x"5b9d0004",  1934 => x"b8603000",
     1935 => x"b8209800",  1936 => x"b8409000",  1937 => x"78010001",
     1938 => x"b880a800",  1939 => x"38211fa0",  1940 => x"ba601000",
     1941 => x"ba401800",  1942 => x"b8c02000",  1943 => x"b8a0a000",
     1944 => x"78110001",  1945 => x"f80023d8",  1946 => x"78100001",
     1947 => x"780f0001",  1948 => x"780e0001",  1949 => x"780d0001",
     1950 => x"b8205800",  1951 => x"340c0000",  1952 => x"3a311fb4",
     1953 => x"3a101fbc",  1954 => x"39ef1c40",  1955 => x"39ce1b1c",
     1956 => x"39ad19b8",  1957 => x"e0000017",  1958 => x"5cc00006",
     1959 => x"ba200800",  1960 => x"ba601000",  1961 => x"ba401800",
     1962 => x"f80023c7",  1963 => x"b5615800",  1964 => x"b6ac1000",
     1965 => x"40420000",  1966 => x"ba000800",  1967 => x"358c0001",
     1968 => x"f80023c1",  1969 => x"21820003",  1970 => x"b42b5800",
     1971 => x"b9e03000",  1972 => x"5c400005",  1973 => x"2181000f",
     1974 => x"b9c03000",  1975 => x"44220002",  1976 => x"b9a03000",
     1977 => x"b8c00800",  1978 => x"f80023b7",  1979 => x"b5615800",
     1980 => x"2186000f",  1981 => x"4a8cffe9",  1982 => x"44c00005",
     1983 => x"78010001",  1984 => x"38211b1c",  1985 => x"f80023b0",
     1986 => x"b42b5800",  1987 => x"b9600800",  1988 => x"2b9d0004",
     1989 => x"2b8b0030",  1990 => x"2b8c002c",  1991 => x"2b8d0028",
     1992 => x"2b8e0024",  1993 => x"2b8f0020",  1994 => x"2b90001c",
     1995 => x"2b910018",  1996 => x"2b920014",  1997 => x"2b930010",
     1998 => x"2b94000c",  1999 => x"2b950008",  2000 => x"379c0030",
     2001 => x"c3a00000",  2002 => x"379cffb8",  2003 => x"5b8b0048",
     2004 => x"5b8c0044",  2005 => x"5b8d0040",  2006 => x"5b8e003c",
     2007 => x"5b8f0038",  2008 => x"5b900034",  2009 => x"5b910030",
     2010 => x"5b92002c",  2011 => x"5b930028",  2012 => x"5b940024",
     2013 => x"5b950020",  2014 => x"5b96001c",  2015 => x"5b970018",
     2016 => x"5b980014",  2017 => x"5b9d0010",  2018 => x"b8608000",
     2019 => x"40430001",  2020 => x"b8206000",  2021 => x"34010002",
     2022 => x"2063000f",  2023 => x"b8406800",  2024 => x"404e0000",
     2025 => x"44610006",  2026 => x"78010001",  2027 => x"b9801000",
     2028 => x"38211fc4",  2029 => x"f8002384",  2030 => x"e000013f",
     2031 => x"40450002",  2032 => x"40460003",  2033 => x"21ce000f",
     2034 => x"3ca50008",  2035 => x"78010001",  2036 => x"b8c52800",
     2037 => x"41a60004",  2038 => x"34030002",  2039 => x"b9c02000",
     2040 => x"344b0022",  2041 => x"38211fe4",  2042 => x"b9801000",
     2043 => x"f8002376",  2044 => x"41a2000c",  2045 => x"41a1000d",
     2046 => x"41a4000e",  2047 => x"41a30006",  2048 => x"3c420018",
     2049 => x"3c210010",  2050 => x"41a60007",  2051 => x"41a5000f",
     2052 => x"3c840008",  2053 => x"b8220800",  2054 => x"3c630008",
     2055 => x"b8812000",  2056 => x"78010001",  2057 => x"b8c31800",
     2058 => x"b8a42000",  2059 => x"b9801000",  2060 => x"38212010",
     2061 => x"f8002364",  2062 => x"78020001",  2063 => x"b9800800",
     2064 => x"38422034",  2065 => x"35a30014",  2066 => x"fbffff54",
     2067 => x"41a3001e",  2068 => x"41a4001f",  2069 => x"41a50021",
     2070 => x"3c630008",  2071 => x"78010001",  2072 => x"b8831800",
     2073 => x"41a40020",  2074 => x"3821203c",  2075 => x"b9801000",
     2076 => x"f8002355",  2077 => x"3401000c",  2078 => x"55c100d1",
     2079 => x"78010001",  2080 => x"3dce0002",  2081 => x"38213dc0",
     2082 => x"b42e0800",  2083 => x"28210000",  2084 => x"c0200000",
     2085 => x"78010001",  2086 => x"b9801000",  2087 => x"38212068",
     2088 => x"f8002349",  2089 => x"41620002",  2090 => x"41610003",
     2091 => x"41640004",  2092 => x"3c420018",  2093 => x"3c210010",
     2094 => x"3c840008",  2095 => x"b8220800",  2096 => x"b8812000",
     2097 => x"41620006",  2098 => x"41610007",  2099 => x"41650008",
     2100 => x"3c420018",  2101 => x"3c210010",  2102 => x"3ca50008",
     2103 => x"b8220800",  2104 => x"b8a12800",  2105 => x"78030001",
     2106 => x"78010001",  2107 => x"41670005",  2108 => x"41660009",
     2109 => x"38212080",  2110 => x"b9801000",  2111 => x"38632090",
     2112 => x"e000001c",  2113 => x"78010001",  2114 => x"b9801000",
     2115 => x"3821209c",  2116 => x"f800232d",  2117 => x"41620002",
     2118 => x"41610003",  2119 => x"41640004",  2120 => x"3c420018",
     2121 => x"3c210010",  2122 => x"3c840008",  2123 => x"b8220800",
     2124 => x"b8812000",  2125 => x"41620006",  2126 => x"41610007",
     2127 => x"41650008",  2128 => x"3c420018",  2129 => x"3c210010",
     2130 => x"3ca50008",  2131 => x"b8220800",  2132 => x"41670005",
     2133 => x"41660009",  2134 => x"b8a12800",  2135 => x"78030001",
     2136 => x"78010001",  2137 => x"38212080",  2138 => x"b9801000",
     2139 => x"386320b8",  2140 => x"b8e42000",  2141 => x"b8c52800",
     2142 => x"f8002313",  2143 => x"e000008e",  2144 => x"78010001",
     2145 => x"b9801000",  2146 => x"382120c8",  2147 => x"f800230e",
     2148 => x"41620002",  2149 => x"41610003",  2150 => x"41640004",
     2151 => x"3c420018",  2152 => x"3c210010",  2153 => x"3c840008",
     2154 => x"b8220800",  2155 => x"b8812000",  2156 => x"41620006",
     2157 => x"41610007",  2158 => x"41650008",  2159 => x"3c420018",
     2160 => x"3c210010",  2161 => x"3ca50008",  2162 => x"b8220800",
     2163 => x"b8a12800",  2164 => x"78030001",  2165 => x"78010001",
     2166 => x"41670005",  2167 => x"41660009",  2168 => x"38212080",
     2169 => x"b9801000",  2170 => x"386320e4",  2171 => x"e3ffffe1",
     2172 => x"78010001",  2173 => x"b9801000",  2174 => x"382120f4",
     2175 => x"f80022f2",  2176 => x"41620002",  2177 => x"41610003",
     2178 => x"41640004",  2179 => x"3c420018",  2180 => x"3c210010",
     2181 => x"3c840008",  2182 => x"b8220800",  2183 => x"b8812000",
     2184 => x"41620006",  2185 => x"41610007",  2186 => x"41650008",
     2187 => x"3c420018",  2188 => x"3c210010",  2189 => x"41670005",
     2190 => x"41660009",  2191 => x"3ca50008",  2192 => x"b8220800",
     2193 => x"780e0001",  2194 => x"39ce2110",  2195 => x"b8a12800",
     2196 => x"78010001",  2197 => x"b9801000",  2198 => x"b9c01800",
     2199 => x"b8e42000",  2200 => x"b8c52800",  2201 => x"38212080",
     2202 => x"f80022d7",  2203 => x"3563000a",  2204 => x"b9800800",
     2205 => x"b9c01000",  2206 => x"fbfffec8",  2207 => x"340b0036",
     2208 => x"e0000080",  2209 => x"78010001",  2210 => x"b9801000",
     2211 => x"38212124",  2212 => x"f80022cd",  2213 => x"41620002",
     2214 => x"41610003",  2215 => x"41640004",  2216 => x"3c420018",
     2217 => x"3c210010",  2218 => x"3c840008",  2219 => x"b8220800",
     2220 => x"b8812000",  2221 => x"41620006",  2222 => x"41610007",
     2223 => x"41650008",  2224 => x"3c420018",  2225 => x"3c210010",
     2226 => x"41670005",  2227 => x"41660009",  2228 => x"3ca50008",
     2229 => x"b8220800",  2230 => x"b8a12800",  2231 => x"78030001",
     2232 => x"78010001",  2233 => x"b8e42000",  2234 => x"b8c52800",
     2235 => x"b9801000",  2236 => x"38632140",  2237 => x"38212080",
     2238 => x"f80022b3",  2239 => x"41660010",  2240 => x"41670011",
     2241 => x"4165000f",  2242 => x"4164000e",  2243 => x"3cc60008",
     2244 => x"78010001",  2245 => x"78030001",  2246 => x"b8e63000",
     2247 => x"b9801000",  2248 => x"3863216c",  2249 => x"38212158",
     2250 => x"f80022a7",  2251 => x"4163000d",  2252 => x"41640012",
     2253 => x"78010001",  2254 => x"b9801000",  2255 => x"38212190",
     2256 => x"f80022a1",  2257 => x"41610018",  2258 => x"41640013",
     2259 => x"41650014",  2260 => x"41660015",  2261 => x"41670016",
     2262 => x"41680017",  2263 => x"5b810004",  2264 => x"41610019",
     2265 => x"78030001",  2266 => x"b9801000",  2267 => x"5b810008",
     2268 => x"4161001a",  2269 => x"386321e8",  2270 => x"340b0040",
     2271 => x"5b81000c",  2272 => x"78010001",  2273 => x"382121b8",
     2274 => x"f800228f",  2275 => x"e000003d",  2276 => x"78010001",
     2277 => x"b9801000",  2278 => x"38212208",  2279 => x"f800228a",
     2280 => x"78020001",  2281 => x"b9800800",  2282 => x"38422224",
     2283 => x"b9601800",  2284 => x"fbfffe7a",  2285 => x"340b002c",
     2286 => x"e0000032",  2287 => x"340b0022",  2288 => x"e0000030",
     2289 => x"55f70009",  2290 => x"78010001",  2291 => x"b9801000",
     2292 => x"ba001800",  2293 => x"b9602000",  2294 => x"b9e02800",
     2295 => x"38212240",  2296 => x"f8002279",  2297 => x"e0000034",
     2298 => x"b5ab7000",  2299 => x"41d60002",  2300 => x"41c10003",
     2301 => x"41c30000",  2302 => x"3ed60008",  2303 => x"41c40001",
     2304 => x"b836b000",  2305 => x"41c10008",  2306 => x"41c50004",
     2307 => x"41c60005",  2308 => x"41c70006",  2309 => x"41c80007",
     2310 => x"5b810004",  2311 => x"41c10009",  2312 => x"3c630008",
     2313 => x"36d10004",  2314 => x"5b810008",  2315 => x"b8831800",
     2316 => x"baa00800",  2317 => x"b9801000",  2318 => x"ba202000",
     2319 => x"f8002262",  2320 => x"4df10007",  2321 => x"ba400800",
     2322 => x"b9801000",  2323 => x"ba201800",  2324 => x"b9e02000",
     2325 => x"f800225c",  2326 => x"e0000008",  2327 => x"b9800800",
     2328 => x"ba801000",  2329 => x"ba601800",  2330 => x"35c4000a",
     2331 => x"36c5fffa",  2332 => x"fbfffe65",  2333 => x"ba207800",
     2334 => x"b56f5800",  2335 => x"e000000b",  2336 => x"78150001",
     2337 => x"78140001",  2338 => x"78130001",  2339 => x"78120001",
     2340 => x"34180002",  2341 => x"34170009",  2342 => x"3ab52264",
     2343 => x"3a9422d0",  2344 => x"3a7322d8",  2345 => x"3a5222a4",
     2346 => x"4d700003",  2347 => x"ca0b7800",  2348 => x"49f8ffc5",
     2349 => x"78020001",  2350 => x"78030001",  2351 => x"b9800800",
     2352 => x"384222e4",  2353 => x"386322ec",  2354 => x"b9a02000",
     2355 => x"ba002800",  2356 => x"fbfffe4d",  2357 => x"2b9d0010",
     2358 => x"2b8b0048",  2359 => x"2b8c0044",  2360 => x"2b8d0040",
     2361 => x"2b8e003c",  2362 => x"2b8f0038",  2363 => x"2b900034",
     2364 => x"2b910030",  2365 => x"2b92002c",  2366 => x"2b930028",
     2367 => x"2b940024",  2368 => x"2b950020",  2369 => x"2b96001c",
     2370 => x"2b970018",  2371 => x"2b980014",  2372 => x"379c0048",
     2373 => x"c3a00000",  2374 => x"379cfff0",  2375 => x"5b8b0010",
     2376 => x"5b8c000c",  2377 => x"5b8d0008",  2378 => x"5b9d0004",
     2379 => x"b8205800",  2380 => x"b8406800",  2381 => x"b8606000",
     2382 => x"4480000f",  2383 => x"2881000c",  2384 => x"78070001",
     2385 => x"28850000",  2386 => x"28860004",  2387 => x"38e73cd4",
     2388 => x"5c200003",  2389 => x"78070001",  2390 => x"38e722f4",
     2391 => x"78010001",  2392 => x"38212300",  2393 => x"b9601000",
     2394 => x"b8a01800",  2395 => x"b8a02000",  2396 => x"f8002215",
     2397 => x"b9600800",  2398 => x"b9a01000",  2399 => x"b9801800",
     2400 => x"fbfffe72",  2401 => x"34010000",  2402 => x"2b9d0004",
     2403 => x"2b8b0010",  2404 => x"2b8c000c",  2405 => x"2b8d0008",
     2406 => x"379c0010",  2407 => x"c3a00000",  2408 => x"379cffe8",
     2409 => x"5b8b0018",  2410 => x"5b8c0014",  2411 => x"5b8d0010",
     2412 => x"5b8e000c",  2413 => x"5b8f0008",  2414 => x"5b9d0004",
     2415 => x"282d0000",  2416 => x"b8207800",  2417 => x"282e0004",
     2418 => x"b8406000",  2419 => x"340b0000",  2420 => x"34010000",
     2421 => x"34040000",  2422 => x"544d0006",  2423 => x"b9a00800",
     2424 => x"f8003a79",  2425 => x"882c1000",  2426 => x"b9602000",
     2427 => x"c9a26800",  2428 => x"34030000",  2429 => x"34020001",
     2430 => x"e000000b",  2431 => x"3d850001",  2432 => x"3d6b0001",
     2433 => x"f5856000",  2434 => x"3c630001",  2435 => x"b58b5800",
     2436 => x"b8a06000",  2437 => x"3c450001",  2438 => x"f4451000",
     2439 => x"b4431800",  2440 => x"b8a01000",  2441 => x"1565001f",
     2442 => x"c8ac3000",  2443 => x"f4c53000",  2444 => x"c8ab2800",
     2445 => x"c8a62800",  2446 => x"00a5001f",  2447 => x"34060001",
     2448 => x"55ab0004",  2449 => x"5dab0002",  2450 => x"55cc0002",
     2451 => x"34060000",  2452 => x"a0a63000",  2453 => x"5cc0ffea",
     2454 => x"556d000d",  2455 => x"5d6d0002",  2456 => x"558e000b",
     2457 => x"c9cc2800",  2458 => x"f4ae7000",  2459 => x"c9ab6800",
     2460 => x"c9ae6800",  2461 => x"b8a07000",  2462 => x"b4822800",
     2463 => x"f4852000",  2464 => x"b4230800",  2465 => x"b4810800",
     2466 => x"b8a02000",  2467 => x"3c65001f",  2468 => x"00420001",
     2469 => x"00630001",  2470 => x"b8a21000",  2471 => x"b8622800",
     2472 => x"44a00006",  2473 => x"3d65001f",  2474 => x"018c0001",
     2475 => x"016b0001",  2476 => x"b8ac6000",  2477 => x"e3ffffe9",
     2478 => x"59e10000",  2479 => x"b9c00800",  2480 => x"59e40004",
     2481 => x"2b9d0004",  2482 => x"2b8b0018",  2483 => x"2b8c0014",
     2484 => x"2b8d0010",  2485 => x"2b8e000c",  2486 => x"2b8f0008",
     2487 => x"379c0018",  2488 => x"c3a00000",  2489 => x"379cfff8",
     2490 => x"5b8b0008",  2491 => x"5b9d0004",  2492 => x"b8405800",
     2493 => x"f80027e6",  2494 => x"b42b0800",  2495 => x"5c200002",
     2496 => x"34010001",  2497 => x"2b9d0004",  2498 => x"2b8b0008",
     2499 => x"379c0008",  2500 => x"c3a00000",  2501 => x"379cfff8",
     2502 => x"5b8b0008",  2503 => x"5b9d0004",  2504 => x"78040001",
     2505 => x"b8405800",  2506 => x"78050001",  2507 => x"34020006",
     2508 => x"34030001",  2509 => x"388423cc",  2510 => x"38a53df4",
     2511 => x"b9603000",  2512 => x"fbfffb53",  2513 => x"45600005",
     2514 => x"1562001f",  2515 => x"34010002",  2516 => x"b9601800",
     2517 => x"f800271f",  2518 => x"34010000",  2519 => x"2b9d0004",
     2520 => x"2b8b0008",  2521 => x"379c0008",  2522 => x"c3a00000",
     2523 => x"379cfff4",  2524 => x"5b8b000c",  2525 => x"5b8c0008",
     2526 => x"5b9d0004",  2527 => x"b8206000",  2528 => x"b8405800",
     2529 => x"b8603000",  2530 => x"44600008",  2531 => x"78040001",
     2532 => x"78050001",  2533 => x"34020006",  2534 => x"34030001",
     2535 => x"388423d8",  2536 => x"38a53e0c",  2537 => x"fbfffb3a",
     2538 => x"b9800800",  2539 => x"b9601000",  2540 => x"fbffffd9",
     2541 => x"2b9d0004",  2542 => x"2b8b000c",  2543 => x"2b8c0008",
     2544 => x"379c000c",  2545 => x"c3a00000",  2546 => x"379cfff0",
     2547 => x"5b8b0010",  2548 => x"5b8c000c",  2549 => x"5b8d0008",
     2550 => x"5b9d0004",  2551 => x"b8206800",  2552 => x"44400012",
     2553 => x"284b0000",  2554 => x"284c0004",  2555 => x"34040003",
     2556 => x"1561001f",  2557 => x"b9601000",  2558 => x"b9801800",
     2559 => x"f8002736",  2560 => x"78040001",  2561 => x"78050001",
     2562 => x"b9a00800",  2563 => x"34020006",  2564 => x"34030001",
     2565 => x"38842404",  2566 => x"38a53e20",  2567 => x"b9603000",
     2568 => x"b9803800",  2569 => x"fbfffb1a",  2570 => x"34010000",
     2571 => x"2b9d0004",  2572 => x"2b8b0010",  2573 => x"2b8c000c",
     2574 => x"2b8d0008",  2575 => x"379c0010",  2576 => x"c3a00000",
     2577 => x"379cffe8",  2578 => x"5b8b000c",  2579 => x"5b8c0008",
     2580 => x"5b9d0004",  2581 => x"b8405800",  2582 => x"b8206000",
     2583 => x"37820018",  2584 => x"37810010",  2585 => x"f800273c",
     2586 => x"78020001",  2587 => x"38424e9c",  2588 => x"2b860014",
     2589 => x"2b870018",  2590 => x"28410000",  2591 => x"59660000",
     2592 => x"59670004",  2593 => x"20210001",  2594 => x"5c200009",
     2595 => x"78040001",  2596 => x"78050001",  2597 => x"b9800800",
     2598 => x"34020006",  2599 => x"34030002",  2600 => x"38842404",
     2601 => x"38a53e30",  2602 => x"fbfffaf9",  2603 => x"34010000",
     2604 => x"2b9d0004",  2605 => x"2b8b000c",  2606 => x"2b8c0008",
     2607 => x"379c0018",  2608 => x"c3a00000",  2609 => x"379cffb4",
     2610 => x"5b8b001c",  2611 => x"5b8c0018",  2612 => x"5b8d0014",
     2613 => x"5b8e0010",  2614 => x"5b8f000c",  2615 => x"5b900008",
     2616 => x"5b9d0004",  2617 => x"28300058",  2618 => x"378c0040",
     2619 => x"b8407800",  2620 => x"b8206800",  2621 => x"78020001",
     2622 => x"340188f7",  2623 => x"b8607000",  2624 => x"0f81004c",
     2625 => x"38423d88",  2626 => x"b9800800",  2627 => x"34030006",
     2628 => x"b8805800",  2629 => x"f8003a0d",  2630 => x"b9801000",
     2631 => x"ba000800",  2632 => x"b9e01800",  2633 => x"b9c02000",
     2634 => x"37850020",  2635 => x"f8001df0",  2636 => x"b8206000",
     2637 => x"45600011",  2638 => x"2b81003c",  2639 => x"2b870024",
     2640 => x"2b880028",  2641 => x"78040001",  2642 => x"78050001",
     2643 => x"5961000c",  2644 => x"59670000",  2645 => x"59680004",
     2646 => x"59600008",  2647 => x"b9a00800",  2648 => x"34020005",
     2649 => x"34030002",  2650 => x"38842414",  2651 => x"38a53e40",
     2652 => x"b9803000",  2653 => x"fbfffac6",  2654 => x"4c0c0010",
     2655 => x"78010001",  2656 => x"38214e9c",  2657 => x"28220000",
     2658 => x"29a10018",  2659 => x"b8410800",  2660 => x"00210014",
     2661 => x"34020001",  2662 => x"2021000f",  2663 => x"50410007",
     2664 => x"78010001",  2665 => x"38212434",  2666 => x"b9e01000",
     2667 => x"b9c01800",  2668 => x"b9602000",  2669 => x"fbfffed9",
     2670 => x"b9800800",  2671 => x"2b9d0004",  2672 => x"2b8b001c",
     2673 => x"2b8c0018",  2674 => x"2b8d0014",  2675 => x"2b8e0010",
     2676 => x"2b8f000c",  2677 => x"2b900008",  2678 => x"379c004c",
     2679 => x"c3a00000",  2680 => x"379cffbc",  2681 => x"5b8b0014",
     2682 => x"5b8c0010",  2683 => x"5b8d000c",  2684 => x"5b8e0008",
     2685 => x"5b9d0004",  2686 => x"b8207000",  2687 => x"28210058",
     2688 => x"b8602800",  2689 => x"b8406800",  2690 => x"b8805800",
     2691 => x"37820038",  2692 => x"b8a02000",  2693 => x"b9a01800",
     2694 => x"37850018",  2695 => x"f8001d1c",  2696 => x"b8206000",
     2697 => x"4560000b",  2698 => x"2b81001c",  2699 => x"59610000",
     2700 => x"2b810020",  2701 => x"59610004",  2702 => x"2b810024",
     2703 => x"59610008",  2704 => x"2b810034",  2705 => x"5961000c",
     2706 => x"2b810030",  2707 => x"59610010",  2708 => x"4c0c0010",
     2709 => x"78040001",  2710 => x"38844e9c",  2711 => x"28820000",
     2712 => x"29c10018",  2713 => x"b8410800",  2714 => x"00210014",
     2715 => x"34020001",  2716 => x"2021000f",  2717 => x"50410007",
     2718 => x"78010001",  2719 => x"3821243c",  2720 => x"b9a01000",
     2721 => x"b9801800",  2722 => x"b9602000",  2723 => x"fbfffea3",
     2724 => x"b9800800",  2725 => x"2b9d0004",  2726 => x"2b8b0014",
     2727 => x"2b8c0010",  2728 => x"2b8d000c",  2729 => x"2b8e0008",
     2730 => x"379c0044",  2731 => x"c3a00000",  2732 => x"379cfffc",
     2733 => x"5b9d0004",  2734 => x"28210058",  2735 => x"f8001ca1",
     2736 => x"34010000",  2737 => x"2b9d0004",  2738 => x"379c0004",
     2739 => x"c3a00000",  2740 => x"379cffd8",  2741 => x"5b8b0010",
     2742 => x"5b8c000c",  2743 => x"5b8d0008",  2744 => x"5b9d0004",
     2745 => x"b8205800",  2746 => x"28210058",  2747 => x"44200002",
     2748 => x"f8001c94",  2749 => x"b9600800",  2750 => x"f8000cfb",
     2751 => x"378c0014",  2752 => x"340188f7",  2753 => x"78020001",
     2754 => x"0f810020",  2755 => x"38423d88",  2756 => x"b9800800",
     2757 => x"34030006",  2758 => x"f800398c",  2759 => x"b9801800",
     2760 => x"34010001",  2761 => x"34020000",  2762 => x"f8001c4e",
     2763 => x"b8206000",  2764 => x"4420000e",  2765 => x"378d0024",
     2766 => x"b9a01000",  2767 => x"f8001c3a",  2768 => x"b9a01000",
     2769 => x"34030006",  2770 => x"35610060",  2771 => x"f800397f",
     2772 => x"3561004c",  2773 => x"596c0058",  2774 => x"b9a01000",
     2775 => x"34030006",  2776 => x"f800397a",  2777 => x"596c0044",
     2778 => x"34010000",  2779 => x"2b9d0004",  2780 => x"2b8b0010",
     2781 => x"2b8c000c",  2782 => x"2b8d0008",  2783 => x"379c0028",
     2784 => x"c3a00000",  2785 => x"379cfff8",  2786 => x"5b8b0008",
     2787 => x"5b9d0004",  2788 => x"78040001",  2789 => x"78050001",
     2790 => x"34020002",  2791 => x"34030002",  2792 => x"38842528",
     2793 => x"38a53ea0",  2794 => x"b8205800",  2795 => x"fbfffa38",
     2796 => x"296302c8",  2797 => x"28610010",  2798 => x"28220064",
     2799 => x"34010000",  2800 => x"44400010",  2801 => x"34010001",
     2802 => x"59610004",  2803 => x"1061000b",  2804 => x"4062000c",
     2805 => x"29640028",  2806 => x"bc411000",  2807 => x"28830018",
     2808 => x"084203e8",  2809 => x"b9600800",  2810 => x"d8600000",
     2811 => x"596102d4",  2812 => x"296102c8",  2813 => x"28210010",
     2814 => x"58200064",  2815 => x"34010001",  2816 => x"2b9d0004",
     2817 => x"2b8b0008",  2818 => x"379c0008",  2819 => x"c3a00000",
     2820 => x"379cfff4",  2821 => x"5b8b000c",  2822 => x"5b8c0008",
     2823 => x"5b9d0004",  2824 => x"78040001",  2825 => x"78050001",
     2826 => x"b8606000",  2827 => x"34020002",  2828 => x"34030002",
     2829 => x"38842528",  2830 => x"38a53eb4",  2831 => x"b8205800",
     2832 => x"fbfffa13",  2833 => x"29820024",  2834 => x"296102c8",
     2835 => x"20430003",  2836 => x"28210010",  2837 => x"7c640000",
     2838 => x"58240038",  2839 => x"20440008",  2840 => x"20420004",
     2841 => x"7c840000",  2842 => x"7c420000",  2843 => x"30230035",
     2844 => x"58220044",  2845 => x"58240040",  2846 => x"29610020",
     2847 => x"28220010",  2848 => x"296102c8",  2849 => x"2c210008",
     2850 => x"0c41002c",  2851 => x"2b9d0004",  2852 => x"2b8b000c",
     2853 => x"2b8c0008",  2854 => x"379c000c",  2855 => x"c3a00000",
     2856 => x"379cfff8",  2857 => x"5b8b0008",  2858 => x"5b9d0004",
     2859 => x"282202c8",  2860 => x"78040001",  2861 => x"78050001",
     2862 => x"284b0010",  2863 => x"34030002",  2864 => x"34020002",
     2865 => x"38842528",  2866 => x"38a53eec",  2867 => x"fbfff9f0",
     2868 => x"34010000",  2869 => x"31600005",  2870 => x"2b9d0004",
     2871 => x"2b8b0008",  2872 => x"379c0008",  2873 => x"c3a00000",
     2874 => x"379cfff8",  2875 => x"5b8b0008",  2876 => x"5b9d0004",
     2877 => x"78040001",  2878 => x"78050001",  2879 => x"b8205800",
     2880 => x"34020002",  2881 => x"34010000",  2882 => x"34030002",
     2883 => x"38842528",  2884 => x"38a53efc",  2885 => x"fbfff9de",
     2886 => x"29610024",  2887 => x"44200006",  2888 => x"34020000",
     2889 => x"34030001",  2890 => x"34040002",  2891 => x"34060003",
     2892 => x"e000001f",  2893 => x"29610000",  2894 => x"29620040",
     2895 => x"58220014",  2896 => x"e000001d",  2897 => x"29650000",
     2898 => x"08410374",  2899 => x"b4a10800",  2900 => x"29650040",
     2901 => x"58250014",  2902 => x"28250368",  2903 => x"5ca30010",
     2904 => x"4025001d",  2905 => x"44a30004",  2906 => x"282102c8",
     2907 => x"5ca40009",  2908 => x"e0000005",  2909 => x"282102c8",
     2910 => x"28210010",  2911 => x"30230004",  2912 => x"e000000a",
     2913 => x"28210010",  2914 => x"30240004",  2915 => x"e0000007",
     2916 => x"28210010",  2917 => x"30260004",  2918 => x"e0000004",
     2919 => x"282102c8",  2920 => x"28210010",  2921 => x"30200004",
     2922 => x"34420001",  2923 => x"29610024",  2924 => x"4822ffe5",
     2925 => x"34010000",  2926 => x"2b9d0004",  2927 => x"2b8b0008",
     2928 => x"379c0008",  2929 => x"c3a00000",  2930 => x"379cfff4",
     2931 => x"5b8b000c",  2932 => x"5b8c0008",  2933 => x"5b9d0004",
     2934 => x"282202c8",  2935 => x"78040001",  2936 => x"78050001",
     2937 => x"284b0010",  2938 => x"34030002",  2939 => x"34020002",
     2940 => x"38842528",  2941 => x"38a53f04",  2942 => x"b8206000",
     2943 => x"fbfff9a4",  2944 => x"41630004",  2945 => x"3401012c",
     2946 => x"59610028",  2947 => x"34020001",  2948 => x"34010bb8",
     2949 => x"59610030",  2950 => x"59600008",  2951 => x"31600035",
     2952 => x"59600040",  2953 => x"59620014",  2954 => x"20630003",
     2955 => x"29610000",  2956 => x"5c620004",  2957 => x"28230034",
     2958 => x"b9800800",  2959 => x"e0000004",  2960 => x"28230034",
     2961 => x"34020000",  2962 => x"b9800800",  2963 => x"d8600000",
     2964 => x"34010000",  2965 => x"2b9d0004",  2966 => x"2b8b000c",
     2967 => x"2b8c0008",  2968 => x"379c000c",  2969 => x"c3a00000",
     2970 => x"379cfff0",  2971 => x"5b8b0010",  2972 => x"5b8c000c",
     2973 => x"5b8d0008",  2974 => x"5b9d0004",  2975 => x"78040001",
     2976 => x"78050001",  2977 => x"2c2d0002",  2978 => x"b8205800",
     2979 => x"b8406000",  2980 => x"34010000",  2981 => x"34020002",
     2982 => x"34030002",  2983 => x"38842528",  2984 => x"38a53e50",
     2985 => x"fbfff97a",  2986 => x"34010040",  2987 => x"4c2d0004",
     2988 => x"b9600800",  2989 => x"b9801000",  2990 => x"f8000466",
     2991 => x"2b9d0004",  2992 => x"2b8b0010",  2993 => x"2b8c000c",
     2994 => x"2b8d0008",  2995 => x"379c0010",  2996 => x"c3a00000",
     2997 => x"379cfff8",  2998 => x"5b8b0008",  2999 => x"5b9d0004",
     3000 => x"78040001",  3001 => x"78050001",  3002 => x"34020002",
     3003 => x"34030002",  3004 => x"38842528",  3005 => x"38a53e64",
     3006 => x"b8205800",  3007 => x"fbfff964",  3008 => x"296102c8",
     3009 => x"34020040",  3010 => x"28210010",  3011 => x"40210004",
     3012 => x"44200006",  3013 => x"34030002",  3014 => x"44230004",
     3015 => x"b9600800",  3016 => x"f8000409",  3017 => x"3402004e",
     3018 => x"b8400800",  3019 => x"2b9d0004",  3020 => x"2b8b0008",
     3021 => x"379c0008",  3022 => x"c3a00000",  3023 => x"379cfff4",
     3024 => x"5b8b000c",  3025 => x"5b8c0008",  3026 => x"5b9d0004",
     3027 => x"78040001",  3028 => x"78050001",  3029 => x"34030002",
     3030 => x"b8406000",  3031 => x"38842528",  3032 => x"34020002",
     3033 => x"38a53e78",  3034 => x"b8205800",  3035 => x"fbfff948",
     3036 => x"296102c8",  3037 => x"34030000",  3038 => x"28210010",
     3039 => x"28210008",  3040 => x"44200007",  3041 => x"35630094",
     3042 => x"59800008",  3043 => x"b9600800",  3044 => x"b9801000",
     3045 => x"f80005c9",  3046 => x"34030001",  3047 => x"b8600800",
     3048 => x"2b9d0004",  3049 => x"2b8b000c",  3050 => x"2b8c0008",
     3051 => x"379c000c",  3052 => x"c3a00000",  3053 => x"379cfff8",
     3054 => x"5b8b0008",  3055 => x"5b9d0004",  3056 => x"78040001",
     3057 => x"78050001",  3058 => x"34020002",  3059 => x"34030002",
     3060 => x"38842528",  3061 => x"38a53e8c",  3062 => x"b8205800",
     3063 => x"fbfff92c",  3064 => x"296102c8",  3065 => x"28220010",
     3066 => x"40410004",  3067 => x"20210002",  3068 => x"4420000b",
     3069 => x"40410035",  3070 => x"20210001",  3071 => x"44200008",
     3072 => x"28410008",  3073 => x"44200003",  3074 => x"28410040",
     3075 => x"5c200004",  3076 => x"b9600800",  3077 => x"34020009",
     3078 => x"f80000a1",  3079 => x"2b9d0004",  3080 => x"2b8b0008",
     3081 => x"379c0008",  3082 => x"c3a00000",  3083 => x"379cffdc",
     3084 => x"5b8b0010",  3085 => x"5b8c000c",  3086 => x"5b8d0008",
     3087 => x"5b9d0004",  3088 => x"28220020",  3089 => x"78040001",
     3090 => x"78050001",  3091 => x"284d0010",  3092 => x"282202c8",
     3093 => x"34030002",  3094 => x"38842528",  3095 => x"284c0010",
     3096 => x"38a53ebc",  3097 => x"34020002",  3098 => x"b8205800",
     3099 => x"fbfff908",  3100 => x"29620318",  3101 => x"2963031c",
     3102 => x"37810014",  3103 => x"f80010b2",  3104 => x"29810008",
     3105 => x"5c200019",  3106 => x"296200a0",  3107 => x"44410003",
     3108 => x"296100b4",  3109 => x"5c200008",  3110 => x"78040001",
     3111 => x"b9600800",  3112 => x"34020004",  3113 => x"34030001",
     3114 => x"38842534",  3115 => x"fbfff8f8",  3116 => x"e0000013",
     3117 => x"b9600800",  3118 => x"f80011a4",  3119 => x"29a20004",
     3120 => x"29810000",  3121 => x"44400005",  3122 => x"28230034",
     3123 => x"34020000",  3124 => x"b9600800",  3125 => x"e0000004",
     3126 => x"28230034",  3127 => x"34020001",  3128 => x"b9600800",
     3129 => x"d8600000",  3130 => x"29620318",  3131 => x"b9600800",
     3132 => x"f800058c",  3133 => x"b9600800",  3134 => x"f80005b4",
     3135 => x"34010000",  3136 => x"2b9d0004",  3137 => x"2b8b0010",
     3138 => x"2b8c000c",  3139 => x"2b8d0008",  3140 => x"379c0024",
     3141 => x"c3a00000",  3142 => x"379cfff8",  3143 => x"5b8b0008",
     3144 => x"5b9d0004",  3145 => x"78040001",  3146 => x"78050001",
     3147 => x"34020002",  3148 => x"34030002",  3149 => x"38842528",
     3150 => x"38a53ecc",  3151 => x"b8205800",  3152 => x"fbfff8d3",
     3153 => x"b9600800",  3154 => x"f8000504",  3155 => x"34010000",
     3156 => x"2b9d0004",  3157 => x"2b8b0008",  3158 => x"379c0008",
     3159 => x"c3a00000",  3160 => x"379cffd8",  3161 => x"5b8b0010",
     3162 => x"5b8c000c",  3163 => x"5b8d0008",  3164 => x"5b9d0004",
     3165 => x"78050001",  3166 => x"b8806000",  3167 => x"78040001",
     3168 => x"b8406800",  3169 => x"34030002",  3170 => x"34020002",
     3171 => x"38842528",  3172 => x"38a53edc",  3173 => x"b8205800",
     3174 => x"fbfff8bd",  3175 => x"34010001",  3176 => x"45810004",
     3177 => x"3401000c",  3178 => x"5d810036",  3179 => x"e0000022",
     3180 => x"296200ec",  3181 => x"5960031c",  3182 => x"37810024",
     3183 => x"4802000c",  3184 => x"1443001f",  3185 => x"00440010",
     3186 => x"3c630010",  3187 => x"3c420010",  3188 => x"b8641800",
     3189 => x"5b820028",  3190 => x"340203e8",  3191 => x"5b830024",
     3192 => x"fbfffcf0",  3193 => x"2b810028",  3194 => x"e000000d",
     3195 => x"c8021000",  3196 => x"1443001f",  3197 => x"00440010",
     3198 => x"3c630010",  3199 => x"3c420010",  3200 => x"b8641800",
     3201 => x"5b820028",  3202 => x"340203e8",  3203 => x"5b830024",
     3204 => x"fbfffce4",  3205 => x"2b810028",  3206 => x"c8010800",
     3207 => x"59610318",  3208 => x"356200e4",  3209 => x"b9600800",
     3210 => x"f8000fe6",  3211 => x"340c0100",  3212 => x"e0000014",
     3213 => x"296102c8",  3214 => x"b9a01000",  3215 => x"37830014",
     3216 => x"28240010",  3217 => x"b9600800",  3218 => x"340c0100",
     3219 => x"3484003c",  3220 => x"f8000416",  3221 => x"296102c8",
     3222 => x"34021000",  3223 => x"28210010",  3224 => x"2c23003c",
     3225 => x"5c620007",  3226 => x"40210004",  3227 => x"20210001",
     3228 => x"44200004",  3229 => x"b9600800",  3230 => x"34020006",
     3231 => x"f8000008",  3232 => x"b9800800",  3233 => x"2b9d0004",
     3234 => x"2b8b0010",  3235 => x"2b8c000c",  3236 => x"2b8d0008",
     3237 => x"379c0028",  3238 => x"c3a00000",  3239 => x"282302c8",
     3240 => x"34040006",  3241 => x"28630010",  3242 => x"44440004",
     3243 => x"34040009",  3244 => x"5c440008",  3245 => x"e0000004",
     3246 => x"34020001",  3247 => x"30620005",  3248 => x"e0000007",
     3249 => x"34020002",  3250 => x"30620005",  3251 => x"e0000006",
     3252 => x"40630005",  3253 => x"34020001",  3254 => x"5c620003",
     3255 => x"34020066",  3256 => x"e0000002",  3257 => x"34020064",
     3258 => x"58220004",  3259 => x"c3a00000",  3260 => x"379cfff4",
     3261 => x"5b8b000c",  3262 => x"5b8c0008",  3263 => x"5b9d0004",
     3264 => x"b8205800",  3265 => x"282102c8",  3266 => x"78050001",
     3267 => x"38a52484",  3268 => x"282c0010",  3269 => x"34010001",
     3270 => x"41820005",  3271 => x"5c410003",  3272 => x"78050001",
     3273 => x"38a5296c",  3274 => x"78040001",  3275 => x"b9600800",
     3276 => x"34020002",  3277 => x"34030001",  3278 => x"3884255c",
     3279 => x"fbfff854",  3280 => x"41820005",  3281 => x"34010001",
     3282 => x"5c410003",  3283 => x"34010006",  3284 => x"e0000002",
     3285 => x"34010009",  3286 => x"59610004",  3287 => x"31800005",
     3288 => x"2b9d0004",  3289 => x"2b8b000c",  3290 => x"2b8c0008",
     3291 => x"379c000c",  3292 => x"c3a00000",  3293 => x"379cfffc",
     3294 => x"5b9d0004",  3295 => x"282202c8",  3296 => x"28420010",
     3297 => x"4043002c",  3298 => x"4460000a",  3299 => x"3463ffff",
     3300 => x"78040001",  3301 => x"3043002c",  3302 => x"38842580",
     3303 => x"34020002",  3304 => x"34030001",  3305 => x"fbfff83a",
     3306 => x"34010001",  3307 => x"e0000003",  3308 => x"fbffffd0",
     3309 => x"34010000",  3310 => x"2b9d0004",  3311 => x"379c0004",
     3312 => x"c3a00000",  3313 => x"379cffd8",  3314 => x"5b8b0018",
     3315 => x"5b8c0014",  3316 => x"5b8d0010",  3317 => x"5b8e000c",
     3318 => x"5b8f0008",  3319 => x"5b9d0004",  3320 => x"b8407000",
     3321 => x"2824000c",  3322 => x"282202c8",  3323 => x"b8205800",
     3324 => x"b8607800",  3325 => x"284d0010",  3326 => x"44800004",
     3327 => x"34010003",  3328 => x"31a1002c",  3329 => x"e000000c",
     3330 => x"282202e0",  3331 => x"44440008",  3332 => x"28220028",
     3333 => x"28440018",  3334 => x"34020000",  3335 => x"d8800000",
     3336 => x"296202e0",  3337 => x"c8220800",  3338 => x"4c20003c",
     3339 => x"340c0000",  3340 => x"e0000015",  3341 => x"29610028",
     3342 => x"340203e8",  3343 => x"28240018",  3344 => x"b9600800",
     3345 => x"d8800000",  3346 => x"596102e0",  3347 => x"296102c8",
     3348 => x"29620028",  3349 => x"4025000c",  3350 => x"1021000b",
     3351 => x"28440018",  3352 => x"bca12800",  3353 => x"b9600800",
     3354 => x"08a203e8",  3355 => x"d8800000",  3356 => x"596102d4",
     3357 => x"34021000",  3358 => x"b9600800",  3359 => x"f80003fb",
     3360 => x"b8206000",  3361 => x"45e0000e",  3362 => x"4162030d",
     3363 => x"3401000c",  3364 => x"5c41000b",  3365 => x"b9600800",
     3366 => x"b9c01000",  3367 => x"3783001c",  3368 => x"35a4003c",
     3369 => x"f8000381",  3370 => x"2da2003c",  3371 => x"34011001",
     3372 => x"5c410003",  3373 => x"34010065",  3374 => x"59610004",
     3375 => x"5d800004",  3376 => x"b9600800",  3377 => x"f8000aae",
     3378 => x"e0000003",  3379 => x"34010002",  3380 => x"59610004",
     3381 => x"29620004",  3382 => x"29610000",  3383 => x"44410002",
     3384 => x"596002d4",  3385 => x"296102c8",  3386 => x"28210010",
     3387 => x"28210028",  3388 => x"59610008",  3389 => x"b9800800",
     3390 => x"2b9d0004",  3391 => x"2b8b0018",  3392 => x"2b8c0014",
     3393 => x"2b8d0010",  3394 => x"2b8e000c",  3395 => x"2b8f0008",
     3396 => x"379c0028",  3397 => x"c3a00000",  3398 => x"b9600800",
     3399 => x"34020005",  3400 => x"f800124e",  3401 => x"b9600800",
     3402 => x"596002e0",  3403 => x"fbffff92",  3404 => x"340c0000",
     3405 => x"5c20ffc0",  3406 => x"e3ffffef",  3407 => x"379cffd8",
     3408 => x"5b8b0018",  3409 => x"5b8c0014",  3410 => x"5b8d0010",
     3411 => x"5b8e000c",  3412 => x"5b8f0008",  3413 => x"5b9d0004",
     3414 => x"b8407000",  3415 => x"2824000c",  3416 => x"282202c8",
     3417 => x"b8205800",  3418 => x"b8607800",  3419 => x"284c0010",
     3420 => x"44800004",  3421 => x"34010003",  3422 => x"3181002c",
     3423 => x"e000000c",  3424 => x"282202e0",  3425 => x"44440008",
     3426 => x"28220028",  3427 => x"28440018",  3428 => x"34020000",
     3429 => x"d8800000",  3430 => x"296202e0",  3431 => x"c8220800",
     3432 => x"4c200029",  3433 => x"340d0000",  3434 => x"e000000b",
     3435 => x"34021001",  3436 => x"b9600800",  3437 => x"f80003ad",
     3438 => x"b8206800",  3439 => x"29610028",  3440 => x"34023a98",
     3441 => x"28240018",  3442 => x"b9600800",  3443 => x"d8800000",
     3444 => x"596102e0",  3445 => x"45e0000e",  3446 => x"4162030d",
     3447 => x"3401000c",  3448 => x"5c41000b",  3449 => x"b9600800",
     3450 => x"b9c01000",  3451 => x"3783001c",  3452 => x"3584003c",
     3453 => x"f800032d",  3454 => x"2d82003c",  3455 => x"34011002",
     3456 => x"5c410003",  3457 => x"34010068",  3458 => x"59610004",
     3459 => x"45a00003",  3460 => x"34010002",  3461 => x"59610004",
     3462 => x"29810028",  3463 => x"59610008",  3464 => x"b9a00800",
     3465 => x"2b9d0004",  3466 => x"2b8b0018",  3467 => x"2b8c0014",
     3468 => x"2b8d0010",  3469 => x"2b8e000c",  3470 => x"2b8f0008",
     3471 => x"379c0028",  3472 => x"c3a00000",  3473 => x"b9600800",
     3474 => x"34020005",  3475 => x"f8001203",  3476 => x"b9600800",
     3477 => x"596002e0",  3478 => x"fbffff47",  3479 => x"340d0000",
     3480 => x"5c20ffd3",  3481 => x"e3ffffef",  3482 => x"379cfff4",
     3483 => x"5b8b000c",  3484 => x"5b8c0008",  3485 => x"5b9d0004",
     3486 => x"282202c8",  3487 => x"b8205800",  3488 => x"284c0010",
     3489 => x"2822000c",  3490 => x"44400004",  3491 => x"34010003",
     3492 => x"3181002c",  3493 => x"e000000b",  3494 => x"282302e0",
     3495 => x"44620013",  3496 => x"28220028",  3497 => x"28430018",
     3498 => x"34020000",  3499 => x"d8600000",  3500 => x"296202e0",
     3501 => x"c8220800",  3502 => x"4c200021",  3503 => x"e000000b",
     3504 => x"29810000",  3505 => x"28220000",  3506 => x"b9600800",
     3507 => x"d8400000",  3508 => x"29610028",  3509 => x"34023a98",
     3510 => x"28230018",  3511 => x"b9600800",  3512 => x"d8600000",
     3513 => x"596102e0",  3514 => x"29810000",  3515 => x"34020000",
     3516 => x"28230004",  3517 => x"b9600800",  3518 => x"d8600000",
     3519 => x"34020001",  3520 => x"5c220007",  3521 => x"34010067",
     3522 => x"59610004",  3523 => x"29810000",  3524 => x"28220008",
     3525 => x"b9600800",  3526 => x"d8400000",  3527 => x"29810028",
     3528 => x"59610008",  3529 => x"34010000",  3530 => x"2b9d0004",
     3531 => x"2b8b000c",  3532 => x"2b8c0008",  3533 => x"379c000c",
     3534 => x"c3a00000",  3535 => x"b9600800",  3536 => x"34020005",
     3537 => x"f80011c5",  3538 => x"29810000",  3539 => x"596002e0",
     3540 => x"28220008",  3541 => x"b9600800",  3542 => x"d8400000",
     3543 => x"b9600800",  3544 => x"fbffff05",  3545 => x"5c20ffd7",
     3546 => x"e3ffffef",  3547 => x"379cffd8",  3548 => x"5b8b0018",
     3549 => x"5b8c0014",  3550 => x"5b8d0010",  3551 => x"5b8e000c",
     3552 => x"5b8f0008",  3553 => x"5b9d0004",  3554 => x"b8407000",
     3555 => x"2824000c",  3556 => x"282202c8",  3557 => x"b8205800",
     3558 => x"b8607800",  3559 => x"284c0010",  3560 => x"44800004",
     3561 => x"34010003",  3562 => x"3181002c",  3563 => x"e000000c",
     3564 => x"282202e0",  3565 => x"44440008",  3566 => x"28220028",
     3567 => x"28440018",  3568 => x"34020000",  3569 => x"d8800000",
     3570 => x"296202e0",  3571 => x"c8220800",  3572 => x"4c200029",
     3573 => x"340d0000",  3574 => x"e000000b",  3575 => x"29610028",
     3576 => x"29820028",  3577 => x"28240018",  3578 => x"b9600800",
     3579 => x"d8800000",  3580 => x"596102e0",  3581 => x"34021002",
     3582 => x"b9600800",  3583 => x"f800031b",  3584 => x"b8206800",
     3585 => x"45e0000e",  3586 => x"4162030d",  3587 => x"3401000c",
     3588 => x"5c41000b",  3589 => x"b9600800",  3590 => x"b9c01000",
     3591 => x"3783001c",  3592 => x"3584003c",  3593 => x"f80002a1",
     3594 => x"2d82003c",  3595 => x"34011003",  3596 => x"5c410003",
     3597 => x"3401006a",  3598 => x"59610004",  3599 => x"45a00003",
     3600 => x"34010002",  3601 => x"59610004",  3602 => x"29810028",
     3603 => x"59610008",  3604 => x"b9a00800",  3605 => x"2b9d0004",
     3606 => x"2b8b0018",  3607 => x"2b8c0014",  3608 => x"2b8d0010",
     3609 => x"2b8e000c",  3610 => x"2b8f0008",  3611 => x"379c0028",
     3612 => x"c3a00000",  3613 => x"b9600800",  3614 => x"34020005",
     3615 => x"f8001177",  3616 => x"b9600800",  3617 => x"596002e0",
     3618 => x"fbfffebb",  3619 => x"340d0000",  3620 => x"5c20ffd3",
     3621 => x"e3ffffef",  3622 => x"379cffec",  3623 => x"5b8b0010",
     3624 => x"5b8c000c",  3625 => x"5b8d0008",  3626 => x"5b9d0004",
     3627 => x"282202c8",  3628 => x"b8206000",  3629 => x"284b0010",
     3630 => x"2822000c",  3631 => x"44400004",  3632 => x"34010003",
     3633 => x"3161002c",  3634 => x"e000000c",  3635 => x"282302e0",
     3636 => x"44620008",  3637 => x"28220028",  3638 => x"28430018",
     3639 => x"34020000",  3640 => x"d8600000",  3641 => x"298202e0",
     3642 => x"c8220800",  3643 => x"4c2000a9",  3644 => x"340d0000",
     3645 => x"e0000011",  3646 => x"29810028",  3647 => x"29620030",
     3648 => x"28230018",  3649 => x"b9800800",  3650 => x"d8600000",
     3651 => x"598102e0",  3652 => x"34021003",  3653 => x"b9800800",
     3654 => x"f80002d4",  3655 => x"b8206800",  3656 => x"3401006c",
     3657 => x"31610010",  3658 => x"29610014",  3659 => x"44200003",
     3660 => x"3401006e",  3661 => x"31610010",  3662 => x"41660010",
     3663 => x"78040001",  3664 => x"78050001",  3665 => x"b9800800",
     3666 => x"34020002",  3667 => x"34030001",  3668 => x"38842594",
     3669 => x"38a53f30",  3670 => x"34c6ff94",  3671 => x"fbfff6cc",
     3672 => x"41620010",  3673 => x"34010008",  3674 => x"3442ff94",
     3675 => x"204200ff",  3676 => x"5441007f",  3677 => x"78010001",
     3678 => x"3c420002",  3679 => x"38213f0c",  3680 => x"b4220800",
     3681 => x"28210000",  3682 => x"c0200000",  3683 => x"29610000",
     3684 => x"34020000",  3685 => x"34030000",  3686 => x"2825002c",
     3687 => x"34040000",  3688 => x"b9800800",  3689 => x"d8a00000",
     3690 => x"5c200071",  3691 => x"3401006d",  3692 => x"31610010",
     3693 => x"29610000",  3694 => x"34020001",  3695 => x"28230024",
     3696 => x"b9800800",  3697 => x"d8600000",  3698 => x"5c200069",
     3699 => x"3401006e",  3700 => x"31610010",  3701 => x"29610000",
     3702 => x"34020001",  3703 => x"37830014",  3704 => x"28240028",
     3705 => x"b9800800",  3706 => x"d8800000",  3707 => x"34020001",
     3708 => x"5c22005f",  3709 => x"2b810014",  3710 => x"78040001",
     3711 => x"34020002",  3712 => x"00250010",  3713 => x"3c210010",
     3714 => x"5965001c",  3715 => x"59610018",  3716 => x"34030001",
     3717 => x"b9800800",  3718 => x"388425a8",  3719 => x"fbfff69c",
     3720 => x"29650018",  3721 => x"78040001",  3722 => x"b9800800",
     3723 => x"34020002",  3724 => x"34030001",  3725 => x"388425cc",
     3726 => x"fbfff695",  3727 => x"3401006f",  3728 => x"31610010",
     3729 => x"29610000",  3730 => x"34020001",  3731 => x"28230020",
     3732 => x"b9800800",  3733 => x"d8600000",  3734 => x"5c200045",
     3735 => x"34010070",  3736 => x"31610010",  3737 => x"29610000",
     3738 => x"28220030",  3739 => x"b9800800",  3740 => x"d8400000",
     3741 => x"5c20003e",  3742 => x"34010071",  3743 => x"31610010",
     3744 => x"29610000",  3745 => x"34020002",  3746 => x"28230024",
     3747 => x"b9800800",  3748 => x"d8600000",  3749 => x"5c200036",
     3750 => x"34010072",  3751 => x"31610010",  3752 => x"29610000",
     3753 => x"34020002",  3754 => x"37830014",  3755 => x"28240028",
     3756 => x"b9800800",  3757 => x"d8800000",  3758 => x"34020001",
     3759 => x"5c22002c",  3760 => x"2b850014",  3761 => x"78040001",
     3762 => x"b9800800",  3763 => x"34020002",  3764 => x"34030001",
     3765 => x"388425f0",  3766 => x"fbfff66d",  3767 => x"2b810014",
     3768 => x"78040001",  3769 => x"34020002",  3770 => x"00250010",
     3771 => x"3c210010",  3772 => x"59650024",  3773 => x"59610020",
     3774 => x"34030001",  3775 => x"b9800800",  3776 => x"38842608",
     3777 => x"fbfff662",  3778 => x"29650020",  3779 => x"78040001",
     3780 => x"b9800800",  3781 => x"34020002",  3782 => x"34030001",
     3783 => x"3884262c",  3784 => x"fbfff65b",  3785 => x"34010073",
     3786 => x"31610010",  3787 => x"29610000",  3788 => x"34020002",
     3789 => x"28230020",  3790 => x"b9800800",  3791 => x"d8600000",
     3792 => x"5c20000b",  3793 => x"34010074",  3794 => x"31610010",
     3795 => x"b9800800",  3796 => x"34021004",  3797 => x"f8000245",
     3798 => x"b8206800",  3799 => x"34010069",  3800 => x"59810004",
     3801 => x"34010001",  3802 => x"59610014",  3803 => x"29610028",
     3804 => x"59810008",  3805 => x"b9a00800",  3806 => x"2b9d0004",
     3807 => x"2b8b0010",  3808 => x"2b8c000c",  3809 => x"2b8d0008",
     3810 => x"379c0014",  3811 => x"c3a00000",  3812 => x"b9800800",
     3813 => x"34020005",  3814 => x"f80010b0",  3815 => x"b9800800",
     3816 => x"598002e0",  3817 => x"fbfffdf4",  3818 => x"340d0000",
     3819 => x"5c20ff53",  3820 => x"e3fffff1",  3821 => x"379cffdc",
     3822 => x"5b8b0014",  3823 => x"5b8c0010",  3824 => x"5b8d000c",
     3825 => x"5b8e0008",  3826 => x"5b9d0004",  3827 => x"b8406800",
     3828 => x"282202c8",  3829 => x"b8205800",  3830 => x"b8607000",
     3831 => x"284c0010",  3832 => x"2822000c",  3833 => x"44400006",
     3834 => x"28220028",  3835 => x"28440018",  3836 => x"29820028",
     3837 => x"d8800000",  3838 => x"596102e0",  3839 => x"296102e0",
     3840 => x"44200009",  3841 => x"29610028",  3842 => x"34020000",
     3843 => x"28240018",  3844 => x"b9600800",  3845 => x"d8800000",
     3846 => x"296202e0",  3847 => x"c8220800",  3848 => x"4c200023",
     3849 => x"45c00018",  3850 => x"4162030d",  3851 => x"3401000c",
     3852 => x"5c410015",  3853 => x"b9600800",  3854 => x"b9a01000",
     3855 => x"37830018",  3856 => x"3584003c",  3857 => x"f8000199",
     3858 => x"2d81003c",  3859 => x"34021003",  3860 => x"5c220006",
     3861 => x"41820005",  3862 => x"34010001",  3863 => x"5c41000a",
     3864 => x"3401006a",  3865 => x"e0000007",  3866 => x"34021005",
     3867 => x"5c220006",  3868 => x"41820005",  3869 => x"34010002",
     3870 => x"5c410003",  3871 => x"3401006b",  3872 => x"59610004",
     3873 => x"29810028",  3874 => x"59610008",  3875 => x"34010000",
     3876 => x"2b9d0004",  3877 => x"2b8b0014",  3878 => x"2b8c0010",
     3879 => x"2b8d000c",  3880 => x"2b8e0008",  3881 => x"379c0024",
     3882 => x"c3a00000",  3883 => x"b9600800",  3884 => x"34020005",
     3885 => x"f8001069",  3886 => x"b9600800",  3887 => x"596002e0",
     3888 => x"fbfffd8c",  3889 => x"e3fffff2",  3890 => x"379cffd4",
     3891 => x"5b8b001c",  3892 => x"5b8c0018",  3893 => x"5b8d0014",
     3894 => x"5b8e0010",  3895 => x"5b8f000c",  3896 => x"5b900008",
     3897 => x"5b9d0004",  3898 => x"b8407000",  3899 => x"282202c8",
     3900 => x"2824000c",  3901 => x"b8205800",  3902 => x"284c0010",
     3903 => x"b8607800",  3904 => x"2d8d0048",  3905 => x"7dad0000",
     3906 => x"44800004",  3907 => x"34010003",  3908 => x"3181002c",
     3909 => x"e0000012",  3910 => x"282202e0",  3911 => x"44440022",
     3912 => x"28220028",  3913 => x"28440018",  3914 => x"34020000",
     3915 => x"d8800000",  3916 => x"296202e0",  3917 => x"c8220800",
     3918 => x"4c20003f",  3919 => x"e000001a",  3920 => x"29810000",
     3921 => x"28240030",  3922 => x"b9600800",  3923 => x"d8800000",
     3924 => x"b9600800",  3925 => x"fbfffd88",  3926 => x"4420002d",
     3927 => x"45a00008",  3928 => x"29810000",  3929 => x"34020000",
     3930 => x"34030000",  3931 => x"2825002c",  3932 => x"34040000",
     3933 => x"b9600800",  3934 => x"d8a00000",  3935 => x"2981004c",
     3936 => x"29700028",  3937 => x"340203e8",  3938 => x"f800348f",
     3939 => x"2a050018",  3940 => x"b8202000",  3941 => x"b8801000",
     3942 => x"b9600800",  3943 => x"d8a00000",  3944 => x"596102e0",
     3945 => x"45e00018",  3946 => x"4162030d",  3947 => x"3401000c",
     3948 => x"5c410015",  3949 => x"b9600800",  3950 => x"b9c01000",
     3951 => x"37830020",  3952 => x"3584003c",  3953 => x"f8000139",
     3954 => x"2d82003c",  3955 => x"34011004",  3956 => x"5c41000d",
     3957 => x"45a00005",  3958 => x"29810000",  3959 => x"28220030",
     3960 => x"b9600800",  3961 => x"d8400000",  3962 => x"41820005",
     3963 => x"34010001",  3964 => x"5c410003",  3965 => x"3401006b",
     3966 => x"e0000002",  3967 => x"34010068",  3968 => x"59610004",
     3969 => x"29810028",  3970 => x"59610008",  3971 => x"34010000",
     3972 => x"2b9d0004",  3973 => x"2b8b001c",  3974 => x"2b8c0018",
     3975 => x"2b8d0014",  3976 => x"2b8e0010",  3977 => x"2b8f000c",
     3978 => x"2b900008",  3979 => x"379c002c",  3980 => x"c3a00000",
     3981 => x"b9600800",  3982 => x"34020005",  3983 => x"f8001007",
     3984 => x"596002e0",  3985 => x"45a0ffc3",  3986 => x"e3ffffbe",
     3987 => x"379cfff0",  3988 => x"5b8b0010",  3989 => x"5b8c000c",
     3990 => x"5b8d0008",  3991 => x"5b9d0004",  3992 => x"282202c8",
     3993 => x"340d0001",  3994 => x"b8206000",  3995 => x"284b0010",
     3996 => x"29620000",  3997 => x"596d0008",  3998 => x"2842000c",
     3999 => x"d8400000",  4000 => x"41610005",  4001 => x"34020000",
     4002 => x"5c2d0005",  4003 => x"34021005",  4004 => x"b9800800",
     4005 => x"f8000175",  4006 => x"b8201000",  4007 => x"34010001",
     4008 => x"59610040",  4009 => x"3401ffff",  4010 => x"5c400009",
     4011 => x"41620005",  4012 => x"34010002",  4013 => x"5c410003",
     4014 => x"34010009",  4015 => x"e0000002",  4016 => x"34010006",
     4017 => x"59810004",  4018 => x"34010000",  4019 => x"2b9d0004",
     4020 => x"2b8b0010",  4021 => x"2b8c000c",  4022 => x"2b8d0008",
     4023 => x"379c0010",  4024 => x"c3a00000",  4025 => x"00430018",
     4026 => x"30220003",  4027 => x"30230000",  4028 => x"00430010",
     4029 => x"30230001",  4030 => x"00430008",  4031 => x"30230002",
     4032 => x"c3a00000",  4033 => x"40220000",  4034 => x"40230003",
     4035 => x"3c420018",  4036 => x"b8621000",  4037 => x"40230001",
     4038 => x"40210002",  4039 => x"3c630010",  4040 => x"3c210008",
     4041 => x"b8431000",  4042 => x"b8410800",  4043 => x"c3a00000",
     4044 => x"40220000",  4045 => x"40210001",  4046 => x"3c420008",
     4047 => x"b8410800",  4048 => x"c3a00000",  4049 => x"379cfff0",
     4050 => x"5b8b0010",  4051 => x"5b8c000c",  4052 => x"5b8d0008",
     4053 => x"5b9d0004",  4054 => x"28230020",  4055 => x"282202c8",
     4056 => x"b8205800",  4057 => x"2863000c",  4058 => x"28420010",
     4059 => x"282c003c",  4060 => x"4064000e",  4061 => x"340300ba",
     4062 => x"48830018",  4063 => x"28420000",  4064 => x"28430004",
     4065 => x"34020001",  4066 => x"d8600000",  4067 => x"ec016800",
     4068 => x"b9600800",  4069 => x"f8000967",  4070 => x"29610020",
     4071 => x"c80d6800",  4072 => x"21ad002e",  4073 => x"2821000c",
     4074 => x"35ad0006",  4075 => x"4021000e",  4076 => x"45a1000a",
     4077 => x"78010001",  4078 => x"b9a01000",  4079 => x"38212650",
     4080 => x"f8001b81",  4081 => x"29610020",  4082 => x"21ad00ff",
     4083 => x"2821000c",  4084 => x"302d000e",  4085 => x"318d0030",
     4086 => x"3401004e",  4087 => x"0d810002",  4088 => x"34010003",
     4089 => x"0d810040",  4090 => x"3401000a",  4091 => x"0d810042",
     4092 => x"34010800",  4093 => x"0d810044",  4094 => x"340130de",
     4095 => x"0d810046",  4096 => x"3401ad01",  4097 => x"0d810048",
     4098 => x"34012000",  4099 => x"0d81004a",  4100 => x"296102c8",
     4101 => x"28220010",  4102 => x"28430014",  4103 => x"40410004",
     4104 => x"44600002",  4105 => x"38210004",  4106 => x"28420008",
     4107 => x"44400002",  4108 => x"38210008",  4109 => x"0d81004c",
     4110 => x"2b9d0004",  4111 => x"2b8b0010",  4112 => x"2b8c000c",
     4113 => x"2b8d0008",  4114 => x"379c0010",  4115 => x"c3a00000",
     4116 => x"379cfff4",  4117 => x"5b8b000c",  4118 => x"5b8c0008",
     4119 => x"5b9d0004",  4120 => x"b8205800",  4121 => x"34210040",
     4122 => x"b8406000",  4123 => x"fbffffb1",  4124 => x"2d650044",
     4125 => x"2d640046",  4126 => x"78070001",  4127 => x"3ca50008",
     4128 => x"00860008",  4129 => x"38e73ce8",  4130 => x"b8a62800",
     4131 => x"28e60000",  4132 => x"64210003",  4133 => x"2d630048",
     4134 => x"e4a62800",  4135 => x"2d62004a",  4136 => x"a0250800",
     4137 => x"44200010",  4138 => x"3c840008",  4139 => x"00610008",
     4140 => x"2084ffff",  4141 => x"b8812000",  4142 => x"206300ff",
     4143 => x"3801dead",  4144 => x"e4812000",  4145 => x"64630001",
     4146 => x"a0831800",  4147 => x"44600006",  4148 => x"34012000",
     4149 => x"5c410004",  4150 => x"3561004c",  4151 => x"fbffff95",
     4152 => x"59810024",  4153 => x"2b9d0004",  4154 => x"2b8b000c",
     4155 => x"2b8c0008",  4156 => x"379c000c",  4157 => x"c3a00000",
     4158 => x"379cfff0",  4159 => x"5b8b0010",  4160 => x"5b8c000c",
     4161 => x"5b8d0008",  4162 => x"5b9d0004",  4163 => x"b8206000",
     4164 => x"282102c8",  4165 => x"204dffff",  4166 => x"28210010",
     4167 => x"40250005",  4168 => x"44a00003",  4169 => x"34012000",
     4170 => x"5da1000a",  4171 => x"78040001",  4172 => x"b9800800",
     4173 => x"34020005",  4174 => x"34030001",  4175 => x"38842668",
     4176 => x"b9a03000",  4177 => x"fbfff4d2",  4178 => x"34010000",
     4179 => x"e0000051",  4180 => x"298b003c",  4181 => x"34030008",
     4182 => x"41610000",  4183 => x"202100f0",  4184 => x"3821000c",
     4185 => x"31610000",  4186 => x"34010005",  4187 => x"31610020",
     4188 => x"29820020",  4189 => x"35610022",  4190 => x"28420014",
     4191 => x"f80033f3",  4192 => x"29810020",  4193 => x"28210014",
     4194 => x"2c210008",  4195 => x"0d6d0036",  4196 => x"00220008",
     4197 => x"3161002b",  4198 => x"34010003",  4199 => x"0d61002c",
     4200 => x"34010800",  4201 => x"0d610030",  4202 => x"340130de",
     4203 => x"0d610032",  4204 => x"3401ad01",  4205 => x"0d610034",
     4206 => x"3162002a",  4207 => x"34011003",  4208 => x"45a10005",
     4209 => x"34011004",  4210 => x"34020008",  4211 => x"5da1002d",
     4212 => x"e0000017",  4213 => x"298102c8",  4214 => x"35620038",
     4215 => x"28210010",  4216 => x"28230014",  4217 => x"44600005",
     4218 => x"40210034",  4219 => x"31610038",  4220 => x"30400001",
     4221 => x"e0000007",  4222 => x"40210034",  4223 => x"3c210008",
     4224 => x"38210001",  4225 => x"00230008",  4226 => x"31630038",
     4227 => x"30410001",  4228 => x"298102c8",  4229 => x"28220010",
     4230 => x"3561003a",  4231 => x"28420030",  4232 => x"fbffff31",
     4233 => x"34020014",  4234 => x"e0000016",  4235 => x"298102c8",
     4236 => x"28220010",  4237 => x"35610038",  4238 => x"2842001c",
     4239 => x"fbffff2a",  4240 => x"298102c8",  4241 => x"28220010",
     4242 => x"3561003c",  4243 => x"28420018",  4244 => x"fbffff25",
     4245 => x"298102c8",  4246 => x"28220010",  4247 => x"35610040",
     4248 => x"28420024",  4249 => x"fbffff20",  4250 => x"298102c8",
     4251 => x"28220010",  4252 => x"35610044",  4253 => x"28420020",
     4254 => x"fbffff1b",  4255 => x"34020018",  4256 => x"34410030",
     4257 => x"31600002",  4258 => x"31610003",  4259 => x"0d62002e",
     4260 => x"2b9d0004",  4261 => x"2b8b0010",  4262 => x"2b8c000c",
     4263 => x"2b8d0008",  4264 => x"379c0010",  4265 => x"c3a00000",
     4266 => x"379cffec",  4267 => x"5b8b0014",  4268 => x"5b8c0010",
     4269 => x"5b8d000c",  4270 => x"5b8e0008",  4271 => x"5b9d0004",
     4272 => x"b8405800",  4273 => x"b8607000",  4274 => x"34420022",
     4275 => x"b8206000",  4276 => x"b8600800",  4277 => x"34030008",
     4278 => x"b8806800",  4279 => x"f800339b",  4280 => x"3561002a",
     4281 => x"fbffff13",  4282 => x"0dc10008",  4283 => x"3561002c",
     4284 => x"fbffff10",  4285 => x"b8202800",  4286 => x"34040003",
     4287 => x"2d630030",  4288 => x"2d620032",  4289 => x"2d610034",
     4290 => x"44a40007",  4291 => x"78040001",  4292 => x"b9800800",
     4293 => x"34020005",  4294 => x"34030001",  4295 => x"3884269c",
     4296 => x"e0000022",  4297 => x"3c650008",  4298 => x"78040001",
     4299 => x"00430008",  4300 => x"38843ce8",  4301 => x"b8a32800",
     4302 => x"28830000",  4303 => x"44a30007",  4304 => x"78040001",
     4305 => x"b9800800",  4306 => x"34020005",  4307 => x"34030001",
     4308 => x"388426ec",  4309 => x"e0000015",  4310 => x"3c450008",
     4311 => x"00230008",  4312 => x"20a5ffff",  4313 => x"b8a32800",
     4314 => x"3802dead",  4315 => x"44a20007",  4316 => x"78040001",
     4317 => x"b9800800",  4318 => x"34020005",  4319 => x"34030001",
     4320 => x"38842724",  4321 => x"e0000009",  4322 => x"202500ff",
     4323 => x"34010001",  4324 => x"44a10008",  4325 => x"78040001",
     4326 => x"b9800800",  4327 => x"34020005",  4328 => x"34030001",
     4329 => x"38842768",  4330 => x"fbfff439",  4331 => x"e0000028",
     4332 => x"2d610036",  4333 => x"45a00002",  4334 => x"0da10000",
     4335 => x"34021003",  4336 => x"44220004",  4337 => x"34021004",
     4338 => x"5c220021",  4339 => x"e0000012",  4340 => x"298102c8",
     4341 => x"356e0038",  4342 => x"282d0010",  4343 => x"b9c00800",
     4344 => x"fbfffed4",  4345 => x"202100ff",  4346 => x"0da10048",
     4347 => x"b9c00800",  4348 => x"fbfffed0",  4349 => x"00210008",
     4350 => x"31a10050",  4351 => x"3561003a",  4352 => x"fbfffec1",
     4353 => x"298202c8",  4354 => x"28420010",  4355 => x"5841004c",
     4356 => x"e000000f",  4357 => x"298102c8",  4358 => x"282c0010",
     4359 => x"35610038",  4360 => x"fbfffeb9",  4361 => x"59810058",
     4362 => x"3561003c",  4363 => x"fbfffeb6",  4364 => x"59810054",
     4365 => x"35610040",  4366 => x"fbfffeb3",  4367 => x"59810060",
     4368 => x"35610044",  4369 => x"fbfffeb0",  4370 => x"5981005c",
     4371 => x"2b9d0004",  4372 => x"2b8b0014",  4373 => x"2b8c0010",
     4374 => x"2b8d000c",  4375 => x"2b8e0008",  4376 => x"379c0014",
     4377 => x"c3a00000",  4378 => x"379cfff4",  4379 => x"5b8b000c",
     4380 => x"5b8c0008",  4381 => x"5b9d0004",  4382 => x"2042ffff",
     4383 => x"b8205800",  4384 => x"fbffff1e",  4385 => x"b8206000",
     4386 => x"29610024",  4387 => x"29630070",  4388 => x"29620034",
     4389 => x"2827000c",  4390 => x"b5831800",  4391 => x"b9600800",
     4392 => x"356400f8",  4393 => x"34050000",  4394 => x"34060000",
     4395 => x"d8e00000",  4396 => x"78080001",  4397 => x"39084a14",
     4398 => x"4c2c000b",  4399 => x"29050030",  4400 => x"78040001",
     4401 => x"b9600800",  4402 => x"34020005",  4403 => x"34030001",
     4404 => x"388427ac",  4405 => x"3406000c",  4406 => x"fbfff3ed",
     4407 => x"3401ffff",  4408 => x"e000000f",  4409 => x"296600f8",
     4410 => x"296700fc",  4411 => x"29080030",  4412 => x"78040001",
     4413 => x"b9600800",  4414 => x"34020005",  4415 => x"34030001",
     4416 => x"388427cc",  4417 => x"b9802800",  4418 => x"fbfff3e1",
     4419 => x"2961036c",  4420 => x"34210001",  4421 => x"5961036c",
     4422 => x"34010000",  4423 => x"2b9d0004",  4424 => x"2b8b000c",
     4425 => x"2b8c0008",  4426 => x"379c000c",  4427 => x"c3a00000",
     4428 => x"78020001",  4429 => x"38424a10",  4430 => x"58410000",
     4431 => x"c3a00000",  4432 => x"78010001",  4433 => x"38215210",
     4434 => x"28210000",  4435 => x"44200002",  4436 => x"58200010",
     4437 => x"c3a00000",  4438 => x"379cffec",  4439 => x"5b8b0014",
     4440 => x"5b8c0010",  4441 => x"5b8d000c",  4442 => x"5b8e0008",
     4443 => x"5b9d0004",  4444 => x"b8206800",  4445 => x"282102c8",
     4446 => x"780e0001",  4447 => x"39ce6db4",  4448 => x"282c0010",
     4449 => x"29c10000",  4450 => x"34020001",  4451 => x"29ab0014",
     4452 => x"fbfff30d",  4453 => x"29810000",  4454 => x"34020000",
     4455 => x"34030000",  4456 => x"2826001c",  4457 => x"35640028",
     4458 => x"b9a00800",  4459 => x"3565002c",  4460 => x"d8c00000",
     4461 => x"3402ffff",  4462 => x"5c200038",  4463 => x"29810000",
     4464 => x"34020000",  4465 => x"28230034",  4466 => x"b9a00800",
     4467 => x"d8600000",  4468 => x"34030010",  4469 => x"35a20358",
     4470 => x"b9600800",  4471 => x"f800345b",  4472 => x"29810000",
     4473 => x"596000a8",  4474 => x"28220018",  4475 => x"34010000",
     4476 => x"d8400000",  4477 => x"34010002",  4478 => x"59610014",
     4479 => x"29810058",  4480 => x"2d820054",  4481 => x"59600088",
     4482 => x"3c210010",  4483 => x"b8220800",  4484 => x"59610018",
     4485 => x"29810060",  4486 => x"2d82005c",  4487 => x"3c210010",
     4488 => x"b8220800",  4489 => x"5961001c",  4490 => x"2981001c",
     4491 => x"2d820018",  4492 => x"3c210010",  4493 => x"b8220800",
     4494 => x"59610020",  4495 => x"29810024",  4496 => x"2d820020",
     4497 => x"3c210010",  4498 => x"b8220800",  4499 => x"78020001",
     4500 => x"59610024",  4501 => x"384227f0",  4502 => x"356100c0",
     4503 => x"f800339b",  4504 => x"78010001",  4505 => x"38215210",
     4506 => x"582b0000",  4507 => x"29610010",  4508 => x"34020000",
     4509 => x"596000b8",  4510 => x"38210001",  4511 => x"59610010",
     4512 => x"78010001",  4513 => x"38215208",  4514 => x"58200000",
     4515 => x"29c10000",  4516 => x"fbfff2cd",  4517 => x"34020000",
     4518 => x"b8400800",  4519 => x"2b9d0004",  4520 => x"2b8b0014",
     4521 => x"2b8c0010",  4522 => x"2b8d000c",  4523 => x"2b8e0008",
     4524 => x"379c0014",  4525 => x"c3a00000",  4526 => x"28460000",
     4527 => x"28450004",  4528 => x"28440008",  4529 => x"28210014",
     4530 => x"28420010",  4531 => x"58260030",  4532 => x"58220040",
     4533 => x"34020001",  4534 => x"58250034",  4535 => x"58240038",
     4536 => x"5822003c",  4537 => x"28670000",  4538 => x"28660004",
     4539 => x"28650008",  4540 => x"2864000c",  4541 => x"28630010",
     4542 => x"58270044",  4543 => x"58260048",  4544 => x"5825004c",
     4545 => x"58240050",  4546 => x"58230054",  4547 => x"78010001",
     4548 => x"38215208",  4549 => x"58220000",  4550 => x"34010000",
     4551 => x"c3a00000",  4552 => x"379cfff8",  4553 => x"5b8b0008",
     4554 => x"5b9d0004",  4555 => x"282500b0",  4556 => x"282400b4",
     4557 => x"282300b8",  4558 => x"282b0014",  4559 => x"282700a8",
     4560 => x"282600ac",  4561 => x"59650060",  4562 => x"59640064",
     4563 => x"282500bc",  4564 => x"282400c0",  4565 => x"59630068",
     4566 => x"282300c4",  4567 => x"282100cc",  4568 => x"59670058",
     4569 => x"59640070",  4570 => x"5961007c",  4571 => x"34010001",
     4572 => x"59610078",  4573 => x"1441001f",  4574 => x"59630074",
     4575 => x"5966005c",  4576 => x"5965006c",  4577 => x"34030000",
     4578 => x"340403e8",  4579 => x"f800319a",  4580 => x"1423001f",
     4581 => x"2063ffff",  4582 => x"b4621000",  4583 => x"f4621800",
     4584 => x"00420010",  4585 => x"b4610800",  4586 => x"3c210010",
     4587 => x"b8221000",  4588 => x"34010000",  4589 => x"59620074",
     4590 => x"2b9d0004",  4591 => x"2b8b0008",  4592 => x"379c0008",
     4593 => x"c3a00000",  4594 => x"379cffbc",  4595 => x"5b8b003c",
     4596 => x"5b8c0038",  4597 => x"5b8d0034",  4598 => x"5b8e0030",
     4599 => x"5b8f002c",  4600 => x"5b900028",  4601 => x"5b910024",
     4602 => x"5b920020",  4603 => x"5b93001c",  4604 => x"5b940018",
     4605 => x"5b950014",  4606 => x"5b960010",  4607 => x"5b97000c",
     4608 => x"5b980008",  4609 => x"5b9d0004",  4610 => x"b8206000",
     4611 => x"282102c8",  4612 => x"298b0014",  4613 => x"282e0010",
     4614 => x"78010001",  4615 => x"38215208",  4616 => x"28210000",
     4617 => x"44200276",  4618 => x"2963003c",  4619 => x"44600007",
     4620 => x"29610050",  4621 => x"44200005",  4622 => x"29610064",
     4623 => x"44200003",  4624 => x"29610078",  4625 => x"5c200011",
     4626 => x"78010001",  4627 => x"3821520c",  4628 => x"28220000",
     4629 => x"34420001",  4630 => x"58220000",  4631 => x"34010005",
     4632 => x"4c220267",  4633 => x"29640050",  4634 => x"29650064",
     4635 => x"29660078",  4636 => x"78010001",  4637 => x"78020001",
     4638 => x"38423f6c",  4639 => x"38212810",  4640 => x"f8001951",
     4641 => x"e000025e",  4642 => x"29c10000",  4643 => x"28230038",
     4644 => x"44600004",  4645 => x"b9600800",  4646 => x"34020000",
     4647 => x"d8600000",  4648 => x"78010001",  4649 => x"38216db4",
     4650 => x"28210000",  4651 => x"34020001",  4652 => x"fbfff245",
     4653 => x"78010001",  4654 => x"3821520c",  4655 => x"58200000",
     4656 => x"296100b8",  4657 => x"29660030",  4658 => x"29670034",
     4659 => x"34210001",  4660 => x"596100b8",  4661 => x"78010001",
     4662 => x"38215208",  4663 => x"58200000",  4664 => x"29680038",
     4665 => x"2965006c",  4666 => x"29640074",  4667 => x"29610070",
     4668 => x"c8a62800",  4669 => x"c8882000",  4670 => x"c8270800",
     4671 => x"e0000002",  4672 => x"348403e8",  4673 => x"b8201800",
     4674 => x"3421ffff",  4675 => x"4804fffd",  4676 => x"b8a00800",
     4677 => x"78050001",  4678 => x"38a53ce0",  4679 => x"28a20000",
     4680 => x"e0000002",  4681 => x"b4621800",  4682 => x"b8205000",
     4683 => x"3421ffff",  4684 => x"4803fffd",  4685 => x"29610044",
     4686 => x"29650058",  4687 => x"29620060",  4688 => x"2969005c",
     4689 => x"c8a12800",  4690 => x"2961004c",  4691 => x"c8410800",
     4692 => x"29620048",  4693 => x"c9224800",  4694 => x"e0000002",
     4695 => x"342103e8",  4696 => x"b9201000",  4697 => x"3529ffff",
     4698 => x"4801fffd",  4699 => x"78090001",  4700 => x"39293ce0",
     4701 => x"292d0000",  4702 => x"e0000002",  4703 => x"b44d1000",
     4704 => x"b8a04800",  4705 => x"34a5ffff",  4706 => x"4802fffd",
     4707 => x"c8810800",  4708 => x"c9495000",  4709 => x"c8622000",
     4710 => x"e0000002",  4711 => x"342103e8",  4712 => x"b8801000",
     4713 => x"3484ffff",  4714 => x"4801fffd",  4715 => x"78040001",
     4716 => x"38843ce0",  4717 => x"b9401800",  4718 => x"28850000",
     4719 => x"e0000002",  4720 => x"b4451000",  4721 => x"b8602000",
     4722 => x"3463ffff",  4723 => x"4802fffd",  4724 => x"59610094",
     4725 => x"78010001",  4726 => x"38214e9c",  4727 => x"59620090",
     4728 => x"28210000",  4729 => x"29820018",  4730 => x"5964008c",
     4731 => x"b8220800",  4732 => x"00210010",  4733 => x"2021000f",
     4734 => x"44200032",  4735 => x"780d0001",  4736 => x"39ad2840",
     4737 => x"78050001",  4738 => x"b9800800",  4739 => x"34020004",
     4740 => x"34030002",  4741 => x"b9a02000",  4742 => x"38a52850",
     4743 => x"fbfff29c",  4744 => x"29660044",  4745 => x"29670048",
     4746 => x"2968004c",  4747 => x"78050001",  4748 => x"b9800800",
     4749 => x"34020004",  4750 => x"34030002",  4751 => x"b9a02000",
     4752 => x"38a5285c",  4753 => x"fbfff292",  4754 => x"29660058",
     4755 => x"2967005c",  4756 => x"29680060",  4757 => x"78050001",
     4758 => x"b9800800",  4759 => x"34020004",  4760 => x"34030002",
     4761 => x"b9a02000",  4762 => x"38a52868",  4763 => x"fbfff288",
     4764 => x"2966006c",  4765 => x"29670070",  4766 => x"29680074",
     4767 => x"78050001",  4768 => x"b9800800",  4769 => x"34020004",
     4770 => x"34030002",  4771 => x"b9a02000",  4772 => x"38a52874",
     4773 => x"fbfff27e",  4774 => x"2966008c",  4775 => x"29670090",
     4776 => x"29680094",  4777 => x"78050001",  4778 => x"b9800800",
     4779 => x"34020004",  4780 => x"34030002",  4781 => x"b9a02000",
     4782 => x"38a52880",  4783 => x"fbfff274",  4784 => x"2962008c",
     4785 => x"78050001",  4786 => x"38a53cec",  4787 => x"28a40000",
     4788 => x"1441001f",  4789 => x"340300e8",  4790 => x"f80030c7",
     4791 => x"b8406800",  4792 => x"29620090",  4793 => x"b8207800",
     4794 => x"34030000",  4795 => x"1441001f",  4796 => x"340403e8",
     4797 => x"f80030c0",  4798 => x"29650094",  4799 => x"b5a21800",
     4800 => x"f5a36800",  4801 => x"14a2001f",  4802 => x"b5e10800",
     4803 => x"b4652800",  4804 => x"b5a10800",  4805 => x"f4651800",
     4806 => x"b4220800",  4807 => x"29640018",  4808 => x"29620020",
     4809 => x"b4611800",  4810 => x"2961001c",  4811 => x"297600a0",
     4812 => x"596300a0",  4813 => x"29630024",  4814 => x"b4821000",
     4815 => x"b4411000",  4816 => x"297400a4",  4817 => x"b4431000",
     4818 => x"596500a4",  4819 => x"1446001f",  4820 => x"4ca20003",
     4821 => x"596600a0",  4822 => x"596200a4",  4823 => x"296500a4",
     4824 => x"296100a0",  4825 => x"1477001f",  4826 => x"c8a21000",
     4827 => x"f4452800",  4828 => x"c8260800",  4829 => x"c8250800",
     4830 => x"1485001f",  4831 => x"b4642000",  4832 => x"f4641800",
     4833 => x"b6e5b800",  4834 => x"b477b800",  4835 => x"004d0001",
     4836 => x"3c23001f",  4837 => x"00250001",  4838 => x"b86d6800",
     4839 => x"b48d6800",  4840 => x"f48d2000",  4841 => x"b6e5b800",
     4842 => x"b497b800",  4843 => x"29640028",  4844 => x"1483001f",
     4845 => x"f8003090",  4846 => x"14350008",  4847 => x"1421001f",
     4848 => x"b5b5a800",  4849 => x"f5b56800",  4850 => x"b6e10800",
     4851 => x"b5a1b800",  4852 => x"29620030",  4853 => x"29610044",
     4854 => x"29720038",  4855 => x"29630034",  4856 => x"c8411000",
     4857 => x"2961004c",  4858 => x"ca419000",  4859 => x"29610048",
     4860 => x"c8611800",  4861 => x"e0000002",  4862 => x"365203e8",
     4863 => x"b8606800",  4864 => x"3463ffff",  4865 => x"4812fffd",
     4866 => x"78090001",  4867 => x"39293ce0",  4868 => x"29210000",
     4869 => x"e0000002",  4870 => x"b5a16800",  4871 => x"b8408800",
     4872 => x"3442ffff",  4873 => x"480dfffd",  4874 => x"378f0040",
     4875 => x"340203e8",  4876 => x"b9e00800",  4877 => x"5b970040",
     4878 => x"5b950044",  4879 => x"fbfff659",  4880 => x"78030001",
     4881 => x"38633ce0",  4882 => x"28620000",  4883 => x"b8208000",
     4884 => x"b9e00800",  4885 => x"fbfff653",  4886 => x"2b820044",
     4887 => x"b42d6800",  4888 => x"b6509000",  4889 => x"b6221000",
     4890 => x"340103e7",  4891 => x"e0000002",  4892 => x"3652fc18",
     4893 => x"b9a08800",  4894 => x"ba408000",  4895 => x"35ad0001",
     4896 => x"4a41fffc",  4897 => x"78040001",  4898 => x"78050001",
     4899 => x"38843cdc",  4900 => x"38a53cf0",  4901 => x"b8400800",
     4902 => x"28830000",  4903 => x"28a20000",  4904 => x"e0000002",
     4905 => x"b6228800",  4906 => x"b8207800",  4907 => x"ba206800",
     4908 => x"34210001",  4909 => x"4a23fffc",  4910 => x"2961002c",
     4911 => x"340203e8",  4912 => x"b9e0c000",  4913 => x"342103e7",
     4914 => x"f8003072",  4915 => x"b8209800",  4916 => x"4c110008",
     4917 => x"ba200800",  4918 => x"ba601000",  4919 => x"f800309a",
     4920 => x"4420000a",  4921 => x"083003e8",  4922 => x"ca216800",
     4923 => x"b6128000",  4924 => x"4da00006",  4925 => x"78090001",
     4926 => x"39293ce0",  4927 => x"29210000",  4928 => x"35efffff",
     4929 => x"b5a16800",  4930 => x"3401ffff",  4931 => x"5de10007",
     4932 => x"4c0d0006",  4933 => x"78020001",  4934 => x"38423cf0",
     4935 => x"28410000",  4936 => x"340f0000",  4937 => x"b5a16800",
     4938 => x"4da00007",  4939 => x"c8130800",  4940 => x"482d0005",
     4941 => x"5de00004",  4942 => x"b5b36800",  4943 => x"0a73fc18",
     4944 => x"b6138000",  4945 => x"78050001",  4946 => x"38a53cec",
     4947 => x"28a40000",  4948 => x"1701001f",  4949 => x"bb001000",
     4950 => x"340300e8",  4951 => x"f8003026",  4952 => x"b820c000",
     4953 => x"1621001f",  4954 => x"b8409800",  4955 => x"34030000",
     4956 => x"340403e8",  4957 => x"ba201000",  4958 => x"f800301f",
     4959 => x"b6621800",  4960 => x"f6639800",  4961 => x"1642001f",
     4962 => x"b7010800",  4963 => x"b4729000",  4964 => x"b6610800",
     4965 => x"b4220800",  4966 => x"f4721800",  4967 => x"78020001",
     4968 => x"38424a10",  4969 => x"b4611800",  4970 => x"28410000",
     4971 => x"596300e8",  4972 => x"34020000",  4973 => x"596100bc",
     4974 => x"29c10000",  4975 => x"597200ec",  4976 => x"597700b0",
     4977 => x"28230004",  4978 => x"597500b4",  4979 => x"b9800800",
     4980 => x"d8600000",  4981 => x"34020001",  4982 => x"4422000c",
     4983 => x"78040001",  4984 => x"b9800800",  4985 => x"34020004",
     4986 => x"34030001",  4987 => x"3884288c",  4988 => x"fbfff1a7",
     4989 => x"29c10000",  4990 => x"34020000",  4991 => x"28230034",
     4992 => x"b9800800",  4993 => x"d8600000",  4994 => x"29c10000",
     4995 => x"28210010",  4996 => x"d8200000",  4997 => x"5c200007",
     4998 => x"29630010",  4999 => x"3402fffd",  5000 => x"a0621000",
     5001 => x"59620010",  5002 => x"5de10009",  5003 => x"e000000a",
     5004 => x"78040001",  5005 => x"b9800800",  5006 => x"34020004",
     5007 => x"34030001",  5008 => x"388428b0",  5009 => x"fbfff192",
     5010 => x"e00000e2",  5011 => x"34010002",  5012 => x"e0000003",
     5013 => x"45af0003",  5014 => x"34010001",  5015 => x"59610014",
     5016 => x"78040001",  5017 => x"b9800800",  5018 => x"34020004",
     5019 => x"b9e02800",  5020 => x"b9a03000",  5021 => x"34030002",
     5022 => x"388428bc",  5023 => x"ba003800",  5024 => x"fbfff183",
     5025 => x"29620014",  5026 => x"78010001",  5027 => x"38213f54",
     5028 => x"3c420002",  5029 => x"78060001",  5030 => x"b4220800",
     5031 => x"28250000",  5032 => x"29610010",  5033 => x"38c63cd4",
     5034 => x"20210002",  5035 => x"44200003",  5036 => x"78060001",
     5037 => x"38c62800",  5038 => x"78040001",  5039 => x"b9800800",
     5040 => x"34020004",  5041 => x"34030001",  5042 => x"388428dc",
     5043 => x"fbfff170",  5044 => x"29620014",  5045 => x"78010001",
     5046 => x"38213f54",  5047 => x"3c420002",  5048 => x"b4221000",
     5049 => x"28420000",  5050 => x"356100c0",  5051 => x"f8003177",
     5052 => x"29620014",  5053 => x"34010004",  5054 => x"3442ffff",
     5055 => x"5441007e",  5056 => x"78010001",  5057 => x"3c420002",
     5058 => x"38213f40",  5059 => x"b4220800",  5060 => x"28210000",
     5061 => x"c0200000",  5062 => x"29c10000",  5063 => x"b9e01000",
     5064 => x"34030000",  5065 => x"28240014",  5066 => x"15e1001f",
     5067 => x"e0000006",  5068 => x"29c10000",  5069 => x"34020000",
     5070 => x"b9a01800",  5071 => x"28240014",  5072 => x"34010000",
     5073 => x"d8800000",  5074 => x"29610010",  5075 => x"38210002",
     5076 => x"59610010",  5077 => x"e0000043",  5078 => x"296500a8",
     5079 => x"78040001",  5080 => x"b9800800",  5081 => x"34020004",
     5082 => x"34030002",  5083 => x"388428f4",  5084 => x"b9a03000",
     5085 => x"ba003800",  5086 => x"fbfff145",  5087 => x"29c20000",
     5088 => x"296100a8",  5089 => x"28420018",  5090 => x"b6010800",
     5091 => x"596100a8",  5092 => x"d8400000",  5093 => x"29610010",
     5094 => x"38210002",  5095 => x"59610010",  5096 => x"34010005",
     5097 => x"59610014",  5098 => x"e0000053",  5099 => x"78090001",
     5100 => x"39293cec",  5101 => x"29240000",  5102 => x"15e1001f",
     5103 => x"b9e01000",  5104 => x"340300e8",  5105 => x"f8002f8c",
     5106 => x"b6027800",  5107 => x"1611001f",  5108 => x"f60f8000",
     5109 => x"b6210800",  5110 => x"b6018000",  5111 => x"15a1001f",
     5112 => x"34030000",  5113 => x"b9a01000",  5114 => x"340403e8",
     5115 => x"f8002f82",  5116 => x"b5e21800",  5117 => x"f5e37800",
     5118 => x"b6010800",  5119 => x"b5e10800",  5120 => x"c8031000",
     5121 => x"48010002",  5122 => x"b8601000",  5123 => x"3401003b",
     5124 => x"4841000d",  5125 => x"29c10000",  5126 => x"34020001",
     5127 => x"28230034",  5128 => x"b9800800",  5129 => x"d8600000",
     5130 => x"296100b0",  5131 => x"59610080",  5132 => x"296100b4",
     5133 => x"59610084",  5134 => x"34010004",  5135 => x"59610014",
     5136 => x"e0000004",  5137 => x"29610088",  5138 => x"34210001",
     5139 => x"59610088",  5140 => x"29620088",  5141 => x"34010009",
     5142 => x"4c220027",  5143 => x"59600088",  5144 => x"34010003",
     5145 => x"e3ffffd0",  5146 => x"296300b4",  5147 => x"29610084",
     5148 => x"296400b0",  5149 => x"29620080",  5150 => x"c8610800",
     5151 => x"f4231800",  5152 => x"596100e4",  5153 => x"78010001",
     5154 => x"38214a10",  5155 => x"c8821000",  5156 => x"28210000",
     5157 => x"c8431000",  5158 => x"596200e0",  5159 => x"44200016",
     5160 => x"1601001f",  5161 => x"29c20000",  5162 => x"0021001e",
     5163 => x"b4308000",  5164 => x"296100a8",  5165 => x"16100002",
     5166 => x"28420018",  5167 => x"b6010800",  5168 => x"596100a8",
     5169 => x"d8400000",  5170 => x"296500a8",  5171 => x"78040001",
     5172 => x"b9800800",  5173 => x"34020006",  5174 => x"34030001",
     5175 => x"38842910",  5176 => x"fbfff0eb",  5177 => x"296100b0",
     5178 => x"59610080",  5179 => x"296100b4",  5180 => x"59610084",
     5181 => x"29620014",  5182 => x"34010004",  5183 => x"44410004",
     5184 => x"296100f0",  5185 => x"34210001",  5186 => x"596100f0",
     5187 => x"296400e8",  5188 => x"296300ec",  5189 => x"1481001f",
     5190 => x"98611800",  5191 => x"c8611000",  5192 => x"98812000",
     5193 => x"f4431800",  5194 => x"c8810800",  5195 => x"c8230800",
     5196 => x"48200005",  5197 => x"5c200007",  5198 => x"340101f4",
     5199 => x"54410002",  5200 => x"e0000004",  5201 => x"296100f4",
     5202 => x"34210001",  5203 => x"596100f4",  5204 => x"296500a4",
     5205 => x"296400a0",  5206 => x"ca851800",  5207 => x"f4740800",
     5208 => x"cac41000",  5209 => x"c8411000",  5210 => x"48020007",
     5211 => x"34010001",  5212 => x"48400013",  5213 => x"5c400011",
     5214 => x"340203e8",  5215 => x"54620010",  5216 => x"e000000e",
     5217 => x"c8140800",  5218 => x"7c220000",  5219 => x"c8161800",
     5220 => x"c8621800",  5221 => x"c8251000",  5222 => x"f4410800",
     5223 => x"c8641800",  5224 => x"c8611800",  5225 => x"34010001",
     5226 => x"48600005",  5227 => x"5c600003",  5228 => x"340303e8",
     5229 => x"54430002",  5230 => x"34010000",  5231 => x"202100ff",
     5232 => x"44200004",  5233 => x"296100f8",  5234 => x"34210001",
     5235 => x"596100f8",  5236 => x"78010001",  5237 => x"38216db4",
     5238 => x"28210000",  5239 => x"34020000",  5240 => x"fbffeff9",
     5241 => x"29c10000",  5242 => x"28230038",  5243 => x"44600004",
     5244 => x"b9600800",  5245 => x"34020001",  5246 => x"d8600000",
     5247 => x"34010000",  5248 => x"2b9d0004",  5249 => x"2b8b003c",
     5250 => x"2b8c0038",  5251 => x"2b8d0034",  5252 => x"2b8e0030",
     5253 => x"2b8f002c",  5254 => x"2b900028",  5255 => x"2b910024",
     5256 => x"2b920020",  5257 => x"2b93001c",  5258 => x"2b940018",
     5259 => x"2b950014",  5260 => x"2b960010",  5261 => x"2b97000c",
     5262 => x"2b980008",  5263 => x"379c0044",  5264 => x"c3a00000",
     5265 => x"379cffe8",  5266 => x"5b8b0018",  5267 => x"5b8c0014",
     5268 => x"5b8d0010",  5269 => x"5b8e000c",  5270 => x"5b8f0008",
     5271 => x"5b9d0004",  5272 => x"b8407800",  5273 => x"28220020",
     5274 => x"b8205800",  5275 => x"b8607000",  5276 => x"284d0008",
     5277 => x"28220024",  5278 => x"282c02c8",  5279 => x"28440000",
     5280 => x"d8800000",  5281 => x"48010058",  5282 => x"29610020",
     5283 => x"34030008",  5284 => x"2824000c",  5285 => x"4161004c",
     5286 => x"30810004",  5287 => x"4161004d",  5288 => x"30810005",
     5289 => x"4161004e",  5290 => x"30810006",  5291 => x"3401ffff",
     5292 => x"30810007",  5293 => x"3401fffe",  5294 => x"30810008",
     5295 => x"4161004f",  5296 => x"30810009",  5297 => x"41610050",
     5298 => x"3081000a",  5299 => x"41610051",  5300 => x"3081000b",
     5301 => x"29610020",  5302 => x"2824000c",  5303 => x"b9800800",
     5304 => x"34820004",  5305 => x"f8002f99",  5306 => x"29610020",
     5307 => x"35620374",  5308 => x"28210000",  5309 => x"3180000a",
     5310 => x"c8410800",  5311 => x"14210002",  5312 => x"0821d775",
     5313 => x"0d810008",  5314 => x"41a10042",  5315 => x"3181000b",
     5316 => x"34010014",  5317 => x"3181000c",  5318 => x"41a10043",
     5319 => x"3181000d",  5320 => x"34010002",  5321 => x"3181000e",
     5322 => x"78010001",  5323 => x"382149dc",  5324 => x"28240000",
     5325 => x"4480000f",  5326 => x"b9600800",  5327 => x"b9e01000",
     5328 => x"b9c01800",  5329 => x"d8800000",  5330 => x"4420000a",
     5331 => x"78040001",  5332 => x"78050001",  5333 => x"b9600800",
     5334 => x"34020002",  5335 => x"34030001",  5336 => x"3884297c",
     5337 => x"38a53f7c",  5338 => x"fbfff049",  5339 => x"e000001e",
     5340 => x"29610020",  5341 => x"78040001",  5342 => x"34020003",
     5343 => x"2825000c",  5344 => x"34030001",  5345 => x"b9600800",
     5346 => x"40a5000e",  5347 => x"38842998",  5348 => x"fbfff03f",
     5349 => x"29610020",  5350 => x"78040001",  5351 => x"34020003",
     5352 => x"2825000c",  5353 => x"34030001",  5354 => x"b9600800",
     5355 => x"40a5000f",  5356 => x"388429ac",  5357 => x"fbfff036",
     5358 => x"2962003c",  5359 => x"b9600800",  5360 => x"f8000634",
     5361 => x"4162001d",  5362 => x"34010001",  5363 => x"44410003",
     5364 => x"34010004",  5365 => x"e0000002",  5366 => x"34010006",
     5367 => x"59610004",  5368 => x"e0000003",  5369 => x"340103e8",
     5370 => x"59610008",  5371 => x"34010000",  5372 => x"2b9d0004",
     5373 => x"2b8b0018",  5374 => x"2b8c0014",  5375 => x"2b8d0010",
     5376 => x"2b8e000c",  5377 => x"2b8f0008",  5378 => x"379c0018",
     5379 => x"c3a00000",  5380 => x"379cfff4",  5381 => x"5b8b000c",
     5382 => x"5b8c0008",  5383 => x"5b9d0004",  5384 => x"2822000c",
     5385 => x"b8205800",  5386 => x"44400006",  5387 => x"28220028",
     5388 => x"28430018",  5389 => x"34020fa0",  5390 => x"d8600000",
     5391 => x"596102dc",  5392 => x"296102dc",  5393 => x"44200009",
     5394 => x"29610028",  5395 => x"34020000",  5396 => x"28230018",
     5397 => x"b9600800",  5398 => x"d8600000",  5399 => x"296202dc",
     5400 => x"c8220800",  5401 => x"4c200014",  5402 => x"296c02dc",
     5403 => x"34010000",  5404 => x"4580000a",  5405 => x"29610028",
     5406 => x"34020000",  5407 => x"28230018",  5408 => x"b9600800",
     5409 => x"d8600000",  5410 => x"c9810800",  5411 => x"a4201000",
     5412 => x"1442001f",  5413 => x"a0220800",  5414 => x"59610008",
     5415 => x"34010000",  5416 => x"2b9d0004",  5417 => x"2b8b000c",
     5418 => x"2b8c0008",  5419 => x"379c000c",  5420 => x"c3a00000",
     5421 => x"b9600800",  5422 => x"34020004",  5423 => x"f8000a67",
     5424 => x"34010001",  5425 => x"59610004",  5426 => x"e3fffff5",
     5427 => x"340203e8",  5428 => x"58220008",  5429 => x"34010000",
     5430 => x"c3a00000",  5431 => x"379cfff0",  5432 => x"5b8b0010",
     5433 => x"5b8c000c",  5434 => x"5b8d0008",  5435 => x"5b9d0004",
     5436 => x"78040001",  5437 => x"388449dc",  5438 => x"2884000c",
     5439 => x"b8205800",  5440 => x"b8406800",  5441 => x"b8606000",
     5442 => x"44800003",  5443 => x"d8800000",  5444 => x"5c20001f",
     5445 => x"2961000c",  5446 => x"4420000b",  5447 => x"296102c8",
     5448 => x"29630028",  5449 => x"4022000c",  5450 => x"1021000b",
     5451 => x"28630018",  5452 => x"bc411000",  5453 => x"b9600800",
     5454 => x"084203e8",  5455 => x"d8600000",  5456 => x"596102d4",
     5457 => x"4580000f",  5458 => x"4161030d",  5459 => x"44200008",
     5460 => x"3402000b",  5461 => x"5c22000b",  5462 => x"b9600800",
     5463 => x"b9a01000",  5464 => x"b9801800",  5465 => x"f8000352",
     5466 => x"e0000005",  5467 => x"b9600800",  5468 => x"b9a01000",
     5469 => x"b9801800",  5470 => x"f8000370",  5471 => x"5c200004",
     5472 => x"b9600800",  5473 => x"f800027e",  5474 => x"44200003",
     5475 => x"34010002",  5476 => x"59610004",  5477 => x"29620004",
     5478 => x"29610000",  5479 => x"44410002",  5480 => x"596002d4",
     5481 => x"296c02d4",  5482 => x"34010000",  5483 => x"4580000a",
     5484 => x"29610028",  5485 => x"34020000",  5486 => x"28230018",
     5487 => x"b9600800",  5488 => x"d8600000",  5489 => x"c9810800",
     5490 => x"a4201000",  5491 => x"1442001f",  5492 => x"a0220800",
     5493 => x"59610008",  5494 => x"34010000",  5495 => x"2b9d0004",
     5496 => x"2b8b0010",  5497 => x"2b8c000c",  5498 => x"2b8d0008",
     5499 => x"379c0010",  5500 => x"c3a00000",  5501 => x"34010000",
     5502 => x"c3a00000",  5503 => x"379cffec",  5504 => x"5b8b0014",
     5505 => x"5b8c0010",  5506 => x"5b8d000c",  5507 => x"5b8e0008",
     5508 => x"5b9d0004",  5509 => x"344b00b2",  5510 => x"3d6b0002",
     5511 => x"b8407000",  5512 => x"b42b5800",  5513 => x"29620004",
     5514 => x"b8206000",  5515 => x"340d0000",  5516 => x"44400008",
     5517 => x"28220028",  5518 => x"28430018",  5519 => x"34020000",
     5520 => x"d8600000",  5521 => x"29620004",  5522 => x"c8220800",
     5523 => x"4c200009",  5524 => x"b9a00800",  5525 => x"2b9d0004",
     5526 => x"2b8b0014",  5527 => x"2b8c0010",  5528 => x"2b8d000c",
     5529 => x"2b8e0008",  5530 => x"379c0014",  5531 => x"c3a00000",
     5532 => x"b9800800",  5533 => x"b9c01000",  5534 => x"f80009f8",
     5535 => x"340d0001",  5536 => x"59600004",  5537 => x"e3fffff3",
     5538 => x"379cffec",  5539 => x"5b8b0014",  5540 => x"5b8c0010",
     5541 => x"5b8d000c",  5542 => x"5b8e0008",  5543 => x"5b9d0004",
     5544 => x"b8407000",  5545 => x"2822000c",  5546 => x"b8205800",
     5547 => x"b8606800",  5548 => x"340c0000",  5549 => x"44400014",
     5550 => x"282302c8",  5551 => x"34020001",  5552 => x"1063000d",
     5553 => x"f80009f4",  5554 => x"296302c8",  5555 => x"b9600800",
     5556 => x"34020003",  5557 => x"1063000b",  5558 => x"f80009ef",
     5559 => x"29630344",  5560 => x"34020001",  5561 => x"34010000",
     5562 => x"5c620002",  5563 => x"29610340",  5564 => x"0d61007e",
     5565 => x"b9600800",  5566 => x"f80005d9",  5567 => x"b8206000",
     5568 => x"48010047",  5569 => x"b9600800",  5570 => x"34020001",
     5571 => x"fbffffbc",  5572 => x"44200010",  5573 => x"296302c8",
     5574 => x"b9600800",  5575 => x"34020001",  5576 => x"1063000d",
     5577 => x"f80009dc",  5578 => x"29630344",  5579 => x"34020001",
     5580 => x"34010000",  5581 => x"5c620002",  5582 => x"29610340",
     5583 => x"0d61007e",  5584 => x"b9600800",  5585 => x"f8000613",
     5586 => x"48010046",  5587 => x"340c0000",  5588 => x"b9600800",
     5589 => x"34020003",  5590 => x"fbffffa9",  5591 => x"44200010",
     5592 => x"29630344",  5593 => x"34020001",  5594 => x"34010000",
     5595 => x"5c620002",  5596 => x"29610340",  5597 => x"0d61007e",
     5598 => x"b9600800",  5599 => x"f80005b8",  5600 => x"48010038",
     5601 => x"296302c8",  5602 => x"b9600800",  5603 => x"34020003",
     5604 => x"1063000b",  5605 => x"340c0000",  5606 => x"f80009bf",
     5607 => x"45a00020",  5608 => x"78010001",  5609 => x"382149dc",
     5610 => x"28250010",  5611 => x"4164030d",  5612 => x"44a00007",
     5613 => x"b9600800",  5614 => x"b9c01000",  5615 => x"b9a01800",
     5616 => x"d8a00000",  5617 => x"b8202000",  5618 => x"48010042",
     5619 => x"34010001",  5620 => x"44810010",  5621 => x"3401000b",
     5622 => x"44810003",  5623 => x"5c800010",  5624 => x"e0000006",
     5625 => x"b9600800",  5626 => x"b9c01000",  5627 => x"b9a01800",
     5628 => x"f80002af",  5629 => x"e0000005",  5630 => x"b9600800",
     5631 => x"b9c01000",  5632 => x"b9a01800",  5633 => x"f80002cd",
     5634 => x"b8206000",  5635 => x"e0000004",  5636 => x"b9600800",
     5637 => x"356200e4",  5638 => x"f800066a",  5639 => x"45800006",
     5640 => x"34010001",  5641 => x"4581000f",  5642 => x"3401ffff",
     5643 => x"5d81000e",  5644 => x"e0000029",  5645 => x"29610020",
     5646 => x"2821000c",  5647 => x"4022000e",  5648 => x"340100ff",
     5649 => x"44410004",  5650 => x"4162001d",  5651 => x"34010002",
     5652 => x"5c410005",  5653 => x"34010004",  5654 => x"59610004",
     5655 => x"e0000002",  5656 => x"340c0000",  5657 => x"296e02d8",
     5658 => x"340d0000",  5659 => x"45c0000a",  5660 => x"29610028",
     5661 => x"34020000",  5662 => x"28230018",  5663 => x"b9600800",
     5664 => x"d8600000",  5665 => x"c9c16800",  5666 => x"a5a00800",
     5667 => x"1421001f",  5668 => x"a1a16800",  5669 => x"296e02d0",
     5670 => x"34010000",  5671 => x"45c0000a",  5672 => x"29610028",
     5673 => x"34020000",  5674 => x"28230018",  5675 => x"b9600800",
     5676 => x"d8600000",  5677 => x"c9c10800",  5678 => x"a4201000",
     5679 => x"1442001f",  5680 => x"a0220800",  5681 => x"4da10007",
     5682 => x"b9a00800",  5683 => x"e0000005",  5684 => x"b8206000",
     5685 => x"34010002",  5686 => x"59610004",  5687 => x"340101f4",
     5688 => x"59610008",  5689 => x"b9800800",  5690 => x"2b9d0004",
     5691 => x"2b8b0014",  5692 => x"2b8c0010",  5693 => x"2b8d000c",
     5694 => x"2b8e0008",  5695 => x"379c0014",  5696 => x"c3a00000",
     5697 => x"379cfff0",  5698 => x"5b8b000c",  5699 => x"5b8c0008",
     5700 => x"5b9d0004",  5701 => x"b8406000",  5702 => x"2822000c",
     5703 => x"b8205800",  5704 => x"4440000c",  5705 => x"282202c8",
     5706 => x"28250028",  5707 => x"4044000c",  5708 => x"1042000b",
     5709 => x"bc821000",  5710 => x"28a40018",  5711 => x"084203e8",
     5712 => x"5b830010",  5713 => x"d8800000",  5714 => x"2b830010",
     5715 => x"596102d4",  5716 => x"4460000d",  5717 => x"4161030d",
     5718 => x"44200007",  5719 => x"3402000b",  5720 => x"5c220009",
     5721 => x"b9600800",  5722 => x"b9801000",  5723 => x"f8000250",
     5724 => x"e0000004",  5725 => x"b9600800",  5726 => x"b9801000",
     5727 => x"f800026f",  5728 => x"5c200004",  5729 => x"b9600800",
     5730 => x"f800017d",  5731 => x"44200003",  5732 => x"34010002",
     5733 => x"59610004",  5734 => x"29620004",  5735 => x"29610000",
     5736 => x"44410002",  5737 => x"596002d4",  5738 => x"340103e8",
     5739 => x"59610008",  5740 => x"34010000",  5741 => x"2b9d0004",
     5742 => x"2b8b000c",  5743 => x"2b8c0008",  5744 => x"379c0010",
     5745 => x"c3a00000",  5746 => x"379cfff8",  5747 => x"5b8b0008",
     5748 => x"5b9d0004",  5749 => x"b8205800",  5750 => x"4460000d",
     5751 => x"4024030d",  5752 => x"44800007",  5753 => x"34050008",
     5754 => x"44850007",  5755 => x"3405000b",  5756 => x"5c850007",
     5757 => x"f8000198",  5758 => x"e0000004",  5759 => x"f80001b1",
     5760 => x"e0000002",  5761 => x"f80001e9",  5762 => x"5c200004",
     5763 => x"b9600800",  5764 => x"f800015b",  5765 => x"44200003",
     5766 => x"34010002",  5767 => x"59610004",  5768 => x"340103e8",
     5769 => x"59610008",  5770 => x"34010000",  5771 => x"2b9d0004",
     5772 => x"2b8b0008",  5773 => x"379c0008",  5774 => x"c3a00000",
     5775 => x"379cffd4",  5776 => x"5b8b0014",  5777 => x"5b8c0010",
     5778 => x"5b8d000c",  5779 => x"5b8e0008",  5780 => x"5b9d0004",
     5781 => x"b8205800",  5782 => x"2821000c",  5783 => x"b8407000",
     5784 => x"b8606800",  5785 => x"44200023",  5786 => x"34020000",
     5787 => x"34030014",  5788 => x"35610080",  5789 => x"f8002e33",
     5790 => x"b9600800",  5791 => x"f80006da",  5792 => x"78010001",
     5793 => x"382149dc",  5794 => x"28240014",  5795 => x"44800007",
     5796 => x"b9600800",  5797 => x"b9c01000",  5798 => x"b9a01800",
     5799 => x"d8800000",  5800 => x"b8206000",  5801 => x"5c20005f",
     5802 => x"4161001c",  5803 => x"29630028",  5804 => x"202100fd",
     5805 => x"3161001c",  5806 => x"296102c8",  5807 => x"28630018",
     5808 => x"4022000c",  5809 => x"1021000b",  5810 => x"bc411000",
     5811 => x"b9600800",  5812 => x"084203e8",  5813 => x"d8600000",
     5814 => x"296302c8",  5815 => x"596102d4",  5816 => x"34020000",
     5817 => x"1063000a",  5818 => x"b9600800",  5819 => x"f80008ea",
     5820 => x"45a00049",  5821 => x"4161030d",  5822 => x"34020008",
     5823 => x"44220012",  5824 => x"54220003",  5825 => x"5c200044",
     5826 => x"e000000a",  5827 => x"34020009",  5828 => x"44220014",
     5829 => x"3402000b",  5830 => x"5c22003f",  5831 => x"b9600800",
     5832 => x"b9c01000",  5833 => x"b9a01800",  5834 => x"f800014b",
     5835 => x"e000000a",  5836 => x"b9600800",  5837 => x"b9c01000",
     5838 => x"b9a01800",  5839 => x"f8000161",  5840 => x"e0000005",
     5841 => x"b9600800",  5842 => x"b9c01000",  5843 => x"b9a01800",
     5844 => x"f8000196",  5845 => x"b8206000",  5846 => x"5c200032",
     5847 => x"e000002e",  5848 => x"34010035",  5849 => x"340c0001",
     5850 => x"4c2d002e",  5851 => x"378c0018",  5852 => x"b9c00800",
     5853 => x"b9801000",  5854 => x"f80004a2",  5855 => x"296102c8",
     5856 => x"37820024",  5857 => x"34030008",  5858 => x"f8002d4f",
     5859 => x"5c20001c",  5860 => x"2d6202f2",  5861 => x"2d61032a",
     5862 => x"5c410019",  5863 => x"296102c8",  5864 => x"2c220008",
     5865 => x"2f81002c",  5866 => x"5c410015",  5867 => x"4161001c",
     5868 => x"20210001",  5869 => x"44200012",  5870 => x"b9801000",
     5871 => x"356100bc",  5872 => x"f8000619",  5873 => x"78010001",
     5874 => x"382149dc",  5875 => x"28220018",  5876 => x"44400006",
     5877 => x"b9600800",  5878 => x"d8400000",  5879 => x"b8206000",
     5880 => x"5c200010",  5881 => x"e0000003",  5882 => x"b9600800",
     5883 => x"f80006d7",  5884 => x"4161032d",  5885 => x"316102ee",
     5886 => x"e0000007",  5887 => x"78040001",  5888 => x"b9600800",
     5889 => x"34020005",  5890 => x"34030002",  5891 => x"388429c4",
     5892 => x"fbffee1f",  5893 => x"b9600800",  5894 => x"f80000d9",
     5895 => x"b8206000",  5896 => x"296102cc",  5897 => x"44200009",
     5898 => x"29610028",  5899 => x"34020000",  5900 => x"28230018",
     5901 => x"b9600800",  5902 => x"d8600000",  5903 => x"296202cc",
     5904 => x"c8220800",  5905 => x"4c200033",  5906 => x"3401ffff",
     5907 => x"45810005",  5908 => x"7d810001",  5909 => x"c8010800",
     5910 => x"a1816000",  5911 => x"e0000003",  5912 => x"34010002",
     5913 => x"59610004",  5914 => x"29620004",  5915 => x"29610000",
     5916 => x"44410005",  5917 => x"596002d4",  5918 => x"596002cc",
     5919 => x"b9600800",  5920 => x"f8000659",  5921 => x"296e02d4",
     5922 => x"340d0000",  5923 => x"45c0000a",  5924 => x"29610028",
     5925 => x"34020000",  5926 => x"28230018",  5927 => x"b9600800",
     5928 => x"d8600000",  5929 => x"c9c16800",  5930 => x"a5a00800",
     5931 => x"1421001f",  5932 => x"a1a16800",  5933 => x"296e02cc",
     5934 => x"b9a00800",  5935 => x"45c0000a",  5936 => x"29610028",
     5937 => x"34020000",  5938 => x"28230018",  5939 => x"b9600800",
     5940 => x"d8600000",  5941 => x"c9c10800",  5942 => x"a4201000",
     5943 => x"1442001f",  5944 => x"a0220800",  5945 => x"4da10002",
     5946 => x"b9a00800",  5947 => x"59610008",  5948 => x"b9800800",
     5949 => x"2b9d0004",  5950 => x"2b8b0014",  5951 => x"2b8c0010",
     5952 => x"2b8d000c",  5953 => x"2b8e0008",  5954 => x"379c002c",
     5955 => x"c3a00000",  5956 => x"b9600800",  5957 => x"34020000",
     5958 => x"f8000850",  5959 => x"b9600800",  5960 => x"596002cc",
     5961 => x"f80004f6",  5962 => x"29630100",  5963 => x"29620104",
     5964 => x"296500f8",  5965 => x"296400fc",  5966 => x"b8206000",
     5967 => x"29610108",  5968 => x"596300b0",  5969 => x"296302c8",
     5970 => x"596200b4",  5971 => x"596100b8",  5972 => x"596500a8",
     5973 => x"596400ac",  5974 => x"1063000a",  5975 => x"b9600800",
     5976 => x"34020000",  5977 => x"f800084c",  5978 => x"29620020",
     5979 => x"356100a8",  5980 => x"28430008",  5981 => x"b8201000",
     5982 => x"34630018",  5983 => x"f80005bd",  5984 => x"e3ffffb2",
     5985 => x"379cfff8",  5986 => x"5b8b0008",  5987 => x"5b9d0004",
     5988 => x"282202c8",  5989 => x"28240028",  5990 => x"b8205800",
     5991 => x"4043000c",  5992 => x"1042000b",  5993 => x"bc621000",
     5994 => x"28830018",  5995 => x"084203e8",  5996 => x"d8600000",
     5997 => x"596102d4",  5998 => x"2b9d0004",  5999 => x"2b8b0008",
     6000 => x"379c0008",  6001 => x"c3a00000",  6002 => x"379cffe4",
     6003 => x"5b8b001c",  6004 => x"5b8c0018",  6005 => x"5b8d0014",
     6006 => x"5b8e0010",  6007 => x"5b8f000c",  6008 => x"5b900008",
     6009 => x"5b9d0004",  6010 => x"340c0000",  6011 => x"b8205800",
     6012 => x"b8407000",  6013 => x"342f030c",  6014 => x"34300320",
     6015 => x"e0000013",  6016 => x"098d0058",  6017 => x"ba000800",
     6018 => x"3403000a",  6019 => x"35a20110",  6020 => x"b5621000",
     6021 => x"f8002cac",  6022 => x"5c20000b",  6023 => x"b56d0800",
     6024 => x"b9e01000",  6025 => x"34030024",  6026 => x"34210144",
     6027 => x"f8002cc7",  6028 => x"b56d5800",  6029 => x"b9c00800",
     6030 => x"3562011c",  6031 => x"f80003be",  6032 => x"e0000020",
     6033 => x"358c0001",  6034 => x"2d63010c",  6035 => x"486cffed",
     6036 => x"34010004",  6037 => x"54610003",  6038 => x"34630001",
     6039 => x"0d63010c",  6040 => x"2d6d010c",  6041 => x"35620320",
     6042 => x"3403000a",  6043 => x"35adffff",  6044 => x"09ac0058",
     6045 => x"35810110",  6046 => x"b5610800",  6047 => x"f8002cb3",
     6048 => x"b56c0800",  6049 => x"34030024",  6050 => x"b9e01000",
     6051 => x"34210144",  6052 => x"f8002cae",  6053 => x"b56c1000",
     6054 => x"b9c00800",  6055 => x"3442011c",  6056 => x"f80003a5",
     6057 => x"78040001",  6058 => x"b9600800",  6059 => x"34020003",
     6060 => x"34030001",  6061 => x"388429f4",  6062 => x"b9a02800",
     6063 => x"fbffed74",  6064 => x"2b9d0004",  6065 => x"2b8b001c",
     6066 => x"2b8c0018",  6067 => x"2b8d0014",  6068 => x"2b8e0010",
     6069 => x"2b8f000c",  6070 => x"2b900008",  6071 => x"379c001c",
     6072 => x"c3a00000",  6073 => x"4022001e",  6074 => x"34030001",
     6075 => x"44430009",  6076 => x"44400008",  6077 => x"34030002",
     6078 => x"5c430008",  6079 => x"34020012",  6080 => x"58220070",
     6081 => x"3402000e",  6082 => x"58220074",  6083 => x"e0000003",
     6084 => x"58200070",  6085 => x"58200074",  6086 => x"28240070",
     6087 => x"2825002c",  6088 => x"34020000",  6089 => x"b4a42800",
     6090 => x"20a30003",  6091 => x"44600003",  6092 => x"34020004",
     6093 => x"c8431000",  6094 => x"b4a22800",  6095 => x"28260030",
     6096 => x"28220074",  6097 => x"5825003c",  6098 => x"34030000",
     6099 => x"b4c23000",  6100 => x"20c70003",  6101 => x"44e00003",
     6102 => x"34030004",  6103 => x"c8671800",  6104 => x"b4c31800",
     6105 => x"c8a42000",  6106 => x"c8621000",  6107 => x"58230040",
     6108 => x"58240034",  6109 => x"58220038",  6110 => x"c3a00000",
     6111 => x"379cfff4",  6112 => x"5b8b000c",  6113 => x"5b8c0008",
     6114 => x"5b9d0004",  6115 => x"78020001",  6116 => x"384249dc",
     6117 => x"28420020",  6118 => x"b8205800",  6119 => x"44400006",
     6120 => x"d8400000",  6121 => x"b8206000",  6122 => x"34010001",
     6123 => x"45810018",  6124 => x"480c0018",  6125 => x"296102d4",
     6126 => x"340c0000",  6127 => x"44200015",  6128 => x"29610028",
     6129 => x"34020000",  6130 => x"28230018",  6131 => x"b9600800",
     6132 => x"d8600000",  6133 => x"296202d4",  6134 => x"c8220800",
     6135 => x"4c200013",  6136 => x"e000000c",  6137 => x"4162001d",
     6138 => x"34010002",  6139 => x"44410004",  6140 => x"34010006",
     6141 => x"59610004",  6142 => x"e0000006",  6143 => x"34010004",
     6144 => x"59610004",  6145 => x"b9600800",  6146 => x"fbffff5f",
     6147 => x"340c0000",  6148 => x"b9800800",  6149 => x"2b9d0004",
     6150 => x"2b8b000c",  6151 => x"2b8c0008",  6152 => x"379c000c",
     6153 => x"c3a00000",  6154 => x"b9600800",  6155 => x"34020002",
     6156 => x"f800078a",  6157 => x"29610020",  6158 => x"596002d4",
     6159 => x"0d60010c",  6160 => x"2821000c",  6161 => x"4022000e",
     6162 => x"340100ff",  6163 => x"5c41ffe6",  6164 => x"e3ffffeb",
     6165 => x"379cfff4",  6166 => x"5b8b000c",  6167 => x"5b8c0008",
     6168 => x"5b9d0004",  6169 => x"3404003f",  6170 => x"b8205800",
     6171 => x"340cffff",  6172 => x"4c83000e",  6173 => x"fbffff55",
     6174 => x"b9600800",  6175 => x"fbffff42",  6176 => x"b9600800",
     6177 => x"f800015a",  6178 => x"59610004",  6179 => x"78010001",
     6180 => x"382149dc",  6181 => x"28220024",  6182 => x"340c0000",
     6183 => x"44400003",  6184 => x"b9600800",  6185 => x"d8400000",
     6186 => x"b9800800",  6187 => x"2b9d0004",  6188 => x"2b8b000c",
     6189 => x"2b8c0008",  6190 => x"379c000c",  6191 => x"c3a00000",
     6192 => x"379cffe0",  6193 => x"5b8b0014",  6194 => x"5b8c0010",
     6195 => x"5b8d000c",  6196 => x"5b8e0008",  6197 => x"5b9d0004",
     6198 => x"b8205800",  6199 => x"3401002b",  6200 => x"b8407000",
     6201 => x"340cffff",  6202 => x"4c230028",  6203 => x"4161001c",
     6204 => x"340c0000",  6205 => x"20210001",  6206 => x"44200024",
     6207 => x"296300ec",  6208 => x"296200f0",  6209 => x"296100f4",
     6210 => x"296500e4",  6211 => x"296400e8",  6212 => x"5963009c",
     6213 => x"596200a0",  6214 => x"2963031c",  6215 => x"29620318",
     6216 => x"596100a4",  6217 => x"59650094",  6218 => x"356100d0",
     6219 => x"59640098",  6220 => x"f8000485",  6221 => x"41610313",
     6222 => x"20210002",  6223 => x"44200007",  6224 => x"4161001c",
     6225 => x"38210002",  6226 => x"3161001c",  6227 => x"2d61032a",
     6228 => x"0d6102ec",  6229 => x"e000000d",  6230 => x"378d0018",
     6231 => x"b9c00800",  6232 => x"b9a01000",  6233 => x"f80002ed",
     6234 => x"4161001c",  6235 => x"b9a01000",  6236 => x"202100fd",
     6237 => x"3161001c",  6238 => x"35610080",  6239 => x"f80004aa",
     6240 => x"b9600800",  6241 => x"f8000551",  6242 => x"b9800800",
     6243 => x"2b9d0004",  6244 => x"2b8b0014",  6245 => x"2b8c0010",
     6246 => x"2b8d000c",  6247 => x"2b8e0008",  6248 => x"379c0020",
     6249 => x"c3a00000",  6250 => x"379cffe4",  6251 => x"5b8b0010",
     6252 => x"5b8c000c",  6253 => x"5b8d0008",  6254 => x"5b9d0004",
     6255 => x"b8205800",  6256 => x"b8400800",  6257 => x"3402002b",
     6258 => x"3404ffff",  6259 => x"4c430031",  6260 => x"4162001c",
     6261 => x"20430001",  6262 => x"5c600004",  6263 => x"78010001",
     6264 => x"38212a14",  6265 => x"e0000005",  6266 => x"20420002",
     6267 => x"5c400007",  6268 => x"78010001",  6269 => x"38212a50",
     6270 => x"78020001",  6271 => x"38423f8c",  6272 => x"f80012f1",
     6273 => x"e0000022",  6274 => x"2d6402ec",  6275 => x"2d63032a",
     6276 => x"44830007",  6277 => x"78010001",  6278 => x"78020001",
     6279 => x"38423f8c",  6280 => x"38212a88",  6281 => x"f80012e8",
     6282 => x"e0000019",  6283 => x"378d0014",  6284 => x"b9a01000",
     6285 => x"f80002ec",  6286 => x"4161001c",  6287 => x"356c0080",
     6288 => x"b9a01000",  6289 => x"202100fd",  6290 => x"3161001c",
     6291 => x"b9800800",  6292 => x"f8000475",  6293 => x"78030001",
     6294 => x"386349dc",  6295 => x"28640028",  6296 => x"44800009",
     6297 => x"b9600800",  6298 => x"b9801000",  6299 => x"356300d0",
     6300 => x"d8800000",  6301 => x"b8202000",  6302 => x"34010001",
     6303 => x"44810004",  6304 => x"48040004",  6305 => x"b9600800",
     6306 => x"f8000510",  6307 => x"34040000",  6308 => x"b8800800",
     6309 => x"2b9d0004",  6310 => x"2b8b0010",  6311 => x"2b8c000c",
     6312 => x"2b8d0008",  6313 => x"379c001c",  6314 => x"c3a00000",
     6315 => x"379cfff0",  6316 => x"5b8b0010",  6317 => x"5b8c000c",
     6318 => x"5b8d0008",  6319 => x"5b9d0004",  6320 => x"b8406800",
     6321 => x"3402003f",  6322 => x"b8205800",  6323 => x"340cffff",
     6324 => x"4c430013",  6325 => x"78040001",  6326 => x"34030002",
     6327 => x"38842ac8",  6328 => x"34020003",  6329 => x"fbffec6a",
     6330 => x"b9a01000",  6331 => x"b9600800",  6332 => x"fbfffeb6",
     6333 => x"b9600800",  6334 => x"f80000bd",  6335 => x"59610004",
     6336 => x"78010001",  6337 => x"382149dc",  6338 => x"28220024",
     6339 => x"340c0000",  6340 => x"44400003",  6341 => x"b9600800",
     6342 => x"d8400000",  6343 => x"b9800800",  6344 => x"2b9d0004",
     6345 => x"2b8b0010",  6346 => x"2b8c000c",  6347 => x"2b8d0008",
     6348 => x"379c0010",  6349 => x"c3a00000",  6350 => x"34010000",
     6351 => x"c3a00000",  6352 => x"379cfffc",  6353 => x"5b9d0004",
     6354 => x"34030008",  6355 => x"f8002b5e",  6356 => x"2b9d0004",
     6357 => x"379c0004",  6358 => x"c3a00000",  6359 => x"379cffe0",
     6360 => x"5b8b0020",  6361 => x"5b8c001c",  6362 => x"5b8d0018",
     6363 => x"5b8e0014",  6364 => x"5b8f0010",  6365 => x"5b90000c",
     6366 => x"5b910008",  6367 => x"5b9d0004",  6368 => x"780e0001",
     6369 => x"39ce3fac",  6370 => x"78040001",  6371 => x"b8406800",
     6372 => x"b8606000",  6373 => x"34020003",  6374 => x"34030002",
     6375 => x"38842e70",  6376 => x"b9c02800",  6377 => x"b8207800",
     6378 => x"35b10021",  6379 => x"fbffec38",  6380 => x"35900021",
     6381 => x"ba200800",  6382 => x"ba001000",  6383 => x"fbffffe1",
     6384 => x"5c200033",  6385 => x"2d81002a",  6386 => x"2dab002a",
     6387 => x"c9615800",  6388 => x"35620001",  6389 => x"34010002",
     6390 => x"54410043",  6391 => x"29e20020",  6392 => x"34030001",
     6393 => x"35a10048",  6394 => x"28420014",  6395 => x"5d63000b",
     6396 => x"fbffffd4",  6397 => x"5c20003c",  6398 => x"78040001",
     6399 => x"b9e00800",  6400 => x"34020003",  6401 => x"34030001",
     6402 => x"38842af8",  6403 => x"b9c02800",  6404 => x"3406008f",
     6405 => x"e000000e",  6406 => x"3403ffff",  6407 => x"358c0048",
     6408 => x"5d63000e",  6409 => x"b9800800",  6410 => x"fbffffc6",
     6411 => x"5c20002e",  6412 => x"78040001",  6413 => x"b9e00800",
     6414 => x"34020003",  6415 => x"34030001",  6416 => x"38842af8",
     6417 => x"b9c02800",  6418 => x"34060098",  6419 => x"fbffec10",
     6420 => x"340b0000",  6421 => x"e0000024",  6422 => x"b9801000",
     6423 => x"fbffffb9",  6424 => x"b8205800",  6425 => x"5c200020",
     6426 => x"78040001",  6427 => x"b9e00800",  6428 => x"34020003",
     6429 => x"34030001",  6430 => x"38842b08",  6431 => x"b9c02800",
     6432 => x"340600a0",  6433 => x"fbffec02",  6434 => x"e0000017",
     6435 => x"41ab001a",  6436 => x"4181001a",  6437 => x"5d61000e",
     6438 => x"41ab001c",  6439 => x"4181001c",  6440 => x"5d61000b",
     6441 => x"41ab001d",  6442 => x"4181001d",  6443 => x"5d610008",
     6444 => x"2da2001e",  6445 => x"2d81001e",  6446 => x"340b0000",
     6447 => x"5c41000a",  6448 => x"41ab0020",  6449 => x"41810020",
     6450 => x"45610003",  6451 => x"c9615800",  6452 => x"e0000005",
     6453 => x"ba200800",  6454 => x"ba001000",  6455 => x"fbffff99",
     6456 => x"b8205800",  6457 => x"b9600800",  6458 => x"2b9d0004",
     6459 => x"2b8b0020",  6460 => x"2b8c001c",  6461 => x"2b8d0018",
     6462 => x"2b8e0014",  6463 => x"2b8f0010",  6464 => x"2b90000c",
     6465 => x"2b910008",  6466 => x"379c0020",  6467 => x"c3a00000",
     6468 => x"379cfffc",  6469 => x"5b9d0004",  6470 => x"34020000",
     6471 => x"34030014",  6472 => x"f8002b88",  6473 => x"2b9d0004",
     6474 => x"379c0004",  6475 => x"c3a00000",  6476 => x"379cfff0",
     6477 => x"5b8b0010",  6478 => x"5b8c000c",  6479 => x"5b8d0008",
     6480 => x"5b9d0004",  6481 => x"b8206800",  6482 => x"28210020",
     6483 => x"282c0014",  6484 => x"282b000c",  6485 => x"28210010",
     6486 => x"0c200000",  6487 => x"34210004",  6488 => x"fbffffec",
     6489 => x"29a10020",  6490 => x"28210010",  6491 => x"34210018",
     6492 => x"fbffffe8",  6493 => x"b9800800",  6494 => x"34020000",
     6495 => x"34030020",  6496 => x"f8002b70",  6497 => x"29610004",
     6498 => x"3402ffa0",  6499 => x"59810000",  6500 => x"29610008",
     6501 => x"59810004",  6502 => x"29610004",  6503 => x"59810010",
     6504 => x"29610008",  6505 => x"59810014",  6506 => x"2d61000e",
     6507 => x"0d810018",  6508 => x"2d610010",  6509 => x"0d81001a",
     6510 => x"41610012",  6511 => x"3181001c",  6512 => x"41610013",
     6513 => x"3181001d",  6514 => x"29a10020",  6515 => x"28210018",
     6516 => x"3022001c",  6517 => x"2b9d0004",  6518 => x"2b8b0010",
     6519 => x"2b8c000c",  6520 => x"2b8d0008",  6521 => x"379c0010",
     6522 => x"c3a00000",  6523 => x"379cff8c",  6524 => x"5b8b0018",
     6525 => x"5b8c0014",  6526 => x"5b8d0010",  6527 => x"5b8e000c",
     6528 => x"5b8f0008",  6529 => x"5b9d0004",  6530 => x"2c22010c",
     6531 => x"b8205800",  6532 => x"340d0000",  6533 => x"340c0001",
     6534 => x"5c400014",  6535 => x"28230000",  6536 => x"b8406800",
     6537 => x"34020006",  6538 => x"5c620010",  6539 => x"fbffffc1",
     6540 => x"29610000",  6541 => x"e0000105",  6542 => x"09820058",
     6543 => x"09a30058",  6544 => x"b9600800",  6545 => x"34420110",
     6546 => x"34630110",  6547 => x"b5621000",  6548 => x"b5631800",
     6549 => x"fbffff42",  6550 => x"48010002",  6551 => x"e0000002",
     6552 => x"b9806800",  6553 => x"358c0001",  6554 => x"2d66010c",
     6555 => x"48ccfff3",  6556 => x"78040001",  6557 => x"b9600800",
     6558 => x"34020003",  6559 => x"34030001",  6560 => x"38842b18",
     6561 => x"b9a02800",  6562 => x"fbffeb81",  6563 => x"1d61010e",
     6564 => x"442d0022",  6565 => x"0d6d010e",  6566 => x"296c0020",
     6567 => x"340f0000",  6568 => x"340e0001",  6569 => x"e0000015",
     6570 => x"29820000",  6571 => x"09c10374",  6572 => x"b4410800",
     6573 => x"2c23010c",  6574 => x"4460000f",  6575 => x"09e40374",
     6576 => x"1c23010e",  6577 => x"b4442000",  6578 => x"1c82010e",
     6579 => x"08630058",  6580 => x"08420058",  6581 => x"34630110",
     6582 => x"b4231800",  6583 => x"34420110",  6584 => x"b4821000",
     6585 => x"fbffff1e",  6586 => x"48010002",  6587 => x"e0000002",
     6588 => x"b9c07800",  6589 => x"35ce0001",  6590 => x"2981000c",
     6591 => x"2c21000c",  6592 => x"482effea",  6593 => x"2981001c",
     6594 => x"442f0004",  6595 => x"34010001",  6596 => x"598f001c",
     6597 => x"59810020",  6598 => x"4162001d",  6599 => x"34010002",
     6600 => x"44410063",  6601 => x"2d61010c",  6602 => x"5c200004",
     6603 => x"29620000",  6604 => x"34010004",  6605 => x"444100c5",
     6606 => x"29610020",  6607 => x"09ac0058",  6608 => x"2821000c",
     6609 => x"4023000a",  6610 => x"4022000b",  6611 => x"40290004",
     6612 => x"40280005",  6613 => x"40270006",  6614 => x"40260007",
     6615 => x"40250008",  6616 => x"40240009",  6617 => x"33830047",
     6618 => x"33890041",  6619 => x"33880042",  6620 => x"33870043",
     6621 => x"33860044",  6622 => x"33850045",  6623 => x"33840046",
     6624 => x"33820048",  6625 => x"2c22000e",  6626 => x"35830110",
     6627 => x"b5631800",  6628 => x"0f82003c",  6629 => x"2c220010",
     6630 => x"0f82003e",  6631 => x"40220012",  6632 => x"3382003a",
     6633 => x"40220013",  6634 => x"0f80004a",  6635 => x"33820040",
     6636 => x"28220004",  6637 => x"5b820068",  6638 => x"28210008",
     6639 => x"37820020",  6640 => x"5b81006c",  6641 => x"b9600800",
     6642 => x"fbfffee5",  6643 => x"4162001d",  6644 => x"34030001",
     6645 => x"44430029",  6646 => x"29620020",  6647 => x"78050001",
     6648 => x"38a53fbc",  6649 => x"2844000c",  6650 => x"1086000e",
     6651 => x"48060004",  6652 => x"48010023",  6653 => x"5c200019",
     6654 => x"e0000006",  6655 => x"48010020",  6656 => x"44200004",
     6657 => x"2c81000c",  6658 => x"5c23000a",  6659 => x"e0000028",
     6660 => x"78040001",  6661 => x"b9600800",  6662 => x"34020003",
     6663 => x"34030001",  6664 => x"38842b38",  6665 => x"fbffeb1a",
     6666 => x"34010002",  6667 => x"e0000087",  6668 => x"29630338",
     6669 => x"2841001c",  6670 => x"4461001d",  6671 => x"b56c1000",
     6672 => x"37810041",  6673 => x"34420131",  6674 => x"5b85001c",
     6675 => x"fbfffebd",  6676 => x"2b85001c",  6677 => x"5c20000c",
     6678 => x"78040001",  6679 => x"b9600800",  6680 => x"34020003",
     6681 => x"34030001",  6682 => x"38842b44",  6683 => x"fbffeb08",
     6684 => x"34010007",  6685 => x"e0000075",  6686 => x"4c200003",
     6687 => x"b9600800",  6688 => x"fbffff2c",  6689 => x"78040001",
     6690 => x"78050001",  6691 => x"b9600800",  6692 => x"34020003",
     6693 => x"34030001",  6694 => x"38842b54",  6695 => x"38a53fbc",
     6696 => x"fbffeafb",  6697 => x"34010006",  6698 => x"e0000068",
     6699 => x"09a30058",  6700 => x"29620020",  6701 => x"b5631800",
     6702 => x"2c64013a",  6703 => x"284c0018",  6704 => x"28410014",
     6705 => x"28420010",  6706 => x"34840001",  6707 => x"0c440000",
     6708 => x"34620150",  6709 => x"28450008",  6710 => x"2844000c",
     6711 => x"58250000",  6712 => x"58240004",  6713 => x"2c420010",
     6714 => x"0c220008",  6715 => x"34620128",  6716 => x"404e0009",
     6717 => x"4045000f",  6718 => x"40440010",  6719 => x"404a000a",
     6720 => x"4049000b",  6721 => x"4048000c",  6722 => x"4047000d",
     6723 => x"4046000e",  6724 => x"302e0010",  6725 => x"30250016",
     6726 => x"302a0011",  6727 => x"30290012",  6728 => x"30280013",
     6729 => x"30270014",  6730 => x"30260015",  6731 => x"30240017",
     6732 => x"28440004",  6733 => x"346e0120",  6734 => x"58240018",
     6735 => x"41c4000a",  6736 => x"3024001c",  6737 => x"40420008",
     6738 => x"3022001d",  6739 => x"4061013c",  6740 => x"3181001c",
     6741 => x"1dc50008",  6742 => x"1d810000",  6743 => x"4425000e",
     6744 => x"78040001",  6745 => x"b9600800",  6746 => x"34020003",
     6747 => x"34030001",  6748 => x"38842b60",  6749 => x"fbffeac6",
     6750 => x"2dc10008",  6751 => x"34020000",  6752 => x"0d810000",
     6753 => x"29610028",  6754 => x"28230004",  6755 => x"b9600800",
     6756 => x"d8600000",  6757 => x"09ad0058",  6758 => x"b56d0800",
     6759 => x"34210141",  6760 => x"4022000b",  6761 => x"20420004",
     6762 => x"7c420000",  6763 => x"59820004",  6764 => x"4022000b",
     6765 => x"20420002",  6766 => x"7c420000",  6767 => x"59820008",
     6768 => x"4022000b",  6769 => x"20420001",  6770 => x"5982000c",
     6771 => x"4022000b",  6772 => x"20420010",  6773 => x"7c420000",
     6774 => x"59820010",  6775 => x"4022000b",  6776 => x"20420020",
     6777 => x"7c420000",  6778 => x"59820014",  6779 => x"4021000b",
     6780 => x"20210008",  6781 => x"7c210000",  6782 => x"59810018",
     6783 => x"78010001",  6784 => x"382149dc",  6785 => x"2824001c",
     6786 => x"44800007",  6787 => x"b56d1000",  6788 => x"b8406800",
     6789 => x"b9600800",  6790 => x"34420144",  6791 => x"35a3011c",
     6792 => x"d8800000",  6793 => x"78040001",  6794 => x"78050001",
     6795 => x"b9600800",  6796 => x"34020003",  6797 => x"34030001",
     6798 => x"38842b74",  6799 => x"38a53fbc",  6800 => x"fbffea93",
     6801 => x"34010009",  6802 => x"2b9d0004",  6803 => x"2b8b0018",
     6804 => x"2b8c0014",  6805 => x"2b8d0010",  6806 => x"2b8e000c",
     6807 => x"2b8f0008",  6808 => x"379c0074",  6809 => x"c3a00000",
     6810 => x"379cffec",  6811 => x"5b8b0014",  6812 => x"5b8c0010",
     6813 => x"5b8d000c",  6814 => x"5b8e0008",  6815 => x"5b9d0004",
     6816 => x"b8406000",  6817 => x"28220024",  6818 => x"b8607000",
     6819 => x"28230070",  6820 => x"2847000c",  6821 => x"28220034",
     6822 => x"b8806800",  6823 => x"b5831800",  6824 => x"342400f8",
     6825 => x"b9a02800",  6826 => x"34060000",  6827 => x"b8205800",
     6828 => x"d8e00000",  6829 => x"78070001",  6830 => x"38e74a14",
     6831 => x"3dc20002",  6832 => x"4c2c000c",  6833 => x"b4e23800",
     6834 => x"28e50000",  6835 => x"78040001",  6836 => x"b9600800",
     6837 => x"34020005",  6838 => x"34030001",  6839 => x"388427ac",
     6840 => x"b9c03000",  6841 => x"fbffea6a",  6842 => x"3401ffff",
     6843 => x"e0000014",  6844 => x"b4e24000",  6845 => x"296600f8",
     6846 => x"296700fc",  6847 => x"29080000",  6848 => x"78040001",
     6849 => x"b9600800",  6850 => x"34020005",  6851 => x"34030001",
     6852 => x"388427cc",  6853 => x"b9802800",  6854 => x"fbffea5d",
     6855 => x"34010001",  6856 => x"5da10003",  6857 => x"29620104",
     6858 => x"44400005",  6859 => x"2961036c",  6860 => x"34210001",
     6861 => x"5961036c",  6862 => x"34010000",  6863 => x"2b9d0004",
     6864 => x"2b8b0014",  6865 => x"2b8c0010",  6866 => x"2b8d000c",
     6867 => x"2b8e0008",  6868 => x"379c0014",  6869 => x"c3a00000",
     6870 => x"379cfff0",  6871 => x"5b8b0010",  6872 => x"5b8c000c",
     6873 => x"5b8d0008",  6874 => x"5b9d0004",  6875 => x"b8205800",
     6876 => x"40410000",  6877 => x"b8406000",  6878 => x"34030002",
     6879 => x"00210004",  6880 => x"356d0320",  6881 => x"3161030c",
     6882 => x"40410000",  6883 => x"2021000f",  6884 => x"3161030d",
     6885 => x"40410001",  6886 => x"2021000f",  6887 => x"3161030e",
     6888 => x"2c410002",  6889 => x"0d610310",  6890 => x"40410004",
     6891 => x"34420006",  6892 => x"31610312",  6893 => x"35610313",
     6894 => x"f8002964",  6895 => x"35820008",  6896 => x"34030004",
     6897 => x"3561031c",  6898 => x"f8002960",  6899 => x"3582000c",
     6900 => x"34030004",  6901 => x"35610318",  6902 => x"f800295c",
     6903 => x"35820014",  6904 => x"34030008",  6905 => x"b9a00800",
     6906 => x"f8002958",  6907 => x"2d81001c",  6908 => x"296202c8",
     6909 => x"34030008",  6910 => x"0d610328",  6911 => x"2d81001e",
     6912 => x"0d61032a",  6913 => x"41810020",  6914 => x"3161032c",
     6915 => x"41810021",  6916 => x"3161032d",  6917 => x"b9a00800",
     6918 => x"f800292b",  6919 => x"3403ffff",  6920 => x"44200015",
     6921 => x"29610020",  6922 => x"28210014",  6923 => x"2c220008",
     6924 => x"4440000a",  6925 => x"b9a01000",  6926 => x"34030008",
     6927 => x"f8002922",  6928 => x"5c200009",  6929 => x"29610020",
     6930 => x"28210014",  6931 => x"2c220008",  6932 => x"2d610328",
     6933 => x"5c410004",  6934 => x"4161001c",  6935 => x"38210001",
     6936 => x"e0000003",  6937 => x"4161001c",  6938 => x"202100fe",
     6939 => x"3161001c",  6940 => x"34030000",  6941 => x"b8600800",
     6942 => x"2b9d0004",  6943 => x"2b8b0010",  6944 => x"2b8c000c",
     6945 => x"2b8d0008",  6946 => x"379c0010",  6947 => x"c3a00000",
     6948 => x"379cfff4",  6949 => x"5b8b000c",  6950 => x"5b8c0008",
     6951 => x"5b9d0004",  6952 => x"30400000",  6953 => x"b8206000",
     6954 => x"282102c8",  6955 => x"b8405800",  6956 => x"34030008",
     6957 => x"4021000e",  6958 => x"30410001",  6959 => x"29810020",
     6960 => x"2821000c",  6961 => x"40210014",  6962 => x"30410004",
     6963 => x"34010002",  6964 => x"30410006",  6965 => x"34410008",
     6966 => x"34020000",  6967 => x"f8002999",  6968 => x"298202c8",
     6969 => x"35610014",  6970 => x"34030008",  6971 => x"f8002917",
     6972 => x"298102c8",  6973 => x"2c210008",  6974 => x"0d61001c",
     6975 => x"3401007f",  6976 => x"31610021",  6977 => x"2b9d0004",
     6978 => x"2b8b000c",  6979 => x"2b8c0008",  6980 => x"379c000c",
     6981 => x"c3a00000",  6982 => x"2c230022",  6983 => x"0c430004",
     6984 => x"28230024",  6985 => x"58430000",  6986 => x"28210028",
     6987 => x"58410008",  6988 => x"c3a00000",  6989 => x"379cfff4",
     6990 => x"5b8b000c",  6991 => x"5b8c0008",  6992 => x"5b9d0004",
     6993 => x"b8205800",  6994 => x"2c210022",  6995 => x"b8406000",
     6996 => x"34030008",  6997 => x"0c410004",  6998 => x"29610024",
     6999 => x"58410000",  7000 => x"29610028",  7001 => x"58410008",
     7002 => x"2d61002c",  7003 => x"0c41000c",  7004 => x"4161002f",
     7005 => x"3041000e",  7006 => x"41610030",  7007 => x"30410010",
     7008 => x"41610031",  7009 => x"30410011",  7010 => x"2d610032",
     7011 => x"0c410012",  7012 => x"41610034",  7013 => x"30410014",
     7014 => x"34410015",  7015 => x"35620035",  7016 => x"f80028ea",
     7017 => x"2d61003d",  7018 => x"0d81001e",  7019 => x"4161003f",
     7020 => x"31810020",  7021 => x"78010001",  7022 => x"382149dc",
     7023 => x"28230030",  7024 => x"44600004",  7025 => x"b9600800",
     7026 => x"b9801000",  7027 => x"d8600000",  7028 => x"2b9d0004",
     7029 => x"2b8b000c",  7030 => x"2b8c0008",  7031 => x"379c000c",
     7032 => x"c3a00000",  7033 => x"2c230022",  7034 => x"0c430004",
     7035 => x"28230024",  7036 => x"58430000",  7037 => x"28210028",
     7038 => x"58410008",  7039 => x"c3a00000",  7040 => x"379cfff4",
     7041 => x"5b8b000c",  7042 => x"5b8c0008",  7043 => x"5b9d0004",
     7044 => x"b8205800",  7045 => x"2c210022",  7046 => x"b8406000",
     7047 => x"34030008",  7048 => x"0c410004",  7049 => x"29610024",
     7050 => x"58410000",  7051 => x"29610028",  7052 => x"58410008",
     7053 => x"3441000c",  7054 => x"3562002c",  7055 => x"f80028c3",
     7056 => x"2d610034",  7057 => x"0d810014",  7058 => x"2b9d0004",
     7059 => x"2b8b000c",  7060 => x"2b8c0008",  7061 => x"379c000c",
     7062 => x"c3a00000",  7063 => x"379cfff4",  7064 => x"5b8b000c",
     7065 => x"5b8c0008",  7066 => x"5b9d0004",  7067 => x"282b003c",
     7068 => x"b8206000",  7069 => x"34020000",  7070 => x"41610000",
     7071 => x"3403000a",  7072 => x"202100f0",  7073 => x"3821000b",
     7074 => x"31610000",  7075 => x"34010040",  7076 => x"0d610002",
     7077 => x"2d810306",  7078 => x"34210001",  7079 => x"2021ffff",
     7080 => x"0d810306",  7081 => x"0d61001e",  7082 => x"34010005",
     7083 => x"31610020",  7084 => x"298102c8",  7085 => x"4021000b",
     7086 => x"31610021",  7087 => x"35610022",  7088 => x"f8002920",
     7089 => x"29810020",  7090 => x"34030008",  7091 => x"28220018",
     7092 => x"28210014",  7093 => x"2c420000",  7094 => x"0d62002c",
     7095 => x"4021001c",  7096 => x"3161002f",  7097 => x"29810020",
     7098 => x"28210014",  7099 => x"40210018",  7100 => x"31610030",
     7101 => x"29810020",  7102 => x"28210014",  7103 => x"40210019",
     7104 => x"31610031",  7105 => x"29810020",  7106 => x"28210014",
     7107 => x"2c22001a",  7108 => x"0d620032",  7109 => x"4021001d",
     7110 => x"31610034",  7111 => x"29810020",  7112 => x"28220014",
     7113 => x"35610035",  7114 => x"34420010",  7115 => x"f8002887",
     7116 => x"29810020",  7117 => x"28220010",  7118 => x"28210018",
     7119 => x"2c420000",  7120 => x"0d62003d",  7121 => x"4021001c",
     7122 => x"34020040",  7123 => x"3161003f",  7124 => x"78010001",
     7125 => x"382149dc",  7126 => x"2823002c",  7127 => x"44600004",
     7128 => x"b9800800",  7129 => x"d8600000",  7130 => x"b8201000",
     7131 => x"b9800800",  7132 => x"3403000b",  7133 => x"34040000",
     7134 => x"fbfffebc",  7135 => x"2b9d0004",  7136 => x"2b8b000c",
     7137 => x"2b8c0008",  7138 => x"379c000c",  7139 => x"c3a00000",
     7140 => x"379cffc8",  7141 => x"5b8b0018",  7142 => x"5b8c0014",
     7143 => x"5b8d0010",  7144 => x"5b8e000c",  7145 => x"5b8f0008",
     7146 => x"5b9d0004",  7147 => x"28220028",  7148 => x"378c001c",
     7149 => x"b8205800",  7150 => x"28430000",  7151 => x"b9801000",
     7152 => x"378f0030",  7153 => x"d8600000",  7154 => x"b9800800",
     7155 => x"b9e01000",  7156 => x"f8000103",  7157 => x"296c003c",
     7158 => x"340efff0",  7159 => x"340d002c",  7160 => x"41810000",
     7161 => x"0d8d0002",  7162 => x"34020000",  7163 => x"a02e0800",
     7164 => x"31810000",  7165 => x"2d6102f0",  7166 => x"34030008",
     7167 => x"34210001",  7168 => x"2021ffff",  7169 => x"0d6102f0",
     7170 => x"31800020",  7171 => x"0d81001e",  7172 => x"296102c8",
     7173 => x"4021000d",  7174 => x"31810021",  7175 => x"35810008",
     7176 => x"f80028c8",  7177 => x"2f810034",  7178 => x"3402002c",
     7179 => x"34030000",  7180 => x"0d810022",  7181 => x"2b810030",
     7182 => x"34040001",  7183 => x"59810024",  7184 => x"2b810038",
     7185 => x"59810028",  7186 => x"b9600800",  7187 => x"fbfffe87",
     7188 => x"5c200023",  7189 => x"29610020",  7190 => x"356c00f8",
     7191 => x"b9801000",  7192 => x"28230008",  7193 => x"b9800800",
     7194 => x"34630018",  7195 => x"f8000101",  7196 => x"b9e01000",
     7197 => x"b9800800",  7198 => x"f80000d9",  7199 => x"2961003c",
     7200 => x"34030008",  7201 => x"34040000",  7202 => x"40220000",
     7203 => x"0c2d0002",  7204 => x"a04e7000",  7205 => x"39ce0008",
     7206 => x"302e0000",  7207 => x"2d6202f0",  7208 => x"0c22001e",
     7209 => x"34020002",  7210 => x"30220020",  7211 => x"296202c8",
     7212 => x"4042000d",  7213 => x"30220021",  7214 => x"2f820034",
     7215 => x"0c220022",  7216 => x"2b820030",  7217 => x"58220024",
     7218 => x"2b820038",  7219 => x"58220028",  7220 => x"b9600800",
     7221 => x"3402002c",  7222 => x"fbfffe64",  7223 => x"2b9d0004",
     7224 => x"2b8b0018",  7225 => x"2b8c0014",  7226 => x"2b8d0010",
     7227 => x"2b8e000c",  7228 => x"2b8f0008",  7229 => x"379c0038",
     7230 => x"c3a00000",  7231 => x"379cffd4",  7232 => x"5b8b000c",
     7233 => x"5b8c0008",  7234 => x"5b9d0004",  7235 => x"28220028",
     7236 => x"378b0010",  7237 => x"b8206000",  7238 => x"28430000",
     7239 => x"b9601000",  7240 => x"d8600000",  7241 => x"37820024",
     7242 => x"b9600800",  7243 => x"f80000ac",  7244 => x"298b003c",
     7245 => x"34020000",  7246 => x"34030008",  7247 => x"41610000",
     7248 => x"202100f0",  7249 => x"38210001",  7250 => x"31610000",
     7251 => x"3401002c",  7252 => x"0d610002",  7253 => x"2d8102f2",
     7254 => x"34210001",  7255 => x"2021ffff",  7256 => x"0d8102f2",
     7257 => x"0d61001e",  7258 => x"34010001",  7259 => x"31610020",
     7260 => x"3401007f",  7261 => x"31610021",  7262 => x"35610008",
     7263 => x"f8002871",  7264 => x"2f810028",  7265 => x"3402002c",
     7266 => x"34030001",  7267 => x"0d610022",  7268 => x"2b810024",
     7269 => x"34040001",  7270 => x"59610024",  7271 => x"2b81002c",
     7272 => x"59610028",  7273 => x"b9800800",  7274 => x"fbfffe30",
     7275 => x"2b9d0004",  7276 => x"2b8b000c",  7277 => x"2b8c0008",
     7278 => x"379c002c",  7279 => x"c3a00000",  7280 => x"379cffe8",
     7281 => x"5b8b000c",  7282 => x"5b8c0008",  7283 => x"5b9d0004",
     7284 => x"b8206000",  7285 => x"b8400800",  7286 => x"37820010",
     7287 => x"f8000080",  7288 => x"298b003c",  7289 => x"34020000",
     7290 => x"34030008",  7291 => x"41610000",  7292 => x"202100f0",
     7293 => x"38210009",  7294 => x"31610000",  7295 => x"34010036",
     7296 => x"0d610002",  7297 => x"41810312",  7298 => x"31610004",
     7299 => x"35610008",  7300 => x"f800284c",  7301 => x"2981031c",
     7302 => x"35820320",  7303 => x"34030008",  7304 => x"59610008",
     7305 => x"29810318",  7306 => x"5961000c",  7307 => x"2d81032a",
     7308 => x"0d61001e",  7309 => x"34010003",  7310 => x"31610020",
     7311 => x"298102c8",  7312 => x"4021000a",  7313 => x"31610021",
     7314 => x"2f810014",  7315 => x"0d610022",  7316 => x"2b810010",
     7317 => x"59610024",  7318 => x"2b810018",  7319 => x"59610028",
     7320 => x"3561002c",  7321 => x"f80027b9",  7322 => x"2d810328",
     7323 => x"34020036",  7324 => x"34030009",  7325 => x"0d610034",
     7326 => x"34040000",  7327 => x"b9800800",  7328 => x"fbfffdfa",
     7329 => x"2b9d0004",  7330 => x"2b8b000c",  7331 => x"2b8c0008",
     7332 => x"379c0018",  7333 => x"c3a00000",  7334 => x"379cfff0",
     7335 => x"5b8b0010",  7336 => x"5b8c000c",  7337 => x"5b8d0008",
     7338 => x"5b9d0004",  7339 => x"78030001",  7340 => x"282d0004",
     7341 => x"38633ce0",  7342 => x"28620000",  7343 => x"b8205800",
     7344 => x"b9a00800",  7345 => x"f80026f3",  7346 => x"78030001",
     7347 => x"296c0000",  7348 => x"38633ce0",  7349 => x"28620000",
     7350 => x"b42c6000",  7351 => x"596c0000",  7352 => x"b9a00800",
     7353 => x"f8002718",  7354 => x"59610004",  7355 => x"4c0c0007",
     7356 => x"4c20000f",  7357 => x"358cffff",  7358 => x"78030001",
     7359 => x"596c0000",  7360 => x"38633ce0",  7361 => x"e0000007",
     7362 => x"45800009",  7363 => x"4c010008",  7364 => x"358c0001",
     7365 => x"78030001",  7366 => x"596c0000",  7367 => x"38633cf0",
     7368 => x"28620000",  7369 => x"b4220800",  7370 => x"59610004",
     7371 => x"2b9d0004",  7372 => x"2b8b0010",  7373 => x"2b8c000c",
     7374 => x"2b8d0008",  7375 => x"379c0010",  7376 => x"c3a00000",
     7377 => x"379cffe8",  7378 => x"5b8b0008",  7379 => x"5b9d0004",
     7380 => x"5b82000c",  7381 => x"5b830010",  7382 => x"5b830014",
     7383 => x"5b820018",  7384 => x"b8205800",  7385 => x"4c600006",
     7386 => x"78010001",  7387 => x"78020001",  7388 => x"38212bf4",
     7389 => x"38423fd0",  7390 => x"f8000e93",  7391 => x"2b810018",
     7392 => x"38028000",  7393 => x"2b830014",  7394 => x"b4221000",
     7395 => x"f4220800",  7396 => x"00420010",  7397 => x"b4230800",
     7398 => x"3c230010",  7399 => x"00210010",  7400 => x"b8431000",
     7401 => x"78030001",  7402 => x"38633ce0",  7403 => x"5b820018",
     7404 => x"28620000",  7405 => x"5b810014",  7406 => x"37810014",
     7407 => x"fbffec79",  7408 => x"59610004",  7409 => x"2b810018",
     7410 => x"59610000",  7411 => x"2b9d0004",  7412 => x"2b8b0008",
     7413 => x"379c0018",  7414 => x"c3a00000",  7415 => x"379cfffc",
     7416 => x"5b9d0004",  7417 => x"28230000",  7418 => x"48030003",
     7419 => x"28210004",  7420 => x"4c200006",  7421 => x"78010001",
     7422 => x"38212c20",  7423 => x"f8000e72",  7424 => x"3401ffff",
     7425 => x"e0000005",  7426 => x"58410008",  7427 => x"58430000",
     7428 => x"0c400004",  7429 => x"34010000",  7430 => x"2b9d0004",
     7431 => x"379c0004",  7432 => x"c3a00000",  7433 => x"379cfffc",
     7434 => x"5b9d0004",  7435 => x"78050001",  7436 => x"38a53cf4",
     7437 => x"28430000",  7438 => x"28a40000",  7439 => x"54640006",
     7440 => x"28420008",  7441 => x"58230000",  7442 => x"58220004",
     7443 => x"34010000",  7444 => x"e0000005",  7445 => x"78010001",
     7446 => x"38212c5c",  7447 => x"f8000e5a",  7448 => x"3401ffff",
     7449 => x"2b9d0004",  7450 => x"379c0004",  7451 => x"c3a00000",
     7452 => x"379cfffc",  7453 => x"5b9d0004",  7454 => x"28660000",
     7455 => x"28450000",  7456 => x"28630004",  7457 => x"28420004",
     7458 => x"b4c52800",  7459 => x"58250000",  7460 => x"b4621000",
     7461 => x"58220004",  7462 => x"fbffff80",  7463 => x"2b9d0004",
     7464 => x"379c0004",  7465 => x"c3a00000",  7466 => x"379cfffc",
     7467 => x"5b9d0004",  7468 => x"28460000",  7469 => x"28650000",
     7470 => x"c8c52800",  7471 => x"58250000",  7472 => x"28450004",
     7473 => x"28620004",  7474 => x"c8a21000",  7475 => x"58220004",
     7476 => x"fbffff72",  7477 => x"2b9d0004",  7478 => x"379c0004",
     7479 => x"c3a00000",  7480 => x"379cfffc",  7481 => x"5b9d0004",
     7482 => x"78040001",  7483 => x"38843cf8",  7484 => x"28230000",
     7485 => x"28820000",  7486 => x"a0621000",  7487 => x"4c400005",
     7488 => x"3442ffff",  7489 => x"3404fffe",  7490 => x"b8441000",
     7491 => x"34420001",  7492 => x"78050001",  7493 => x"38a53ce0",
     7494 => x"28a40000",  7495 => x"88441000",  7496 => x"28240004",
     7497 => x"b4441000",  7498 => x"0064001f",  7499 => x"b4831800",
     7500 => x"14630001",  7501 => x"58230000",  7502 => x"0043001f",
     7503 => x"b4621000",  7504 => x"14420001",  7505 => x"58220004",
     7506 => x"fbffff54",  7507 => x"2b9d0004",  7508 => x"379c0004",
     7509 => x"c3a00000",  7510 => x"379cfff8",  7511 => x"5b8b0008",
     7512 => x"5b9d0004",  7513 => x"28250000",  7514 => x"78030001",
     7515 => x"b8201000",  7516 => x"38632cac",  7517 => x"4805000a",
     7518 => x"78030001",  7519 => x"38631c40",  7520 => x"5ca00007",
     7521 => x"28210004",  7522 => x"78030001",  7523 => x"38632cac",
     7524 => x"48a10003",  7525 => x"78030001",  7526 => x"38631c40",
     7527 => x"28410004",  7528 => x"14a4001f",  7529 => x"780b0001",
     7530 => x"1426001f",  7531 => x"98853800",  7532 => x"396b5214",
     7533 => x"98c12800",  7534 => x"78020001",  7535 => x"b9600800",
     7536 => x"38422cb0",  7537 => x"c8e42000",  7538 => x"c8a62800",
     7539 => x"f8000df0",  7540 => x"b9600800",  7541 => x"2b9d0004",
     7542 => x"2b8b0008",  7543 => x"379c0008",  7544 => x"c3a00000",
     7545 => x"379cfff8",  7546 => x"5b8b0008",  7547 => x"5b9d0004",
     7548 => x"28220020",  7549 => x"28240028",  7550 => x"b8205800",
     7551 => x"28430004",  7552 => x"58600038",  7553 => x"28430014",
     7554 => x"0c20010c",  7555 => x"0c600008",  7556 => x"28830014",
     7557 => x"44600013",  7558 => x"d8600000",  7559 => x"3402ffff",
     7560 => x"5c220008",  7561 => x"78040001",  7562 => x"b9600800",
     7563 => x"34020004",  7564 => x"34030001",  7565 => x"38842cbc",
     7566 => x"fbffe795",  7567 => x"34010000",  7568 => x"29620020",
     7569 => x"c8010800",  7570 => x"3c21000a",  7571 => x"28420004",
     7572 => x"1423001f",  7573 => x"5841002c",  7574 => x"58430028",
     7575 => x"e000000d",  7576 => x"28420008",  7577 => x"28420038",
     7578 => x"20420001",  7579 => x"5c430005",  7580 => x"28840008",
     7581 => x"34020000",  7582 => x"34030000",  7583 => x"d8800000",
     7584 => x"29610020",  7585 => x"28210004",  7586 => x"58200028",
     7587 => x"5820002c",  7588 => x"29610020",  7589 => x"78040001",
     7590 => x"34020004",  7591 => x"28260004",  7592 => x"34030001",
     7593 => x"b9600800",  7594 => x"28c50028",  7595 => x"28c6002c",
     7596 => x"38842cd8",  7597 => x"fbffe776",  7598 => x"2b9d0004",
     7599 => x"2b8b0008",  7600 => x"379c0008",  7601 => x"c3a00000",
     7602 => x"379cfff0",  7603 => x"5b8b0010",  7604 => x"5b8c000c",
     7605 => x"5b8d0008",  7606 => x"5b9d0004",  7607 => x"b8205800",
     7608 => x"28210020",  7609 => x"35620094",  7610 => x"35630080",
     7611 => x"282d0004",  7612 => x"356c00d0",  7613 => x"b9a00800",
     7614 => x"fbffff6c",  7615 => x"b9a01000",  7616 => x"b9801800",
     7617 => x"b9a00800",  7618 => x"fbffff68",  7619 => x"b9800800",
     7620 => x"fbffff92",  7621 => x"78040001",  7622 => x"b8202800",
     7623 => x"34020004",  7624 => x"b9600800",  7625 => x"34030003",
     7626 => x"38842cf8",  7627 => x"fbffe758",  7628 => x"2b9d0004",
     7629 => x"2b8b0010",  7630 => x"2b8c000c",  7631 => x"2b8d0008",
     7632 => x"379c0010",  7633 => x"c3a00000",  7634 => x"379cffb8",
     7635 => x"5b8b0024",  7636 => x"5b8c0020",  7637 => x"5b8d001c",
     7638 => x"5b8e0018",  7639 => x"5b8f0014",  7640 => x"5b900010",
     7641 => x"5b91000c",  7642 => x"5b920008",  7643 => x"5b9d0004",
     7644 => x"28220020",  7645 => x"b8205800",  7646 => x"284d0004",
     7647 => x"284c0010",  7648 => x"28220080",  7649 => x"5c400008",
     7650 => x"28230084",  7651 => x"5c620006",  7652 => x"78040001",
     7653 => x"34020004",  7654 => x"34030002",  7655 => x"38842d10",
     7656 => x"e000006e",  7657 => x"35af0014",  7658 => x"357000bc",
     7659 => x"357100a8",  7660 => x"b9e00800",  7661 => x"ba001000",
     7662 => x"ba201800",  7663 => x"fbffff3b",  7664 => x"357200d0",
     7665 => x"b9e01000",  7666 => x"ba401800",  7667 => x"b9e00800",
     7668 => x"fbffff36",  7669 => x"ba400800",  7670 => x"fbffff60",
     7671 => x"78040001",  7672 => x"b8202800",  7673 => x"34020004",
     7674 => x"34030003",  7675 => x"38842d30",  7676 => x"b9600800",
     7677 => x"fbffe726",  7678 => x"35610080",  7679 => x"fbffff57",
     7680 => x"78040001",  7681 => x"b8202800",  7682 => x"34020004",
     7683 => x"34030002",  7684 => x"38842d48",  7685 => x"b9600800",
     7686 => x"fbffe71d",  7687 => x"35610094",  7688 => x"fbffff4e",
     7689 => x"78040001",  7690 => x"b8202800",  7691 => x"34020004",
     7692 => x"34030002",  7693 => x"38842d50",  7694 => x"b9600800",
     7695 => x"fbffe714",  7696 => x"ba200800",  7697 => x"fbffff45",
     7698 => x"78040001",  7699 => x"b8202800",  7700 => x"34020004",
     7701 => x"34030002",  7702 => x"38842d58",  7703 => x"b9600800",
     7704 => x"fbffe70b",  7705 => x"ba000800",  7706 => x"fbffff3c",
     7707 => x"78040001",  7708 => x"b8202800",  7709 => x"34020004",
     7710 => x"34030002",  7711 => x"38842d60",  7712 => x"b9600800",
     7713 => x"fbffe702",  7714 => x"b9a00800",  7715 => x"fbffff33",
     7716 => x"78040001",  7717 => x"b8202800",  7718 => x"34020004",
     7719 => x"34030001",  7720 => x"38842d68",  7721 => x"b9600800",
     7722 => x"fbffe6f9",  7723 => x"b9e00800",  7724 => x"fbffff2a",
     7725 => x"78040001",  7726 => x"b8202800",  7727 => x"38842d80",
     7728 => x"b9600800",  7729 => x"34020004",  7730 => x"34030001",
     7731 => x"fbffe6f0",  7732 => x"29610020",  7733 => x"358e0018",
     7734 => x"28220004",  7735 => x"b9c00800",  7736 => x"34430014",
     7737 => x"fbfffee3",  7738 => x"b9c00800",  7739 => x"fbfffefd",
     7740 => x"b9c00800",  7741 => x"fbffff19",  7742 => x"78040001",
     7743 => x"b8202800",  7744 => x"34020004",  7745 => x"b9600800",
     7746 => x"34030001",  7747 => x"38842d98",  7748 => x"fbffe6df",
     7749 => x"29610020",  7750 => x"28220010",  7751 => x"28260004",
     7752 => x"28420018",  7753 => x"5c400142",  7754 => x"28210008",
     7755 => x"28270030",  7756 => x"44e2013c",  7757 => x"28c20000",
     7758 => x"5c400003",  7759 => x"28c30014",  7760 => x"44620008",
     7761 => x"78040001",  7762 => x"b9600800",  7763 => x"34020004",
     7764 => x"34030001",  7765 => x"38842dac",  7766 => x"fbffe6cd",
     7767 => x"e0000134",  7768 => x"28c50004",  7769 => x"48a70003",
     7770 => x"28c20018",  7771 => x"4ce2012d",  7772 => x"28c60018",
     7773 => x"78040001",  7774 => x"b9600800",  7775 => x"34020004",
     7776 => x"34030001",  7777 => x"38842dd8",  7778 => x"fbffe6c1",
     7779 => x"e0000128",  7780 => x"2982001c",  7781 => x"59a20034",
     7782 => x"1c220040",  7783 => x"29a10034",  7784 => x"3444ffff",
     7785 => x"1423001f",  7786 => x"98612800",  7787 => x"c8a32800",
     7788 => x"3403001f",  7789 => x"c8621800",  7790 => x"94a33800",
     7791 => x"34820001",  7792 => x"34630001",  7793 => x"3484ffff",
     7794 => x"5ce0fffc",  7795 => x"34030001",  7796 => x"bc621000",
     7797 => x"4c460002",  7798 => x"59a20038",  7799 => x"29a30038",
     7800 => x"4c620003",  7801 => x"34630001",  7802 => x"59a30038",
     7803 => x"2982001c",  7804 => x"4c400002",  7805 => x"5981001c",
     7806 => x"2982001c",  7807 => x"4c400002",  7808 => x"5980001c",
     7809 => x"2985001c",  7810 => x"08210003",  7811 => x"4c25000d",
     7812 => x"78040001",  7813 => x"b9600800",  7814 => x"34020004",
     7815 => x"34030001",  7816 => x"38842e1c",  7817 => x"fbffe69a",
     7818 => x"29a10034",  7819 => x"29a20038",  7820 => x"3c210001",
     7821 => x"34420001",  7822 => x"b4410800",  7823 => x"5981001c",
     7824 => x"29af0038",  7825 => x"29a20034",  7826 => x"35900004",
     7827 => x"35e1ffff",  7828 => x"88220800",  7829 => x"2982001c",
     7830 => x"b4220800",  7831 => x"b9e01000",  7832 => x"f800250c",
     7833 => x"59a10034",  7834 => x"78040001",  7835 => x"b8203000",
     7836 => x"b9e02800",  7837 => x"38842e34",  7838 => x"5981001c",
     7839 => x"34020004",  7840 => x"b9600800",  7841 => x"34030001",
     7842 => x"fbffe681",  7843 => x"b9a01000",  7844 => x"b9c01800",
     7845 => x"ba000800",  7846 => x"fbfffe84",  7847 => x"ba000800",
     7848 => x"fbfffeae",  7849 => x"78040001",  7850 => x"b8202800",
     7851 => x"34020004",  7852 => x"b9600800",  7853 => x"34030001",
     7854 => x"38842e58",  7855 => x"fbffe674",  7856 => x"296f0020",
     7857 => x"29e10008",  7858 => x"2825002c",  7859 => x"44a00011",
     7860 => x"29820004",  7861 => x"44400007",  7862 => x"78040001",
     7863 => x"b9600800",  7864 => x"34020004",  7865 => x"34030001",
     7866 => x"38842e74",  7867 => x"e3ffff9b",  7868 => x"29820008",
     7869 => x"4ca20007",  7870 => x"78040001",  7871 => x"b9600800",
     7872 => x"34020004",  7873 => x"34030001",  7874 => x"38842ea4",
     7875 => x"e00000c3",  7876 => x"29820004",  7877 => x"44400031",
     7878 => x"28220038",  7879 => x"20410001",  7880 => x"5c2000c3",
     7881 => x"20420002",  7882 => x"5c410019",  7883 => x"296300c4",
     7884 => x"296200c8",  7885 => x"296100cc",  7886 => x"5b830030",
     7887 => x"29e30010",  7888 => x"296500bc",  7889 => x"296400c0",
     7890 => x"378c0028",  7891 => x"5b820034",  7892 => x"5b810038",
     7893 => x"b9801000",  7894 => x"b9800800",  7895 => x"34630018",
     7896 => x"5b850028",  7897 => x"5b84002c",  7898 => x"fbfffe42",
     7899 => x"29610028",  7900 => x"b9801000",  7901 => x"28230004",
     7902 => x"b9600800",  7903 => x"d8600000",  7904 => x"b9600800",
     7905 => x"fbfffe98",  7906 => x"e00000a9",  7907 => x"29820008",
     7908 => x"78030001",  7909 => x"38633cfc",  7910 => x"28610000",
     7911 => x"ec021000",  7912 => x"78050001",  7913 => x"c8021000",
     7914 => x"38a53d00",  7915 => x"a0411000",  7916 => x"28a10000",
     7917 => x"b4411000",  7918 => x"29610028",  7919 => x"c8021000",
     7920 => x"28230010",  7921 => x"5c600002",  7922 => x"2823000c",
     7923 => x"b9600800",  7924 => x"d8600000",  7925 => x"e0000096",
     7926 => x"29830008",  7927 => x"29ed0004",  7928 => x"78050001",
     7929 => x"1462001f",  7930 => x"29b0002c",  7931 => x"00640016",
     7932 => x"3c63000a",  7933 => x"29ae0028",  7934 => x"3c42000a",
     7935 => x"b4708000",  7936 => x"b8821000",  7937 => x"f4701800",
     7938 => x"b44e1000",  7939 => x"b4627000",  7940 => x"1c22003e",
     7941 => x"38a53d00",  7942 => x"28a40000",  7943 => x"1441001f",
     7944 => x"34030000",  7945 => x"59ae0028",  7946 => x"59b0002c",
     7947 => x"f8002472",  7948 => x"00430016",  7949 => x"3c21000a",
     7950 => x"3c42000a",  7951 => x"b8610800",  7952 => x"49c1000b",
     7953 => x"5dc10002",  7954 => x"56020009",  7955 => x"c8021000",
     7956 => x"7c430000",  7957 => x"c8010800",  7958 => x"c8230800",
     7959 => x"482e0004",  7960 => x"5c2e0005",  7961 => x"54500002",
     7962 => x"e0000003",  7963 => x"59a10028",  7964 => x"59a2002c",
     7965 => x"29a10028",  7966 => x"29a2002c",  7967 => x"48200003",
     7968 => x"5c200004",  7969 => x"44410003",  7970 => x"340d0000",
     7971 => x"e0000002",  7972 => x"340dffff",  7973 => x"5b810044",
     7974 => x"5b820048",  7975 => x"45a00007",  7976 => x"c8021000",
     7977 => x"7c430000",  7978 => x"c8010800",  7979 => x"c8230800",
     7980 => x"5b810044",  7981 => x"5b820048",  7982 => x"29e20008",
     7983 => x"37810044",  7984 => x"1c42003e",  7985 => x"fbffea37",
     7986 => x"45a00009",  7987 => x"2b810048",  7988 => x"2b820044",
     7989 => x"c8010800",  7990 => x"7c230000",  7991 => x"c8021000",
     7992 => x"c8431000",  7993 => x"5b820044",  7994 => x"5b810048",
     7995 => x"29820008",  7996 => x"1441001f",  7997 => x"00430016",
     7998 => x"3c21000a",  7999 => x"ec026000",  8000 => x"3c42000a",
     8001 => x"b8610800",  8002 => x"c80c6000",  8003 => x"5b81003c",
     8004 => x"5b820040",  8005 => x"45800007",  8006 => x"c8021000",
     8007 => x"7c430000",  8008 => x"c8010800",  8009 => x"c8230800",
     8010 => x"5b81003c",  8011 => x"5b820040",  8012 => x"29610020",
     8013 => x"28220008",  8014 => x"3781003c",  8015 => x"1c42003c",
     8016 => x"fbffea18",  8017 => x"45800009",  8018 => x"2b810040",
     8019 => x"2b82003c",  8020 => x"c8010800",  8021 => x"7c230000",
     8022 => x"c8021000",  8023 => x"c8431000",  8024 => x"5b82003c",
     8025 => x"5b810040",  8026 => x"2b830048",  8027 => x"2b820040",
     8028 => x"2b81003c",  8029 => x"2b840044",  8030 => x"b4621000",
     8031 => x"f4621800",  8032 => x"b4810800",  8033 => x"b4610800",
     8034 => x"48200003",  8035 => x"5c200006",  8036 => x"44410005",
     8037 => x"3c210016",  8038 => x"0042000a",  8039 => x"b8221000",
     8040 => x"e0000009",  8041 => x"c8021000",  8042 => x"7c430000",
     8043 => x"c8010800",  8044 => x"c8230800",  8045 => x"3c210016",
     8046 => x"0042000a",  8047 => x"b8221000",  8048 => x"c8021000",
     8049 => x"29610020",  8050 => x"28210008",  8051 => x"28250038",
     8052 => x"20a50001",  8053 => x"5ca00008",  8054 => x"29640028",
     8055 => x"c8021000",  8056 => x"28830010",  8057 => x"5c650002",
     8058 => x"2883000c",  8059 => x"b9600800",  8060 => x"d8600000",
     8061 => x"29610020",  8062 => x"78040001",  8063 => x"34020004",
     8064 => x"28210004",  8065 => x"34030002",  8066 => x"38842ee0",
     8067 => x"2825002c",  8068 => x"b9600800",  8069 => x"14a5000a",
     8070 => x"fbffe59d",  8071 => x"e0000004",  8072 => x"29a60038",
     8073 => x"4c06fedb",  8074 => x"e3fffedc",  8075 => x"2b9d0004",
     8076 => x"2b8b0024",  8077 => x"2b8c0020",  8078 => x"2b8d001c",
     8079 => x"2b8e0018",  8080 => x"2b8f0014",  8081 => x"2b900010",
     8082 => x"2b91000c",  8083 => x"2b920008",  8084 => x"379c0048",
     8085 => x"c3a00000",  8086 => x"379cfffc",  8087 => x"5b9d0004",
     8088 => x"78030001",  8089 => x"3c420002",  8090 => x"38634a54",
     8091 => x"b4622800",  8092 => x"28a50000",  8093 => x"78040001",
     8094 => x"34020006",  8095 => x"34030001",  8096 => x"38842ef8",
     8097 => x"fbffe582",  8098 => x"2b9d0004",  8099 => x"379c0004",
     8100 => x"c3a00000",  8101 => x"379cfff0",  8102 => x"5b8b0010",
     8103 => x"5b8c000c",  8104 => x"5b8d0008",  8105 => x"5b9d0004",
     8106 => x"b8205800",  8107 => x"78010001",  8108 => x"3821522c",
     8109 => x"b8406800",  8110 => x"28220000",  8111 => x"5c400005",
     8112 => x"29620020",  8113 => x"2844000c",  8114 => x"28820008",
     8115 => x"58220000",  8116 => x"78040001",  8117 => x"78010001",
     8118 => x"3884522c",  8119 => x"38213d04",  8120 => x"28260000",
     8121 => x"28850000",  8122 => x"340c0190",  8123 => x"bd836000",
     8124 => x"88a62800",  8125 => x"b9801000",  8126 => x"34a53039",
     8127 => x"00a10010",  8128 => x"88a62800",  8129 => x"202107ff",
     8130 => x"34a53039",  8131 => x"58850000",  8132 => x"00a50010",
     8133 => x"3c24000a",  8134 => x"20a103ff",  8135 => x"b8240800",
     8136 => x"f8002439",  8137 => x"3d820001",  8138 => x"b4221000",
     8139 => x"29610028",  8140 => x"28230018",  8141 => x"b9600800",
     8142 => x"d8600000",  8143 => x"35a200b2",  8144 => x"3c420002",
     8145 => x"b5625800",  8146 => x"59610004",  8147 => x"2b9d0004",
     8148 => x"2b8b0010",  8149 => x"2b8c000c",  8150 => x"2b8d0008",
     8151 => x"379c0010",  8152 => x"c3a00000",  8153 => x"379cfff0",
     8154 => x"5b8b0010",  8155 => x"5b8c000c",  8156 => x"5b8d0008",
     8157 => x"5b9d0004",  8158 => x"282b000c",  8159 => x"b8206000",
     8160 => x"34010001",  8161 => x"59610000",  8162 => x"29810024",
     8163 => x"48200002",  8164 => x"34010001",  8165 => x"0d61000c",
     8166 => x"29810008",  8167 => x"5c200002",  8168 => x"59820008",
     8169 => x"298d0008",  8170 => x"3561000e",  8171 => x"34030004",
     8172 => x"b9a01000",  8173 => x"f8002465",  8174 => x"2d62000c",
     8175 => x"34010001",  8176 => x"5c410004",  8177 => x"29810000",
     8178 => x"4021001d",  8179 => x"64210002",  8180 => x"59610018",
     8181 => x"41a10044",  8182 => x"2d67000c",  8183 => x"34060002",
     8184 => x"31610012",  8185 => x"41a10045",  8186 => x"34050001",
     8187 => x"3404ffff",  8188 => x"31610013",  8189 => x"41a10046",
     8190 => x"31610014",  8191 => x"34010000",  8192 => x"e000000c",
     8193 => x"08220374",  8194 => x"29880000",  8195 => x"b5021000",
     8196 => x"44600004",  8197 => x"4043001d",  8198 => x"44660002",
     8199 => x"59600018",  8200 => x"58410338",  8201 => x"58450000",
     8202 => x"0c44010e",  8203 => x"34210001",  8204 => x"29630018",
     8205 => x"48e1fff4",  8206 => x"44600006",  8207 => x"78010001",
     8208 => x"38212f88",  8209 => x"f8000b60",  8210 => x"3401ffff",
     8211 => x"3161000e",  8212 => x"78010001",  8213 => x"382149dc",
     8214 => x"28230004",  8215 => x"34010000",  8216 => x"44600004",
     8217 => x"b9800800",  8218 => x"b9a01000",  8219 => x"d8600000",
     8220 => x"2b9d0004",  8221 => x"2b8b0010",  8222 => x"2b8c000c",
     8223 => x"2b8d0008",  8224 => x"379c0010",  8225 => x"c3a00000",
     8226 => x"379cfffc",  8227 => x"5b9d0004",  8228 => x"78020001",
     8229 => x"384249dc",  8230 => x"28430008",  8231 => x"34020000",
     8232 => x"44600003",  8233 => x"d8600000",  8234 => x"b8201000",
     8235 => x"b8400800",  8236 => x"2b9d0004",  8237 => x"379c0004",
     8238 => x"c3a00000",  8239 => x"379cfffc",  8240 => x"5b9d0004",
     8241 => x"b8201000",  8242 => x"78010001",  8243 => x"38212fac",
     8244 => x"f8000b3d",  8245 => x"2b9d0004",  8246 => x"379c0004",
     8247 => x"c3a00000",  8248 => x"379cffcc",  8249 => x"5b8b0010",
     8250 => x"5b8c000c",  8251 => x"5b8d0008",  8252 => x"5b9d0004",
     8253 => x"378b0014",  8254 => x"34020000",  8255 => x"34030024",
     8256 => x"b9600800",  8257 => x"f800248f",  8258 => x"78030001",
     8259 => x"b9600800",  8260 => x"34040000",  8261 => x"34020000",
     8262 => x"38635230",  8263 => x"34080020",  8264 => x"34070008",
     8265 => x"e0000004",  8266 => x"34840001",  8267 => x"34210004",
     8268 => x"44870017",  8269 => x"b4432800",  8270 => x"e0000004",
     8271 => x"30a00000",  8272 => x"34420001",  8273 => x"34a50001",
     8274 => x"40a60000",  8275 => x"44c8fffc",  8276 => x"44c0000d",
     8277 => x"b4432800",  8278 => x"58250000",  8279 => x"e0000002",
     8280 => x"34420001",  8281 => x"b4432800",  8282 => x"40a50000",
     8283 => x"7ca90000",  8284 => x"7ca60020",  8285 => x"a1263000",
     8286 => x"5cc0fffa",  8287 => x"5ca6ffeb",  8288 => x"e0000003",
     8289 => x"340c0000",  8290 => x"448c0021",  8291 => x"2b810014",
     8292 => x"340c0000",  8293 => x"40220000",  8294 => x"34010023",
     8295 => x"4441001c",  8296 => x"780b0001",  8297 => x"780c0001",
     8298 => x"396b4dc8",  8299 => x"398c4e68",  8300 => x"e0000011",
     8301 => x"29610000",  8302 => x"f80024a3",  8303 => x"b8206800",
     8304 => x"5c20000c",  8305 => x"29620004",  8306 => x"37810018",
     8307 => x"d8400000",  8308 => x"b8206000",  8309 => x"4c2d000e",
     8310 => x"29620000",  8311 => x"78010001",  8312 => x"b9801800",
     8313 => x"38212fb4",  8314 => x"f8000af7",  8315 => x"e0000008",
     8316 => x"356b0008",  8317 => x"2b820014",  8318 => x"558bffef",
     8319 => x"78010001",  8320 => x"38212fcc",  8321 => x"f8000af0",
     8322 => x"340cffea",  8323 => x"b9800800",  8324 => x"2b9d0004",
     8325 => x"2b8b0010",  8326 => x"2b8c000c",  8327 => x"2b8d0008",
     8328 => x"379c0034",  8329 => x"c3a00000",  8330 => x"379cfff8",
     8331 => x"5b8b0008",  8332 => x"5b9d0004",  8333 => x"780b0001",
     8334 => x"396b5284",  8335 => x"29650000",  8336 => x"78020001",
     8337 => x"34240001",  8338 => x"b8201800",  8339 => x"38425230",
     8340 => x"b4220800",  8341 => x"c8a31800",  8342 => x"b4821000",
     8343 => x"f80023f4",  8344 => x"29610000",  8345 => x"3421ffff",
     8346 => x"59610000",  8347 => x"2b9d0004",  8348 => x"2b8b0008",
     8349 => x"379c0008",  8350 => x"c3a00000",  8351 => x"78010001",
     8352 => x"3821528c",  8353 => x"58200000",  8354 => x"78010001",
     8355 => x"38215284",  8356 => x"58200000",  8357 => x"78010001",
     8358 => x"38215288",  8359 => x"58200000",  8360 => x"c3a00000",
     8361 => x"379cfff4",  8362 => x"5b8b000c",  8363 => x"5b8c0008",
     8364 => x"5b9d0004",  8365 => x"780b0001",  8366 => x"396b5288",
     8367 => x"29610000",  8368 => x"340c0001",  8369 => x"442c000f",
     8370 => x"34020002",  8371 => x"44220099",  8372 => x"5c2000a1",
     8373 => x"78010001",  8374 => x"38212fe8",  8375 => x"f8000aba",
     8376 => x"78010001",  8377 => x"3821528c",  8378 => x"58200000",
     8379 => x"78010001",  8380 => x"38215284",  8381 => x"58200000",
     8382 => x"596c0000",  8383 => x"e0000096",  8384 => x"f800194d",
     8385 => x"48010094",  8386 => x"3402001b",  8387 => x"44220008",
     8388 => x"78020001",  8389 => x"38425290",  8390 => x"28430000",
     8391 => x"6424005b",  8392 => x"00650010",  8393 => x"a0a42000",
     8394 => x"44800006",  8395 => x"78010001",  8396 => x"38215290",
     8397 => x"78020001",  8398 => x"58220000",  8399 => x"e0000003",
     8400 => x"b8230800",  8401 => x"58410000",  8402 => x"78010001",
     8403 => x"38215290",  8404 => x"282b0000",  8405 => x"216100ff",
     8406 => x"4420007f",  8407 => x"3401007e",  8408 => x"4561002e",
     8409 => x"49610006",  8410 => x"34010009",  8411 => x"4561006d",
     8412 => x"3401000d",  8413 => x"5d610042",  8414 => x"e0000020",
     8415 => x"78020001",  8416 => x"38423d08",  8417 => x"28410000",
     8418 => x"45610010",  8419 => x"78020001",  8420 => x"38423d0c",
     8421 => x"28410000",  8422 => x"45610004",  8423 => x"3401007f",
     8424 => x"5d610037",  8425 => x"e0000027",  8426 => x"78010001",
     8427 => x"3821528c",  8428 => x"28220000",  8429 => x"4c02005b",
     8430 => x"3442ffff",  8431 => x"58220000",  8432 => x"34010044",
     8433 => x"e000000b",  8434 => x"78010001",  8435 => x"78020001",
     8436 => x"3821528c",  8437 => x"38425284",  8438 => x"28230000",
     8439 => x"28420000",  8440 => x"4c620050",  8441 => x"34630001",
     8442 => x"58230000",  8443 => x"34010043",  8444 => x"fbffff33",
     8445 => x"e000004b",  8446 => x"78010001",  8447 => x"38211b1c",
     8448 => x"f8000a71",  8449 => x"78010001",  8450 => x"38215288",
     8451 => x"34020002",  8452 => x"58220000",  8453 => x"e0000043",
     8454 => x"78010001",  8455 => x"78020001",  8456 => x"3821528c",
     8457 => x"38425284",  8458 => x"28210000",  8459 => x"28420000",
     8460 => x"4422003c",  8461 => x"fbffff7d",  8462 => x"34010050",
     8463 => x"e3ffffed",  8464 => x"780b0001",  8465 => x"396b528c",
     8466 => x"29610000",  8467 => x"4c010035",  8468 => x"34010044",
     8469 => x"fbffff1a",  8470 => x"34010050",  8471 => x"fbffff18",
     8472 => x"29610000",  8473 => x"3421ffff",  8474 => x"fbffff70",
     8475 => x"29610000",  8476 => x"3421ffff",  8477 => x"59610000",
     8478 => x"e000002a",  8479 => x"78010001",  8480 => x"a1610800",
     8481 => x"5c200027",  8482 => x"78010001",  8483 => x"38215284",
     8484 => x"28240000",  8485 => x"3401004f",  8486 => x"48810022",
     8487 => x"78010001",  8488 => x"3821528c",  8489 => x"28230000",
     8490 => x"44640008",  8491 => x"78020001",  8492 => x"34610001",
     8493 => x"38425230",  8494 => x"b4220800",  8495 => x"b4621000",
     8496 => x"c8831800",  8497 => x"f800235a",  8498 => x"78010001",
     8499 => x"3821528c",  8500 => x"28230000",  8501 => x"78020001",
     8502 => x"38425230",  8503 => x"b4431000",  8504 => x"304b0000",
     8505 => x"34620001",  8506 => x"58220000",  8507 => x"78010001",
     8508 => x"38215284",  8509 => x"28220000",  8510 => x"34420001",
     8511 => x"58220000",  8512 => x"34010040",  8513 => x"fbfffeee",
     8514 => x"78020001",  8515 => x"38425290",  8516 => x"28420000",
     8517 => x"78010001",  8518 => x"38212ff0",  8519 => x"f8000a2a",
     8520 => x"78010001",  8521 => x"38215290",  8522 => x"58200000",
     8523 => x"e000000a",  8524 => x"78020001",  8525 => x"38425284",
     8526 => x"28420000",  8527 => x"78010001",  8528 => x"38215230",
     8529 => x"b4220800",  8530 => x"30200000",  8531 => x"fbfffee5",
     8532 => x"59600000",  8533 => x"2b9d0004",  8534 => x"2b8b000c",
     8535 => x"2b8c0008",  8536 => x"379c000c",  8537 => x"c3a00000",
     8538 => x"34030000",  8539 => x"34070009",  8540 => x"34050005",
     8541 => x"e0000014",  8542 => x"3486ffd0",  8543 => x"20c800ff",
     8544 => x"55070004",  8545 => x"3c630004",  8546 => x"b4c31800",
     8547 => x"e000000d",  8548 => x"3486ffbf",  8549 => x"20c600ff",
     8550 => x"54c50004",  8551 => x"3c630004",  8552 => x"3484ffc9",
     8553 => x"e0000006",  8554 => x"3486ff9f",  8555 => x"20c600ff",
     8556 => x"54c50007",  8557 => x"3c630004",  8558 => x"3484ffa9",
     8559 => x"b4831800",  8560 => x"34210001",  8561 => x"40240000",
     8562 => x"5c80ffec",  8563 => x"58430000",  8564 => x"c3a00000",
     8565 => x"34030000",  8566 => x"34050009",  8567 => x"e0000007",
     8568 => x"3484ffd0",  8569 => x"208600ff",  8570 => x"54c50006",
     8571 => x"0863000a",  8572 => x"34210001",  8573 => x"b4831800",
     8574 => x"40240000",  8575 => x"5c80fff9",  8576 => x"58430000",
     8577 => x"c3a00000",  8578 => x"379cffec",  8579 => x"5b8b0014",
     8580 => x"5b8c0010",  8581 => x"5b8d000c",  8582 => x"5b8e0008",
     8583 => x"5b9d0004",  8584 => x"78010001",  8585 => x"38216a58",
     8586 => x"40210000",  8587 => x"340bffff",  8588 => x"4420001c",
     8589 => x"780b0001",  8590 => x"780e0001",  8591 => x"780d0001",
     8592 => x"340c0000",  8593 => x"396b5230",  8594 => x"39ce5284",
     8595 => x"39ad300c",  8596 => x"b9600800",  8597 => x"34020050",
     8598 => x"b9801800",  8599 => x"f800149d",  8600 => x"59c10000",
     8601 => x"48200007",  8602 => x"340b0000",  8603 => x"5d80000d",
     8604 => x"78010001",  8605 => x"38212ff4",  8606 => x"f80009d3",
     8607 => x"e0000009",  8608 => x"b5610800",  8609 => x"3020ffff",
     8610 => x"b9601000",  8611 => x"b9a00800",  8612 => x"f80009cd",
     8613 => x"fbfffe93",  8614 => x"340c0001",  8615 => x"e3ffffed",
     8616 => x"b9600800",  8617 => x"2b9d0004",  8618 => x"2b8b0014",
     8619 => x"2b8c0010",  8620 => x"2b8d000c",  8621 => x"2b8e0008",
     8622 => x"379c0014",  8623 => x"c3a00000",  8624 => x"379cfff8",
     8625 => x"5b8b0008",  8626 => x"5b9d0004",  8627 => x"78010001",
     8628 => x"38216db8",  8629 => x"28210000",  8630 => x"78030001",
     8631 => x"386343d8",  8632 => x"28620000",  8633 => x"282b000c",
     8634 => x"78030001",  8635 => x"78010001",  8636 => x"38633034",
     8637 => x"3821301c",  8638 => x"f80009b3",  8639 => x"78040001",
     8640 => x"78030001",  8641 => x"388443dc",  8642 => x"386343e0",
     8643 => x"28820000",  8644 => x"28630000",  8645 => x"78010001",
     8646 => x"38213054",  8647 => x"f80009aa",  8648 => x"216b000f",
     8649 => x"356b0001",  8650 => x"78010001",  8651 => x"34020080",
     8652 => x"3d6b0004",  8653 => x"38213064",  8654 => x"34030800",
     8655 => x"f80009a2",  8656 => x"3561ff80",  8657 => x"3402000f",
     8658 => x"50410006",  8659 => x"78010001",  8660 => x"3821308c",
     8661 => x"b9601000",  8662 => x"35630010",  8663 => x"f800099a",
     8664 => x"34010000",  8665 => x"2b9d0004",  8666 => x"2b8b0008",
     8667 => x"379c0008",  8668 => x"c3a00000",  8669 => x"379cffe8",
     8670 => x"5b8b0010",  8671 => x"5b8c000c",  8672 => x"5b8d0008",
     8673 => x"5b9d0004",  8674 => x"b8205800",  8675 => x"28210000",
     8676 => x"78020001",  8677 => x"384230bc",  8678 => x"f800232b",
     8679 => x"5c200011",  8680 => x"2963000c",  8681 => x"3402ffea",
     8682 => x"44610086",  8683 => x"29610004",  8684 => x"f80004b9",
     8685 => x"b8206800",  8686 => x"29610008",  8687 => x"f80004b6",
     8688 => x"b8206000",  8689 => x"2961000c",  8690 => x"f80004b3",
     8691 => x"b8201800",  8692 => x"b9801000",  8693 => x"b9a00800",
     8694 => x"f8001d6d",  8695 => x"e0000078",  8696 => x"29610000",
     8697 => x"78020001",  8698 => x"384230c4",  8699 => x"f8002316",
     8700 => x"b8201800",  8701 => x"5c200007",  8702 => x"29610004",
     8703 => x"3402ffea",  8704 => x"44230070",  8705 => x"f80004a4",
     8706 => x"f8001e46",  8707 => x"e0000060",  8708 => x"29610000",
     8709 => x"78020001",  8710 => x"384230c8",  8711 => x"f800230a",
     8712 => x"5c200003",  8713 => x"f8001ed8",  8714 => x"e0000065",
     8715 => x"29610000",  8716 => x"78020001",  8717 => x"384230d0",
     8718 => x"f8002303",  8719 => x"5c20000d",  8720 => x"29630008",
     8721 => x"3402ffea",  8722 => x"4461005e",  8723 => x"29610004",
     8724 => x"f8000491",  8725 => x"b8206000",  8726 => x"29610008",
     8727 => x"f800048e",  8728 => x"b8201000",  8729 => x"b9800800",
     8730 => x"f8001e3f",  8731 => x"e0000054",  8732 => x"29610000",
     8733 => x"78020001",  8734 => x"384230d4",  8735 => x"f80022f2",
     8736 => x"b8201800",  8737 => x"5c20000e",  8738 => x"29610004",
     8739 => x"3402ffea",  8740 => x"4423004c",  8741 => x"f8000480",
     8742 => x"37820018",  8743 => x"37830014",  8744 => x"f8001e59",
     8745 => x"2b820018",  8746 => x"2b830014",  8747 => x"78010001",
     8748 => x"382130d8",  8749 => x"f8000944",  8750 => x"e0000041",
     8751 => x"29610000",  8752 => x"78020001",  8753 => x"384230e0",
     8754 => x"f80022df",  8755 => x"b8201800",  8756 => x"5c200007",
     8757 => x"29610004",  8758 => x"3402ffea",  8759 => x"44230039",
     8760 => x"f800046d",  8761 => x"f8001deb",  8762 => x"e0000035",
     8763 => x"29610000",  8764 => x"78020001",  8765 => x"384230e8",
     8766 => x"f80022d3",  8767 => x"b8201800",  8768 => x"5c200007",
     8769 => x"29610004",  8770 => x"3402ffea",  8771 => x"4423002d",
     8772 => x"f8000461",  8773 => x"f8001df6",  8774 => x"e0000029",
     8775 => x"29610000",  8776 => x"78020001",  8777 => x"384230f0",
     8778 => x"f80022c7",  8779 => x"5c20000d",  8780 => x"29630008",
     8781 => x"3402ffea",  8782 => x"44610022",  8783 => x"29610004",
     8784 => x"f8000455",  8785 => x"b8206000",  8786 => x"29610008",
     8787 => x"f8000452",  8788 => x"b8201000",  8789 => x"b9800800",
     8790 => x"f8001f05",  8791 => x"e0000018",  8792 => x"29610000",
     8793 => x"78020001",  8794 => x"384230f8",  8795 => x"f80022b6",
     8796 => x"b8201800",  8797 => x"5c20000b",  8798 => x"29610004",
     8799 => x"3402ffea",  8800 => x"44230010",  8801 => x"f8000444",
     8802 => x"f8001eea",  8803 => x"b8201000",  8804 => x"78010001",
     8805 => x"382138d8",  8806 => x"f800090b",  8807 => x"e0000008",
     8808 => x"29610000",  8809 => x"78020001",  8810 => x"38423100",
     8811 => x"f80022a6",  8812 => x"3402ffea",  8813 => x"5c200003",
     8814 => x"f8001fa0",  8815 => x"34020000",  8816 => x"b8400800",
     8817 => x"2b9d0004",  8818 => x"2b8b0010",  8819 => x"2b8c000c",
     8820 => x"2b8d0008",  8821 => x"379c0018",  8822 => x"c3a00000",
     8823 => x"379cffb4",  8824 => x"5b8b002c",  8825 => x"5b8c0028",
     8826 => x"5b8d0024",  8827 => x"5b8e0020",  8828 => x"5b8f001c",
     8829 => x"5b900018",  8830 => x"5b910014",  8831 => x"5b920010",
     8832 => x"5b93000c",  8833 => x"5b940008",  8834 => x"5b9d0004",
     8835 => x"b8205800",  8836 => x"28210000",  8837 => x"44200015",
     8838 => x"78020001",  8839 => x"38423110",  8840 => x"f8002289",
     8841 => x"b8206000",  8842 => x"5c200010",  8843 => x"f8000f26",
     8844 => x"5c2c0005",  8845 => x"78010001",  8846 => x"38213118",
     8847 => x"f80008e2",  8848 => x"e0000004",  8849 => x"78010001",
     8850 => x"38214ac0",  8851 => x"f8000f25",  8852 => x"78020001",
     8853 => x"38424ac0",  8854 => x"78010001",  8855 => x"30400010",
     8856 => x"38212e70",  8857 => x"e000004d",  8858 => x"29610000",
     8859 => x"78020001",  8860 => x"38423124",  8861 => x"f8002274",
     8862 => x"5c200009",  8863 => x"f80011ca",  8864 => x"3402ffff",
     8865 => x"340c0000",  8866 => x"5c2200b3",  8867 => x"78010001",
     8868 => x"3821312c",  8869 => x"f80008cc",  8870 => x"e00000af",
     8871 => x"29610010",  8872 => x"44200040",  8873 => x"29610000",
     8874 => x"78020001",  8875 => x"38423140",  8876 => x"f8002265",
     8877 => x"5c20003b",  8878 => x"29610004",  8879 => x"356c0004",
     8880 => x"f80022a6",  8881 => x"34020010",  8882 => x"54220005",
     8883 => x"29610004",  8884 => x"f80022a2",  8885 => x"3c220018",
     8886 => x"14420018",  8887 => x"34030000",  8888 => x"37840030",
     8889 => x"e0000007",  8890 => x"29810000",  8891 => x"b4832800",
     8892 => x"b4230800",  8893 => x"40210000",  8894 => x"34630001",
     8895 => x"30a10000",  8896 => x"b0600800",  8897 => x"4841fff9",
     8898 => x"b4811000",  8899 => x"34030020",  8900 => x"3404000f",
     8901 => x"e0000005",  8902 => x"34210001",  8903 => x"30430000",
     8904 => x"b0200800",  8905 => x"34420001",  8906 => x"4c81fffc",
     8907 => x"29610008",  8908 => x"f80003d9",  8909 => x"5b810044",
     8910 => x"2961000c",  8911 => x"f80003d6",  8912 => x"5b810048",
     8913 => x"29610010",  8914 => x"f80003d3",  8915 => x"5b810040",
     8916 => x"34020001",  8917 => x"37810030",  8918 => x"34030000",
     8919 => x"f80011a7",  8920 => x"3c220018",  8921 => x"3401fffe",
     8922 => x"14420018",  8923 => x"5c410004",  8924 => x"78010001",
     8925 => x"38213144",  8926 => x"e0000067",  8927 => x"3401ffff",
     8928 => x"5c410004",  8929 => x"78010001",  8930 => x"38213154",
     8931 => x"e0000062",  8932 => x"78010001",  8933 => x"38213160",
     8934 => x"f800088b",  8935 => x"e000006d",  8936 => x"29610000",
     8937 => x"44200033",  8938 => x"78020001",  8939 => x"38423170",
     8940 => x"f8002225",  8941 => x"5c20002f",  8942 => x"78100001",
     8943 => x"780f0001",  8944 => x"780e0001",  8945 => x"340c0000",
     8946 => x"340b0000",  8947 => x"34120001",  8948 => x"37910030",
     8949 => x"3414ffff",  8950 => x"3a1031ac",  8951 => x"37930040",
     8952 => x"39ef2ff0",  8953 => x"39ce31b4",  8954 => x"ba200800",
     8955 => x"34020000",  8956 => x"b9801800",  8957 => x"f8001181",
     8958 => x"5d60000b",  8959 => x"b0201000",  8960 => x"5c4b0004",
     8961 => x"78010001",  8962 => x"38213178",  8963 => x"e0000042",
     8964 => x"5c540004",  8965 => x"78010001",  8966 => x"38213190",
     8967 => x"e000003e",  8968 => x"b8409000",  8969 => x"358c0001",
     8970 => x"ba000800",  8971 => x"b9801000",  8972 => x"f8000865",
     8973 => x"ba206800",  8974 => x"41a20000",  8975 => x"b9e00800",
     8976 => x"35ad0001",  8977 => x"f8000860",  8978 => x"5db3fffc",
     8979 => x"2b820044",  8980 => x"2b830048",  8981 => x"2b840040",
     8982 => x"356b0001",  8983 => x"b9c00800",  8984 => x"b1605800",
     8985 => x"f8000858",  8986 => x"4a4bffe0",  8987 => x"e0000039",
     8988 => x"29610000",  8989 => x"4420002a",  8990 => x"78020001",
     8991 => x"384231d4",  8992 => x"f80021f1",  8993 => x"5c200026",
     8994 => x"78020001",  8995 => x"38424ac0",  8996 => x"40430000",
     8997 => x"5c610004",  8998 => x"78010001",  8999 => x"382131dc",
     9000 => x"e000001d",  9001 => x"378b0030",  9002 => x"b9600800",
     9003 => x"34030010",  9004 => x"f80022a6",  9005 => x"b9600800",
     9006 => x"f80011c0",  9007 => x"4c010014",  9008 => x"2b820044",
     9009 => x"2b830048",  9010 => x"2b840040",  9011 => x"78010001",
     9012 => x"382131f4",  9013 => x"f800083c",  9014 => x"2b820044",
     9015 => x"78010001",  9016 => x"38214e6c",  9017 => x"58220000",
     9018 => x"2b820048",  9019 => x"78010001",  9020 => x"38214e70",
     9021 => x"58220000",  9022 => x"2b820040",  9023 => x"78010001",
     9024 => x"382143ec",  9025 => x"58220000",  9026 => x"e0000012",
     9027 => x"78010001",  9028 => x"3821321c",  9029 => x"f800082c",
     9030 => x"e000000e",  9031 => x"29610000",  9032 => x"340c0000",
     9033 => x"4420000c",  9034 => x"78020001",  9035 => x"38423234",
     9036 => x"f80021c5",  9037 => x"b8201000",  9038 => x"5c200007",
     9039 => x"29610004",  9040 => x"340cffea",  9041 => x"44220004",
     9042 => x"f8000353",  9043 => x"f80009dc",  9044 => x"340c0000",
     9045 => x"b9800800",  9046 => x"2b9d0004",  9047 => x"2b8b002c",
     9048 => x"2b8c0028",  9049 => x"2b8d0024",  9050 => x"2b8e0020",
     9051 => x"2b8f001c",  9052 => x"2b900018",  9053 => x"2b910014",
     9054 => x"2b920010",  9055 => x"2b93000c",  9056 => x"2b940008",
     9057 => x"379c004c",  9058 => x"c3a00000",  9059 => x"379cfff8",
     9060 => x"5b8b0008",  9061 => x"5b9d0004",  9062 => x"b8205800",
     9063 => x"28210000",  9064 => x"5c200011",  9065 => x"78010001",
     9066 => x"38216dac",  9067 => x"28220000",  9068 => x"340b0000",
     9069 => x"64420000",  9070 => x"58220000",  9071 => x"78010001",
     9072 => x"38216d04",  9073 => x"28230000",  9074 => x"3463ffff",
     9075 => x"58230000",  9076 => x"5c4b002b",  9077 => x"78010001",
     9078 => x"3821323c",  9079 => x"f80007fa",  9080 => x"e0000027",
     9081 => x"78020001",  9082 => x"38423250",  9083 => x"f8002196",
     9084 => x"5c200007",  9085 => x"f8000965",  9086 => x"b8201000",
     9087 => x"78010001",  9088 => x"3821371c",  9089 => x"f80007f0",
     9090 => x"e000001c",  9091 => x"29610000",  9092 => x"78020001",
     9093 => x"38422524",  9094 => x"f800218b",  9095 => x"5c20000b",
     9096 => x"78010001",  9097 => x"38216dac",  9098 => x"34020001",
     9099 => x"58220000",  9100 => x"78010001",  9101 => x"38216d04",
     9102 => x"28220000",  9103 => x"3442ffff",  9104 => x"58220000",
     9105 => x"e000000d",  9106 => x"29610000",  9107 => x"78020001",
     9108 => x"38423254",  9109 => x"f800217c",  9110 => x"340bffea",
     9111 => x"5c200008",  9112 => x"78010001",  9113 => x"38216dac",
     9114 => x"58200000",  9115 => x"78010001",  9116 => x"3821323c",
     9117 => x"f80007d4",  9118 => x"340b0000",  9119 => x"b9600800",
     9120 => x"2b9d0004",  9121 => x"2b8b0008",  9122 => x"379c0008",
     9123 => x"c3a00000",  9124 => x"379cfff8",  9125 => x"5b8b0008",
     9126 => x"5b9d0004",  9127 => x"b8205800",  9128 => x"28210000",
     9129 => x"78020001",  9130 => x"384230e0",  9131 => x"f8002166",
     9132 => x"5c200003",  9133 => x"fbffe2a3",  9134 => x"e0000008",
     9135 => x"29610000",  9136 => x"78020001",  9137 => x"384230e8",
     9138 => x"f800215f",  9139 => x"3402ffea",  9140 => x"5c200003",
     9141 => x"fbffe2bd",  9142 => x"b8201000",  9143 => x"b8400800",
     9144 => x"2b9d0004",  9145 => x"2b8b0008",  9146 => x"379c0008",
     9147 => x"c3a00000",  9148 => x"379cfff8",  9149 => x"5b8b0008",
     9150 => x"5b9d0004",  9151 => x"b8205800",  9152 => x"28210000",
     9153 => x"78020001",  9154 => x"3842325c",  9155 => x"f800214e",
     9156 => x"34020001",  9157 => x"44200018",  9158 => x"29610000",
     9159 => x"78020001",  9160 => x"3842296c",  9161 => x"f8002148",
     9162 => x"34020002",  9163 => x"44200012",  9164 => x"29610000",
     9165 => x"78020001",  9166 => x"38422484",  9167 => x"f8002142",
     9168 => x"34020003",  9169 => x"4420000c",  9170 => x"fbffe27a",
     9171 => x"3c210002",  9172 => x"78020001",  9173 => x"38423fe8",
     9174 => x"b4411000",  9175 => x"28420000",  9176 => x"78010001",
     9177 => x"38212e70",  9178 => x"f8000797",  9179 => x"34010000",
     9180 => x"e0000003",  9181 => x"b8400800",  9182 => x"fbffe2b6",
     9183 => x"2b9d0004",  9184 => x"2b8b0008",  9185 => x"379c0008",
     9186 => x"c3a00000",  9187 => x"379cfff0",  9188 => x"5b8b000c",
     9189 => x"5b8c0008",  9190 => x"5b9d0004",  9191 => x"b8205800",
     9192 => x"28210000",  9193 => x"4420000b",  9194 => x"78020001",
     9195 => x"38423274",  9196 => x"f8002125",  9197 => x"b8206000",
     9198 => x"5c200006",  9199 => x"37810010",  9200 => x"f8000f2f",
     9201 => x"340bffff",  9202 => x"49810021",  9203 => x"e000001c",
     9204 => x"29610000",  9205 => x"340b0000",  9206 => x"5c20001d",
     9207 => x"37810010",  9208 => x"34020000",  9209 => x"f8001136",
     9210 => x"4d61000a",  9211 => x"2b820010",  9212 => x"78010001",
     9213 => x"3821327c",  9214 => x"f8000773",  9215 => x"2b820010",
     9216 => x"78010001",  9217 => x"382143f0",  9218 => x"58220000",
     9219 => x"e0000010",  9220 => x"78010001",  9221 => x"382132a4",
     9222 => x"f800076b",  9223 => x"37810010",  9224 => x"f8000f17",
     9225 => x"340bffff",  9226 => x"48010009",  9227 => x"2b820010",
     9228 => x"78010001",  9229 => x"382143f0",  9230 => x"58220000",
     9231 => x"37810010",  9232 => x"34020001",  9233 => x"f800111e",
     9234 => x"b8205800",  9235 => x"b9600800",  9236 => x"2b9d0004",
     9237 => x"2b8b000c",  9238 => x"2b8c0008",  9239 => x"379c0010",
     9240 => x"c3a00000",  9241 => x"379cffe8",  9242 => x"5b8b000c",
     9243 => x"5b8c0008",  9244 => x"5b9d0004",  9245 => x"b8205800",
     9246 => x"37820018",  9247 => x"37810010",  9248 => x"f8000d35",
     9249 => x"29610008",  9250 => x"44200014",  9251 => x"29610000",
     9252 => x"78020001",  9253 => x"384232d8",  9254 => x"f80020eb",
     9255 => x"5c20000f",  9256 => x"fbffe224",  9257 => x"34030003",
     9258 => x"3402fff0",  9259 => x"4423003f",  9260 => x"29610004",
     9261 => x"f8000278",  9262 => x"b8206000",  9263 => x"29610008",
     9264 => x"f8000275",  9265 => x"b8201800",  9266 => x"b9801000",
     9267 => x"1581001f",  9268 => x"34040003",  9269 => x"e0000020",
     9270 => x"29610000",  9271 => x"4420000f",  9272 => x"78020001",
     9273 => x"384232dc",  9274 => x"f80020d7",  9275 => x"5c20000b",
     9276 => x"fbffe210",  9277 => x"34020003",  9278 => x"44220023",
     9279 => x"29610004",  9280 => x"f8000265",  9281 => x"b8201000",
     9282 => x"34030000",  9283 => x"1421001f",  9284 => x"34040001",
     9285 => x"e0000010",  9286 => x"29610000",  9287 => x"44200010",
     9288 => x"78020001",  9289 => x"384232e4",  9290 => x"f80020c7",
     9291 => x"5c20000c",  9292 => x"fbffe200",  9293 => x"34020003",
     9294 => x"44220013",  9295 => x"29610004",  9296 => x"f8000255",
     9297 => x"b8201800",  9298 => x"34020000",  9299 => x"34010000",
     9300 => x"34040002",  9301 => x"f8000ce0",  9302 => x"e0000013",
     9303 => x"29610000",  9304 => x"44200009",  9305 => x"78020001",
     9306 => x"384232ec",  9307 => x"f80020b6",  9308 => x"5c200005",
     9309 => x"78010001",  9310 => x"382130d8",  9311 => x"2b820014",
     9312 => x"e0000007",  9313 => x"2b820014",  9314 => x"2b810010",
     9315 => x"f8000169",  9316 => x"b8201000",  9317 => x"78010001",
     9318 => x"382132f0",  9319 => x"2b830018",  9320 => x"f8000709",
     9321 => x"34020000",  9322 => x"b8400800",  9323 => x"2b9d0004",
     9324 => x"2b8b000c",  9325 => x"2b8c0008",  9326 => x"379c0018",
     9327 => x"c3a00000",  9328 => x"78010001",  9329 => x"38214e68",
     9330 => x"34020001",  9331 => x"58220000",  9332 => x"34010000",
     9333 => x"c3a00000",  9334 => x"379cfffc",  9335 => x"5b9d0004",
     9336 => x"f8000d86",  9337 => x"34010000",  9338 => x"2b9d0004",
     9339 => x"379c0004",  9340 => x"c3a00000",  9341 => x"379cffec",
     9342 => x"5b8b0010",  9343 => x"5b8c000c",  9344 => x"5b8d0008",
     9345 => x"5b9d0004",  9346 => x"340b0000",  9347 => x"b8406800",
     9348 => x"340c0006",  9349 => x"37820014",  9350 => x"fbfffcd4",
     9351 => x"2b830014",  9352 => x"b5ab1000",  9353 => x"356b0001",
     9354 => x"30430000",  9355 => x"40220000",  9356 => x"6442003a",
     9357 => x"b4220800",  9358 => x"5d6cfff7",  9359 => x"2b9d0004",
     9360 => x"2b8b0010",  9361 => x"2b8c000c",  9362 => x"2b8d0008",
     9363 => x"379c0014",  9364 => x"c3a00000",  9365 => x"379cfff0",
     9366 => x"5b8b0008",  9367 => x"5b9d0004",  9368 => x"b8205800",
     9369 => x"28210000",  9370 => x"44200005",  9371 => x"78020001",
     9372 => x"38423318",  9373 => x"f8002074",  9374 => x"5c200004",
     9375 => x"3781000c",  9376 => x"f80007d9",  9377 => x"e000002b",
     9378 => x"29610000",  9379 => x"78020001",  9380 => x"3842331c",
     9381 => x"f800206c",  9382 => x"5c200008",  9383 => x"378b000c",
     9384 => x"b9600800",  9385 => x"f80007d0",  9386 => x"b9601000",
     9387 => x"34010000",  9388 => x"f80011e3",  9389 => x"e000001f",
     9390 => x"29610000",  9391 => x"78020001",  9392 => x"384232d8",
     9393 => x"f8002060",  9394 => x"5c20000b",  9395 => x"29630004",
     9396 => x"44610009",  9397 => x"378b000c",  9398 => x"b8600800",
     9399 => x"b9601000",  9400 => x"fbffffc5",  9401 => x"b9600800",
     9402 => x"f80007ab",  9403 => x"f80008a6",  9404 => x"e0000010",
     9405 => x"29610000",  9406 => x"78020001",  9407 => x"38423324",
     9408 => x"f8002051",  9409 => x"b8201800",  9410 => x"3402ffea",
     9411 => x"5c200013",  9412 => x"29610004",  9413 => x"44230011",
     9414 => x"378b000c",  9415 => x"b9601000",  9416 => x"fbffffb5",
     9417 => x"34010000",  9418 => x"b9601000",  9419 => x"f80011bb",
     9420 => x"4382000c",  9421 => x"4383000d",  9422 => x"4384000e",
     9423 => x"4385000f",  9424 => x"43860010",  9425 => x"43870011",
     9426 => x"78010001",  9427 => x"3821332c",  9428 => x"f800069d",
     9429 => x"34020000",  9430 => x"b8400800",  9431 => x"2b9d0004",
     9432 => x"2b8b0008",  9433 => x"379c0010",  9434 => x"c3a00000",
     9435 => x"379cfff4",  9436 => x"5b8b000c",  9437 => x"5b8c0008",
     9438 => x"5b9d0004",  9439 => x"34020050",  9440 => x"b8205800",
     9441 => x"34010000",  9442 => x"f80009ef",  9443 => x"5c200006",
     9444 => x"78010001",  9445 => x"3821335c",  9446 => x"f800068b",
     9447 => x"340bffff",  9448 => x"e0000031",  9449 => x"29610000",
     9450 => x"4420000c",  9451 => x"78020001",  9452 => x"38423124",
     9453 => x"f8002024",  9454 => x"5c200008",  9455 => x"f8001075",
     9456 => x"340b0000",  9457 => x"4c2b0028",  9458 => x"78010001",
     9459 => x"38213370",  9460 => x"f800067d",  9461 => x"e0000024",
     9462 => x"29610004",  9463 => x"44200012",  9464 => x"29610000",
     9465 => x"78020001",  9466 => x"38423140",  9467 => x"f8002016",
     9468 => x"b8206000",  9469 => x"5c20000c",  9470 => x"b9600800",
     9471 => x"f800107a",  9472 => x"4c2c0004",  9473 => x"78010001",
     9474 => x"38213390",  9475 => x"e0000003",  9476 => x"78010001",
     9477 => x"382133ac",  9478 => x"f800066b",  9479 => x"340b0000",
     9480 => x"e0000011",  9481 => x"29610000",  9482 => x"44200007",
     9483 => x"78020001",  9484 => x"38423170",  9485 => x"f8002004",
     9486 => x"5c200003",  9487 => x"f80010e4",  9488 => x"e3fffff7",
     9489 => x"29610000",  9490 => x"340b0000",  9491 => x"44200006",
     9492 => x"78020001",  9493 => x"384233b4",  9494 => x"f8001ffb",
     9495 => x"5c200002",  9496 => x"fbfffc6a",  9497 => x"b9600800",
     9498 => x"2b9d0004",  9499 => x"2b8b000c",  9500 => x"2b8c0008",
     9501 => x"379c000c",  9502 => x"c3a00000",  9503 => x"379cfff8",
     9504 => x"5b8b0008",  9505 => x"5b9d0004",  9506 => x"b8205800",
     9507 => x"28210000",  9508 => x"4420000c",  9509 => x"78020001",
     9510 => x"384233c4",  9511 => x"f8001fea",  9512 => x"5c200008",
     9513 => x"34010001",  9514 => x"fbffec22",  9515 => x"78010001",
     9516 => x"382143e8",  9517 => x"34020001",  9518 => x"58220000",
     9519 => x"e000000b",  9520 => x"29610000",  9521 => x"44200009",
     9522 => x"78020001",  9523 => x"384233cc",  9524 => x"f8001fdd",
     9525 => x"5c200005",  9526 => x"fbffec16",  9527 => x"78010001",
     9528 => x"382143e8",  9529 => x"58200000",  9530 => x"78010001",
     9531 => x"382143e8",  9532 => x"28210000",  9533 => x"78020001",
     9534 => x"384233c0",  9535 => x"44200003",  9536 => x"78020001",
     9537 => x"384233bc",  9538 => x"78010001",  9539 => x"382133d4",
     9540 => x"f800062d",  9541 => x"34010000",  9542 => x"2b9d0004",
     9543 => x"2b8b0008",  9544 => x"379c0008",  9545 => x"c3a00000",
     9546 => x"379cfff0",  9547 => x"5b8b0010",  9548 => x"5b8c000c",
     9549 => x"5b8d0008",  9550 => x"5b9d0004",  9551 => x"78010001",
     9552 => x"382133f0",  9553 => x"780b0001",  9554 => x"780d0001",
     9555 => x"780c0001",  9556 => x"f800061d",  9557 => x"396b4dc8",
     9558 => x"39ad4e68",  9559 => x"398c3408",  9560 => x"e0000005",
     9561 => x"29620000",  9562 => x"b9800800",  9563 => x"356b0008",
     9564 => x"f8000615",  9565 => x"55abfffc",  9566 => x"34010000",
     9567 => x"2b9d0004",  9568 => x"2b8b0010",  9569 => x"2b8c000c",
     9570 => x"2b8d0008",  9571 => x"379c0010",  9572 => x"c3a00000",
     9573 => x"379cfff8",  9574 => x"5b9d0004",  9575 => x"b8201000",
     9576 => x"28210000",  9577 => x"4420000d",  9578 => x"28420004",
     9579 => x"5c40000b",  9580 => x"37820008",  9581 => x"fbfffc08",
     9582 => x"2b820008",  9583 => x"78010001",  9584 => x"382143e4",
     9585 => x"084203e8",  9586 => x"58220000",  9587 => x"78010001",
     9588 => x"38211b1c",  9589 => x"e0000003",  9590 => x"78010001",
     9591 => x"38213418",  9592 => x"f80005f9",  9593 => x"34010000",
     9594 => x"2b9d0004",  9595 => x"379c0008",  9596 => x"c3a00000",
     9597 => x"379cffe8",  9598 => x"5b8b0010",  9599 => x"5b8c000c",
     9600 => x"5b9b0008",  9601 => x"5b9d0004",  9602 => x"b820d800",
     9603 => x"28210000",  9604 => x"44200005",  9605 => x"78020001",
     9606 => x"38423318",  9607 => x"f8001f8a",  9608 => x"5c200004",
     9609 => x"37810018",  9610 => x"f80004ca",  9611 => x"e0000018",
     9612 => x"2b610000",  9613 => x"78020001",  9614 => x"384232d8",
     9615 => x"f8001f82",  9616 => x"b8201800",  9617 => x"3402ffea",
     9618 => x"5c200021",  9619 => x"2b610004",  9620 => x"4423001f",
     9621 => x"379b0018",  9622 => x"378c001c",  9623 => x"378b0014",
     9624 => x"b9601000",  9625 => x"fbfffbdc",  9626 => x"2b820014",
     9627 => x"33620000",  9628 => x"40220000",  9629 => x"377b0001",
     9630 => x"6442002e",  9631 => x"b4220800",  9632 => x"5f6cfff8",
     9633 => x"37810018",  9634 => x"f80004bb",  9635 => x"78010001",
     9636 => x"38215d6c",  9637 => x"28210000",  9638 => x"44200005",
     9639 => x"78010001",  9640 => x"3821343c",  9641 => x"f80005c8",
     9642 => x"e0000008",  9643 => x"43820018",  9644 => x"43830019",
     9645 => x"4384001a",  9646 => x"4385001b",  9647 => x"78010001",
     9648 => x"38213458",  9649 => x"f80005c0",  9650 => x"34020000",
     9651 => x"b8400800",  9652 => x"2b9d0004",  9653 => x"2b8b0010",
     9654 => x"2b8c000c",  9655 => x"2b9b0008",  9656 => x"379c0018",
     9657 => x"c3a00000",  9658 => x"379cfffc",  9659 => x"5b9d0004",
     9660 => x"28210000",  9661 => x"44200005",  9662 => x"fbffdf97",
     9663 => x"78020001",  9664 => x"38424e9c",  9665 => x"58410000",
     9666 => x"78020001",  9667 => x"38424e9c",  9668 => x"28420000",
     9669 => x"78010001",  9670 => x"38213478",  9671 => x"f80005aa",
     9672 => x"34010000",  9673 => x"2b9d0004",  9674 => x"379c0004",
     9675 => x"c3a00000",  9676 => x"379cffd8",  9677 => x"5b8b0028",
     9678 => x"5b8c0024",  9679 => x"5b8d0020",  9680 => x"5b8e001c",
     9681 => x"5b8f0018",  9682 => x"5b900014",  9683 => x"5b910010",
     9684 => x"5b92000c",  9685 => x"5b9d0008",  9686 => x"78030001",
     9687 => x"38633d10",  9688 => x"b8406000",  9689 => x"b8400800",
     9690 => x"28620000",  9691 => x"f8001e26",  9692 => x"78030001",
     9693 => x"38633d10",  9694 => x"28620000",  9695 => x"b8205800",
     9696 => x"b9800800",  9697 => x"f8001e10",  9698 => x"b8206000",
     9699 => x"3402003c",  9700 => x"b9600800",  9701 => x"f8001e1c",
     9702 => x"34020e10",  9703 => x"b8208800",  9704 => x"b9600800",
     9705 => x"f8001e18",  9706 => x"3402003c",  9707 => x"f8001e06",
     9708 => x"34020e10",  9709 => x"b8207800",  9710 => x"b9600800",
     9711 => x"f8001e02",  9712 => x"b8208000",  9713 => x"34020007",
     9714 => x"35810004",  9715 => x"f8001e0e",  9716 => x"b8209000",
     9717 => x"340b07b2",  9718 => x"e000000f",  9719 => x"3402016d",
     9720 => x"5da0000b",  9721 => x"34020064",  9722 => x"b9600800",
     9723 => x"f8001dd6",  9724 => x"3402016e",  9725 => x"5c2d0006",
     9726 => x"34020190",  9727 => x"b9600800",  9728 => x"f8001dd1",
     9729 => x"64220000",  9730 => x"3442016d",  9731 => x"c9826000",
     9732 => x"356b0001",  9733 => x"216d0003",  9734 => x"3402016d",
     9735 => x"5da0000b",  9736 => x"34020064",  9737 => x"b9600800",
     9738 => x"f8001dc7",  9739 => x"3402016e",  9740 => x"5c2d0006",
     9741 => x"34020190",  9742 => x"b9600800",  9743 => x"f8001dc2",
     9744 => x"64220000",  9745 => x"3442016d",  9746 => x"5182ffe5",
     9747 => x"34020064",  9748 => x"b9600800",  9749 => x"f8001dbc",
     9750 => x"34020190",  9751 => x"b8207000",  9752 => x"b9600800",
     9753 => x"f8001db8",  9754 => x"78030001",  9755 => x"34020000",
     9756 => x"64250000",  9757 => x"38633ff8",  9758 => x"e000000d",
     9759 => x"34040000",  9760 => x"5da00004",  9761 => x"34040001",
     9762 => x"5dcd0002",  9763 => x"b8a02000",  9764 => x"0884000c",
     9765 => x"b4822000",  9766 => x"3c840002",  9767 => x"34420001",
     9768 => x"b4642000",  9769 => x"28810000",  9770 => x"c9816000",
     9771 => x"34040000",  9772 => x"5da00004",  9773 => x"34040001",
     9774 => x"5dcd0002",  9775 => x"b8a02000",  9776 => x"0884000c",
     9777 => x"b4822000",  9778 => x"3c840002",  9779 => x"b4642000",
     9780 => x"28810000",  9781 => x"5181ffea",  9782 => x"3e450002",
     9783 => x"78030001",  9784 => x"38634058",  9785 => x"b4652800",
     9786 => x"3c420002",  9787 => x"78030001",  9788 => x"38634074",
     9789 => x"b4622000",  9790 => x"28840000",  9791 => x"28a30000",
     9792 => x"780d0001",  9793 => x"39ad5294",  9794 => x"78020001",
     9795 => x"b9a00800",  9796 => x"38423498",  9797 => x"35850001",
     9798 => x"b9603000",  9799 => x"ba003800",  9800 => x"b9e04000",
     9801 => x"5b910004",  9802 => x"f8000519",  9803 => x"b9a00800",
     9804 => x"2b9d0008",  9805 => x"2b8b0028",  9806 => x"2b8c0024",
     9807 => x"2b8d0020",  9808 => x"2b8e001c",  9809 => x"2b8f0018",
     9810 => x"2b900014",  9811 => x"2b910010",  9812 => x"2b92000c",
     9813 => x"379c0028",  9814 => x"c3a00000",  9815 => x"379cffdc",
     9816 => x"5b8b0008",  9817 => x"5b9d0004",  9818 => x"5b840014",
     9819 => x"20240080",  9820 => x"64840000",  9821 => x"5b830010",
     9822 => x"78030001",  9823 => x"b8204800",  9824 => x"b8600800",
     9825 => x"34030002",  9826 => x"5b82000c",  9827 => x"b8405800",
     9828 => x"382134b8",  9829 => x"c8641000",  9830 => x"2123007f",
     9831 => x"5b850018",  9832 => x"5b86001c",  9833 => x"5b870020",
     9834 => x"5b880024",  9835 => x"f8000506",  9836 => x"37820010",
     9837 => x"b9600800",  9838 => x"f80004e1",  9839 => x"78010001",
     9840 => x"382134c4",  9841 => x"f8000500",  9842 => x"2b9d0004",
     9843 => x"2b8b0008",  9844 => x"379c0024",  9845 => x"c3a00000",
     9846 => x"379cffe0",  9847 => x"5b8b000c",  9848 => x"5b8c0008",
     9849 => x"5b9d0004",  9850 => x"b8404800",  9851 => x"78020001",
     9852 => x"b8205000",  9853 => x"b8400800",  9854 => x"b8605800",
     9855 => x"b9401000",  9856 => x"b9201800",  9857 => x"382134c8",
     9858 => x"b8806000",  9859 => x"5b840010",  9860 => x"5b850014",
     9861 => x"5b860018",  9862 => x"5b87001c",  9863 => x"5b880020",
     9864 => x"f80004e9",  9865 => x"21620080",  9866 => x"78030001",
     9867 => x"64420000",  9868 => x"b8600800",  9869 => x"34030002",
     9870 => x"c8621000",  9871 => x"382134b8",  9872 => x"2163007f",
     9873 => x"f80004e0",  9874 => x"37820014",  9875 => x"b9800800",
     9876 => x"f80004bb",  9877 => x"78010001",  9878 => x"382134c4",
     9879 => x"f80004da",  9880 => x"2b9d0004",  9881 => x"2b8b000c",
     9882 => x"2b8c0008",  9883 => x"379c0020",  9884 => x"c3a00000",
     9885 => x"379cfffc",  9886 => x"5b9d0004",  9887 => x"78010001",
     9888 => x"382134d4",  9889 => x"f80004d0",  9890 => x"2b9d0004",
     9891 => x"379c0004",  9892 => x"c3a00000",  9893 => x"40240000",
     9894 => x"3402002d",  9895 => x"34030001",  9896 => x"5c820003",
     9897 => x"34210001",  9898 => x"3403ffff",  9899 => x"34020000",
     9900 => x"34050009",  9901 => x"e0000004",  9902 => x"0842000a",
     9903 => x"34210001",  9904 => x"b4821000",  9905 => x"40240000",
     9906 => x"3484ffd0",  9907 => x"208600ff",  9908 => x"50a6fffa",
     9909 => x"88430800",  9910 => x"c3a00000",  9911 => x"379cfff4",
     9912 => x"5b8b000c",  9913 => x"5b8c0008",  9914 => x"5b9d0004",
     9915 => x"b8206000",  9916 => x"f8000ae7",  9917 => x"342b0001",
     9918 => x"f8000ae5",  9919 => x"5c2bffff",  9920 => x"b9800800",
     9921 => x"e0000002",  9922 => x"3421ffff",  9923 => x"4820ffff",
     9924 => x"f8000adf",  9925 => x"c82b0800",  9926 => x"2b9d0004",
     9927 => x"2b8b000c",  9928 => x"2b8c0008",  9929 => x"379c000c",
     9930 => x"c3a00000",  9931 => x"379cfff0",  9932 => x"5b8b0010",
     9933 => x"5b8c000c",  9934 => x"5b8d0008",  9935 => x"5b9d0004",
     9936 => x"340b0400",  9937 => x"340c0400",  9938 => x"e0000003",
     9939 => x"b58b6000",  9940 => x"3d6b0001",  9941 => x"b9800800",
     9942 => x"fbffffe1",  9943 => x"4420fffc",  9944 => x"158c0001",
     9945 => x"156b0002",  9946 => x"e0000009",  9947 => x"b56c6800",
     9948 => x"b9a00800",  9949 => x"fbffffda",  9950 => x"5c200002",
     9951 => x"b9a06000",  9952 => x"0161001f",  9953 => x"b42b5800",
     9954 => x"156b0001",  9955 => x"5d60fff8",  9956 => x"78010001",
     9957 => x"382152d4",  9958 => x"582c0000",  9959 => x"78010001",
     9960 => x"b9801000",  9961 => x"3821352c",  9962 => x"f8000487",
     9963 => x"2b9d0004",  9964 => x"2b8b0010",  9965 => x"2b8c000c",
     9966 => x"2b8d0008",  9967 => x"379c0010",  9968 => x"c3a00000",
     9969 => x"379cfffc",  9970 => x"5b9d0004",  9971 => x"78020001",
     9972 => x"384252d4",  9973 => x"28430000",  9974 => x"34042710",
     9975 => x"0865000a",  9976 => x"e0000004",  9977 => x"3442ffff",
     9978 => x"4840ffff",  9979 => x"3421d8f0",  9980 => x"50810003",
     9981 => x"b8a01000",  9982 => x"e3fffffc",  9983 => x"88230800",
     9984 => x"340203e8",  9985 => x"f8001cf0",  9986 => x"e0000002",
     9987 => x"3421ffff",  9988 => x"4820ffff",  9989 => x"34010000",
     9990 => x"2b9d0004",  9991 => x"379c0004",  9992 => x"c3a00000",
     9993 => x"379cfffc",  9994 => x"5b9d0004",  9995 => x"b8400800",
     9996 => x"f800056d",  9997 => x"34010000",  9998 => x"2b9d0004",
     9999 => x"379c0004", 10000 => x"c3a00000", 10001 => x"78020001",
    10002 => x"384252d8", 10003 => x"58410018", 10004 => x"58410240",
    10005 => x"58410468", 10006 => x"58410690", 10007 => x"c3a00000",
    10008 => x"379cff24", 10009 => x"5b8b0014", 10010 => x"5b8c0010",
    10011 => x"5b8d000c", 10012 => x"5b8e0008", 10013 => x"5b9d0004",
    10014 => x"78010001", 10015 => x"b8607000", 10016 => x"382152d8",
    10017 => x"340c0000", 10018 => x"34020004", 10019 => x"28230000",
    10020 => x"5c600009", 10021 => x"78040001", 10022 => x"b8801000",
    10023 => x"37810018", 10024 => x"38423544", 10025 => x"fbffdd12",
    10026 => x"340b0000", 10027 => x"4961001d", 10028 => x"e0000006",
    10029 => x"358c0001", 10030 => x"34210228", 10031 => x"5d82fff4",
    10032 => x"340b0000", 10033 => x"e0000017", 10034 => x"098d0228",
    10035 => x"780c0001", 10036 => x"398c52d8", 10037 => x"b5ac5800",
    10038 => x"b9c01000", 10039 => x"3403000e", 10040 => x"35610004",
    10041 => x"f8001d19", 10042 => x"35610012", 10043 => x"f800053e",
    10044 => x"2b8100d0", 10045 => x"34020200", 10046 => x"0d600220",
    10047 => x"59610018", 10048 => x"2b8100b8", 10049 => x"5961001c",
    10050 => x"35610220", 10051 => x"0c200002", 10052 => x"0c220004",
    10053 => x"0c200006", 10054 => x"34010001", 10055 => x"59610000",
    10056 => x"b9600800", 10057 => x"2b9d0004", 10058 => x"2b8b0014",
    10059 => x"2b8c0010", 10060 => x"2b8d000c", 10061 => x"2b8e0008",
    10062 => x"379c00dc", 10063 => x"c3a00000", 10064 => x"44200002",
    10065 => x"58200000", 10066 => x"34010000", 10067 => x"c3a00000",
    10068 => x"379cffe8", 10069 => x"5b8b0018", 10070 => x"5b8c0014",
    10071 => x"5b8d0010", 10072 => x"5b8e000c", 10073 => x"5b8f0008",
    10074 => x"5b9d0004", 10075 => x"b8205800", 10076 => x"59620010",
    10077 => x"b8407000", 10078 => x"b8807800", 10079 => x"b8a06000",
    10080 => x"282d0008", 10081 => x"44600005", 10082 => x"b8a00800",
    10083 => x"3402fc18", 10084 => x"f8001c40", 10085 => x"b42d6800",
    10086 => x"c9cf2000", 10087 => x"b8801800", 10088 => x"4c800002",
    10089 => x"b48c1800", 10090 => x"0181001f", 10091 => x"b42c0800",
    10092 => x"14210001", 10093 => x"b4242000", 10094 => x"4c800002",
    10095 => x"b48c2000", 10096 => x"49840002", 10097 => x"c88c2000",
    10098 => x"09820003", 10099 => x"1445001f", 10100 => x"00a5001e",
    10101 => x"b4a21000", 10102 => x"14420002", 10103 => x"48620006",
    10104 => x"1582001f", 10105 => x"0042001e", 10106 => x"b44c1000",
    10107 => x"14420002", 10108 => x"4c62000d", 10109 => x"b4812000",
    10110 => x"596d0008", 10111 => x"5964000c", 10112 => x"4984000a",
    10113 => x"c88c2000", 10114 => x"5964000c", 10115 => x"b9800800",
    10116 => x"340203e8", 10117 => x"f8001c1f", 10118 => x"b5a10800",
    10119 => x"59610008", 10120 => x"e0000002", 10121 => x"5963000c",
    10122 => x"78030001", 10123 => x"38633cdc", 10124 => x"29610008",
    10125 => x"28620000", 10126 => x"4c41000d", 10127 => x"78030001",
    10128 => x"38633cf0", 10129 => x"28620000", 10130 => x"29630000",
    10131 => x"b4220800", 10132 => x"29620004", 10133 => x"59610008",
    10134 => x"34410001", 10135 => x"f4411000", 10136 => x"59610004",
    10137 => x"b4431000", 10138 => x"59620000", 10139 => x"2b9d0004",
    10140 => x"2b8b0018", 10141 => x"2b8c0014", 10142 => x"2b8d0010",
    10143 => x"2b8e000c", 10144 => x"2b8f0008", 10145 => x"379c0018",
    10146 => x"c3a00000", 10147 => x"379cffb8", 10148 => x"5b8b0020",
    10149 => x"5b8c001c", 10150 => x"5b8d0018", 10151 => x"5b8e0014",
    10152 => x"5b8f0010", 10153 => x"5b90000c", 10154 => x"5b910008",
    10155 => x"5b9d0004", 10156 => x"b8407800", 10157 => x"2c220226",
    10158 => x"b8205800", 10159 => x"b8806800", 10160 => x"b8a06000",
    10161 => x"34010000", 10162 => x"4440007f", 10163 => x"2d610222",
    10164 => x"3442ffff", 10165 => x"0d620226", 10166 => x"b5612000",
    10167 => x"40840020", 10168 => x"34210001", 10169 => x"2021ffff",
    10170 => x"3384004a", 10171 => x"0d610222", 10172 => x"34040200",
    10173 => x"2d620224", 10174 => x"5c240002", 10175 => x"0d600222",
    10176 => x"2d610222", 10177 => x"b5612000", 10178 => x"40840020",
    10179 => x"34210001", 10180 => x"2021ffff", 10181 => x"3384004b",
    10182 => x"0d610222", 10183 => x"34040200", 10184 => x"5c240002",
    10185 => x"0d600222", 10186 => x"34420002", 10187 => x"2042ffff",
    10188 => x"0d620224", 10189 => x"3787004a", 10190 => x"3785003c",
    10191 => x"34060200", 10192 => x"e000000b", 10193 => x"2d610222",
    10194 => x"b5612000", 10195 => x"40840020", 10196 => x"34210001",
    10197 => x"2021ffff", 10198 => x"30a40000", 10199 => x"0d610222",
    10200 => x"34a50001", 10201 => x"5c260002", 10202 => x"0d600222",
    10203 => x"5ca7fff6", 10204 => x"3442000e", 10205 => x"2042ffff",
    10206 => x"0d620224", 10207 => x"3787003c", 10208 => x"37850024",
    10209 => x"34060200", 10210 => x"e000000b", 10211 => x"2d610222",
    10212 => x"b5612000", 10213 => x"40840020", 10214 => x"34210001",
    10215 => x"2021ffff", 10216 => x"30a40000", 10217 => x"0d610222",
    10218 => x"34a50001", 10219 => x"5c260002", 10220 => x"0d600222",
    10221 => x"5ca7fff6", 10222 => x"34420018", 10223 => x"2f8e004a",
    10224 => x"2042ffff", 10225 => x"0d620224", 10226 => x"b9a00800",
    10227 => x"51cd0002", 10228 => x"b9c00800", 10229 => x"b4613000",
    10230 => x"34050200", 10231 => x"e000000c", 10232 => x"2d640222",
    10233 => x"b5642000", 10234 => x"40840020", 10235 => x"30640000",
    10236 => x"2d640222", 10237 => x"34630001", 10238 => x"34840001",
    10239 => x"2084ffff", 10240 => x"0d640222", 10241 => x"5c850002",
    10242 => x"0d600222", 10243 => x"5c66fff5", 10244 => x"b4410800",
    10245 => x"0d610224", 10246 => x"2f810048", 10247 => x"37820042",
    10248 => x"34030006", 10249 => x"0de1000c", 10250 => x"b9e00800",
    10251 => x"f8001c47", 10252 => x"35e10006", 10253 => x"3782003c",
    10254 => x"34030006", 10255 => x"f8001c43", 10256 => x"4580001d",
    10257 => x"2b900034", 10258 => x"2b8f0028", 10259 => x"34010000",
    10260 => x"59900014", 10261 => x"598f0018", 10262 => x"f80018ed",
    10263 => x"b8208800", 10264 => x"35820010", 10265 => x"34030000",
    10266 => x"34010000", 10267 => x"f8001892", 10268 => x"2b81002c",
    10269 => x"43820024", 10270 => x"29640018", 10271 => x"59810000",
    10272 => x"2b810030", 10273 => x"59900008", 10274 => x"5980000c",
    10275 => x"59810004", 10276 => x"222100ff", 10277 => x"64210000",
    10278 => x"b9e01800", 10279 => x"a0220800", 10280 => x"29820010",
    10281 => x"5981001c", 10282 => x"34051f40", 10283 => x"b9800800",
    10284 => x"fbffff28", 10285 => x"35cefff2", 10286 => x"b9a00800",
    10287 => x"51cd0002", 10288 => x"b9c00800", 10289 => x"2b9d0004",
    10290 => x"2b8b0020", 10291 => x"2b8c001c", 10292 => x"2b8d0018",
    10293 => x"2b8e0014", 10294 => x"2b8f0010", 10295 => x"2b90000c",
    10296 => x"2b910008", 10297 => x"379c0048", 10298 => x"c3a00000",
    10299 => x"379cffbc", 10300 => x"5b8b001c", 10301 => x"5b8c0018",
    10302 => x"5b8d0014", 10303 => x"5b8e0010", 10304 => x"5b8f000c",
    10305 => x"5b900008", 10306 => x"5b9d0004", 10307 => x"378c0038",
    10308 => x"b8208000", 10309 => x"b8607800", 10310 => x"b9800800",
    10311 => x"34030006", 10312 => x"b8807000", 10313 => x"b8406800",
    10314 => x"b8a05800", 10315 => x"f8001c07", 10316 => x"36020012",
    10317 => x"34030006", 10318 => x"3781003e", 10319 => x"f8001c03",
    10320 => x"2da1000c", 10321 => x"b9e01000", 10322 => x"35c3000e",
    10323 => x"0f810044", 10324 => x"37840020", 10325 => x"b9800800",
    10326 => x"f80007d8", 10327 => x"4560000a", 10328 => x"2b820028",
    10329 => x"5960000c", 10330 => x"59620000", 10331 => x"2b82002c",
    10332 => x"59620004", 10333 => x"2b820030", 10334 => x"59620008",
    10335 => x"43820020", 10336 => x"5962001c", 10337 => x"2b9d0004",
    10338 => x"2b8b001c", 10339 => x"2b8c0018", 10340 => x"2b8d0014",
    10341 => x"2b8e0010", 10342 => x"2b8f000c", 10343 => x"2b900008",
    10344 => x"379c0044", 10345 => x"c3a00000", 10346 => x"379cffc4",
    10347 => x"5b8b0020", 10348 => x"5b8c001c", 10349 => x"5b8d0018",
    10350 => x"5b8e0014", 10351 => x"5b8f0010", 10352 => x"5b90000c",
    10353 => x"5b9b0008", 10354 => x"5b9d0004", 10355 => x"780b0001",
    10356 => x"396b5d58", 10357 => x"78020001", 10358 => x"b9600800",
    10359 => x"38425b78", 10360 => x"340301e0", 10361 => x"37840024",
    10362 => x"f8000708", 10363 => x"b8207000", 10364 => x"4c01006d",
    10365 => x"780c0001", 10366 => x"398c52d8", 10367 => x"340d0000",
    10368 => x"b9808000", 10369 => x"b9607800", 10370 => x"341b0004",
    10371 => x"09ab0228", 10372 => x"29810000", 10373 => x"b5705800",
    10374 => x"44200009", 10375 => x"b9e00800", 10376 => x"35620004",
    10377 => x"34030006", 10378 => x"f8001ba7", 10379 => x"5c200004",
    10380 => x"2de2000c", 10381 => x"2d810010", 10382 => x"44410005",
    10383 => x"35ad0001", 10384 => x"358c0228", 10385 => x"5dbbfff2",
    10386 => x"e0000057", 10387 => x"2d630224", 10388 => x"35c10028",
    10389 => x"48230054", 10390 => x"2d620220", 10391 => x"21c1ffff",
    10392 => x"00250008", 10393 => x"b5622000", 10394 => x"34420001",
    10395 => x"0f81003e", 10396 => x"2042ffff", 10397 => x"30850020",
    10398 => x"0d620220", 10399 => x"34040200", 10400 => x"5c440002",
    10401 => x"0d600220", 10402 => x"2d620220", 10403 => x"4385003f",
    10404 => x"b5622000", 10405 => x"34420001", 10406 => x"2042ffff",
    10407 => x"30850020", 10408 => x"0d620220", 10409 => x"34040200",
    10410 => x"5c440002", 10411 => x"0d600220", 10412 => x"3463fffe",
    10413 => x"78020001", 10414 => x"2063ffff", 10415 => x"38425d58",
    10416 => x"0d630224", 10417 => x"3446000e", 10418 => x"34050200",
    10419 => x"e000000b", 10420 => x"2d640220", 10421 => x"40480000",
    10422 => x"34420001", 10423 => x"b5643800", 10424 => x"34840001",
    10425 => x"2084ffff", 10426 => x"30e80020", 10427 => x"0d640220",
    10428 => x"5c850002", 10429 => x"0d600220", 10430 => x"5c46fff6",
    10431 => x"3463fff2", 10432 => x"2063ffff", 10433 => x"0d630224",
    10434 => x"379b003c", 10435 => x"37820024", 10436 => x"34050200",
    10437 => x"e000000b", 10438 => x"2d640220", 10439 => x"40470000",
    10440 => x"34420001", 10441 => x"b5643000", 10442 => x"34840001",
    10443 => x"2084ffff", 10444 => x"30c70020", 10445 => x"0d640220",
    10446 => x"5c850002", 10447 => x"0d600220", 10448 => x"5c5bfff6",
    10449 => x"3463ffe8", 10450 => x"78020001", 10451 => x"2063ffff",
    10452 => x"38425b78", 10453 => x"0d630224", 10454 => x"b4223000",
    10455 => x"34050200", 10456 => x"e000000b", 10457 => x"2d640220",
    10458 => x"40480000", 10459 => x"34420001", 10460 => x"b5643800",
    10461 => x"34840001", 10462 => x"2084ffff", 10463 => x"30e80020",
    10464 => x"0d640220", 10465 => x"5c850002", 10466 => x"0d600220",
    10467 => x"5c46fff6", 10468 => x"c8610800", 10469 => x"0d610224",
    10470 => x"2d610226", 10471 => x"34210001", 10472 => x"0d610226",
    10473 => x"2b9d0004", 10474 => x"2b8b0020", 10475 => x"2b8c001c",
    10476 => x"2b8d0018", 10477 => x"2b8e0014", 10478 => x"2b8f0010",
    10479 => x"2b90000c", 10480 => x"2b9b0008", 10481 => x"379c003c",
    10482 => x"c3a00000", 10483 => x"379cffe8", 10484 => x"5b8b0008",
    10485 => x"5b9d0004", 10486 => x"378b000c", 10487 => x"b9600800",
    10488 => x"34020000", 10489 => x"3403000e", 10490 => x"f8001bd6",
    10491 => x"b9600800", 10492 => x"340200ff", 10493 => x"34030006",
    10494 => x"f8001bd2", 10495 => x"34010806", 10496 => x"0f810018",
    10497 => x"34020000", 10498 => x"b9601800", 10499 => x"34010000",
    10500 => x"fbfffe14", 10501 => x"78020001", 10502 => x"38425d68",
    10503 => x"58410000", 10504 => x"2b9d0004", 10505 => x"2b8b0008",
    10506 => x"379c0018", 10507 => x"c3a00000", 10508 => x"379cff38",
    10509 => x"5b8b0028", 10510 => x"5b8c0024", 10511 => x"5b8d0020",
    10512 => x"5b8e001c", 10513 => x"5b8f0018", 10514 => x"5b900014",
    10515 => x"5b910010", 10516 => x"5b92000c", 10517 => x"5b930008",
    10518 => x"5b9d0004", 10519 => x"78010001", 10520 => x"38215d6c",
    10521 => x"282c0000", 10522 => x"5d800047", 10523 => x"780b0001",
    10524 => x"396b5d68", 10525 => x"29610000", 10526 => x"378e00ac",
    10527 => x"378d002c", 10528 => x"b9c01000", 10529 => x"b9a01800",
    10530 => x"34040080", 10531 => x"34050000", 10532 => x"fbfffe7f",
    10533 => x"4d81003c", 10534 => x"3402001b", 10535 => x"4c41003a",
    10536 => x"378c00c4", 10537 => x"b9800800", 10538 => x"f800012a",
    10539 => x"43810032", 10540 => x"5c200035", 10541 => x"43930033",
    10542 => x"34010001", 10543 => x"5e610032", 10544 => x"378f0044",
    10545 => x"b9e00800", 10546 => x"b9801000", 10547 => x"34030004",
    10548 => x"f8001afd", 10549 => x"5c20002c", 10550 => x"379000bc",
    10551 => x"37920034", 10552 => x"ba401000", 10553 => x"34030006",
    10554 => x"ba000800", 10555 => x"f8001b17", 10556 => x"3791003a",
    10557 => x"ba201000", 10558 => x"34030004", 10559 => x"378100c8",
    10560 => x"f8001b12", 10561 => x"34010008", 10562 => x"3381002e",
    10563 => x"34010006", 10564 => x"33810030", 10565 => x"34010004",
    10566 => x"33810031", 10567 => x"34010002", 10568 => x"33810033",
    10569 => x"ba400800", 10570 => x"3380002c", 10571 => x"3393002d",
    10572 => x"3380002f", 10573 => x"33800032", 10574 => x"f800032b",
    10575 => x"b9801000", 10576 => x"34030004", 10577 => x"ba200800",
    10578 => x"f8001b00", 10579 => x"ba001000", 10580 => x"34030006",
    10581 => x"3781003e", 10582 => x"f8001afc", 10583 => x"378200c8",
    10584 => x"34030004", 10585 => x"b9e00800", 10586 => x"f8001af8",
    10587 => x"29610000", 10588 => x"b9c01000", 10589 => x"b9a01800",
    10590 => x"3404001c", 10591 => x"34050000", 10592 => x"fbfffedb",
    10593 => x"2b9d0004", 10594 => x"2b8b0028", 10595 => x"2b8c0024",
    10596 => x"2b8d0020", 10597 => x"2b8e001c", 10598 => x"2b8f0018",
    10599 => x"2b900014", 10600 => x"2b910010", 10601 => x"2b92000c",
    10602 => x"2b930008", 10603 => x"379c00c8", 10604 => x"c3a00000",
    10605 => x"379cffe0", 10606 => x"5b8b0018", 10607 => x"5b8c0014",
    10608 => x"5b8d0010", 10609 => x"5b8e000c", 10610 => x"5b8f0008",
    10611 => x"5b9d0004", 10612 => x"378d001c", 10613 => x"b8205800",
    10614 => x"b9a00800", 10615 => x"f80000dd", 10616 => x"41620000",
    10617 => x"34010045", 10618 => x"340c0000", 10619 => x"5c41004a",
    10620 => x"356e0010", 10621 => x"b9a01000", 10622 => x"b9c00800",
    10623 => x"34030004", 10624 => x"f8001ab1", 10625 => x"b8201000",
    10626 => x"5c200043", 10627 => x"41640009", 10628 => x"34030001",
    10629 => x"416d0002", 10630 => x"41610003", 10631 => x"b8406000",
    10632 => x"5c83003d", 10633 => x"41630014", 10634 => x"34020008",
    10635 => x"5c62003a", 10636 => x"3dad0008", 10637 => x"b9a16800",
    10638 => x"35adffe8", 10639 => x"34010040", 10640 => x"4c2d0002",
    10641 => x"340d0040", 10642 => x"356f000c", 10643 => x"b9e01000",
    10644 => x"34030004", 10645 => x"37810020", 10646 => x"f8001abc",
    10647 => x"35ac0018", 10648 => x"34010045", 10649 => x"31610000",
    10650 => x"15810008", 10651 => x"3782001c", 10652 => x"31610002",
    10653 => x"3401003f", 10654 => x"31610008", 10655 => x"34010001",
    10656 => x"31610009", 10657 => x"34030004", 10658 => x"31600001",
    10659 => x"316c0003", 10660 => x"31600004", 10661 => x"31600005",
    10662 => x"31600006", 10663 => x"31600007", 10664 => x"3160000a",
    10665 => x"3160000b", 10666 => x"b9e00800", 10667 => x"f8001aa7",
    10668 => x"34030004", 10669 => x"37820020", 10670 => x"b9c00800",
    10671 => x"f8001aa3", 10672 => x"35ad0005", 10673 => x"01a1001f",
    10674 => x"31600014", 10675 => x"b42d6800", 10676 => x"15a20001",
    10677 => x"31600015", 10678 => x"31600016", 10679 => x"31600017",
    10680 => x"35610014", 10681 => x"f8000015", 10682 => x"2021ffff",
    10683 => x"00220008", 10684 => x"31610017", 10685 => x"31620016",
    10686 => x"b9600800", 10687 => x"3402000a", 10688 => x"f800000e",
    10689 => x"2021ffff", 10690 => x"00220008", 10691 => x"3161000b",
    10692 => x"3162000a", 10693 => x"b9800800", 10694 => x"2b9d0004",
    10695 => x"2b8b0018", 10696 => x"2b8c0014", 10697 => x"2b8d0010",
    10698 => x"2b8e000c", 10699 => x"2b8f0008", 10700 => x"379c0020",
    10701 => x"c3a00000", 10702 => x"34030000", 10703 => x"34040000",
    10704 => x"e0000005", 10705 => x"2c250000", 10706 => x"34840001",
    10707 => x"34210002", 10708 => x"b4651800", 10709 => x"4844fffc",
    10710 => x"00610010", 10711 => x"2063ffff", 10712 => x"b4611800",
    10713 => x"00610010", 10714 => x"b4231800", 10715 => x"a4600800",
    10716 => x"2021ffff", 10717 => x"c3a00000", 10718 => x"379cffe8",
    10719 => x"5b8b0008", 10720 => x"5b9d0004", 10721 => x"78010001",
    10722 => x"378b000c", 10723 => x"38215d6c", 10724 => x"34020000",
    10725 => x"3403000e", 10726 => x"58200000", 10727 => x"b9600800",
    10728 => x"f8001ae8", 10729 => x"b9600800", 10730 => x"f800028f",
    10731 => x"34010800", 10732 => x"0f810018", 10733 => x"34020000",
    10734 => x"b9601800", 10735 => x"34010000", 10736 => x"fbfffd28",
    10737 => x"78020001", 10738 => x"38425d74", 10739 => x"58410000",
    10740 => x"2b9d0004", 10741 => x"2b8b0008", 10742 => x"379c0018",
    10743 => x"c3a00000", 10744 => x"379cfe50", 10745 => x"5b8b0010",
    10746 => x"5b8c000c", 10747 => x"5b8d0008", 10748 => x"5b9d0004",
    10749 => x"78020001", 10750 => x"38425d74", 10751 => x"28410000",
    10752 => x"378c0014", 10753 => x"378201a4", 10754 => x"b9801800",
    10755 => x"34040190", 10756 => x"34050000", 10757 => x"fbfffd9e",
    10758 => x"b8205800", 10759 => x"4c010019", 10760 => x"78020001",
    10761 => x"38425d6c", 10762 => x"28410000", 10763 => x"44200004",
    10764 => x"b9800800", 10765 => x"b9601000", 10766 => x"f800010a",
    10767 => x"78010001", 10768 => x"38215d6c", 10769 => x"282d0000",
    10770 => x"5da0000e", 10771 => x"378c0014", 10772 => x"b9800800",
    10773 => x"b9601000", 10774 => x"fbffff57", 10775 => x"b8202000",
    10776 => x"4da10008", 10777 => x"78020001", 10778 => x"38425d74",
    10779 => x"28410000", 10780 => x"b9801800", 10781 => x"378201a4",
    10782 => x"34050000", 10783 => x"fbfffe1c", 10784 => x"78010001",
    10785 => x"38215d6c", 10786 => x"28210000", 10787 => x"4420001d",
    10788 => x"78010001", 10789 => x"38215d78", 10790 => x"28210000",
    10791 => x"5c200019", 10792 => x"78010001", 10793 => x"38215d7c",
    10794 => x"28220000", 10795 => x"378b0014", 10796 => x"378c01a4",
    10797 => x"34420001", 10798 => x"58220000", 10799 => x"b9600800",
    10800 => x"f8000052", 10801 => x"b8206800", 10802 => x"340200ff",
    10803 => x"34030006", 10804 => x"b9800800", 10805 => x"f8001a9b",
    10806 => x"78050001", 10807 => x"34010800", 10808 => x"38a55d74",
    10809 => x"0f8101b0", 10810 => x"28a10000", 10811 => x"b9801000",
    10812 => x"b9601800", 10813 => x"b9a02000", 10814 => x"34050000",
    10815 => x"fbfffdfc", 10816 => x"78010001", 10817 => x"38215d6c",
    10818 => x"28210000", 10819 => x"4420000b", 10820 => x"78010001",
    10821 => x"38215d78", 10822 => x"28220000", 10823 => x"78040001",
    10824 => x"38843d14", 10825 => x"28830000", 10826 => x"34420001",
    10827 => x"58220000", 10828 => x"5c430002", 10829 => x"58200000",
    10830 => x"2b9d0004", 10831 => x"2b8b0010", 10832 => x"2b8c000c",
    10833 => x"2b8d0008", 10834 => x"379c01b0", 10835 => x"c3a00000",
    10836 => x"379cfffc", 10837 => x"5b9d0004", 10838 => x"78020001",
    10839 => x"38425d70", 10840 => x"34030004", 10841 => x"f80019f9",
    10842 => x"2b9d0004", 10843 => x"379c0004", 10844 => x"c3a00000",
    10845 => x"379cfff0", 10846 => x"5b8b0010", 10847 => x"5b8c000c",
    10848 => x"5b8d0008", 10849 => x"5b9d0004", 10850 => x"78030001",
    10851 => x"780b0001", 10852 => x"396b5d70", 10853 => x"b8206000",
    10854 => x"38636dc8", 10855 => x"286d0000", 10856 => x"b9801000",
    10857 => x"34030004", 10858 => x"b9600800", 10859 => x"f80019e7",
    10860 => x"41620000", 10861 => x"41610001", 10862 => x"3c420018",
    10863 => x"3c210010", 10864 => x"b8410800", 10865 => x"41620003",
    10866 => x"b8220800", 10867 => x"41620002", 10868 => x"3c420008",
    10869 => x"b8220800", 10870 => x"59a10018", 10871 => x"b9800800",
    10872 => x"f8000926", 10873 => x"78010001", 10874 => x"38215d6c",
    10875 => x"58200000", 10876 => x"2b9d0004", 10877 => x"2b8b0010",
    10878 => x"2b8c000c", 10879 => x"2b8d0008", 10880 => x"379c0010",
    10881 => x"c3a00000", 10882 => x"379cffe8", 10883 => x"5b8b0018",
    10884 => x"5b8c0014", 10885 => x"5b8d0010", 10886 => x"5b8e000c",
    10887 => x"5b8f0008", 10888 => x"5b9d0004", 10889 => x"340c0001",
    10890 => x"b8205800", 10891 => x"302c001c", 10892 => x"302c001d",
    10893 => x"34010006", 10894 => x"3161001e", 10895 => x"3160001f",
    10896 => x"35610020", 10897 => x"b8406800", 10898 => x"f80001e7",
    10899 => x"41620024", 10900 => x"41610020", 10901 => x"34030002",
    10902 => x"356e0008", 10903 => x"98410800", 10904 => x"31610020",
    10905 => x"41620025", 10906 => x"41610021", 10907 => x"316d0025",
    10908 => x"356f0010", 10909 => x"98410800", 10910 => x"41620022",
    10911 => x"31610021", 10912 => x"15a10008", 10913 => x"98221000",
    10914 => x"31620022", 10915 => x"41620023", 10916 => x"31610024",
    10917 => x"35610026", 10918 => x"984d1000", 10919 => x"31620023",
    10920 => x"34020000", 10921 => x"f8001a27", 10922 => x"34020000",
    10923 => x"34030004", 10924 => x"35610028", 10925 => x"f8001a23",
    10926 => x"34020000", 10927 => x"34030004", 10928 => x"3561002c",
    10929 => x"f8001a1f", 10930 => x"34020000", 10931 => x"34030004",
    10932 => x"35610030", 10933 => x"f8001a1b", 10934 => x"34020000",
    10935 => x"34030004", 10936 => x"35610034", 10937 => x"f8001a17",
    10938 => x"356d0038", 10939 => x"34020000", 10940 => x"34030010",
    10941 => x"b9a00800", 10942 => x"f8001a12", 10943 => x"b9a00800",
    10944 => x"f80001b9", 10945 => x"34020000", 10946 => x"34030040",
    10947 => x"35610048", 10948 => x"f8001a0c", 10949 => x"34020000",
    10950 => x"34030080", 10951 => x"35610088", 10952 => x"f8001a08",
    10953 => x"34020000", 10954 => x"34030040", 10955 => x"35610108",
    10956 => x"f8001a04", 10957 => x"34020000", 10958 => x"34030004",
    10959 => x"b9c00800", 10960 => x"f8001a00", 10961 => x"356d000c",
    10962 => x"340200ff", 10963 => x"34030004", 10964 => x"b9a00800",
    10965 => x"f80019fb", 10966 => x"34010011", 10967 => x"31610011",
    10968 => x"34010044", 10969 => x"34020034", 10970 => x"31610015",
    10971 => x"34010043", 10972 => x"31620013", 10973 => x"31610017",
    10974 => x"31620019", 10975 => x"31600010", 10976 => x"340200a0",
    10977 => x"316c0012", 10978 => x"31600014", 10979 => x"31600016",
    10980 => x"316c0018", 10981 => x"3160001a", 10982 => x"3160001b",
    10983 => x"b9c00800", 10984 => x"fbfffee6", 10985 => x"2022ffff",
    10986 => x"5c400002", 10987 => x"3802ffff", 10988 => x"00410008",
    10989 => x"3162001b", 10990 => x"3161001a", 10991 => x"34010045",
    10992 => x"31610000", 10993 => x"34010001", 10994 => x"31610002",
    10995 => x"34010048", 10996 => x"31610003", 10997 => x"3401003f",
    10998 => x"31610008", 10999 => x"34010011", 11000 => x"31610009",
    11001 => x"31600001", 11002 => x"31600004", 11003 => x"31600005",
    11004 => x"31600006", 11005 => x"31600007", 11006 => x"3160000a",
    11007 => x"3160000b", 11008 => x"b9a00800", 11009 => x"34020000",
    11010 => x"34030004", 11011 => x"f80019cd", 11012 => x"34030004",
    11013 => x"b9e00800", 11014 => x"340200ff", 11015 => x"f80019c9",
    11016 => x"b9600800", 11017 => x"3402000a", 11018 => x"fbfffec4",
    11019 => x"2021ffff", 11020 => x"00220008", 11021 => x"3161000b",
    11022 => x"34010148", 11023 => x"3162000a", 11024 => x"2b9d0004",
    11025 => x"2b8b0018", 11026 => x"2b8c0014", 11027 => x"2b8d0010",
    11028 => x"2b8e000c", 11029 => x"2b8f0008", 11030 => x"379c0018",
    11031 => x"c3a00000", 11032 => x"379cffe0", 11033 => x"5b8b0014",
    11034 => x"5b8c0010", 11035 => x"5b8d000c", 11036 => x"5b8e0008",
    11037 => x"5b9d0004", 11038 => x"378d0018", 11039 => x"b8205800",
    11040 => x"b9a00800", 11041 => x"b8407000", 11042 => x"f8000157",
    11043 => x"34010148", 11044 => x"340c0000", 11045 => x"5dc10022",
    11046 => x"41620000", 11047 => x"34010045", 11048 => x"5c41001f",
    11049 => x"41620009", 11050 => x"34010011", 11051 => x"5c41001c",
    11052 => x"41610016", 11053 => x"5c20001a", 11054 => x"41620017",
    11055 => x"34010044", 11056 => x"5c410017", 11057 => x"41610014",
    11058 => x"5c200015", 11059 => x"41620015", 11060 => x"34010043",
    11061 => x"5c410012", 11062 => x"35610038", 11063 => x"b9a01000",
    11064 => x"34030006", 11065 => x"f80018f8", 11066 => x"5c20000d",
    11067 => x"3561002c", 11068 => x"fbffff21", 11069 => x"37810020",
    11070 => x"fbffff16", 11071 => x"43820020", 11072 => x"43830021",
    11073 => x"43840022", 11074 => x"43850023", 11075 => x"78010001",
    11076 => x"38213548", 11077 => x"f800002c", 11078 => x"340c0001",
    11079 => x"b9800800", 11080 => x"2b9d0004", 11081 => x"2b8b0014",
    11082 => x"2b8c0010", 11083 => x"2b8d000c", 11084 => x"2b8e0008",
    11085 => x"379c0020", 11086 => x"c3a00000", 11087 => x"379cfff4",
    11088 => x"5b8b000c", 11089 => x"5b8c0008", 11090 => x"5b9d0004",
    11091 => x"780b0001", 11092 => x"b8202000", 11093 => x"396b5d80",
    11094 => x"b8401800", 11095 => x"b9600800", 11096 => x"b8801000",
    11097 => x"f8000027", 11098 => x"b8206000", 11099 => x"b9600800",
    11100 => x"f8000e9f", 11101 => x"b9800800", 11102 => x"2b9d0004",
    11103 => x"2b8b000c", 11104 => x"2b8c0008", 11105 => x"379c000c",
    11106 => x"c3a00000", 11107 => x"379cffe0", 11108 => x"5b9d0004",
    11109 => x"5b83000c", 11110 => x"3783000c", 11111 => x"5b820008",
    11112 => x"5b840010", 11113 => x"5b850014", 11114 => x"5b860018",
    11115 => x"5b87001c", 11116 => x"5b880020", 11117 => x"f8000013",
    11118 => x"2b9d0004", 11119 => x"379c0020", 11120 => x"c3a00000",
    11121 => x"379cffdc", 11122 => x"5b9d0004", 11123 => x"5b82000c",
    11124 => x"3782000c", 11125 => x"5b810008", 11126 => x"5b830010",
    11127 => x"5b840014", 11128 => x"5b850018", 11129 => x"5b86001c",
    11130 => x"5b870020", 11131 => x"5b880024", 11132 => x"fbffffd3",
    11133 => x"2b9d0004", 11134 => x"379c0024", 11135 => x"c3a00000",
    11136 => x"379cff94", 11137 => x"5b8b0044", 11138 => x"5b8c0040",
    11139 => x"5b8d003c", 11140 => x"5b8e0038", 11141 => x"5b8f0034",
    11142 => x"5b900030", 11143 => x"5b91002c", 11144 => x"5b920028",
    11145 => x"5b930024", 11146 => x"5b940020", 11147 => x"5b95001c",
    11148 => x"5b960018", 11149 => x"5b970014", 11150 => x"5b980010",
    11151 => x"5b99000c", 11152 => x"5b9b0008", 11153 => x"5b9d0004",
    11154 => x"78160001", 11155 => x"b820c800", 11156 => x"b840a000",
    11157 => x"b8209800", 11158 => x"34180025", 11159 => x"34090069",
    11160 => x"34080070", 11161 => x"34070058", 11162 => x"34060063",
    11163 => x"34050064", 11164 => x"341b002a", 11165 => x"340a0030",
    11166 => x"34170010", 11167 => x"37950060", 11168 => x"3ad63570",
    11169 => x"e0000093", 11170 => x"34110001", 11171 => x"34100020",
    11172 => x"340e000a", 11173 => x"44380004", 11174 => x"32610000",
    11175 => x"e0000038", 11176 => x"34100030", 11177 => x"36940001",
    11178 => x"42810000", 11179 => x"4429003c", 11180 => x"5429000d",
    11181 => x"44270037", 11182 => x"54270008", 11183 => x"443b0018",
    11184 => x"543b0004", 11185 => x"44200085", 11186 => x"5c380017",
    11187 => x"e000002b", 11188 => x"5c2a0015", 11189 => x"e3fffff3",
    11190 => x"44260019", 11191 => x"5c250012", 11192 => x"e000002f",
    11193 => x"4428002b", 11194 => x"54280006", 11195 => x"3402006e",
    11196 => x"44220077", 11197 => x"3404006f", 11198 => x"5c24000b",
    11199 => x"e0000022", 11200 => x"34020075", 11201 => x"44220026",
    11202 => x"34040078", 11203 => x"44240021", 11204 => x"34020073",
    11205 => x"5c220004", 11206 => x"e000000e", 11207 => x"286e0000",
    11208 => x"34630004", 11209 => x"3422ffcf", 11210 => x"204200ff",
    11211 => x"34040008", 11212 => x"5444ffdd", 11213 => x"3431ffd0",
    11214 => x"e3ffffdb", 11215 => x"28610000", 11216 => x"34630004",
    11217 => x"32610000", 11218 => x"36730001", 11219 => x"e0000060",
    11220 => x"b8600800", 11221 => x"28210000", 11222 => x"34630004",
    11223 => x"e0000004", 11224 => x"32620000", 11225 => x"34210001",
    11226 => x"36730001", 11227 => x"40220000", 11228 => x"5c40fffc",
    11229 => x"e0000056", 11230 => x"32780000", 11231 => x"36730001",
    11232 => x"e0000053", 11233 => x"3401000a", 11234 => x"45c10004",
    11235 => x"e0000004", 11236 => x"340e0010", 11237 => x"e0000002",
    11238 => x"340e0008", 11239 => x"286d0000", 11240 => x"34720004",
    11241 => x"65c3000a", 11242 => x"01a4001f", 11243 => x"340f0000",
    11244 => x"a0831800", 11245 => x"44600003", 11246 => x"c80d6800",
    11247 => x"340f0001", 11248 => x"340c0010", 11249 => x"e0000019",
    11250 => x"b9a00800", 11251 => x"b9c01000", 11252 => x"5b85004c",
    11253 => x"5b860050", 11254 => x"5b870054", 11255 => x"5b880058",
    11256 => x"5b89005c", 11257 => x"5b8a0048", 11258 => x"f8001807",
    11259 => x"b6c11800", 11260 => x"40630000", 11261 => x"358cffff",
    11262 => x"b6ac5800", 11263 => x"b9a00800", 11264 => x"31630000",
    11265 => x"b9c01000", 11266 => x"f80017ef", 11267 => x"2b8a0048",
    11268 => x"2b89005c", 11269 => x"2b880058", 11270 => x"2b870054",
    11271 => x"2b860050", 11272 => x"2b85004c", 11273 => x"b8206800",
    11274 => x"7d840000", 11275 => x"7da30000", 11276 => x"a0831800",
    11277 => x"5c60ffe5", 11278 => x"5d970004", 11279 => x"34020030",
    11280 => x"3382006f", 11281 => x"340c000f", 11282 => x"66020020",
    11283 => x"a1e21000", 11284 => x"4440000b", 11285 => x"358cffff",
    11286 => x"b6ac1000", 11287 => x"3403002d", 11288 => x"30430000",
    11289 => x"340f0000", 11290 => x"e0000005", 11291 => x"358cffff",
    11292 => x"b6ac1000", 11293 => x"30500000", 11294 => x"e0000003",
    11295 => x"caf10800", 11296 => x"b42f0800", 11297 => x"4981fffa",
    11298 => x"45e00005", 11299 => x"358cffff", 11300 => x"b6ac0800",
    11301 => x"3402002d", 11302 => x"30220000", 11303 => x"caec1800",
    11304 => x"ba600800", 11305 => x"3404000f", 11306 => x"e0000006",
    11307 => x"b6ac1000", 11308 => x"40420000", 11309 => x"358c0001",
    11310 => x"30220000", 11311 => x"34210001", 11312 => x"4c8cfffb",
    11313 => x"b6639800", 11314 => x"ba401800", 11315 => x"36940001",
    11316 => x"42810000", 11317 => x"5c20ff6d", 11318 => x"ca790800",
    11319 => x"32600000", 11320 => x"2b9d0004", 11321 => x"2b8b0044",
    11322 => x"2b8c0040", 11323 => x"2b8d003c", 11324 => x"2b8e0038",
    11325 => x"2b8f0034", 11326 => x"2b900030", 11327 => x"2b91002c",
    11328 => x"2b920028", 11329 => x"2b930024", 11330 => x"2b940020",
    11331 => x"2b95001c", 11332 => x"2b960018", 11333 => x"2b970014",
    11334 => x"2b980010", 11335 => x"2b99000c", 11336 => x"2b9b0008",
    11337 => x"379c006c", 11338 => x"c3a00000", 11339 => x"78020001",
    11340 => x"14210002", 11341 => x"38426dbc", 11342 => x"28420000",
    11343 => x"202100ff", 11344 => x"3c210010", 11345 => x"5841002c",
    11346 => x"28410030", 11347 => x"4c20ffff", 11348 => x"28410030",
    11349 => x"2021ffff", 11350 => x"c3a00000", 11351 => x"14210002",
    11352 => x"78030001", 11353 => x"38636dbc", 11354 => x"202100ff",
    11355 => x"28630000", 11356 => x"2042ffff", 11357 => x"78048000",
    11358 => x"3c210010", 11359 => x"b8441000", 11360 => x"b8411000",
    11361 => x"5862002c", 11362 => x"28610030", 11363 => x"4c20ffff",
    11364 => x"c3a00000", 11365 => x"40240002", 11366 => x"40230003",
    11367 => x"78020001", 11368 => x"3c840018", 11369 => x"3c630010",
    11370 => x"38426dbc", 11371 => x"b8831800", 11372 => x"40240005",
    11373 => x"28420000", 11374 => x"b8641800", 11375 => x"40240004",
    11376 => x"3c840008", 11377 => x"b8641800", 11378 => x"58430028",
    11379 => x"40230001", 11380 => x"40210000", 11381 => x"3c210008",
    11382 => x"b8610800", 11383 => x"58410024", 11384 => x"c3a00000",
    11385 => x"78020001", 11386 => x"38426dbc", 11387 => x"28430000",
    11388 => x"28630028", 11389 => x"30230005", 11390 => x"28430000",
    11391 => x"28630028", 11392 => x"00630008", 11393 => x"30230004",
    11394 => x"28430000", 11395 => x"28630028", 11396 => x"00630010",
    11397 => x"30230003", 11398 => x"28430000", 11399 => x"28630028",
    11400 => x"00630018", 11401 => x"30230002", 11402 => x"28430000",
    11403 => x"28630024", 11404 => x"30230001", 11405 => x"28420000",
    11406 => x"28420024", 11407 => x"00420008", 11408 => x"30220000",
    11409 => x"c3a00000", 11410 => x"379cfff4", 11411 => x"5b8b000c",
    11412 => x"5b8c0008", 11413 => x"5b9d0004", 11414 => x"780b0001",
    11415 => x"b8406000", 11416 => x"396b6dbc", 11417 => x"5c200004",
    11418 => x"29610000", 11419 => x"58200000", 11420 => x"e0000022",
    11421 => x"29610000", 11422 => x"58200000", 11423 => x"28220034",
    11424 => x"78010001", 11425 => x"38213584", 11426 => x"fbfffecf",
    11427 => x"f80000be", 11428 => x"29610000", 11429 => x"340200e0",
    11430 => x"58220000", 11431 => x"78010001", 11432 => x"38215e00",
    11433 => x"34020800", 11434 => x"582c0000", 11435 => x"34010000",
    11436 => x"fbffffab", 11437 => x"340100c8", 11438 => x"f80004fa",
    11439 => x"34010000", 11440 => x"38028000", 11441 => x"fbffffa6",
    11442 => x"34010000", 11443 => x"34020000", 11444 => x"fbffffa3",
    11445 => x"34010010", 11446 => x"34020000", 11447 => x"fbffffa0",
    11448 => x"7d820000", 11449 => x"34010000", 11450 => x"c8021000",
    11451 => x"20421200", 11452 => x"34420140", 11453 => x"fbffff9a",
    11454 => x"34010000", 11455 => x"2b9d0004", 11456 => x"2b8b000c",
    11457 => x"2b8c0008", 11458 => x"379c000c", 11459 => x"c3a00000",
    11460 => x"379cfff0", 11461 => x"5b8b000c", 11462 => x"5b8c0008",
    11463 => x"5b9d0004", 11464 => x"78020001", 11465 => x"38425e00",
    11466 => x"284b0000", 11467 => x"b8206000", 11468 => x"34010004",
    11469 => x"fbffff7e", 11470 => x"7d6b0000", 11471 => x"0f810012",
    11472 => x"34010004", 11473 => x"c80b5800", 11474 => x"fbffff79",
    11475 => x"216b0020", 11476 => x"0f810012", 11477 => x"356b0004",
    11478 => x"45800004", 11479 => x"34010014", 11480 => x"fbffff73",
    11481 => x"0d810000", 11482 => x"2f810012", 11483 => x"a1610800",
    11484 => x"e42b0800", 11485 => x"2b9d0004", 11486 => x"2b8b000c",
    11487 => x"2b8c0008", 11488 => x"379c0010", 11489 => x"c3a00000",
    11490 => x"379cfffc", 11491 => x"5b9d0004", 11492 => x"34010040",
    11493 => x"fbffff66", 11494 => x"00210004", 11495 => x"2021001f",
    11496 => x"08210320", 11497 => x"2b9d0004", 11498 => x"379c0004",
    11499 => x"c3a00000", 11500 => x"379cfff4", 11501 => x"5b8b000c",
    11502 => x"5b8c0008", 11503 => x"5b9d0004", 11504 => x"78030001",
    11505 => x"38634e6c", 11506 => x"b8405800", 11507 => x"28620000",
    11508 => x"58220000", 11509 => x"78010001", 11510 => x"38214e70",
    11511 => x"282c0000", 11512 => x"34010040", 11513 => x"fbffff52",
    11514 => x"00210004", 11515 => x"2021001f", 11516 => x"08210320",
    11517 => x"b42c0800", 11518 => x"59610000", 11519 => x"34010000",
    11520 => x"2b9d0004", 11521 => x"2b8b000c", 11522 => x"2b8c0008",
    11523 => x"379c000c", 11524 => x"c3a00000", 11525 => x"379cfffc",
    11526 => x"5b9d0004", 11527 => x"34010040", 11528 => x"fbffff43",
    11529 => x"38220001", 11530 => x"34010040", 11531 => x"fbffff4c",
    11532 => x"34010000", 11533 => x"2b9d0004", 11534 => x"379c0004",
    11535 => x"c3a00000", 11536 => x"379cfffc", 11537 => x"5b9d0004",
    11538 => x"34010040", 11539 => x"fbffff38", 11540 => x"3402fffe",
    11541 => x"a0221000", 11542 => x"34010040", 11543 => x"fbffff40",
    11544 => x"34010000", 11545 => x"2b9d0004", 11546 => x"379c0004",
    11547 => x"c3a00000", 11548 => x"379cfff8", 11549 => x"5b8b0008",
    11550 => x"5b9d0004", 11551 => x"780b0001", 11552 => x"396b6dbc",
    11553 => x"29610000", 11554 => x"28220004", 11555 => x"38420010",
    11556 => x"58220004", 11557 => x"34010001", 11558 => x"f8000482",
    11559 => x"29610000", 11560 => x"28210004", 11561 => x"20210020",
    11562 => x"7c210000", 11563 => x"2b9d0004", 11564 => x"2b8b0008",
    11565 => x"379c0008", 11566 => x"c3a00000", 11567 => x"379cfff8",
    11568 => x"5b8b0008", 11569 => x"5b9d0004", 11570 => x"b8205800",
    11571 => x"34010044", 11572 => x"fbffff17", 11573 => x"38220020",
    11574 => x"45600003", 11575 => x"3402ffdf", 11576 => x"a0221000",
    11577 => x"34010044", 11578 => x"fbffff1d", 11579 => x"34010000",
    11580 => x"2b9d0004", 11581 => x"2b8b0008", 11582 => x"379c0008",
    11583 => x"c3a00000", 11584 => x"379cfff8", 11585 => x"5b8b0008",
    11586 => x"5b9d0004", 11587 => x"78020001", 11588 => x"38426d00",
    11589 => x"28420000", 11590 => x"780b0001", 11591 => x"396b6dbc",
    11592 => x"59620000", 11593 => x"fbffff1c", 11594 => x"34010001",
    11595 => x"fbffffe4", 11596 => x"78020001", 11597 => x"38423d18",
    11598 => x"28410000", 11599 => x"78040001", 11600 => x"38843d1c",
    11601 => x"58200000", 11602 => x"29610000", 11603 => x"28830000",
    11604 => x"34020003", 11605 => x"58200000", 11606 => x"5822000c",
    11607 => x"58230008", 11608 => x"78030001", 11609 => x"38633d20",
    11610 => x"58220004", 11611 => x"28620000", 11612 => x"5822003c",
    11613 => x"2b9d0004", 11614 => x"2b8b0008", 11615 => x"379c0008",
    11616 => x"c3a00000", 11617 => x"379cfffc", 11618 => x"5b9d0004",
    11619 => x"78010001", 11620 => x"78040001", 11621 => x"38214ad4",
    11622 => x"38843d24", 11623 => x"28220000", 11624 => x"28830000",
    11625 => x"44430012", 11626 => x"78030001", 11627 => x"38634ba0",
    11628 => x"780500ff", 11629 => x"e000000d", 11630 => x"28240000",
    11631 => x"3c870018", 11632 => x"00860018", 11633 => x"b8e63000",
    11634 => x"a0853800", 11635 => x"00e70008", 11636 => x"2084ff00",
    11637 => x"3c840008", 11638 => x"b8c73000", 11639 => x"b8c42000",
    11640 => x"58240000", 11641 => x"34210004", 11642 => x"5461fff4",
    11643 => x"78010001", 11644 => x"78050001", 11645 => x"38214ad4",
    11646 => x"38a53d24", 11647 => x"28240000", 11648 => x"28a30000",
    11649 => x"44830005", 11650 => x"78010001", 11651 => x"3821358c",
    11652 => x"fbfffded", 11653 => x"e000004f", 11654 => x"78020001",
    11655 => x"38425e04", 11656 => x"28430000", 11657 => x"5c600016",
    11658 => x"2824000c", 11659 => x"34031234", 11660 => x"0084000d",
    11661 => x"2084ffff", 11662 => x"5c83000b", 11663 => x"28240014",
    11664 => x"34035678", 11665 => x"0084000d", 11666 => x"2084ffff",
    11667 => x"5c830006", 11668 => x"2823001c", 11669 => x"38019abc",
    11670 => x"0063000d", 11671 => x"2063ffff", 11672 => x"44610005",
    11673 => x"78010001", 11674 => x"382135b4", 11675 => x"fbfffdd6",
    11676 => x"e0000038", 11677 => x"34010001", 11678 => x"58410000",
    11679 => x"78020001", 11680 => x"38423d28", 11681 => x"28430000",
    11682 => x"78020001", 11683 => x"38426dbc", 11684 => x"28420000",
    11685 => x"78010001", 11686 => x"38214ad4", 11687 => x"28460024",
    11688 => x"28250014", 11689 => x"2824001c", 11690 => x"2827000c",
    11691 => x"20c6ffff", 11692 => x"3cc6000d", 11693 => x"a0832000",
    11694 => x"a0a32800", 11695 => x"a0e31800", 11696 => x"b8c31800",
    11697 => x"5823000c", 11698 => x"28430028", 11699 => x"00630010",
    11700 => x"3c63000d", 11701 => x"b8651800", 11702 => x"58230014",
    11703 => x"28430028", 11704 => x"2063ffff", 11705 => x"3c63000d",
    11706 => x"b8641800", 11707 => x"5823001c", 11708 => x"78010001",
    11709 => x"78030001", 11710 => x"58400014", 11711 => x"34040000",
    11712 => x"38214ad8", 11713 => x"38634ba0", 11714 => x"e000000f",
    11715 => x"28250000", 11716 => x"28270004", 11717 => x"34210008",
    11718 => x"20a60fff", 11719 => x"3ce70014", 11720 => x"00a5000c",
    11721 => x"58460018", 11722 => x"b8e52800", 11723 => x"3ca50008",
    11724 => x"2087003f", 11725 => x"38a50040", 11726 => x"b8a72800",
    11727 => x"58450014", 11728 => x"34840001", 11729 => x"5461fff2",
    11730 => x"34010080", 11731 => x"58410014", 11732 => x"2b9d0004",
    11733 => x"379c0004", 11734 => x"c3a00000", 11735 => x"78030001",
    11736 => x"38636db8", 11737 => x"44400004", 11738 => x"28620000",
    11739 => x"58410004", 11740 => x"c3a00000", 11741 => x"28620000",
    11742 => x"58410008", 11743 => x"c3a00000", 11744 => x"78030001",
    11745 => x"38636db8", 11746 => x"44400004", 11747 => x"28620000",
    11748 => x"58410004", 11749 => x"c3a00000", 11750 => x"28620000",
    11751 => x"58410008", 11752 => x"c3a00000", 11753 => x"3401012c",
    11754 => x"34000000", 11755 => x"3421ffff", 11756 => x"5c20fffe",
    11757 => x"c3a00000", 11758 => x"379cfff8", 11759 => x"5b8b0008",
    11760 => x"5b9d0004", 11761 => x"202100ff", 11762 => x"3c2b0003",
    11763 => x"78020001", 11764 => x"38424ba0", 11765 => x"b44b5800",
    11766 => x"29610004", 11767 => x"34020000", 11768 => x"fbffffdf",
    11769 => x"fbfffff0", 11770 => x"29610000", 11771 => x"34020000",
    11772 => x"fbffffdb", 11773 => x"fbffffec", 11774 => x"2b9d0004",
    11775 => x"2b8b0008", 11776 => x"379c0008", 11777 => x"c3a00000",
    11778 => x"379cfff8", 11779 => x"5b8b0008", 11780 => x"5b9d0004",
    11781 => x"202100ff", 11782 => x"3c2b0003", 11783 => x"78020001",
    11784 => x"38424ba0", 11785 => x"b44b5800", 11786 => x"29610004",
    11787 => x"34020001", 11788 => x"fbffffcb", 11789 => x"fbffffdc",
    11790 => x"29610000", 11791 => x"34020001", 11792 => x"fbffffc7",
    11793 => x"fbffffd8", 11794 => x"29610004", 11795 => x"34020000",
    11796 => x"fbffffc3", 11797 => x"fbffffd4", 11798 => x"29610000",
    11799 => x"34020000", 11800 => x"fbffffbf", 11801 => x"fbffffd0",
    11802 => x"2b9d0004", 11803 => x"2b8b0008", 11804 => x"379c0008",
    11805 => x"c3a00000", 11806 => x"379cfff8", 11807 => x"5b8b0008",
    11808 => x"5b9d0004", 11809 => x"202100ff", 11810 => x"3c2b0003",
    11811 => x"78020001", 11812 => x"38424ba0", 11813 => x"b44b5800",
    11814 => x"29610004", 11815 => x"34020000", 11816 => x"fbffffaf",
    11817 => x"fbffffc0", 11818 => x"29610000", 11819 => x"34020001",
    11820 => x"fbffffab", 11821 => x"fbffffbc", 11822 => x"29610004",
    11823 => x"34020001", 11824 => x"fbffffa7", 11825 => x"fbffffb8",
    11826 => x"2b9d0004", 11827 => x"2b8b0008", 11828 => x"379c0008",
    11829 => x"c3a00000", 11830 => x"379cffec", 11831 => x"5b8b0014",
    11832 => x"5b8c0010", 11833 => x"5b8d000c", 11834 => x"5b8e0008",
    11835 => x"5b9d0004", 11836 => x"202100ff", 11837 => x"78030001",
    11838 => x"3c2b0003", 11839 => x"38634ba0", 11840 => x"204e00ff",
    11841 => x"340d0008", 11842 => x"b46b5800", 11843 => x"29610004",
    11844 => x"21c20080", 11845 => x"35adffff", 11846 => x"fbffff91",
    11847 => x"fbffffa2", 11848 => x"29610000", 11849 => x"34020001",
    11850 => x"3dce0001", 11851 => x"fbffff8c", 11852 => x"fbffff9d",
    11853 => x"29610000", 11854 => x"34020000", 11855 => x"21ad00ff",
    11856 => x"fbffff87", 11857 => x"356c0004", 11858 => x"fbffff97",
    11859 => x"21ce00ff", 11860 => x"5da0ffef", 11861 => x"29810000",
    11862 => x"34020001", 11863 => x"fbffff80", 11864 => x"fbffff91",
    11865 => x"29610000", 11866 => x"34020001", 11867 => x"fbffff7c",
    11868 => x"fbffff8d", 11869 => x"78010001", 11870 => x"38216db8",
    11871 => x"28210000", 11872 => x"298d0000", 11873 => x"34020000",
    11874 => x"28210004", 11875 => x"a02d6800", 11876 => x"29610000",
    11877 => x"fbffff72", 11878 => x"fbffff83", 11879 => x"29810000",
    11880 => x"34020000", 11881 => x"fbffff6e", 11882 => x"fbffff7f",
    11883 => x"7da10000", 11884 => x"2b9d0004", 11885 => x"2b8b0014",
    11886 => x"2b8c0010", 11887 => x"2b8d000c", 11888 => x"2b8e0008",
    11889 => x"379c0014", 11890 => x"c3a00000", 11891 => x"379cffe0",
    11892 => x"5b8b0020", 11893 => x"5b8c001c", 11894 => x"5b8d0018",
    11895 => x"5b8e0014", 11896 => x"5b8f0010", 11897 => x"5b90000c",
    11898 => x"5b910008", 11899 => x"5b9d0004", 11900 => x"202100ff",
    11901 => x"3c2b0003", 11902 => x"78040001", 11903 => x"38844ba0",
    11904 => x"b48b5800", 11905 => x"29610004", 11906 => x"b8407800",
    11907 => x"34020001", 11908 => x"207000ff", 11909 => x"fbffff52",
    11910 => x"fbffff63", 11911 => x"29610000", 11912 => x"34020000",
    11913 => x"780d0001", 11914 => x"fbffff4d", 11915 => x"340c0000",
    11916 => x"fbffff5d", 11917 => x"340e0000", 11918 => x"39ad6db8",
    11919 => x"34110008", 11920 => x"29610000", 11921 => x"34020001",
    11922 => x"3d8c0001", 11923 => x"fbffff44", 11924 => x"fbffff55",
    11925 => x"29a10000", 11926 => x"29620004", 11927 => x"218c00ff",
    11928 => x"28210004", 11929 => x"a0220800", 11930 => x"44200002",
    11931 => x"398c0001", 11932 => x"29610000", 11933 => x"34020000",
    11934 => x"35ce0001", 11935 => x"fbffff38", 11936 => x"fbffff49",
    11937 => x"5dd1ffef", 11938 => x"46000004", 11939 => x"29610004",
    11940 => x"34020001", 11941 => x"e0000003", 11942 => x"29610004",
    11943 => x"34020000", 11944 => x"fbffff2f", 11945 => x"fbffff40",
    11946 => x"29610000", 11947 => x"34020001", 11948 => x"fbffff2b",
    11949 => x"fbffff3c", 11950 => x"29610000", 11951 => x"34020000",
    11952 => x"fbffff27", 11953 => x"fbffff38", 11954 => x"31ec0000",
    11955 => x"2b9d0004", 11956 => x"2b8b0020", 11957 => x"2b8c001c",
    11958 => x"2b8d0018", 11959 => x"2b8e0014", 11960 => x"2b8f0010",
    11961 => x"2b90000c", 11962 => x"2b910008", 11963 => x"379c0020",
    11964 => x"c3a00000", 11965 => x"379cfff8", 11966 => x"5b8b0008",
    11967 => x"5b9d0004", 11968 => x"202100ff", 11969 => x"3c2b0003",
    11970 => x"78020001", 11971 => x"38424ba0", 11972 => x"b44b5800",
    11973 => x"29610000", 11974 => x"34020001", 11975 => x"fbffff10",
    11976 => x"fbffff21", 11977 => x"29610004", 11978 => x"34020001",
    11979 => x"fbffff0c", 11980 => x"fbffff1d", 11981 => x"2b9d0004",
    11982 => x"2b8b0008", 11983 => x"379c0008", 11984 => x"c3a00000",
    11985 => x"379cfff4", 11986 => x"5b8b000c", 11987 => x"5b8c0008",
    11988 => x"5b9d0004", 11989 => x"202b00ff", 11990 => x"b9600800",
    11991 => x"204c00ff", 11992 => x"fbffff16", 11993 => x"3d820001",
    11994 => x"b9600800", 11995 => x"204200fe", 11996 => x"fbffff5a",
    11997 => x"b8206000", 11998 => x"b9600800", 11999 => x"fbffff3f",
    12000 => x"65810000", 12001 => x"2b9d0004", 12002 => x"2b8b000c",
    12003 => x"2b8c0008", 12004 => x"379c000c", 12005 => x"c3a00000",
    12006 => x"379cffe8", 12007 => x"5b8b0018", 12008 => x"5b8c0014",
    12009 => x"5b8d0010", 12010 => x"5b8e000c", 12011 => x"5b8f0008",
    12012 => x"5b9d0004", 12013 => x"780b0001", 12014 => x"396b5e08",
    12015 => x"296d000c", 12016 => x"296f0004", 12017 => x"b8206000",
    12018 => x"3dad0002", 12019 => x"c84f0800", 12020 => x"b9a01000",
    12021 => x"b8607000", 12022 => x"f800150b", 12023 => x"b42f1000",
    12024 => x"b5af6800", 12025 => x"b44e0800", 12026 => x"542d0006",
    12027 => x"b9800800", 12028 => x"b9c01800", 12029 => x"f8001555",
    12030 => x"b8206000", 12031 => x"e0000009", 12032 => x"c9a26800",
    12033 => x"b9a01800", 12034 => x"b9800800", 12035 => x"f800154f",
    12036 => x"29620004", 12037 => x"b58d0800", 12038 => x"c9cd1800",
    12039 => x"f800154b", 12040 => x"b9800800", 12041 => x"2b9d0004",
    12042 => x"2b8b0018", 12043 => x"2b8c0014", 12044 => x"2b8d0010",
    12045 => x"2b8e000c", 12046 => x"2b8f0008", 12047 => x"379c0018",
    12048 => x"c3a00000", 12049 => x"379cffe8", 12050 => x"5b8b0018",
    12051 => x"5b8c0014", 12052 => x"5b8d0010", 12053 => x"5b8e000c",
    12054 => x"5b8f0008", 12055 => x"5b9d0004", 12056 => x"780b0001",
    12057 => x"396b5e08", 12058 => x"296f000c", 12059 => x"296e0004",
    12060 => x"b8406800", 12061 => x"3def0002", 12062 => x"c82e0800",
    12063 => x"b9e01000", 12064 => x"f80014e1", 12065 => x"b42e6000",
    12066 => x"b58d0800", 12067 => x"b5ee7000", 12068 => x"542e0006",
    12069 => x"b9800800", 12070 => x"34020000", 12071 => x"b9a01800",
    12072 => x"f80015a8", 12073 => x"e000000b", 12074 => x"c9cc7000",
    12075 => x"34020000", 12076 => x"b9c01800", 12077 => x"b9800800",
    12078 => x"f80015a2", 12079 => x"29610004", 12080 => x"34020000",
    12081 => x"c9ae1800", 12082 => x"f800159e", 12083 => x"b9800800",
    12084 => x"2b9d0004", 12085 => x"2b8b0018", 12086 => x"2b8c0014",
    12087 => x"2b8d0010", 12088 => x"2b8e000c", 12089 => x"2b8f0008",
    12090 => x"379c0018", 12091 => x"c3a00000", 12092 => x"379cfff4",
    12093 => x"5b8b000c", 12094 => x"5b8c0008", 12095 => x"5b9d0004",
    12096 => x"780c0001", 12097 => x"398c6dcc", 12098 => x"29810000",
    12099 => x"780b0001", 12100 => x"396b5e08", 12101 => x"58200000",
    12102 => x"34020200", 12103 => x"78010001", 12104 => x"38216230",
    12105 => x"5962000c", 12106 => x"34020800", 12107 => x"59610004",
    12108 => x"59610000", 12109 => x"fbffffc4", 12110 => x"29620004",
    12111 => x"29810000", 12112 => x"58220008", 12113 => x"2962000c",
    12114 => x"5822000c", 12115 => x"34020002", 12116 => x"5822004c",
    12117 => x"34020400", 12118 => x"58220000", 12119 => x"2b9d0004",
    12120 => x"2b8b000c", 12121 => x"2b8c0008", 12122 => x"379c000c",
    12123 => x"c3a00000", 12124 => x"379cfff4", 12125 => x"5b8b000c",
    12126 => x"5b8c0008", 12127 => x"5b9d0004", 12128 => x"780b0001",
    12129 => x"396b6dcc", 12130 => x"29630000", 12131 => x"340c0002",
    12132 => x"78010001", 12133 => x"586c0040", 12134 => x"78020001",
    12135 => x"586c004c", 12136 => x"38215e08", 12137 => x"38426230",
    12138 => x"58220004", 12139 => x"00420002", 12140 => x"34040800",
    12141 => x"5824000c", 12142 => x"344401ff", 12143 => x"3c840010",
    12144 => x"2042ffff", 12145 => x"b8821000", 12146 => x"58620020",
    12147 => x"78020001", 12148 => x"38425e30", 12149 => x"58220014",
    12150 => x"34020100", 12151 => x"5822001c", 12152 => x"58200020",
    12153 => x"58200024", 12154 => x"fbffffc2", 12155 => x"29610000",
    12156 => x"582c0044", 12157 => x"2b9d0004", 12158 => x"2b8b000c",
    12159 => x"2b8c0008", 12160 => x"379c000c", 12161 => x"c3a00000",
    12162 => x"379cffc4", 12163 => x"5b8b0028", 12164 => x"5b8c0024",
    12165 => x"5b8d0020", 12166 => x"5b8e001c", 12167 => x"5b8f0018",
    12168 => x"5b900014", 12169 => x"5b910010", 12170 => x"5b92000c",
    12171 => x"5b930008", 12172 => x"5b9d0004", 12173 => x"b8805800",
    12174 => x"78040001", 12175 => x"38846dcc", 12176 => x"28840000",
    12177 => x"b8209000", 12178 => x"b8408800", 12179 => x"2881004c",
    12180 => x"b8608000", 12181 => x"340c0000", 12182 => x"20210002",
    12183 => x"4420008a", 12184 => x"780e0001", 12185 => x"39ce5e08",
    12186 => x"29c20000", 12187 => x"28430000", 12188 => x"48030009",
    12189 => x"28810000", 12190 => x"20210200", 12191 => x"5c200004",
    12192 => x"78010001", 12193 => x"382135dc", 12194 => x"fbfffbcf",
    12195 => x"fbffff99", 12196 => x"e000007d", 12197 => x"20610001",
    12198 => x"206d0ffe", 12199 => x"c9a16800", 12200 => x"35af0003",
    12201 => x"01ef0002", 12202 => x"78044000", 12203 => x"a0642000",
    12204 => x"35ef0001", 12205 => x"340cffff", 12206 => x"5c800054",
    12207 => x"7d610000", 12208 => x"0063001d", 12209 => x"a0611800",
    12210 => x"4464003e", 12211 => x"b44d1000", 12212 => x"34030004",
    12213 => x"37810038", 12214 => x"fbffff30", 12215 => x"29c30000",
    12216 => x"35b3fffa", 12217 => x"35adfffe", 12218 => x"b46d1000",
    12219 => x"3781003e", 12220 => x"34030002", 12221 => x"fbffff29",
    12222 => x"78010001", 12223 => x"38213d2c", 12224 => x"282c0000",
    12225 => x"37820034", 12226 => x"3781002c", 12227 => x"2b8d0038",
    12228 => x"f8000191", 12229 => x"78020001", 12230 => x"38423d30",
    12231 => x"28410000", 12232 => x"a1ac6000", 12233 => x"01ad001c",
    12234 => x"502c000e", 12235 => x"78030001", 12236 => x"38633d34",
    12237 => x"2b820034", 12238 => x"28610000", 12239 => x"54410009",
    12240 => x"2b820030", 12241 => x"2b81002c", 12242 => x"3444ffff",
    12243 => x"f4441000", 12244 => x"3421ffff", 12245 => x"b4410800",
    12246 => x"5b81002c", 12247 => x"5b840030", 12248 => x"78020001",
    12249 => x"38423d38", 12250 => x"28410000", 12251 => x"2b820030",
    12252 => x"2183000f", 12253 => x"c86d1800", 12254 => x"a0410800",
    12255 => x"5961000c", 12256 => x"6461fff1", 12257 => x"64630001",
    12258 => x"59600008", 12259 => x"b8231800", 12260 => x"44600004",
    12261 => x"34010001", 12262 => x"59610004", 12263 => x"e0000002",
    12264 => x"59600004", 12265 => x"2f81003e", 12266 => x"3d8c0003",
    12267 => x"ba606800", 12268 => x"20210800", 12269 => x"64210000",
    12270 => x"596c0010", 12271 => x"31610000", 12272 => x"b9a06000",
    12273 => x"520d0002", 12274 => x"ba006000", 12275 => x"780b0001",
    12276 => x"396b5e08", 12277 => x"29610024", 12278 => x"29620000",
    12279 => x"3403000e", 12280 => x"34210001", 12281 => x"59610024",
    12282 => x"34420004", 12283 => x"ba400800", 12284 => x"fbfffeea",
    12285 => x"29630000", 12286 => x"ba200800", 12287 => x"34620012",
    12288 => x"3583fff2", 12289 => x"fbfffee5", 12290 => x"780b0001",
    12291 => x"396b5e08", 12292 => x"3dee0002", 12293 => x"29610000",
    12294 => x"b9c01000", 12295 => x"fbffff0a", 12296 => x"78030001",
    12297 => x"38636dcc", 12298 => x"286d0000", 12299 => x"29610000",
    12300 => x"59af0010", 12301 => x"2962000c", 12302 => x"296f0004",
    12303 => x"3c420002", 12304 => x"c82f0800", 12305 => x"b42e0800",
    12306 => x"f80013ef", 12307 => x"b42f0800", 12308 => x"59610000",
    12309 => x"29a20010", 12310 => x"28210000", 12311 => x"4801000a",
    12312 => x"29a10000", 12313 => x"20210200", 12314 => x"44200002",
    12315 => x"fbffff21", 12316 => x"78010001", 12317 => x"38216dcc",
    12318 => x"28210000", 12319 => x"34020002", 12320 => x"5822004c",
    12321 => x"b9800800", 12322 => x"2b9d0004", 12323 => x"2b8b0028",
    12324 => x"2b8c0024", 12325 => x"2b8d0020", 12326 => x"2b8e001c",
    12327 => x"2b8f0018", 12328 => x"2b900014", 12329 => x"2b910010",
    12330 => x"2b92000c", 12331 => x"2b930008", 12332 => x"379c003c",
    12333 => x"c3a00000", 12334 => x"379cffd8", 12335 => x"5b8b001c",
    12336 => x"5b8c0018", 12337 => x"5b8d0014", 12338 => x"5b8e0010",
    12339 => x"5b8f000c", 12340 => x"5b900008", 12341 => x"5b9d0004",
    12342 => x"780d0001", 12343 => x"39ad5e08", 12344 => x"b8605800",
    12345 => x"34030100", 12346 => x"59a3001c", 12347 => x"59a30018",
    12348 => x"78030001", 12349 => x"38636dcc", 12350 => x"b8207800",
    12351 => x"b8407000", 12352 => x"78010001", 12353 => x"28620000",
    12354 => x"38215e30", 12355 => x"59a10014", 12356 => x"59a10010",
    12357 => x"58410004", 12358 => x"35630010", 12359 => x"34020000",
    12360 => x"b8806000", 12361 => x"f8001487", 12362 => x"29a10010",
    12363 => x"3402003c", 12364 => x"b9601800", 12365 => x"34210004",
    12366 => x"51620002", 12367 => x"3403003c", 12368 => x"34020000",
    12369 => x"780d0001", 12370 => x"f800147e", 12371 => x"39ad5e08",
    12372 => x"29a10010", 12373 => x"b9e01000", 12374 => x"3403000e",
    12375 => x"34210004", 12376 => x"f80013fa", 12377 => x"29a10010",
    12378 => x"b9c01000", 12379 => x"3563fff2", 12380 => x"34210012",
    12381 => x"f80013f5", 12382 => x"3401003b", 12383 => x"502b0002",
    12384 => x"e0000002", 12385 => x"340b003c", 12386 => x"35630001",
    12387 => x"7d810000", 12388 => x"00630001", 12389 => x"3c21001e",
    12390 => x"78048000", 12391 => x"b8642000", 12392 => x"b8812000",
    12393 => x"78010001", 12394 => x"38215e08", 12395 => x"28220010",
    12396 => x"3c630002", 12397 => x"78010001", 12398 => x"58440000",
    12399 => x"38216dcc", 12400 => x"b4431000", 12401 => x"58400000",
    12402 => x"28220000", 12403 => x"340d0000", 12404 => x"b8207800",
    12405 => x"28430000", 12406 => x"341003e8", 12407 => x"38630001",
    12408 => x"58430000", 12409 => x"29e10000", 12410 => x"282e0000",
    12411 => x"21c10002", 12412 => x"5c200009", 12413 => x"34010001",
    12414 => x"35ad0001", 12415 => x"f8000129", 12416 => x"5db0fff9",
    12417 => x"78010001", 12418 => x"382135fc", 12419 => x"b9c01000",
    12420 => x"fbfffaed", 12421 => x"45800046", 12422 => x"780d0001",
    12423 => x"340e0000", 12424 => x"39ad6dcc", 12425 => x"340f0064",
    12426 => x"29a10000", 12427 => x"28220000", 12428 => x"20420800",
    12429 => x"5c40000a", 12430 => x"34010001", 12431 => x"35ce0001",
    12432 => x"f8000118", 12433 => x"5dcffff9", 12434 => x"78010001",
    12435 => x"3821362c", 12436 => x"fbfffadd", 12437 => x"340e0000",
    12438 => x"e0000003", 12439 => x"282e0014", 12440 => x"21ce0001",
    12441 => x"78010001", 12442 => x"38216dcc", 12443 => x"28210000",
    12444 => x"282d0018", 12445 => x"28230014", 12446 => x"00630006",
    12447 => x"2063ffff", 12448 => x"44600006", 12449 => x"78020001",
    12450 => x"34010000", 12451 => x"3842365c", 12452 => x"34040000",
    12453 => x"fbffcfe0", 12454 => x"78020001", 12455 => x"38423d2c",
    12456 => x"28410000", 12457 => x"37820028", 12458 => x"a1a16800",
    12459 => x"37810020", 12460 => x"f80000a9", 12461 => x"78030001",
    12462 => x"38633d30", 12463 => x"28610000", 12464 => x"502d000e",
    12465 => x"78030001", 12466 => x"38633d34", 12467 => x"2b820028",
    12468 => x"28610000", 12469 => x"54410009", 12470 => x"2b830024",
    12471 => x"2b820020", 12472 => x"3461ffff", 12473 => x"f4611800",
    12474 => x"3442ffff", 12475 => x"b4621000", 12476 => x"5b820020",
    12477 => x"5b810024", 12478 => x"2b810020", 12479 => x"318e0000",
    12480 => x"3dad0003", 12481 => x"59810008", 12482 => x"2b810024",
    12483 => x"59800004", 12484 => x"598d0010", 12485 => x"5981000c",
    12486 => x"78010001", 12487 => x"38215e08", 12488 => x"28220020",
    12489 => x"34420001", 12490 => x"58220020", 12491 => x"b9600800",
    12492 => x"2b9d0004", 12493 => x"2b8b001c", 12494 => x"2b8c0018",
    12495 => x"2b8d0014", 12496 => x"2b8e0010", 12497 => x"2b8f000c",
    12498 => x"2b900008", 12499 => x"379c0028", 12500 => x"c3a00000",
    12501 => x"78030001", 12502 => x"38635e08", 12503 => x"28640020",
    12504 => x"58240000", 12505 => x"28610024", 12506 => x"58410000",
    12507 => x"c3a00000", 12508 => x"78010001", 12509 => x"38216d10",
    12510 => x"28210000", 12511 => x"28220008", 12512 => x"2821000c",
    12513 => x"202100ff", 12514 => x"c3a00000", 12515 => x"78010001",
    12516 => x"78030001", 12517 => x"38633d3c", 12518 => x"38216d10",
    12519 => x"28210000", 12520 => x"28620000", 12521 => x"78040001",
    12522 => x"38843d40", 12523 => x"58220000", 12524 => x"58200014",
    12525 => x"28830000", 12526 => x"58200018", 12527 => x"58200010",
    12528 => x"58230000", 12529 => x"58220000", 12530 => x"5820001c",
    12531 => x"c3a00000", 12532 => x"379cffe8", 12533 => x"5b8b0018",
    12534 => x"5b8c0014", 12535 => x"5b8d0010", 12536 => x"5b8e000c",
    12537 => x"5b8f0008", 12538 => x"5b9d0004", 12539 => x"780b0001",
    12540 => x"b8207800", 12541 => x"34010001", 12542 => x"b8406800",
    12543 => x"b8607000", 12544 => x"396b3684", 12545 => x"5de10003",
    12546 => x"780b0001", 12547 => x"396b3688", 12548 => x"15ac001f",
    12549 => x"b9c00800", 12550 => x"f8001327", 12551 => x"218c0002",
    12552 => x"358c002b", 12553 => x"78020001", 12554 => x"b8202800",
    12555 => x"38423690", 12556 => x"34010000", 12557 => x"b9601800",
    12558 => x"b9802000", 12559 => x"fbffcf76", 12560 => x"78020001",
    12561 => x"34010002", 12562 => x"38426d10", 12563 => x"5de1000e",
    12564 => x"28410000", 12565 => x"15a2001f", 12566 => x"20420007",
    12567 => x"b44e7000", 12568 => x"f44e1000", 12569 => x"01ce0003",
    12570 => x"b44d6800", 12571 => x"3dad001d", 12572 => x"58200014",
    12573 => x"58200018", 12574 => x"b9ae7000", 12575 => x"582e0010",
    12576 => x"e0000006", 12577 => x"28420000", 12578 => x"21ad00ff",
    12579 => x"584e0014", 12580 => x"584d0018", 12581 => x"58400010",
    12582 => x"78010001", 12583 => x"38216d10", 12584 => x"28210000",
    12585 => x"28220000", 12586 => x"38420004", 12587 => x"58220000",
    12588 => x"34010000", 12589 => x"2b9d0004", 12590 => x"2b8b0018",
    12591 => x"2b8c0014", 12592 => x"2b8d0010", 12593 => x"2b8e000c",
    12594 => x"2b8f0008", 12595 => x"379c0018", 12596 => x"c3a00000",
    12597 => x"78050001", 12598 => x"38a56d10", 12599 => x"28a50000",
    12600 => x"202100ff", 12601 => x"00630003", 12602 => x"58a20014",
    12603 => x"58a10018", 12604 => x"58a30010", 12605 => x"34010003",
    12606 => x"5c810007", 12607 => x"28a20000", 12608 => x"3401fff3",
    12609 => x"a0410800", 12610 => x"38210008", 12611 => x"58a10000",
    12612 => x"c3a00000", 12613 => x"34010001", 12614 => x"5c810007",
    12615 => x"28a2001c", 12616 => x"3401ffe7", 12617 => x"a0410800",
    12618 => x"38210008", 12619 => x"58a1001c", 12620 => x"c3a00000",
    12621 => x"34010002", 12622 => x"5c810006", 12623 => x"28a2001c",
    12624 => x"3401ffe7", 12625 => x"a0410800", 12626 => x"38210010",
    12627 => x"58a1001c", 12628 => x"c3a00000", 12629 => x"379cffe0",
    12630 => x"5b8b0020", 12631 => x"5b8c001c", 12632 => x"5b8d0018",
    12633 => x"5b8e0014", 12634 => x"5b8f0010", 12635 => x"5b90000c",
    12636 => x"5b910008", 12637 => x"5b9d0004", 12638 => x"b8206000",
    12639 => x"78010001", 12640 => x"38213d2c", 12641 => x"282f0000",
    12642 => x"780b0001", 12643 => x"b8406800", 12644 => x"396b6d10",
    12645 => x"fbffff77", 12646 => x"b8208800", 12647 => x"29610000",
    12648 => x"b8408000", 12649 => x"282e0004", 12650 => x"a1cf7000",
    12651 => x"fbffff71", 12652 => x"5c31fff9", 12653 => x"5c50fff8",
    12654 => x"45800003", 12655 => x"59810000", 12656 => x"59820004",
    12657 => x"45a00003", 12658 => x"3dc10003", 12659 => x"59a10000",
    12660 => x"2b9d0004", 12661 => x"2b8b0020", 12662 => x"2b8c001c",
    12663 => x"2b8d0018", 12664 => x"2b8e0014", 12665 => x"2b8f0010",
    12666 => x"2b90000c", 12667 => x"2b910008", 12668 => x"379c0020",
    12669 => x"c3a00000", 12670 => x"78010001", 12671 => x"38216d10",
    12672 => x"28210000", 12673 => x"28210000", 12674 => x"20210004",
    12675 => x"64210000", 12676 => x"c3a00000", 12677 => x"78020001",
    12678 => x"38426d10", 12679 => x"28420000", 12680 => x"2843001c",
    12681 => x"44200003", 12682 => x"38630006", 12683 => x"e0000003",
    12684 => x"3401fff9", 12685 => x"a0611800", 12686 => x"5843001c",
    12687 => x"34010000", 12688 => x"c3a00000", 12689 => x"78020001",
    12690 => x"38426dd0", 12691 => x"28420000", 12692 => x"78030001",
    12693 => x"38636db8", 12694 => x"58620000", 12695 => x"44200005",
    12696 => x"28430010", 12697 => x"78018000", 12698 => x"b8610800",
    12699 => x"e0000006", 12700 => x"78040001", 12701 => x"38843d38",
    12702 => x"28430010", 12703 => x"28810000", 12704 => x"a0610800",
    12705 => x"58410010", 12706 => x"c3a00000", 12707 => x"78010001",
    12708 => x"38216db8", 12709 => x"28210000", 12710 => x"28210014",
    12711 => x"c3a00000", 12712 => x"78020001", 12713 => x"38426db8",
    12714 => x"28420000", 12715 => x"28430014", 12716 => x"b4230800",
    12717 => x"28430014", 12718 => x"c8611800", 12719 => x"4803fffe",
    12720 => x"c3a00000", 12721 => x"78010001", 12722 => x"38216db8",
    12723 => x"28210000", 12724 => x"28210004", 12725 => x"20210080",
    12726 => x"64210000", 12727 => x"c3a00000", 12728 => x"379cffe0",
    12729 => x"5b8b001c", 12730 => x"5b8c0018", 12731 => x"5b8d0014",
    12732 => x"5b8e0010", 12733 => x"5b8f000c", 12734 => x"5b900008",
    12735 => x"5b9d0004", 12736 => x"b8208000", 12737 => x"34010001",
    12738 => x"fbfffcfb", 12739 => x"34010001", 12740 => x"fbfffc2a",
    12741 => x"340200a0", 12742 => x"34010001", 12743 => x"fbfffc6f",
    12744 => x"34020000", 12745 => x"34010001", 12746 => x"fbfffc6c",
    12747 => x"34010001", 12748 => x"fbfffc36", 12749 => x"340200a1",
    12750 => x"34010001", 12751 => x"fbfffc67", 12752 => x"378d0023",
    12753 => x"b9a01000", 12754 => x"34030001", 12755 => x"34010001",
    12756 => x"fbfffc9f", 12757 => x"34010001", 12758 => x"fbfffc48",
    12759 => x"34010001", 12760 => x"438c0023", 12761 => x"fbfffc15",
    12762 => x"34010001", 12763 => x"340200a1", 12764 => x"fbfffc5a",
    12765 => x"340bffd9", 12766 => x"340f000f", 12767 => x"340e0017",
    12768 => x"34030000", 12769 => x"34010001", 12770 => x"b9a01000",
    12771 => x"fbfffc90", 12772 => x"43830023", 12773 => x"b5836000",
    12774 => x"218c00ff", 12775 => x"556f0003", 12776 => x"b60b0800",
    12777 => x"30230000", 12778 => x"356b0001", 12779 => x"5d6efff5",
    12780 => x"37820023", 12781 => x"34030001", 12782 => x"34010001",
    12783 => x"fbfffc84", 12784 => x"34010001", 12785 => x"fbfffc2d",
    12786 => x"43810023", 12787 => x"fc2c6000", 12788 => x"c80c0800",
    12789 => x"2b9d0004", 12790 => x"2b8b001c", 12791 => x"2b8c0018",
    12792 => x"2b8d0014", 12793 => x"2b8e0010", 12794 => x"2b8f000c",
    12795 => x"2b900008", 12796 => x"379c0020", 12797 => x"c3a00000",
    12798 => x"379cffe0", 12799 => x"5b9b0008", 12800 => x"341b0020",
    12801 => x"b77cd800", 12802 => x"5b8b0020", 12803 => x"5b8c001c",
    12804 => x"5b8d0018", 12805 => x"5b8e0014", 12806 => x"5b8f0010",
    12807 => x"5b90000c", 12808 => x"5b9d0004", 12809 => x"780b0001",
    12810 => x"780c0001", 12811 => x"bb807800", 12812 => x"34020001",
    12813 => x"396b4c88", 12814 => x"398c36b0", 12815 => x"e0000012",
    12816 => x"bb808000", 12817 => x"379cffe4", 12818 => x"378e000b",
    12819 => x"01ce0003", 12820 => x"35a2002c", 12821 => x"3dce0003",
    12822 => x"34030014", 12823 => x"b9c00800", 12824 => x"f800123a",
    12825 => x"31c00013", 12826 => x"29a20020", 12827 => x"29630074",
    12828 => x"b9800800", 12829 => x"b9c02000", 12830 => x"fbfff953",
    12831 => x"34020000", 12832 => x"ba00e000", 12833 => x"b9600800",
    12834 => x"f8001099", 12835 => x"b8206800", 12836 => x"5c20ffec",
    12837 => x"b9e0e000", 12838 => x"2b9d0004", 12839 => x"2b8b0020",
    12840 => x"2b8c001c", 12841 => x"2b8d0018", 12842 => x"2b8e0014",
    12843 => x"2b8f0010", 12844 => x"2b90000c", 12845 => x"2b9b0008",
    12846 => x"379c0020", 12847 => x"c3a00000", 12848 => x"379cffec",
    12849 => x"5b8b0014", 12850 => x"5b8c0010", 12851 => x"5b8d000c",
    12852 => x"5b8e0008", 12853 => x"5b9d0004", 12854 => x"780b0001",
    12855 => x"396b6a30", 12856 => x"29610000", 12857 => x"5c200007",
    12858 => x"78010001", 12859 => x"38214c88", 12860 => x"f800105d",
    12861 => x"29610000", 12862 => x"34210001", 12863 => x"59610000",
    12864 => x"780b0001", 12865 => x"396b4bb0", 12866 => x"780c0001",
    12867 => x"356d00d8", 12868 => x"398c4c88", 12869 => x"e0000009",
    12870 => x"29620008", 12871 => x"2963000c", 12872 => x"29640010",
    12873 => x"296e0000", 12874 => x"b9800800", 12875 => x"f8001122",
    12876 => x"59c10000", 12877 => x"356b0018", 12878 => x"5d6dfff8",
    12879 => x"2b9d0004", 12880 => x"2b8b0014", 12881 => x"2b8c0010",
    12882 => x"2b8d000c", 12883 => x"2b8e0008", 12884 => x"379c0014",
    12885 => x"c3a00000", 12886 => x"379cfff4", 12887 => x"5b8b000c",
    12888 => x"5b8c0008", 12889 => x"5b9d0004", 12890 => x"34020000",
    12891 => x"b8206000", 12892 => x"f80002d3", 12893 => x"b8205800",
    12894 => x"4c200005", 12895 => x"78010001", 12896 => x"382136d8",
    12897 => x"b9601000", 12898 => x"e0000004", 12899 => x"29820000",
    12900 => x"78010001", 12901 => x"38213704", 12902 => x"fbfff90b",
    12903 => x"b9600800", 12904 => x"2b9d0004", 12905 => x"2b8b000c",
    12906 => x"2b8c0008", 12907 => x"379c000c", 12908 => x"c3a00000",
    12909 => x"379cfffc", 12910 => x"5b9d0004", 12911 => x"78010001",
    12912 => x"38216a34", 12913 => x"58200000", 12914 => x"78020001",
    12915 => x"78010001", 12916 => x"38216a48", 12917 => x"38426a38",
    12918 => x"3403ffff", 12919 => x"58230000", 12920 => x"58430000",
    12921 => x"58200008", 12922 => x"58400008", 12923 => x"58400004",
    12924 => x"58200004", 12925 => x"5840000c", 12926 => x"5820000c",
    12927 => x"34020000", 12928 => x"34010000", 12929 => x"f8000dd8",
    12930 => x"2b9d0004", 12931 => x"379c0004", 12932 => x"c3a00000",
    12933 => x"379cfff4", 12934 => x"5b8b000c", 12935 => x"5b8c0008",
    12936 => x"5b9d0004", 12937 => x"b8206000", 12938 => x"34010000",
    12939 => x"f8000e78", 12940 => x"b8205800", 12941 => x"34020000",
    12942 => x"5c20008b", 12943 => x"fbfffa8d", 12944 => x"78030001",
    12945 => x"38636a38", 12946 => x"28650008", 12947 => x"78020001",
    12948 => x"38426a34", 12949 => x"b8202000", 12950 => x"28420000",
    12951 => x"44ab0004", 12952 => x"34010001", 12953 => x"5ca1001d",
    12954 => x"e0000010", 12955 => x"34010001", 12956 => x"44810005",
    12957 => x"28610004", 12958 => x"34210001", 12959 => x"58610004",
    12960 => x"e0000002", 12961 => x"58600004", 12962 => x"78030001",
    12963 => x"38636a38", 12964 => x"28650004", 12965 => x"34010004",
    12966 => x"4c250010", 12967 => x"34010001", 12968 => x"58610008",
    12969 => x"e0000002", 12970 => x"44850003", 12971 => x"58600004",
    12972 => x"e000000a", 12973 => x"28650004", 12974 => x"34010004",
    12975 => x"34a50001", 12976 => x"58650004", 12977 => x"4c250005",
    12978 => x"34010002", 12979 => x"58610008", 12980 => x"3441fe0c",
    12981 => x"5861000c", 12982 => x"78030001", 12983 => x"38636a48",
    12984 => x"28650008", 12985 => x"44a00004", 12986 => x"34010001",
    12987 => x"5ca1001c", 12988 => x"e000000f", 12989 => x"44850005",
    12990 => x"28610004", 12991 => x"34210001", 12992 => x"58610004",
    12993 => x"e0000002", 12994 => x"58600004", 12995 => x"78030001",
    12996 => x"38636a48", 12997 => x"28640004", 12998 => x"34010004",
    12999 => x"4c240010", 13000 => x"34010001", 13001 => x"58610008",
    13002 => x"e0000002", 13003 => x"44800003", 13004 => x"58600004",
    13005 => x"e000000a", 13006 => x"28640004", 13007 => x"34010004",
    13008 => x"34840001", 13009 => x"58640004", 13010 => x"4c240005",
    13011 => x"34010002", 13012 => x"58610008", 13013 => x"3441fe0c",
    13014 => x"5861000c", 13015 => x"3401251b", 13016 => x"4c22003a",
    13017 => x"78020001", 13018 => x"38426a38", 13019 => x"28430008",
    13020 => x"34010002", 13021 => x"5c610008", 13022 => x"78020001",
    13023 => x"38426a48", 13024 => x"28410008", 13025 => x"5c230004",
    13026 => x"2844000c", 13027 => x"34011f3f", 13028 => x"e0000008",
    13029 => x"78020001", 13030 => x"38423724", 13031 => x"34010000",
    13032 => x"fbffcd9d", 13033 => x"3402ffff", 13034 => x"e000002f",
    13035 => x"3484e0c0", 13036 => x"4881ffff", 13037 => x"78020001",
    13038 => x"38426a48", 13039 => x"5844000c", 13040 => x"78020001",
    13041 => x"38426a38", 13042 => x"2843000c", 13043 => x"34011f3f",
    13044 => x"e0000002", 13045 => x"3463e0c0", 13046 => x"4861ffff",
    13047 => x"78020001", 13048 => x"38426a38", 13049 => x"5843000c",
    13050 => x"4c640003", 13051 => x"348bf060", 13052 => x"e0000004",
    13053 => x"340b0000", 13054 => x"4c830002", 13055 => x"348b0fa0",
    13056 => x"b5635800", 13057 => x"0161001f", 13058 => x"b42b5800",
    13059 => x"156b0001", 13060 => x"4d600003", 13061 => x"356b1f40",
    13062 => x"e0000004", 13063 => x"34011f3f", 13064 => x"4c2b0002",
    13065 => x"356be0c0", 13066 => x"78020001", 13067 => x"38423740",
    13068 => x"34010000", 13069 => x"b9602800", 13070 => x"fbffcd77",
    13071 => x"34020001", 13072 => x"598b0000", 13073 => x"e0000008",
    13074 => x"78010001", 13075 => x"34420064", 13076 => x"38216a34",
    13077 => x"58220000", 13078 => x"34010000", 13079 => x"f8000d42",
    13080 => x"34020000", 13081 => x"b8400800", 13082 => x"2b9d0004",
    13083 => x"2b8b000c", 13084 => x"2b8c0008", 13085 => x"379c000c",
    13086 => x"c3a00000", 13087 => x"379cfff8", 13088 => x"5b8b0008",
    13089 => x"5b9d0004", 13090 => x"78020001", 13091 => x"b8205800",
    13092 => x"b8400800", 13093 => x"38213774", 13094 => x"fbfff84b",
    13095 => x"e0000003", 13096 => x"34010064", 13097 => x"fbfffe7f",
    13098 => x"34010000", 13099 => x"fbfff999", 13100 => x"4420fffc",
    13101 => x"34010003", 13102 => x"34020000", 13103 => x"34030001",
    13104 => x"f8000c33", 13105 => x"78020001", 13106 => x"b8400800",
    13107 => x"3821378c", 13108 => x"fbfff83d", 13109 => x"e0000003",
    13110 => x"34010064", 13111 => x"fbfffe71", 13112 => x"34010000",
    13113 => x"f8000d0f", 13114 => x"4420fffc", 13115 => x"78020001",
    13116 => x"b8400800", 13117 => x"38211b1c", 13118 => x"fbfff833",
    13119 => x"78020001", 13120 => x"b8400800", 13121 => x"3821379c",
    13122 => x"fbfff82f", 13123 => x"fbffff2a", 13124 => x"b9600800",
    13125 => x"fbffff40", 13126 => x"4420fffe", 13127 => x"2b9d0004",
    13128 => x"2b8b0008", 13129 => x"379c0008", 13130 => x"c3a00000",
    13131 => x"379cfff0", 13132 => x"5b8b000c", 13133 => x"5b8c0008",
    13134 => x"5b9d0004", 13135 => x"b8405800", 13136 => x"34020003",
    13137 => x"5c220020", 13138 => x"fbffff1b", 13139 => x"b9600800",
    13140 => x"fbffff31", 13141 => x"4420fffe", 13142 => x"4c200002",
    13143 => x"e000001a", 13144 => x"37810010", 13145 => x"34020000",
    13146 => x"f80001d5", 13147 => x"b8206000", 13148 => x"48010007",
    13149 => x"29620000", 13150 => x"2b810010", 13151 => x"3443ff38",
    13152 => x"54610003", 13153 => x"344200c8", 13154 => x"50410012",
    13155 => x"34020001", 13156 => x"b9600800", 13157 => x"f80001ca",
    13158 => x"78030001", 13159 => x"b8206000", 13160 => x"29620000",
    13161 => x"386337c4", 13162 => x"4c200003", 13163 => x"78030001",
    13164 => x"386337bc", 13165 => x"78010001", 13166 => x"382137cc",
    13167 => x"fbfff802", 13168 => x"e0000004", 13169 => x"b9600800",
    13170 => x"fbfffee4", 13171 => x"b8206000", 13172 => x"29610000",
    13173 => x"fbfff39c", 13174 => x"b9800800", 13175 => x"2b9d0004",
    13176 => x"2b8b000c", 13177 => x"2b8c0008", 13178 => x"379c0010",
    13179 => x"c3a00000", 13180 => x"379cfffc", 13181 => x"5b9d0004",
    13182 => x"34010800", 13183 => x"34020001", 13184 => x"fbfffa60",
    13185 => x"34010400", 13186 => x"34020000", 13187 => x"fbfffa5d",
    13188 => x"34011000", 13189 => x"34020000", 13190 => x"fbfffa5a",
    13191 => x"2b9d0004", 13192 => x"379c0004", 13193 => x"c3a00000",
    13194 => x"40230000", 13195 => x"78020001", 13196 => x"40240001",
    13197 => x"38426dc0", 13198 => x"28420000", 13199 => x"3c630008",
    13200 => x"b8831800", 13201 => x"58430010", 13202 => x"40240002",
    13203 => x"40230003", 13204 => x"3c840018", 13205 => x"3c630010",
    13206 => x"b8832000", 13207 => x"40230005", 13208 => x"b8832000",
    13209 => x"40230004", 13210 => x"3c630008", 13211 => x"b8830800",
    13212 => x"58410014", 13213 => x"c3a00000", 13214 => x"40230000",
    13215 => x"40240003", 13216 => x"78020001", 13217 => x"3c630018",
    13218 => x"38426dc0", 13219 => x"b8831800", 13220 => x"40240001",
    13221 => x"40210002", 13222 => x"28420000", 13223 => x"3c840010",
    13224 => x"3c210008", 13225 => x"b8641800", 13226 => x"b8611800",
    13227 => x"3401ff00", 13228 => x"58430018", 13229 => x"a0611800",
    13230 => x"34630001", 13231 => x"58410020", 13232 => x"3801ea60",
    13233 => x"5843001c", 13234 => x"58410024", 13235 => x"78030001",
    13236 => x"34210001", 13237 => x"38633d44", 13238 => x"58410028",
    13239 => x"34210001", 13240 => x"5841002c", 13241 => x"28610000",
    13242 => x"78030001", 13243 => x"38633d48", 13244 => x"58410030",
    13245 => x"38018cae", 13246 => x"58410034", 13247 => x"28610000",
    13248 => x"58410038", 13249 => x"34011f40", 13250 => x"5841003c",
    13251 => x"c3a00000", 13252 => x"379cffe0", 13253 => x"5b8b001c",
    13254 => x"5b8c0018", 13255 => x"5b8d0014", 13256 => x"5b8e0010",
    13257 => x"5b8f000c", 13258 => x"5b900008", 13259 => x"5b9d0004",
    13260 => x"b8205800", 13261 => x"78010001", 13262 => x"38216a58",
    13263 => x"b8406000", 13264 => x"40220000", 13265 => x"b8607000",
    13266 => x"b8807800", 13267 => x"b8a06800", 13268 => x"3401ffff",
    13269 => x"4440002b", 13270 => x"3d8c0001", 13271 => x"b9600800",
    13272 => x"fbfffa16", 13273 => x"218200fe", 13274 => x"b9600800",
    13275 => x"fbfffa5b", 13276 => x"01c20008", 13277 => x"b9600800",
    13278 => x"204200ff", 13279 => x"fbfffa57", 13280 => x"21c200ff",
    13281 => x"b9600800", 13282 => x"fbfffa54", 13283 => x"b9600800",
    13284 => x"fbfffa1e", 13285 => x"39820001", 13286 => x"b9600800",
    13287 => x"204200ff", 13288 => x"fbfffa4e", 13289 => x"340c0000",
    13290 => x"35aeffff", 13291 => x"37900023", 13292 => x"e0000009",
    13293 => x"b9600800", 13294 => x"ba001000", 13295 => x"34030000",
    13296 => x"fbfffa83", 13297 => x"43820023", 13298 => x"b5ec0800",
    13299 => x"358c0001", 13300 => x"30220000", 13301 => x"55ccfff8",
    13302 => x"b9600800", 13303 => x"ba001000", 13304 => x"34030001",
    13305 => x"fbfffa7a", 13306 => x"43810023", 13307 => x"b5ee7000",
    13308 => x"31c10000", 13309 => x"b9600800", 13310 => x"fbfffa20",
    13311 => x"b9a00800", 13312 => x"2b9d0004", 13313 => x"2b8b001c",
    13314 => x"2b8c0018", 13315 => x"2b8d0014", 13316 => x"2b8e0010",
    13317 => x"2b8f000c", 13318 => x"2b900008", 13319 => x"379c0020",
    13320 => x"c3a00000", 13321 => x"379cffe0", 13322 => x"5b8b0020",
    13323 => x"5b8c001c", 13324 => x"5b8d0018", 13325 => x"5b8e0014",
    13326 => x"5b8f0010", 13327 => x"5b90000c", 13328 => x"5b910008",
    13329 => x"5b9d0004", 13330 => x"b8205800", 13331 => x"78010001",
    13332 => x"38216a58", 13333 => x"b8606800", 13334 => x"40230000",
    13335 => x"3c4f0001", 13336 => x"b8808000", 13337 => x"b8a07000",
    13338 => x"3401ffff", 13339 => x"21ef00ff", 13340 => x"340c0000",
    13341 => x"5c60001f", 13342 => x"e0000020", 13343 => x"b9600800",
    13344 => x"fbfff9ce", 13345 => x"b9e01000", 13346 => x"b9600800",
    13347 => x"fbfffa13", 13348 => x"01a20008", 13349 => x"b9600800",
    13350 => x"204200ff", 13351 => x"fbfffa0f", 13352 => x"21a200ff",
    13353 => x"b9600800", 13354 => x"fbfffa0c", 13355 => x"b60c1000",
    13356 => x"40420000", 13357 => x"b9600800", 13358 => x"35ad0001",
    13359 => x"fbfffa07", 13360 => x"b9600800", 13361 => x"fbfff9ed",
    13362 => x"b9600800", 13363 => x"fbfff9bb", 13364 => x"b9600800",
    13365 => x"b9e01000", 13366 => x"fbfffa00", 13367 => x"b8208800",
    13368 => x"b9600800", 13369 => x"fbfff9e5", 13370 => x"5e20fff8",
    13371 => x"358c0001", 13372 => x"55ccffe3", 13373 => x"b9c00800",
    13374 => x"2b9d0004", 13375 => x"2b8b0020", 13376 => x"2b8c001c",
    13377 => x"2b8d0018", 13378 => x"2b8e0014", 13379 => x"2b8f0010",
    13380 => x"2b90000c", 13381 => x"2b910008", 13382 => x"379c0020",
    13383 => x"c3a00000", 13384 => x"379cffec", 13385 => x"5b8b0014",
    13386 => x"5b8c0010", 13387 => x"5b8d000c", 13388 => x"5b8e0008",
    13389 => x"5b9d0004", 13390 => x"780d0001", 13391 => x"780c0001",
    13392 => x"39ad6a5c", 13393 => x"398c6a60", 13394 => x"780b0001",
    13395 => x"59a10000", 13396 => x"59820000", 13397 => x"34030001",
    13398 => x"396b6a58", 13399 => x"202100ff", 13400 => x"204200ff",
    13401 => x"31630000", 13402 => x"fbfffa77", 13403 => x"b8207000",
    13404 => x"5c200006", 13405 => x"41a10003", 13406 => x"41820003",
    13407 => x"fbfffa72", 13408 => x"5c2e0002", 13409 => x"31600000",
    13410 => x"2b9d0004", 13411 => x"2b8b0014", 13412 => x"2b8c0010",
    13413 => x"2b8d000c", 13414 => x"2b8e0008", 13415 => x"379c0014",
    13416 => x"c3a00000", 13417 => x"379cfff8", 13418 => x"5b9d0004",
    13419 => x"78010001", 13420 => x"78020001", 13421 => x"38216a5c",
    13422 => x"38426a60", 13423 => x"40420003", 13424 => x"40210003",
    13425 => x"34031004", 13426 => x"3784000b", 13427 => x"34050001",
    13428 => x"3380000b", 13429 => x"fbffff94", 13430 => x"34030001",
    13431 => x"3402ffff", 13432 => x"5c230002", 13433 => x"4382000b",
    13434 => x"b8400800", 13435 => x"2b9d0004", 13436 => x"379c0008",
    13437 => x"c3a00000", 13438 => x"379cffec", 13439 => x"5b8b0014",
    13440 => x"5b8c0010", 13441 => x"5b8d000c", 13442 => x"5b8e0008",
    13443 => x"5b9d0004", 13444 => x"b8205800", 13445 => x"206d00ff",
    13446 => x"34010003", 13447 => x"204c00ff", 13448 => x"3405fffc",
    13449 => x"55a1005d", 13450 => x"5da0000f", 13451 => x"78010001",
    13452 => x"78020001", 13453 => x"38216a5c", 13454 => x"38426a60",
    13455 => x"40420003", 13456 => x"40210003", 13457 => x"78040001",
    13458 => x"34050001", 13459 => x"34031004", 13460 => x"38846a68",
    13461 => x"fbffff2f", 13462 => x"34020001", 13463 => x"3405ffff",
    13464 => x"5c22004e", 13465 => x"45800007", 13466 => x"78010001",
    13467 => x"38216a68", 13468 => x"40220000", 13469 => x"34010004",
    13470 => x"3405fffe", 13471 => x"44410047", 13472 => x"b9ac0800",
    13473 => x"5c200007", 13474 => x"78010001", 13475 => x"38216a68",
    13476 => x"40210000", 13477 => x"34050000", 13478 => x"5c250006",
    13479 => x"e000003f", 13480 => x"3562001c", 13481 => x"b9600800",
    13482 => x"34030000", 13483 => x"5d80001b", 13484 => x"78010001",
    13485 => x"78020001", 13486 => x"38216a5c", 13487 => x"38426a60",
    13488 => x"09a3001d", 13489 => x"40420003", 13490 => x"40210003",
    13491 => x"3405001d", 13492 => x"34631005", 13493 => x"b9602000",
    13494 => x"fbffff0e", 13495 => x"3402001d", 13496 => x"b9606000",
    13497 => x"3405ffff", 13498 => x"5c22002c", 13499 => x"3562001c",
    13500 => x"34010000", 13501 => x"41830000", 13502 => x"358c0001",
    13503 => x"b4230800", 13504 => x"202100ff", 13505 => x"5d82fffc",
    13506 => x"4162001c", 13507 => x"3405fffd", 13508 => x"5c410022",
    13509 => x"e000001e", 13510 => x"40240000", 13511 => x"34210001",
    13512 => x"b4641800", 13513 => x"206300ff", 13514 => x"5c22fffc",
    13515 => x"780c0001", 13516 => x"3163001c", 13517 => x"398c6a68",
    13518 => x"41830000", 13519 => x"780e0001", 13520 => x"780d0001",
    13521 => x"39ce6a5c", 13522 => x"39ad6a60", 13523 => x"0863001d",
    13524 => x"41a20003", 13525 => x"41c10003", 13526 => x"34631005",
    13527 => x"b9602000", 13528 => x"3405001d", 13529 => x"fbffff30",
    13530 => x"41810000", 13531 => x"41a20003", 13532 => x"34031004",
    13533 => x"34210001", 13534 => x"31810000", 13535 => x"41c10003",
    13536 => x"b9802000", 13537 => x"34050001", 13538 => x"fbffff27",
    13539 => x"78010001", 13540 => x"38216a68", 13541 => x"40250000",
    13542 => x"b8a00800", 13543 => x"2b9d0004", 13544 => x"2b8b0014",
    13545 => x"2b8c0010", 13546 => x"2b8d000c", 13547 => x"2b8e0008",
    13548 => x"379c0014", 13549 => x"c3a00000", 13550 => x"379cffc8",
    13551 => x"5b8b0018", 13552 => x"5b8c0014", 13553 => x"5b8d0010",
    13554 => x"5b8e000c", 13555 => x"5b8f0008", 13556 => x"5b9d0004",
    13557 => x"340c0000", 13558 => x"b8205800", 13559 => x"340d0001",
    13560 => x"378e001c", 13561 => x"340f00fd", 13562 => x"e000002b",
    13563 => x"34020000", 13564 => x"b9c00800", 13565 => x"b9801800",
    13566 => x"fbffff80", 13567 => x"b1801000", 13568 => x"5c400005",
    13569 => x"202d00ff", 13570 => x"35a1ffff", 13571 => x"202100ff",
    13572 => x"542f0022", 13573 => x"b9c00800", 13574 => x"b9601000",
    13575 => x"34030010", 13576 => x"f800107d", 13577 => x"358c0001",
    13578 => x"5c20001b", 13579 => x"2b810030", 13580 => x"00220018",
    13581 => x"31610017", 13582 => x"31620014", 13583 => x"00220010",
    13584 => x"31620015", 13585 => x"00220008", 13586 => x"2b810034",
    13587 => x"31620016", 13588 => x"00220018", 13589 => x"3161001b",
    13590 => x"31620018", 13591 => x"00220010", 13592 => x"31620019",
    13593 => x"00220008", 13594 => x"2b81002c", 13595 => x"3162001a",
    13596 => x"00220018", 13597 => x"31610013", 13598 => x"31620010",
    13599 => x"00220010", 13600 => x"31620011", 13601 => x"00220008",
    13602 => x"34010001", 13603 => x"31620012", 13604 => x"e0000003",
    13605 => x"49acffd6", 13606 => x"34010000", 13607 => x"2b9d0004",
    13608 => x"2b8b0018", 13609 => x"2b8c0014", 13610 => x"2b8d0010",
    13611 => x"2b8e000c", 13612 => x"2b8f0008", 13613 => x"379c0038",
    13614 => x"c3a00000", 13615 => x"379cfff8", 13616 => x"5b8b0008",
    13617 => x"5b9d0004", 13618 => x"78030001", 13619 => x"b8205800",
    13620 => x"204200ff", 13621 => x"78010001", 13622 => x"38216a5c",
    13623 => x"38636a60", 13624 => x"44400015", 13625 => x"29640000",
    13626 => x"78028000", 13627 => x"34050004", 13628 => x"b8821000",
    13629 => x"59620000", 13630 => x"40620003", 13631 => x"40210003",
    13632 => x"34031000", 13633 => x"b9602000", 13634 => x"fbfffec7",
    13635 => x"7c210004", 13636 => x"78040001", 13637 => x"38843d38",
    13638 => x"c8011000", 13639 => x"29630000", 13640 => x"28810000",
    13641 => x"38420001", 13642 => x"a0610800", 13643 => x"59610000",
    13644 => x"e0000013", 13645 => x"40620003", 13646 => x"40210003",
    13647 => x"34031000", 13648 => x"b9602000", 13649 => x"34050004",
    13650 => x"fbfffe72", 13651 => x"34030004", 13652 => x"3402ffff",
    13653 => x"5c23000a", 13654 => x"29610000", 13655 => x"34020000",
    13656 => x"4c200007", 13657 => x"78030001", 13658 => x"38633d38",
    13659 => x"28620000", 13660 => x"a0220800", 13661 => x"59610000",
    13662 => x"34020001", 13663 => x"b8400800", 13664 => x"2b9d0004",
    13665 => x"2b8b0008", 13666 => x"379c0008", 13667 => x"c3a00000",
    13668 => x"379cfff8", 13669 => x"5b9d0004", 13670 => x"78010001",
    13671 => x"78020001", 13672 => x"38216a5c", 13673 => x"38426a60",
    13674 => x"40420003", 13675 => x"40210003", 13676 => x"34031074",
    13677 => x"3784000a", 13678 => x"34050002", 13679 => x"0f80000a",
    13680 => x"fbfffe99", 13681 => x"34030002", 13682 => x"3402ffff",
    13683 => x"5c230002", 13684 => x"2f82000a", 13685 => x"b8400800",
    13686 => x"2b9d0004", 13687 => x"379c0008", 13688 => x"c3a00000",
    13689 => x"379cffcc", 13690 => x"5b8b002c", 13691 => x"5b8c0028",
    13692 => x"5b8d0024", 13693 => x"5b8e0020", 13694 => x"5b8f001c",
    13695 => x"5b900018", 13696 => x"5b910014", 13697 => x"5b920010",
    13698 => x"5b93000c", 13699 => x"5b940008", 13700 => x"5b9d0004",
    13701 => x"78030001", 13702 => x"78020001", 13703 => x"38636a5c",
    13704 => x"b8208800", 13705 => x"38426a60", 13706 => x"34010020",
    13707 => x"33810037", 13708 => x"40420003", 13709 => x"40610003",
    13710 => x"37840034", 13711 => x"34031074", 13712 => x"34050002",
    13713 => x"fbfffe33", 13714 => x"34020002", 13715 => x"340bffff",
    13716 => x"5c220051", 13717 => x"2f820034", 13718 => x"3801ffff",
    13719 => x"5c410002", 13720 => x"0f800034", 13721 => x"780d0001",
    13722 => x"780c0001", 13723 => x"340b0001", 13724 => x"39ad6a5c",
    13725 => x"398c6a60", 13726 => x"37900037", 13727 => x"e0000023",
    13728 => x"41b40003", 13729 => x"41930003", 13730 => x"b9c00800",
    13731 => x"34721076", 13732 => x"f8000fb2", 13733 => x"b8202800",
    13734 => x"b9c02000", 13735 => x"ba800800", 13736 => x"ba601000",
    13737 => x"ba401800", 13738 => x"fbfffe5f", 13739 => x"b8207000",
    13740 => x"29e10000", 13741 => x"f8000fa9", 13742 => x"5dc10036",
    13743 => x"29e10000", 13744 => x"2f8e0034", 13745 => x"f8000fa5",
    13746 => x"b5c11800", 13747 => x"41820003", 13748 => x"41a10003",
    13749 => x"2063ffff", 13750 => x"0f830034", 13751 => x"ba002000",
    13752 => x"34631076", 13753 => x"34050001", 13754 => x"fbfffe4f",
    13755 => x"34020001", 13756 => x"5c220028", 13757 => x"2f810034",
    13758 => x"356b0001", 13759 => x"216b00ff", 13760 => x"34210001",
    13761 => x"0f810034", 13762 => x"3d6f0002", 13763 => x"2f830034",
    13764 => x"b62f7800", 13765 => x"29ee0000", 13766 => x"5dc0ffda",
    13767 => x"3401000a", 13768 => x"33810037", 13769 => x"41820003",
    13770 => x"41a10003", 13771 => x"34631075", 13772 => x"37840037",
    13773 => x"34050001", 13774 => x"fbfffe3b", 13775 => x"34020001",
    13776 => x"340bffff", 13777 => x"5c220014", 13778 => x"41a10003",
    13779 => x"41820003", 13780 => x"34031074", 13781 => x"37840034",
    13782 => x"34050002", 13783 => x"fbfffe32", 13784 => x"b8207000",
    13785 => x"34010002", 13786 => x"5dc1000b", 13787 => x"41a10003",
    13788 => x"41820003", 13789 => x"34031074", 13790 => x"37840032",
    13791 => x"34050002", 13792 => x"fbfffde4", 13793 => x"e42e5800",
    13794 => x"356bffff", 13795 => x"e0000002", 13796 => x"340bffff",
    13797 => x"b9600800", 13798 => x"2b9d0004", 13799 => x"2b8b002c",
    13800 => x"2b8c0028", 13801 => x"2b8d0024", 13802 => x"2b8e0020",
    13803 => x"2b8f001c", 13804 => x"2b900018", 13805 => x"2b910014",
    13806 => x"2b920010", 13807 => x"2b93000c", 13808 => x"2b940008",
    13809 => x"379c0034", 13810 => x"c3a00000", 13811 => x"379cffe4",
    13812 => x"5b8b0018", 13813 => x"5b8c0014", 13814 => x"5b8d0010",
    13815 => x"5b8e000c", 13816 => x"5b8f0008", 13817 => x"5b9d0004",
    13818 => x"78010001", 13819 => x"78020001", 13820 => x"38216a5c",
    13821 => x"38426a60", 13822 => x"40420003", 13823 => x"40210003",
    13824 => x"34031074", 13825 => x"3784001c", 13826 => x"34050002",
    13827 => x"fbfffdc1", 13828 => x"34030002", 13829 => x"3402ffff",
    13830 => x"5c230025", 13831 => x"2f81001c", 13832 => x"3802fffd",
    13833 => x"3421ffff", 13834 => x"2021ffff", 13835 => x"50410005",
    13836 => x"78010001", 13837 => x"38212ff4", 13838 => x"0f80001c",
    13839 => x"fbfff562", 13840 => x"780e0001", 13841 => x"780d0001",
    13842 => x"780c0001", 13843 => x"340b0000", 13844 => x"39ce6a5c",
    13845 => x"39ad6a60", 13846 => x"378f001f", 13847 => x"398c2ff0",
    13848 => x"e000000e", 13849 => x"41a20003", 13850 => x"41c10003",
    13851 => x"35631076", 13852 => x"b9e02000", 13853 => x"34050001",
    13854 => x"fbfffda6", 13855 => x"34020001", 13856 => x"5c22000a",
    13857 => x"4382001f", 13858 => x"b9800800", 13859 => x"356b0001",
    13860 => x"fbfff54d", 13861 => x"216bffff", 13862 => x"2f81001c",
    13863 => x"542bfff2", 13864 => x"34020000", 13865 => x"e0000002",
    13866 => x"3402ffff", 13867 => x"b8400800", 13868 => x"2b9d0004",
    13869 => x"2b8b0018", 13870 => x"2b8c0014", 13871 => x"2b8d0010",
    13872 => x"2b8e000c", 13873 => x"2b8f0008", 13874 => x"379c001c",
    13875 => x"c3a00000", 13876 => x"379cffdc", 13877 => x"5b8b0024",
    13878 => x"5b8c0020", 13879 => x"5b8d001c", 13880 => x"5b8e0018",
    13881 => x"5b8f0014", 13882 => x"5b900010", 13883 => x"5b91000c",
    13884 => x"5b920008", 13885 => x"5b9d0004", 13886 => x"206300ff",
    13887 => x"b8208800", 13888 => x"205200ff", 13889 => x"5c600012",
    13890 => x"78040001", 13891 => x"78030001", 13892 => x"38846a5c",
    13893 => x"38636a60", 13894 => x"40620003", 13895 => x"40810003",
    13896 => x"78040001", 13897 => x"34031074", 13898 => x"38846a64",
    13899 => x"34050002", 13900 => x"fbfffd78", 13901 => x"34020002",
    13902 => x"3403ffff", 13903 => x"5c22002b", 13904 => x"78030001",
    13905 => x"38636a66", 13906 => x"0c610000", 13907 => x"78040001",
    13908 => x"38846a66", 13909 => x"78030001", 13910 => x"38636a64",
    13911 => x"2c820000", 13912 => x"2c610000", 13913 => x"34030000",
    13914 => x"3442fffe", 13915 => x"5041001f", 13916 => x"780d0001",
    13917 => x"780c0001", 13918 => x"340b0000", 13919 => x"b8807000",
    13920 => x"39ad6a5c", 13921 => x"398c6a60", 13922 => x"3410000a",
    13923 => x"2dc30000", 13924 => x"3461fffe", 13925 => x"54320012",
    13926 => x"41820003", 13927 => x"41a10003", 13928 => x"34640001",
    13929 => x"b62b7800", 13930 => x"0dc40000", 13931 => x"34631074",
    13932 => x"b9e02000", 13933 => x"34050001", 13934 => x"fbfffd56",
    13935 => x"34020001", 13936 => x"5c220009", 13937 => x"41e10000",
    13938 => x"356b0001", 13939 => x"216b00ff", 13940 => x"5c30ffef",
    13941 => x"b9601800", 13942 => x"e0000004", 13943 => x"3403fffd",
    13944 => x"e0000002", 13945 => x"3403ffff", 13946 => x"b8600800",
    13947 => x"2b9d0004", 13948 => x"2b8b0024", 13949 => x"2b8c0020",
    13950 => x"2b8d001c", 13951 => x"2b8e0018", 13952 => x"2b8f0014",
    13953 => x"2b900010", 13954 => x"2b91000c", 13955 => x"2b920008",
    13956 => x"379c0024", 13957 => x"c3a00000", 13958 => x"379cfffc",
    13959 => x"5b9d0004", 13960 => x"78010001", 13961 => x"382137f0",
    13962 => x"fbfff4e7", 13963 => x"3401ffff", 13964 => x"2b9d0004",
    13965 => x"379c0004", 13966 => x"c3a00000", 13967 => x"379cfff8",
    13968 => x"5b8b0008", 13969 => x"5b9d0004", 13970 => x"78010001",
    13971 => x"b8405800", 13972 => x"78020001", 13973 => x"384240a4",
    13974 => x"38213814", 13975 => x"fbfff4da", 13976 => x"78020001",
    13977 => x"78010001", 13978 => x"38426d18", 13979 => x"38216d28",
    13980 => x"34460090", 13981 => x"34050022", 13982 => x"34040033",
    13983 => x"28220004", 13984 => x"204300ff", 13985 => x"7c670042",
    13986 => x"7c630028", 13987 => x"a0e31800", 13988 => x"5c60000b",
    13989 => x"28230000", 13990 => x"31650000", 13991 => x"31640001",
    13992 => x"31630002", 13993 => x"00430018", 13994 => x"31630003",
    13995 => x"00430010", 13996 => x"00420008", 13997 => x"31630004",
    13998 => x"31620005", 13999 => x"34210010", 14000 => x"5c26ffef",
    14001 => x"34010000", 14002 => x"2b9d0004", 14003 => x"2b8b0008",
    14004 => x"379c0008", 14005 => x"c3a00000", 14006 => x"379cffe8",
    14007 => x"5b8b0018", 14008 => x"5b8c0014", 14009 => x"5b8d0010",
    14010 => x"5b8e000c", 14011 => x"5b8f0008", 14012 => x"5b9d0004",
    14013 => x"780b0001", 14014 => x"b8207800", 14015 => x"b8407000",
    14016 => x"340d0008", 14017 => x"340c0001", 14018 => x"396b4d40",
    14019 => x"a18e1800", 14020 => x"29640008", 14021 => x"7c620000",
    14022 => x"b9e00800", 14023 => x"35adffff", 14024 => x"d8800000",
    14025 => x"3d8c0001", 14026 => x"5da0fff9", 14027 => x"2b9d0004",
    14028 => x"2b8b0018", 14029 => x"2b8c0014", 14030 => x"2b8d0010",
    14031 => x"2b8e000c", 14032 => x"2b8f0008", 14033 => x"379c0018",
    14034 => x"c3a00000", 14035 => x"379cffe8", 14036 => x"5b8b0018",
    14037 => x"5b8c0014", 14038 => x"5b8d0010", 14039 => x"5b8e000c",
    14040 => x"5b8f0008", 14041 => x"5b9d0004", 14042 => x"780b0001",
    14043 => x"b8207800", 14044 => x"340e0008", 14045 => x"340c0000",
    14046 => x"340d0001", 14047 => x"396b4d40", 14048 => x"29620004",
    14049 => x"b9e00800", 14050 => x"35ceffff", 14051 => x"d8400000",
    14052 => x"7c220000", 14053 => x"c8021000", 14054 => x"a1a21000",
    14055 => x"b9826000", 14056 => x"3dad0001", 14057 => x"5dc0fff7",
    14058 => x"34010064", 14059 => x"fbfff006", 14060 => x"b9800800",
    14061 => x"2b9d0004", 14062 => x"2b8b0018", 14063 => x"2b8c0014",
    14064 => x"2b8d0010", 14065 => x"2b8e000c", 14066 => x"2b8f0008",
    14067 => x"379c0018", 14068 => x"c3a00000", 14069 => x"379cffc0",
    14070 => x"5b8b0040", 14071 => x"5b8c003c", 14072 => x"5b8d0038",
    14073 => x"5b8e0034", 14074 => x"5b8f0030", 14075 => x"5b90002c",
    14076 => x"5b910028", 14077 => x"5b920024", 14078 => x"5b930020",
    14079 => x"5b94001c", 14080 => x"5b950018", 14081 => x"5b960014",
    14082 => x"5b970010", 14083 => x"5b98000c", 14084 => x"5b990008",
    14085 => x"5b9d0004", 14086 => x"34020000", 14087 => x"b8206000",
    14088 => x"34030080", 14089 => x"34210008", 14090 => x"780d0001",
    14091 => x"f8000dc5", 14092 => x"39ad4d40", 14093 => x"29a10000",
    14094 => x"340f0000", 14095 => x"44200061", 14096 => x"b9805800",
    14097 => x"34120000", 14098 => x"34110000", 14099 => x"78194000",
    14100 => x"34160001", 14101 => x"34180008", 14102 => x"596c0008",
    14103 => x"45e00022", 14104 => x"29610000", 14105 => x"78028000",
    14106 => x"34030000", 14107 => x"59610010", 14108 => x"29610004",
    14109 => x"59610014", 14110 => x"a0590800", 14111 => x"44200003",
    14112 => x"78024000", 14113 => x"34030000", 14114 => x"a0710800",
    14115 => x"a0522800", 14116 => x"b8a12800", 14117 => x"29640010",
    14118 => x"29610014", 14119 => x"5ca0000e", 14120 => x"a4603000",
    14121 => x"a0260800", 14122 => x"59610014", 14123 => x"00630001",
    14124 => x"3c41001f", 14125 => x"a4403800", 14126 => x"00420001",
    14127 => x"a0872000", 14128 => x"b8231800", 14129 => x"59640010",
    14130 => x"b8430800", 14131 => x"5c25ffeb", 14132 => x"e000003c",
    14133 => x"b8821000", 14134 => x"b8231800", 14135 => x"59620010",
    14136 => x"59630014", 14137 => x"35ee0001", 14138 => x"29a20000",
    14139 => x"3dce0004", 14140 => x"b9800800", 14141 => x"b58e7000",
    14142 => x"d8400000", 14143 => x"5c360031", 14144 => x"b9800800",
    14145 => x"340200f0", 14146 => x"fbffff74", 14147 => x"34140040",
    14148 => x"34130000", 14149 => x"34100001", 14150 => x"34120000",
    14151 => x"34110000", 14152 => x"29a20004", 14153 => x"b9800800",
    14154 => x"29d70004", 14155 => x"d8400000", 14156 => x"29a20004",
    14157 => x"b820a800", 14158 => x"b9800800", 14159 => x"a2f0b800",
    14160 => x"d8400000", 14161 => x"46a10008", 14162 => x"29a30008",
    14163 => x"baa01000", 14164 => x"7eb50000", 14165 => x"b9800800",
    14166 => x"d8600000", 14167 => x"5eb60011", 14168 => x"e0000007",
    14169 => x"29a30008", 14170 => x"b9800800", 14171 => x"bae01000",
    14172 => x"d8600000", 14173 => x"46e00009", 14174 => x"e000000a",
    14175 => x"29c10000", 14176 => x"b8330800", 14177 => x"59c10000",
    14178 => x"29c10004", 14179 => x"b8300800", 14180 => x"59c10004",
    14181 => x"e0000003", 14182 => x"ba539000", 14183 => x"ba308800",
    14184 => x"3e010001", 14185 => x"3e730001", 14186 => x"f6018000",
    14187 => x"3694ffff", 14188 => x"b6139800", 14189 => x"b8208000",
    14190 => x"5e80ffda", 14191 => x"e0000014", 14192 => x"b9e00800",
    14193 => x"2b9d0004", 14194 => x"2b8b0040", 14195 => x"2b8c003c",
    14196 => x"2b8d0038", 14197 => x"2b8e0034", 14198 => x"2b8f0030",
    14199 => x"2b90002c", 14200 => x"2b910028", 14201 => x"2b920024",
    14202 => x"2b930020", 14203 => x"2b94001c", 14204 => x"2b950018",
    14205 => x"2b960014", 14206 => x"2b970010", 14207 => x"2b98000c",
    14208 => x"2b990008", 14209 => x"379c0040", 14210 => x"c3a00000",
    14211 => x"35ef0001", 14212 => x"356b0010", 14213 => x"5df8ff91",
    14214 => x"e3ffffea", 14215 => x"379cfff0", 14216 => x"5b8b0010",
    14217 => x"5b8c000c", 14218 => x"5b8d0008", 14219 => x"5b9d0004",
    14220 => x"b8205800", 14221 => x"78010001", 14222 => x"38214d40",
    14223 => x"28220000", 14224 => x"29610000", 14225 => x"340c0000",
    14226 => x"340d0040", 14227 => x"d8400000", 14228 => x"29610000",
    14229 => x"34020055", 14230 => x"fbffff20", 14231 => x"29610008",
    14232 => x"2962000c", 14233 => x"b9801800", 14234 => x"358c0008",
    14235 => x"f8000bfa", 14236 => x"29610000", 14237 => x"fbffff19",
    14238 => x"5d8dfff9", 14239 => x"2b9d0004", 14240 => x"2b8b0010",
    14241 => x"2b8c000c", 14242 => x"2b8d0008", 14243 => x"379c0010",
    14244 => x"c3a00000", 14245 => x"28210000", 14246 => x"78020001",
    14247 => x"38426da0", 14248 => x"28420000", 14249 => x"3c210008",
    14250 => x"3821000a", 14251 => x"58410000", 14252 => x"28410000",
    14253 => x"20230008", 14254 => x"5c60fffe", 14255 => x"20210001",
    14256 => x"18210001", 14257 => x"c3a00000", 14258 => x"28210000",
    14259 => x"78020001", 14260 => x"38426da0", 14261 => x"28420000",
    14262 => x"3c210008", 14263 => x"38210009", 14264 => x"58410000",
    14265 => x"28410000", 14266 => x"20230008", 14267 => x"5c60fffe",
    14268 => x"20210001", 14269 => x"c3a00000", 14270 => x"28210000",
    14271 => x"78030001", 14272 => x"38636da0", 14273 => x"3c210008",
    14274 => x"28630000", 14275 => x"7c420000", 14276 => x"38210008",
    14277 => x"b8221000", 14278 => x"58620000", 14279 => x"28610000",
    14280 => x"20210008", 14281 => x"5c20fffe", 14282 => x"c3a00000",
    14283 => x"78010001", 14284 => x"78030001", 14285 => x"38216da0",
    14286 => x"38633d4c", 14287 => x"28210000", 14288 => x"28620000",
    14289 => x"58220004", 14290 => x"c3a00000", 14291 => x"379cffc4",
    14292 => x"5b8b001c", 14293 => x"5b8c0018", 14294 => x"5b8d0014",
    14295 => x"5b8e0010", 14296 => x"5b8f000c", 14297 => x"5b900008",
    14298 => x"5b9d0004", 14299 => x"b8206000", 14300 => x"28210000",
    14301 => x"340bffff", 14302 => x"4420002a", 14303 => x"29820004",
    14304 => x"44400028", 14305 => x"fbffeec4", 14306 => x"780e0001",
    14307 => x"b8206800", 14308 => x"340b0000", 14309 => x"3410001f",
    14310 => x"378f0020", 14311 => x"39ce3830", 14312 => x"e000000b",
    14313 => x"fbffeebc", 14314 => x"202400ff", 14315 => x"b56d1000",
    14316 => x"b5eb0800", 14317 => x"30240000", 14318 => x"b8401800",
    14319 => x"b9c00800", 14320 => x"b8802800", 14321 => x"fbfff380",
    14322 => x"356b0001", 14323 => x"29810004", 14324 => x"ee0b1800",
    14325 => x"358c0004", 14326 => x"7c220000", 14327 => x"a0621000",
    14328 => x"5c40fff1", 14329 => x"78010001", 14330 => x"b9602000",
    14331 => x"b9a01000", 14332 => x"b9e01800", 14333 => x"38216d18",
    14334 => x"f80001cc", 14335 => x"b8206000", 14336 => x"b9601800",
    14337 => x"78010001", 14338 => x"fd8b5800", 14339 => x"38213854",
    14340 => x"b9a01000", 14341 => x"b9802000", 14342 => x"fbfff36b",
    14343 => x"c80b5800", 14344 => x"b9600800", 14345 => x"2b9d0004",
    14346 => x"2b8b001c", 14347 => x"2b8c0018", 14348 => x"2b8d0014",
    14349 => x"2b8e0010", 14350 => x"2b8f000c", 14351 => x"2b900008",
    14352 => x"379c003c", 14353 => x"c3a00000", 14354 => x"379cffc8",
    14355 => x"5b8b0018", 14356 => x"5b8c0014", 14357 => x"5b8d0010",
    14358 => x"5b8e000c", 14359 => x"5b8f0008", 14360 => x"5b9d0004",
    14361 => x"b8205800", 14362 => x"28210000", 14363 => x"3405ffff",
    14364 => x"4420002c", 14365 => x"29620004", 14366 => x"4440002a",
    14367 => x"fbffee86", 14368 => x"b8207000", 14369 => x"29610004",
    14370 => x"fbffee83", 14371 => x"b8205800", 14372 => x"34010020",
    14373 => x"4c2b0002", 14374 => x"340b0020", 14375 => x"378d001c",
    14376 => x"78010001", 14377 => x"b9602000", 14378 => x"b9c01000",
    14379 => x"b9a01800", 14380 => x"38216d18", 14381 => x"f8000189",
    14382 => x"b8206000", 14383 => x"78010001", 14384 => x"b9601800",
    14385 => x"38213874", 14386 => x"b9c01000", 14387 => x"b9802000",
    14388 => x"fbfff33d", 14389 => x"e98b5800", 14390 => x"ec0c0800",
    14391 => x"3405ffff", 14392 => x"b9615800", 14393 => x"5d60000f",
    14394 => x"b9a07800", 14395 => x"780d0001", 14396 => x"39ad3830",
    14397 => x"b5eb0800", 14398 => x"40240000", 14399 => x"b56e1000",
    14400 => x"b9a00800", 14401 => x"b8401800", 14402 => x"b8802800",
    14403 => x"356b0001", 14404 => x"fbfff32d", 14405 => x"498bfff8",
    14406 => x"fd8b2800", 14407 => x"c8052800", 14408 => x"b8a00800",
    14409 => x"2b9d0004", 14410 => x"2b8b0018", 14411 => x"2b8c0014",
    14412 => x"2b8d0010", 14413 => x"2b8e000c", 14414 => x"2b8f0008",
    14415 => x"379c0038", 14416 => x"c3a00000", 14417 => x"379cffe4",
    14418 => x"5b8b001c", 14419 => x"5b8c0018", 14420 => x"5b8d0014",
    14421 => x"5b8e0010", 14422 => x"5b8f000c", 14423 => x"5b900008",
    14424 => x"5b9d0004", 14425 => x"780d0001", 14426 => x"39ad6d18",
    14427 => x"b9a00800", 14428 => x"780b0001", 14429 => x"780f0001",
    14430 => x"780e0001", 14431 => x"fbfffe96", 14432 => x"396b6d28",
    14433 => x"340c0000", 14434 => x"39ef3894", 14435 => x"39ce38ac",
    14436 => x"34100008", 14437 => x"29630000", 14438 => x"29640004",
    14439 => x"b8640800", 14440 => x"44200010", 14441 => x"b9801000",
    14442 => x"b9e00800", 14443 => x"fbfff306", 14444 => x"3d810004",
    14445 => x"34020000", 14446 => x"34210008", 14447 => x"b5a10800",
    14448 => x"f8000015", 14449 => x"2023ffff", 14450 => x"08632710",
    14451 => x"b8201000", 14452 => x"14420010", 14453 => x"14630010",
    14454 => x"b9c00800", 14455 => x"fbfff2fa", 14456 => x"358c0001",
    14457 => x"356b0010", 14458 => x"5d90ffeb", 14459 => x"34010000",
    14460 => x"2b9d0004", 14461 => x"2b8b001c", 14462 => x"2b8c0018",
    14463 => x"2b8d0014", 14464 => x"2b8e0010", 14465 => x"2b8f000c",
    14466 => x"2b900008", 14467 => x"379c001c", 14468 => x"c3a00000",
    14469 => x"379cffec", 14470 => x"5b8b0014", 14471 => x"5b8c0010",
    14472 => x"5b8d000c", 14473 => x"5b8e0008", 14474 => x"5b9d0004",
    14475 => x"402d000f", 14476 => x"b8206000", 14477 => x"34010028",
    14478 => x"b8407000", 14479 => x"45a10005", 14480 => x"34010042",
    14481 => x"45a10003", 14482 => x"34010010", 14483 => x"5da10034",
    14484 => x"21cb0002", 14485 => x"5d60000f", 14486 => x"b9800800",
    14487 => x"fbfffef0", 14488 => x"29810000", 14489 => x"34020044",
    14490 => x"21ce0001", 14491 => x"fbfffe1b", 14492 => x"34010000",
    14493 => x"5dcb002d", 14494 => x"780b0001", 14495 => x"396b4d40",
    14496 => x"29620004", 14497 => x"29810000", 14498 => x"d8400000",
    14499 => x"4420fffd", 14500 => x"b9800800", 14501 => x"fbfffee2",
    14502 => x"29810000", 14503 => x"780b0001", 14504 => x"340200be",
    14505 => x"396b6a6c", 14506 => x"fbfffe0c", 14507 => x"356e0008",
    14508 => x"e0000005", 14509 => x"29810000", 14510 => x"fbfffe25",
    14511 => x"31610000", 14512 => x"356b0001", 14513 => x"5d6efffc",
    14514 => x"78020001", 14515 => x"38426a6c", 14516 => x"40410001",
    14517 => x"40430000", 14518 => x"3c210008", 14519 => x"b8230800",
    14520 => x"34030028", 14521 => x"dc200800", 14522 => x"45a3000b",
    14523 => x"34030042", 14524 => x"45a30009", 14525 => x"34030010",
    14526 => x"5da3000b", 14527 => x"40420006", 14528 => x"3c21000f",
    14529 => x"3c42000c", 14530 => x"3421c000", 14531 => x"b8220800",
    14532 => x"e0000006", 14533 => x"3c21000c", 14534 => x"e0000004",
    14535 => x"78018000", 14536 => x"e0000002", 14537 => x"34010000",
    14538 => x"2b9d0004", 14539 => x"2b8b0014", 14540 => x"2b8c0010",
    14541 => x"2b8d000c", 14542 => x"2b8e0008", 14543 => x"379c0014",
    14544 => x"c3a00000", 14545 => x"379cfffc", 14546 => x"5b9d0004",
    14547 => x"34030000", 14548 => x"b8202000", 14549 => x"34090028",
    14550 => x"34080042", 14551 => x"34070010", 14552 => x"34060008",
    14553 => x"40850017", 14554 => x"44a90003", 14555 => x"44a80002",
    14556 => x"5ca70006", 14557 => x"3c630004", 14558 => x"34630008",
    14559 => x"b4230800", 14560 => x"fbffffa5", 14561 => x"e0000005",
    14562 => x"34630001", 14563 => x"34840010", 14564 => x"5c66fff5",
    14565 => x"78018000", 14566 => x"2b9d0004", 14567 => x"379c0004",
    14568 => x"c3a00000", 14569 => x"379cffe0", 14570 => x"5b8b0020",
    14571 => x"5b8c001c", 14572 => x"5b8d0018", 14573 => x"5b8e0014",
    14574 => x"5b8f0010", 14575 => x"5b90000c", 14576 => x"5b910008",
    14577 => x"5b9d0004", 14578 => x"b8205800", 14579 => x"b8408800",
    14580 => x"b8608000", 14581 => x"b8806000", 14582 => x"fbfffe91",
    14583 => x"29610000", 14584 => x"3402000f", 14585 => x"222e00ff",
    14586 => x"fbfffdbc", 14587 => x"29610000", 14588 => x"b9c01000",
    14589 => x"2231ff00", 14590 => x"fbfffdb8", 14591 => x"16310008",
    14592 => x"29610000", 14593 => x"ba201000", 14594 => x"340d0000",
    14595 => x"fbfffdb3", 14596 => x"e0000006", 14597 => x"b60d1000",
    14598 => x"29610000", 14599 => x"40420000", 14600 => x"35ad0001",
    14601 => x"fbfffdad", 14602 => x"498dfffb", 14603 => x"b9600800",
    14604 => x"fbfffe7b", 14605 => x"29610000", 14606 => x"340200aa",
    14607 => x"fbfffda7", 14608 => x"29610000", 14609 => x"fbfffdc2",
    14610 => x"b8207800", 14611 => x"5c2e0022", 14612 => x"29610000",
    14613 => x"fbfffdbe", 14614 => x"b8207000", 14615 => x"5c310020",
    14616 => x"29610000", 14617 => x"340d0000", 14618 => x"fbfffdb9",
    14619 => x"b8208800", 14620 => x"e0000007", 14621 => x"29610000",
    14622 => x"fbfffdb5", 14623 => x"b60d1000", 14624 => x"40420000",
    14625 => x"5c220018", 14626 => x"35ad0001", 14627 => x"498dfffa",
    14628 => x"b9600800", 14629 => x"fbfffe62", 14630 => x"29610000",
    14631 => x"34020055", 14632 => x"fbfffd8e", 14633 => x"29610000",
    14634 => x"b9e01000", 14635 => x"fbfffd8b", 14636 => x"29610000",
    14637 => x"b9c01000", 14638 => x"fbfffd88", 14639 => x"29610000",
    14640 => x"ba201000", 14641 => x"fbfffd85", 14642 => x"34012710",
    14643 => x"fbffedbe", 14644 => x"e0000006", 14645 => x"340cffff",
    14646 => x"e0000004", 14647 => x"340cfffe", 14648 => x"e0000002",
    14649 => x"340cfffd", 14650 => x"b9800800", 14651 => x"2b9d0004",
    14652 => x"2b8b0020", 14653 => x"2b8c001c", 14654 => x"2b8d0018",
    14655 => x"2b8e0014", 14656 => x"2b8f0010", 14657 => x"2b90000c",
    14658 => x"2b910008", 14659 => x"379c0020", 14660 => x"c3a00000",
    14661 => x"379cffe4", 14662 => x"5b8b001c", 14663 => x"5b8c0018",
    14664 => x"5b8d0014", 14665 => x"5b8e0010", 14666 => x"5b8f000c",
    14667 => x"5b900008", 14668 => x"5b9d0004", 14669 => x"b8208000",
    14670 => x"2041001f", 14671 => x"b8405800", 14672 => x"b8607000",
    14673 => x"b8806000", 14674 => x"340d0000", 14675 => x"44200030",
    14676 => x"3441ffff", 14677 => x"b4240800", 14678 => x"1422001f",
    14679 => x"b8807800", 14680 => x"0042001b", 14681 => x"b4410800",
    14682 => x"1562001f", 14683 => x"14210005", 14684 => x"0042001b",
    14685 => x"b44b1000", 14686 => x"14420005", 14687 => x"4422000c",
    14688 => x"78010001", 14689 => x"38213d50", 14690 => x"28220000",
    14691 => x"a1621000", 14692 => x"4c400005", 14693 => x"3442ffff",
    14694 => x"3401ffe0", 14695 => x"b8411000", 14696 => x"34420001",
    14697 => x"340f0020", 14698 => x"c9e27800", 14699 => x"ba000800",
    14700 => x"b9601000", 14701 => x"b9c01800", 14702 => x"b9e02000",
    14703 => x"fbffff7a", 14704 => x"b8206800", 14705 => x"48010016",
    14706 => x"b5cf7000", 14707 => x"b56f5800", 14708 => x"c98f6000",
    14709 => x"e000000e", 14710 => x"b9802000", 14711 => x"4dec0002",
    14712 => x"34040020", 14713 => x"ba000800", 14714 => x"b9601000",
    14715 => x"b9c01800", 14716 => x"fbffff6d", 14717 => x"48010009",
    14718 => x"b5a16800", 14719 => x"35ce0020", 14720 => x"356b0020",
    14721 => x"358cffe0", 14722 => x"e0000002", 14723 => x"340f0020",
    14724 => x"4980fff2", 14725 => x"e0000002", 14726 => x"b8206800",
    14727 => x"b9a00800", 14728 => x"2b9d0004", 14729 => x"2b8b001c",
    14730 => x"2b8c0018", 14731 => x"2b8d0014", 14732 => x"2b8e0010",
    14733 => x"2b8f000c", 14734 => x"2b900008", 14735 => x"379c001c",
    14736 => x"c3a00000", 14737 => x"379cffec", 14738 => x"5b8b0014",
    14739 => x"5b8c0010", 14740 => x"5b8d000c", 14741 => x"5b8e0008",
    14742 => x"5b9d0004", 14743 => x"b8405800", 14744 => x"b8206000",
    14745 => x"b8607000", 14746 => x"b8806800", 14747 => x"fbfffdec",
    14748 => x"29810000", 14749 => x"340200f0", 14750 => x"fbfffd18",
    14751 => x"29810000", 14752 => x"216200ff", 14753 => x"fbfffd15",
    14754 => x"2162ff00", 14755 => x"29810000", 14756 => x"00420008",
    14757 => x"340b0000", 14758 => x"fbfffd10", 14759 => x"e0000006",
    14760 => x"29810000", 14761 => x"fbfffd2a", 14762 => x"b5cb1000",
    14763 => x"30410000", 14764 => x"356b0001", 14765 => x"49abfffb",
    14766 => x"b9a00800", 14767 => x"2b9d0004", 14768 => x"2b8b0014",
    14769 => x"2b8c0010", 14770 => x"2b8d000c", 14771 => x"2b8e0008",
    14772 => x"379c0014", 14773 => x"c3a00000", 14774 => x"379cfffc",
    14775 => x"5b9d0004", 14776 => x"34050000", 14777 => x"b8203000",
    14778 => x"34080043", 14779 => x"34070008", 14780 => x"40c90017",
    14781 => x"5d280006", 14782 => x"3ca50004", 14783 => x"34a50008",
    14784 => x"b4250800", 14785 => x"fbffffd0", 14786 => x"e0000005",
    14787 => x"34a50001", 14788 => x"34c60010", 14789 => x"5ca7fff7",
    14790 => x"3401ffff", 14791 => x"2b9d0004", 14792 => x"379c0004",
    14793 => x"c3a00000", 14794 => x"379cfffc", 14795 => x"5b9d0004",
    14796 => x"34050000", 14797 => x"b8203000", 14798 => x"34080043",
    14799 => x"34070008", 14800 => x"40c90017", 14801 => x"5d280006",
    14802 => x"3ca50004", 14803 => x"34a50008", 14804 => x"b4250800",
    14805 => x"fbffff70", 14806 => x"e0000005", 14807 => x"34a50001",
    14808 => x"34c60010", 14809 => x"5ca7fff7", 14810 => x"3401ffff",
    14811 => x"2b9d0004", 14812 => x"379c0004", 14813 => x"c3a00000",
    14814 => x"78010001", 14815 => x"38216da4", 14816 => x"28220000",
    14817 => x"78010001", 14818 => x"38216dc4", 14819 => x"58220000",
    14820 => x"340103c6", 14821 => x"58410004", 14822 => x"c3a00000",
    14823 => x"c3a00000", 14824 => x"379cfff8", 14825 => x"5b8b0008",
    14826 => x"5b9d0004", 14827 => x"b8205800", 14828 => x"3401000a",
    14829 => x"5d610003", 14830 => x"3401000d", 14831 => x"fbfffff9",
    14832 => x"78020001", 14833 => x"38426dc4", 14834 => x"28420000",
    14835 => x"28410000", 14836 => x"20210001", 14837 => x"5c20fffe",
    14838 => x"584b0008", 14839 => x"2b9d0004", 14840 => x"2b8b0008",
    14841 => x"379c0008", 14842 => x"c3a00000", 14843 => x"379cfff4",
    14844 => x"5b8b000c", 14845 => x"5b8c0008", 14846 => x"5b9d0004",
    14847 => x"b8206000", 14848 => x"b8205800", 14849 => x"e0000004",
    14850 => x"b8400800", 14851 => x"356b0001", 14852 => x"fbffffe4",
    14853 => x"41620000", 14854 => x"5c40fffc", 14855 => x"c96c0800",
    14856 => x"2b9d0004", 14857 => x"2b8b000c", 14858 => x"2b8c0008",
    14859 => x"379c000c", 14860 => x"c3a00000", 14861 => x"78010001",
    14862 => x"38216dc4", 14863 => x"28220000", 14864 => x"3401ffff",
    14865 => x"28430000", 14866 => x"20630002", 14867 => x"44600003",
    14868 => x"2841000c", 14869 => x"202100ff", 14870 => x"c3a00000",
    14871 => x"28250008", 14872 => x"28240000", 14873 => x"28260004",
    14874 => x"b4451800", 14875 => x"88642000", 14876 => x"5822001c",
    14877 => x"88461000", 14878 => x"b4821000", 14879 => x"2824000c",
    14880 => x"1442000c", 14881 => x"b4442000", 14882 => x"28220014",
    14883 => x"4c820005", 14884 => x"28240010", 14885 => x"44800008",
    14886 => x"4ca3000b", 14887 => x"e0000006", 14888 => x"28220018",
    14889 => x"4c440006", 14890 => x"28240010", 14891 => x"44800002",
    14892 => x"4c650005", 14893 => x"58230008", 14894 => x"e0000003",
    14895 => x"58230008", 14896 => x"b8801000", 14897 => x"58220020",
    14898 => x"b8400800", 14899 => x"c3a00000", 14900 => x"2822000c",
    14901 => x"58200008", 14902 => x"58220020", 14903 => x"c3a00000",
    14904 => x"379cfff8", 14905 => x"5b8b0008", 14906 => x"5b9d0004",
    14907 => x"b8205800", 14908 => x"58200014", 14909 => x"b8400800",
    14910 => x"f80009ef", 14911 => x"2963000c", 14912 => x"29620000",
    14913 => x"4823000b", 14914 => x"29610004", 14915 => x"4c410003",
    14916 => x"34420001", 14917 => x"59620000", 14918 => x"29620000",
    14919 => x"5c410011", 14920 => x"34010001", 14921 => x"59610014",
    14922 => x"59610010", 14923 => x"e000000e", 14924 => x"29610008",
    14925 => x"4c220003", 14926 => x"3442ffff", 14927 => x"59620000",
    14928 => x"29620000", 14929 => x"5c410007", 14930 => x"34010001",
    14931 => x"59610014", 14932 => x"59600000", 14933 => x"59600010",
    14934 => x"3401ffff", 14935 => x"e0000002", 14936 => x"29610010",
    14937 => x"2b9d0004", 14938 => x"2b8b0008", 14939 => x"379c0008",
    14940 => x"c3a00000", 14941 => x"58200010", 14942 => x"58200000",
    14943 => x"58200014", 14944 => x"c3a00000", 14945 => x"379cfff4",
    14946 => x"5b8b000c", 14947 => x"5b8c0008", 14948 => x"5b9d0004",
    14949 => x"b8205800", 14950 => x"b8406000", 14951 => x"78020001",
    14952 => x"34010000", 14953 => x"384238c8", 14954 => x"b9601800",
    14955 => x"b9802000", 14956 => x"fbffc619", 14957 => x"78010001",
    14958 => x"38216db0", 14959 => x"28220000", 14960 => x"484b0013",
    14961 => x"78050001", 14962 => x"38a56d08", 14963 => x"c9621000",
    14964 => x"45800007", 14965 => x"28a10000", 14966 => x"34040001",
    14967 => x"bc821000", 14968 => x"28230028", 14969 => x"b8431000",
    14970 => x"e0000007", 14971 => x"28a10000", 14972 => x"34040001",
    14973 => x"bc821000", 14974 => x"28230028", 14975 => x"a4401000",
    14976 => x"a0431000", 14977 => x"58220028", 14978 => x"e0000011",
    14979 => x"78050001", 14980 => x"38a56d08", 14981 => x"45800007",
    14982 => x"28a10000", 14983 => x"34020001", 14984 => x"bc4b1000",
    14985 => x"28230024", 14986 => x"b8431000", 14987 => x"e0000007",
    14988 => x"28a10000", 14989 => x"34020001", 14990 => x"bc4b1000",
    14991 => x"28230024", 14992 => x"a4401000", 14993 => x"a0431000",
    14994 => x"58220024", 14995 => x"78010001", 14996 => x"38216d08",
    14997 => x"28210000", 14998 => x"78020001", 14999 => x"78030001",
    15000 => x"28250028", 15001 => x"28260024", 15002 => x"384238dc",
    15003 => x"34010000", 15004 => x"386340b8", 15005 => x"b9602000",
    15006 => x"fbffc5e7", 15007 => x"2b9d0004", 15008 => x"2b8b000c",
    15009 => x"2b8c0008", 15010 => x"379c000c", 15011 => x"c3a00000",
    15012 => x"379cfff0", 15013 => x"5b8b0010", 15014 => x"5b8c000c",
    15015 => x"5b8d0008", 15016 => x"5b9d0004", 15017 => x"b8406800",
    15018 => x"b8606000", 15019 => x"34020000", 15020 => x"34030028",
    15021 => x"b8205800", 15022 => x"f8000a22", 15023 => x"b9600800",
    15024 => x"b9a01000", 15025 => x"34030014", 15026 => x"f80009a0",
    15027 => x"596c0014", 15028 => x"2b9d0004", 15029 => x"2b8b0010",
    15030 => x"2b8c000c", 15031 => x"2b8d0008", 15032 => x"379c0010",
    15033 => x"c3a00000", 15034 => x"b8201800", 15035 => x"e0000004",
    15036 => x"28840000", 15037 => x"34630008", 15038 => x"44820006",
    15039 => x"28610004", 15040 => x"b8602000", 15041 => x"5c20fffb",
    15042 => x"78010001", 15043 => x"38213900", 15044 => x"c3a00000",
    15045 => x"78020001", 15046 => x"38426d08", 15047 => x"28420000",
    15048 => x"b8201800", 15049 => x"34010000", 15050 => x"28440008",
    15051 => x"20840002", 15052 => x"4480000c", 15053 => x"34040002",
    15054 => x"58440008", 15055 => x"78060001", 15056 => x"28420010",
    15057 => x"38c63d54", 15058 => x"28c40000", 15059 => x"3445ff9b",
    15060 => x"54a40004", 15061 => x"08420064", 15062 => x"34010001",
    15063 => x"58620000", 15064 => x"c3a00000", 15065 => x"379cfff0",
    15066 => x"5b8b0010", 15067 => x"5b8c000c", 15068 => x"5b8d0008",
    15069 => x"5b9d0004", 15070 => x"780b0001", 15071 => x"b8206000",
    15072 => x"78010001", 15073 => x"396b6db0", 15074 => x"38216da8",
    15075 => x"28210000", 15076 => x"296d0000", 15077 => x"b42d6800",
    15078 => x"29810000", 15079 => x"b9a01000", 15080 => x"f8000116",
    15081 => x"29810004", 15082 => x"29630000", 15083 => x"b9a01000",
    15084 => x"f800019b", 15085 => x"5980000c", 15086 => x"59800008",
    15087 => x"2b9d0004", 15088 => x"2b8b0010", 15089 => x"2b8c000c",
    15090 => x"2b8d0008", 15091 => x"379c0010", 15092 => x"c3a00000",
    15093 => x"379cfff8", 15094 => x"5b8b0008", 15095 => x"5b9d0004",
    15096 => x"b8205800", 15097 => x"28210000", 15098 => x"f800016e",
    15099 => x"78010001", 15100 => x"38216d08", 15101 => x"28210000",
    15102 => x"34020001", 15103 => x"34030009", 15104 => x"58220004",
    15105 => x"5963000c", 15106 => x"78030001", 15107 => x"38633d58",
    15108 => x"59620008", 15109 => x"28620000", 15110 => x"5822004c",
    15111 => x"2b9d0004", 15112 => x"2b8b0008", 15113 => x"379c0008",
    15114 => x"c3a00000", 15115 => x"b8201000", 15116 => x"28210000",
    15117 => x"2823004c", 15118 => x"34010000", 15119 => x"44600016",
    15120 => x"28430004", 15121 => x"28630038", 15122 => x"44600013",
    15123 => x"78030001", 15124 => x"38636d08", 15125 => x"28630000",
    15126 => x"28640004", 15127 => x"20840004", 15128 => x"4480000d",
    15129 => x"28630004", 15130 => x"20630008", 15131 => x"5c60000a",
    15132 => x"2842000c", 15133 => x"3403000a", 15134 => x"34010001",
    15135 => x"54430006", 15136 => x"78010001", 15137 => x"3c420002",
    15138 => x"382140f4", 15139 => x"b4220800", 15140 => x"28210000",
    15141 => x"c3a00000", 15142 => x"379cfff0", 15143 => x"5b8b000c",
    15144 => x"5b8c0008", 15145 => x"5b9d0004", 15146 => x"2822000c",
    15147 => x"b8205800", 15148 => x"34010009", 15149 => x"3442ffff",
    15150 => x"544100a9", 15151 => x"78010001", 15152 => x"3c420002",
    15153 => x"382140cc", 15154 => x"b4220800", 15155 => x"28210000",
    15156 => x"c0200000", 15157 => x"78010001", 15158 => x"38216d08",
    15159 => x"28210000", 15160 => x"28220004", 15161 => x"20420008",
    15162 => x"5c40009d", 15163 => x"28230004", 15164 => x"78028000",
    15165 => x"b8621000", 15166 => x"58220004", 15167 => x"3401000a",
    15168 => x"e0000096", 15169 => x"78010001", 15170 => x"38216d08",
    15171 => x"28210000", 15172 => x"78040001", 15173 => x"38843d38",
    15174 => x"28230004", 15175 => x"28820000", 15176 => x"a0621000",
    15177 => x"58220004", 15178 => x"28220004", 15179 => x"20420008",
    15180 => x"5c400089", 15181 => x"28210004", 15182 => x"20210004",
    15183 => x"44220088", 15184 => x"34010001", 15185 => x"e0000085",
    15186 => x"29610000", 15187 => x"2821004c", 15188 => x"44200083",
    15189 => x"fbffc51d", 15190 => x"29610004", 15191 => x"f800015e",
    15192 => x"fbffc523", 15193 => x"34010008", 15194 => x"e000007c",
    15195 => x"78010001", 15196 => x"38216d08", 15197 => x"28210000",
    15198 => x"34020002", 15199 => x"58220008", 15200 => x"29610000",
    15201 => x"2821004c", 15202 => x"44200075", 15203 => x"29610004",
    15204 => x"28210038", 15205 => x"44200072", 15206 => x"78010001",
    15207 => x"38216d0c", 15208 => x"28210000", 15209 => x"340300a2",
    15210 => x"58230000", 15211 => x"34030003", 15212 => x"58230010",
    15213 => x"34030001", 15214 => x"5823001c", 15215 => x"5962000c",
    15216 => x"78020001", 15217 => x"34010000", 15218 => x"3842390c",
    15219 => x"e0000017", 15220 => x"78010001", 15221 => x"38216d0c",
    15222 => x"28210000", 15223 => x"2822001c", 15224 => x"20420001",
    15225 => x"4440005e", 15226 => x"34020002", 15227 => x"5822001c",
    15228 => x"fbfff627", 15229 => x"342107d0", 15230 => x"59610010",
    15231 => x"34010003", 15232 => x"e0000056", 15233 => x"fbfff622",
    15234 => x"29620010", 15235 => x"54410054", 15236 => x"34010007",
    15237 => x"5961000c", 15238 => x"78020001", 15239 => x"5960001c",
    15240 => x"34010000", 15241 => x"38423920", 15242 => x"fbffc4fb",
    15243 => x"e000004c", 15244 => x"37810010", 15245 => x"fbffff38",
    15246 => x"44200049", 15247 => x"78030001", 15248 => x"38633d14",
    15249 => x"2b810010", 15250 => x"28620000", 15251 => x"f800083e",
    15252 => x"3802c34f", 15253 => x"e8221000", 15254 => x"5b810010",
    15255 => x"64210000", 15256 => x"b8410800", 15257 => x"44200005",
    15258 => x"34010064", 15259 => x"59610014", 15260 => x"3401ff9c",
    15261 => x"e0000003", 15262 => x"59600014", 15263 => x"34010064",
    15264 => x"59610018", 15265 => x"29630014", 15266 => x"29640018",
    15267 => x"78020001", 15268 => x"34010000", 15269 => x"38423938",
    15270 => x"fbffc4df", 15271 => x"34010004", 15272 => x"e000002e",
    15273 => x"29610004", 15274 => x"f80001e9", 15275 => x"b8206000",
    15276 => x"5c20002b", 15277 => x"37810010", 15278 => x"fbffff17",
    15279 => x"442c0028", 15280 => x"78040001", 15281 => x"38843d14",
    15282 => x"2b810010", 15283 => x"28820000", 15284 => x"f800081d",
    15285 => x"29620014", 15286 => x"5b810010", 15287 => x"44220009",
    15288 => x"2961001c", 15289 => x"29620018", 15290 => x"b4410800",
    15291 => x"5961001c", 15292 => x"29610004", 15293 => x"2962001c",
    15294 => x"f80001b3", 15295 => x"e0000018", 15296 => x"29620014",
    15297 => x"5c220016", 15298 => x"2961001c", 15299 => x"34217530",
    15300 => x"5961001c", 15301 => x"29610004", 15302 => x"2962001c",
    15303 => x"f80001aa", 15304 => x"34010005", 15305 => x"e000000d",
    15306 => x"29610004", 15307 => x"f80001c8", 15308 => x"5c20000b",
    15309 => x"78020001", 15310 => x"38423958", 15311 => x"fbffc4b6",
    15312 => x"34010006", 15313 => x"e0000005", 15314 => x"b9600800",
    15315 => x"fbffff38", 15316 => x"5c200003", 15317 => x"34010009",
    15318 => x"5961000c", 15319 => x"2b9d0004", 15320 => x"2b8b000c",
    15321 => x"2b8c0008", 15322 => x"379c0010", 15323 => x"c3a00000",
    15324 => x"78040001", 15325 => x"64630000", 15326 => x"38846d08",
    15327 => x"28850000", 15328 => x"c8031800", 15329 => x"78048000",
    15330 => x"78060001", 15331 => x"a0641800", 15332 => x"38c63d5c",
    15333 => x"b4641800", 15334 => x"28c40000", 15335 => x"3c210018",
    15336 => x"a0441000", 15337 => x"b8410800", 15338 => x"b8231800",
    15339 => x"58a3004c", 15340 => x"c3a00000", 15341 => x"78040001",
    15342 => x"64630000", 15343 => x"38846d08", 15344 => x"28850000",
    15345 => x"c8031800", 15346 => x"78048000", 15347 => x"78060001",
    15348 => x"a0641800", 15349 => x"38c63d5c", 15350 => x"b4641800",
    15351 => x"28c40000", 15352 => x"3c210018", 15353 => x"a0441000",
    15354 => x"b8410800", 15355 => x"b8231800", 15356 => x"58a3004c",
    15357 => x"c3a00000", 15358 => x"34030005", 15359 => x"5823002c",
    15360 => x"3803fffb", 15361 => x"58230030", 15362 => x"3403ff6a",
    15363 => x"5823001c", 15364 => x"3403fffe", 15365 => x"58230018",
    15366 => x"34030001", 15367 => x"58230028", 15368 => x"340300c8",
    15369 => x"58230048", 15370 => x"34032710", 15371 => x"58230040",
    15372 => x"34030064", 15373 => x"58230044", 15374 => x"5822000c",
    15375 => x"58200014", 15376 => x"c3a00000", 15377 => x"379cfff0",
    15378 => x"5b8b0010", 15379 => x"5b8c000c", 15380 => x"5b8d0008",
    15381 => x"5b9d0004", 15382 => x"b8205800", 15383 => x"2821000c",
    15384 => x"b8406800", 15385 => x"340c0000", 15386 => x"5c610047",
    15387 => x"34010022", 15388 => x"34030000", 15389 => x"fbffffbf",
    15390 => x"29620004", 15391 => x"34010025", 15392 => x"34030000",
    15393 => x"fbffffbb", 15394 => x"29610008", 15395 => x"4c200004",
    15396 => x"596d0004", 15397 => x"596d0008", 15398 => x"e000003b",
    15399 => x"4da10005", 15400 => x"29620000", 15401 => x"78010040",
    15402 => x"b4410800", 15403 => x"59610000", 15404 => x"29630000",
    15405 => x"78050001", 15406 => x"29620004", 15407 => x"38a53d60",
    15408 => x"28a10000", 15409 => x"b5a32000", 15410 => x"c8826000",
    15411 => x"482c0006", 15412 => x"78050001", 15413 => x"38a53d64",
    15414 => x"28a10000", 15415 => x"49810002", 15416 => x"e0000002",
    15417 => x"b8206000", 15418 => x"78050001", 15419 => x"38a53d68",
    15420 => x"28a10000", 15421 => x"4c240006", 15422 => x"4c220005",
    15423 => x"c8611800", 15424 => x"c8410800", 15425 => x"59630000",
    15426 => x"59610004", 15427 => x"29610004", 15428 => x"b9801000",
    15429 => x"596d0008", 15430 => x"34214000", 15431 => x"59610004",
    15432 => x"35610018", 15433 => x"fbfffdce", 15434 => x"78030001",
    15435 => x"38636d08", 15436 => x"29620010", 15437 => x"b8206800",
    15438 => x"28610000", 15439 => x"34030000", 15440 => x"582d0040",
    15441 => x"34410001", 15442 => x"59610010", 15443 => x"34010026",
    15444 => x"fbffff88", 15445 => x"34010020", 15446 => x"b9a01000",
    15447 => x"34030000", 15448 => x"fbffff84", 15449 => x"b9801000",
    15450 => x"34010021", 15451 => x"34030001", 15452 => x"fbffff80",
    15453 => x"b9801000", 15454 => x"3561003c", 15455 => x"fbfffdd9",
    15456 => x"7c2c0000", 15457 => x"b9800800", 15458 => x"2b9d0004",
    15459 => x"2b8b0010", 15460 => x"2b8c000c", 15461 => x"2b8d0008",
    15462 => x"379c0010", 15463 => x"c3a00000", 15464 => x"379cfff8",
    15465 => x"5b8b0008", 15466 => x"5b9d0004", 15467 => x"b8205800",
    15468 => x"2821002c", 15469 => x"59600004", 15470 => x"59600000",
    15471 => x"59610024", 15472 => x"3401ffff", 15473 => x"59610008",
    15474 => x"59600010", 15475 => x"35610018", 15476 => x"fbfffdc0",
    15477 => x"3561003c", 15478 => x"fbfffde7", 15479 => x"78020001",
    15480 => x"35610054", 15481 => x"34030010", 15482 => x"38424120",
    15483 => x"fbfffe29", 15484 => x"2961000c", 15485 => x"34020001",
    15486 => x"fbfffde3", 15487 => x"34010024", 15488 => x"34020001",
    15489 => x"34030001", 15490 => x"fbffff5a", 15491 => x"2b9d0004",
    15492 => x"2b8b0008", 15493 => x"379c0008", 15494 => x"c3a00000",
    15495 => x"379cfff8", 15496 => x"5b8b0008", 15497 => x"5b9d0004",
    15498 => x"b8205800", 15499 => x"34010005", 15500 => x"59610018",
    15501 => x"3801fffa", 15502 => x"5961001c", 15503 => x"34010001",
    15504 => x"59610014", 15505 => x"34017530", 15506 => x"59610010",
    15507 => x"3401fbb4", 15508 => x"59610008", 15509 => x"3401ffe2",
    15510 => x"59610004", 15511 => x"340104b0", 15512 => x"59610034",
    15513 => x"340103e8", 15514 => x"5961002c", 15515 => x"34010064",
    15516 => x"59610030", 15517 => x"78010001", 15518 => x"38216db0",
    15519 => x"28250000", 15520 => x"b8403000", 15521 => x"59620070",
    15522 => x"c8652800", 15523 => x"78020001", 15524 => x"b8602000",
    15525 => x"59650080", 15526 => x"3842396c", 15527 => x"59630074",
    15528 => x"5960007c", 15529 => x"b8c01800", 15530 => x"59600084",
    15531 => x"34010000", 15532 => x"fbffc3d9", 15533 => x"35610004",
    15534 => x"fbfffd86", 15535 => x"35610028", 15536 => x"fbfffdad",
    15537 => x"2b9d0004", 15538 => x"2b8b0008", 15539 => x"379c0008",
    15540 => x"c3a00000", 15541 => x"379cfff8", 15542 => x"5b8b0008",
    15543 => x"5b9d0004", 15544 => x"b8205800", 15545 => x"29630080",
    15546 => x"78020001", 15547 => x"38423984", 15548 => x"34010000",
    15549 => x"fbffc3c8", 15550 => x"3401ffff", 15551 => x"59610048",
    15552 => x"5961004c", 15553 => x"59610050", 15554 => x"59610054",
    15555 => x"34010001", 15556 => x"59610084", 15557 => x"59600044",
    15558 => x"35610004", 15559 => x"59600040", 15560 => x"59600058",
    15561 => x"5960005c", 15562 => x"59600060", 15563 => x"59600068",
    15564 => x"5960006c", 15565 => x"59600078", 15566 => x"fbfffd66",
    15567 => x"35610028", 15568 => x"fbfffd8d", 15569 => x"29610070",
    15570 => x"34020001", 15571 => x"fbfffd8e", 15572 => x"29610074",
    15573 => x"34020001", 15574 => x"fbfffd8b", 15575 => x"34010004",
    15576 => x"34020001", 15577 => x"34030001", 15578 => x"fbffff13",
    15579 => x"2b9d0004", 15580 => x"2b8b0008", 15581 => x"379c0008",
    15582 => x"c3a00000", 15583 => x"379cfff8", 15584 => x"5b8b0008",
    15585 => x"5b9d0004", 15586 => x"b8205800", 15587 => x"28210074",
    15588 => x"34020000", 15589 => x"fbfffd7c", 15590 => x"59600084",
    15591 => x"2b9d0004", 15592 => x"2b8b0008", 15593 => x"379c0008",
    15594 => x"c3a00000", 15595 => x"379cfff0", 15596 => x"5b8b0010",
    15597 => x"5b8c000c", 15598 => x"5b8d0008", 15599 => x"5b9d0004",
    15600 => x"28240084", 15601 => x"b8205800", 15602 => x"34010001",
    15603 => x"44800078", 15604 => x"29610070", 15605 => x"5c610002",
    15606 => x"59620048", 15607 => x"29610074", 15608 => x"5c610002",
    15609 => x"5962004c", 15610 => x"29610048", 15611 => x"48010009",
    15612 => x"29620050", 15613 => x"48020006", 15614 => x"4c220005",
    15615 => x"29630040", 15616 => x"78020040", 15617 => x"b4621000",
    15618 => x"59620040", 15619 => x"59610050", 15620 => x"2961004c",
    15621 => x"48010009", 15622 => x"29620054", 15623 => x"48020006",
    15624 => x"4c220005", 15625 => x"29630044", 15626 => x"78020040",
    15627 => x"b4621000", 15628 => x"59620044", 15629 => x"59610054",
    15630 => x"29630048", 15631 => x"34010000", 15632 => x"4803005b",
    15633 => x"2962004c", 15634 => x"48020059", 15635 => x"296c0040",
    15636 => x"29610038", 15637 => x"b46c1800", 15638 => x"296c0044",
    15639 => x"c8621000", 15640 => x"c84c6000", 15641 => x"44200006",
    15642 => x"218c3fff", 15643 => x"21812000", 15644 => x"44200003",
    15645 => x"3401c000", 15646 => x"b9816000", 15647 => x"b9801000",
    15648 => x"35610004", 15649 => x"fbfffcf6", 15650 => x"29620080",
    15651 => x"78030001", 15652 => x"38636d08", 15653 => x"2042000f",
    15654 => x"b8206800", 15655 => x"3c420010", 15656 => x"28610000",
    15657 => x"21a3ffff", 15658 => x"b8621000", 15659 => x"58220044",
    15660 => x"29630040", 15661 => x"29620048", 15662 => x"34010005",
    15663 => x"b4621000", 15664 => x"34030000", 15665 => x"fbfffebc",
    15666 => x"29630044", 15667 => x"2962004c", 15668 => x"34010002",
    15669 => x"b4621000", 15670 => x"34030000", 15671 => x"fbfffeb6",
    15672 => x"34010001", 15673 => x"b9801000", 15674 => x"34030000",
    15675 => x"fbfffeb2", 15676 => x"29620078", 15677 => x"34030000",
    15678 => x"34410001", 15679 => x"59610078", 15680 => x"34010006",
    15681 => x"fbfffeac", 15682 => x"34010000", 15683 => x"b9a01000",
    15684 => x"34030001", 15685 => x"fbfffea8", 15686 => x"78020001",
    15687 => x"3401ffff", 15688 => x"38423d6c", 15689 => x"5961004c",
    15690 => x"59610048", 15691 => x"29630040", 15692 => x"28410000",
    15693 => x"4c23000a", 15694 => x"29620044", 15695 => x"4c220008",
    15696 => x"78040001", 15697 => x"38843d70", 15698 => x"28810000",
    15699 => x"b4611800", 15700 => x"b4410800", 15701 => x"59630040",
    15702 => x"59610044", 15703 => x"29610038", 15704 => x"4420000f",
    15705 => x"2961006c", 15706 => x"29620068", 15707 => x"4c220006",
    15708 => x"34210001", 15709 => x"5961006c", 15710 => x"29610040",
    15711 => x"3421ffff", 15712 => x"e0000006", 15713 => x"4c410006",
    15714 => x"3421ffff", 15715 => x"5961006c", 15716 => x"29610040",
    15717 => x"34210001", 15718 => x"59610040", 15719 => x"35610028",
    15720 => x"b9801000", 15721 => x"fbfffccf", 15722 => x"7c210000",
    15723 => x"2b9d0004", 15724 => x"2b8b0010", 15725 => x"2b8c000c",
    15726 => x"2b8d0008", 15727 => x"379c0010", 15728 => x"c3a00000",
    15729 => x"379cfff0", 15730 => x"5b8b0008", 15731 => x"5b9d0004",
    15732 => x"b8205800", 15733 => x"1443001f", 15734 => x"3781000c",
    15735 => x"4802000b", 15736 => x"00440012", 15737 => x"3c63000e",
    15738 => x"3c42000e", 15739 => x"b8641800", 15740 => x"5b820010",
    15741 => x"34021f40", 15742 => x"5b83000c", 15743 => x"fbffcbe9",
    15744 => x"2b820010", 15745 => x"e0000009", 15746 => x"0842c000",
    15747 => x"5b820010", 15748 => x"1442001f", 15749 => x"5b82000c",
    15750 => x"34021f40", 15751 => x"fbffcbe1", 15752 => x"2b820010",
    15753 => x"c8021000", 15754 => x"0041001f", 15755 => x"b4221000",
    15756 => x"14420001", 15757 => x"34010000", 15758 => x"59620068",
    15759 => x"2b9d0004", 15760 => x"2b8b0008", 15761 => x"379c0010",
    15762 => x"c3a00000", 15763 => x"28220068", 15764 => x"2821006c",
    15765 => x"fc410800", 15766 => x"c3a00000", 15767 => x"58220004",
    15768 => x"5820001c", 15769 => x"58230008", 15770 => x"5820000c",
    15771 => x"58200010", 15772 => x"58200000", 15773 => x"c3a00000",
    15774 => x"379cfffc", 15775 => x"5b9d0004", 15776 => x"34020001",
    15777 => x"58220000", 15778 => x"58200014", 15779 => x"5820001c",
    15780 => x"5820000c", 15781 => x"58200010", 15782 => x"28210004",
    15783 => x"fbfffcba", 15784 => x"78010001", 15785 => x"38216db0",
    15786 => x"28210000", 15787 => x"34020001", 15788 => x"fbfffcb5",
    15789 => x"2b9d0004", 15790 => x"379c0004", 15791 => x"c3a00000",
    15792 => x"379cffb0", 15793 => x"5b8b0010", 15794 => x"5b8c000c",
    15795 => x"5b8d0008", 15796 => x"5b9d0004", 15797 => x"b8205800",
    15798 => x"b8406000", 15799 => x"b8606800", 15800 => x"37810014",
    15801 => x"34020000", 15802 => x"34030040", 15803 => x"f8000715",
    15804 => x"3401c000", 15805 => x"78040001", 15806 => x"5b810020",
    15807 => x"38846db0", 15808 => x"34014000", 15809 => x"5b810044",
    15810 => x"28810000", 15811 => x"5da10005", 15812 => x"78030001",
    15813 => x"38634d4c", 15814 => x"586c0000", 15815 => x"e0000027",
    15816 => x"3dad0005", 15817 => x"b56d5800", 15818 => x"29610000",
    15819 => x"44200023", 15820 => x"78030001", 15821 => x"38634d4c",
    15822 => x"28610000", 15823 => x"29620010", 15824 => x"c9810800",
    15825 => x"20213fff", 15826 => x"1423000c", 15827 => x"5c400007",
    15828 => x"3c630002", 15829 => x"5961000c", 15830 => x"34010001",
    15831 => x"59630014", 15832 => x"59610010", 15833 => x"e0000015",
    15834 => x"2964000c", 15835 => x"34420001", 15836 => x"b4240800",
    15837 => x"29640014", 15838 => x"b4641800", 15839 => x"3c630002",
    15840 => x"37840050", 15841 => x"b4831800", 15842 => x"2863ffc4",
    15843 => x"59620010", 15844 => x"b4230800", 15845 => x"29630008",
    15846 => x"5961000c", 15847 => x"5c430007", 15848 => x"f80005bc",
    15849 => x"59610018", 15850 => x"34010001", 15851 => x"5961001c",
    15852 => x"5960000c", 15853 => x"59600010", 15854 => x"34010000",
    15855 => x"2b9d0004", 15856 => x"2b8b0010", 15857 => x"2b8c000c",
    15858 => x"2b8d0008", 15859 => x"379c0050", 15860 => x"c3a00000",
    15861 => x"78030001", 15862 => x"38636d08", 15863 => x"5c40000a",
    15864 => x"34040001", 15865 => x"28620000", 15866 => x"bc810800",
    15867 => x"202100ff", 15868 => x"28430020", 15869 => x"3c210010",
    15870 => x"a4200800", 15871 => x"a0230800", 15872 => x"e0000008",
    15873 => x"28620000", 15874 => x"34040001", 15875 => x"bc810800",
    15876 => x"28430020", 15877 => x"202100ff", 15878 => x"3c210010",
    15879 => x"b8230800", 15880 => x"58410020", 15881 => x"c3a00000",
    15882 => x"379cffe0", 15883 => x"5b8b0010", 15884 => x"5b8c000c",
    15885 => x"5b8d0008", 15886 => x"5b9d0004", 15887 => x"b8406000",
    15888 => x"c8231000", 15889 => x"1441001f", 15890 => x"b8605800",
    15891 => x"48010002", 15892 => x"e0000020", 15893 => x"c9836000",
    15894 => x"1583001f", 15895 => x"5c60001d", 15896 => x"4583001c",
    15897 => x"78050001", 15898 => x"38a53d74", 15899 => x"28a40000",
    15900 => x"3403ffff", 15901 => x"f8000560", 15902 => x"5b81001c",
    15903 => x"5b820020", 15904 => x"3781001c", 15905 => x"b9601000",
    15906 => x"fbffcb46", 15907 => x"78050001", 15908 => x"38a53ce4",
    15909 => x"28a40000", 15910 => x"34030000", 15911 => x"34010000",
    15912 => x"b9801000", 15913 => x"f8000554", 15914 => x"5b810014",
    15915 => x"5b820018", 15916 => x"37810014", 15917 => x"b9601000",
    15918 => x"2b8d0020", 15919 => x"fbffcb39", 15920 => x"2b810018",
    15921 => x"4da10004", 15922 => x"b9a00800", 15923 => x"e0000002",
    15924 => x"3401ffff", 15925 => x"2b9d0004", 15926 => x"2b8b0010",
    15927 => x"2b8c000c", 15928 => x"2b8d0008", 15929 => x"379c0020",
    15930 => x"c3a00000", 15931 => x"379cfff8", 15932 => x"5b8b0008",
    15933 => x"5b9d0004", 15934 => x"34020001", 15935 => x"44220009",
    15936 => x"34020002", 15937 => x"4422000c", 15938 => x"5c200017",
    15939 => x"78010001", 15940 => x"38216d08", 15941 => x"282b0000",
    15942 => x"356b0018", 15943 => x"e000000a", 15944 => x"78010001",
    15945 => x"38216d08", 15946 => x"282b0000", 15947 => x"356b0014",
    15948 => x"e0000005", 15949 => x"78010001", 15950 => x"38216d08",
    15951 => x"282b0000", 15952 => x"356b001c", 15953 => x"340107d0",
    15954 => x"fbfff356", 15955 => x"78030001", 15956 => x"38633d2c",
    15957 => x"29620000", 15958 => x"28610000", 15959 => x"a0410800",
    15960 => x"e0000002", 15961 => x"34010000", 15962 => x"2b9d0004",
    15963 => x"2b8b0008", 15964 => x"379c0008", 15965 => x"c3a00000",
    15966 => x"379cfff8", 15967 => x"5b8b0008", 15968 => x"5b9d0004",
    15969 => x"78030001", 15970 => x"b8405800", 15971 => x"38636b2c",
    15972 => x"44200007", 15973 => x"3421ffff", 15974 => x"08230090",
    15975 => x"78010001", 15976 => x"38216a78", 15977 => x"b4610800",
    15978 => x"34230144", 15979 => x"b8600800", 15980 => x"b9601000",
    15981 => x"fbffff04", 15982 => x"78010001", 15983 => x"38216a78",
    15984 => x"582b0014", 15985 => x"2b9d0004", 15986 => x"2b8b0008",
    15987 => x"379c0008", 15988 => x"c3a00000", 15989 => x"379cffec",
    15990 => x"5b8b0014", 15991 => x"5b8c0010", 15992 => x"5b8d000c",
    15993 => x"5b8e0008", 15994 => x"5b9d0004", 15995 => x"780c0001",
    15996 => x"780d0001", 15997 => x"b8207000", 15998 => x"340b0000",
    15999 => x"398c6db0", 16000 => x"39ad6cf4", 16001 => x"e000000a",
    16002 => x"29a10000", 16003 => x"942b0800", 16004 => x"20210001",
    16005 => x"44200005", 16006 => x"3d620005", 16007 => x"b5c21000",
    16008 => x"3441025c", 16009 => x"fbffff15", 16010 => x"356b0001",
    16011 => x"29810000", 16012 => x"482bfff6", 16013 => x"2b9d0004",
    16014 => x"2b8b0014", 16015 => x"2b8c0010", 16016 => x"2b8d000c",
    16017 => x"2b8e0008", 16018 => x"379c0014", 16019 => x"c3a00000",
    16020 => x"379cffb8", 16021 => x"5b8b0044", 16022 => x"5b8c0040",
    16023 => x"5b8d003c", 16024 => x"5b8e0038", 16025 => x"5b8f0034",
    16026 => x"5b900030", 16027 => x"5b91002c", 16028 => x"5b920028",
    16029 => x"5b930024", 16030 => x"5b940020", 16031 => x"5b95001c",
    16032 => x"5b960018", 16033 => x"5b970014", 16034 => x"5b980010",
    16035 => x"5b99000c", 16036 => x"5b9b0008", 16037 => x"5b9d0004",
    16038 => x"78010001", 16039 => x"78190001", 16040 => x"38213d5c",
    16041 => x"780b0001", 16042 => x"78180001", 16043 => x"780d0001",
    16044 => x"78110001", 16045 => x"78100001", 16046 => x"780c0001",
    16047 => x"78160001", 16048 => x"780f0001", 16049 => x"3b396d08",
    16050 => x"283b0000", 16051 => x"396b6a78", 16052 => x"34130009",
    16053 => x"3b184134", 16054 => x"34170001", 16055 => x"34120003",
    16056 => x"39ad6b0c", 16057 => x"3a316b2c", 16058 => x"3a106a90",
    16059 => x"398c6db0", 16060 => x"3ad66cd4", 16061 => x"39ef6da8",
    16062 => x"e000007b", 16063 => x"2861007c", 16064 => x"5b810048",
    16065 => x"2b8e0048", 16066 => x"2b940048", 16067 => x"29610004",
    16068 => x"01ce0018", 16069 => x"a29ba000", 16070 => x"3421ffff",
    16071 => x"21ce007f", 16072 => x"54330050", 16073 => x"3c210002",
    16074 => x"b7010800", 16075 => x"28210000", 16076 => x"c0200000",
    16077 => x"29610048", 16078 => x"58610040", 16079 => x"296100d0",
    16080 => x"296200cc", 16081 => x"b4410800", 16082 => x"0022001f",
    16083 => x"b4410800", 16084 => x"14210001", 16085 => x"34020001",
    16086 => x"58610044", 16087 => x"29810000", 16088 => x"fbfffb89",
    16089 => x"fbfff2ca", 16090 => x"34210032", 16091 => x"59610008",
    16092 => x"3401000a", 16093 => x"e0000011", 16094 => x"29750008",
    16095 => x"fbfff2c4", 16096 => x"caa10800", 16097 => x"4c200037",
    16098 => x"29610000", 16099 => x"5c370003", 16100 => x"59770004",
    16101 => x"e0000033", 16102 => x"59720004", 16103 => x"e0000031",
    16104 => x"29810000", 16105 => x"34020000", 16106 => x"fbfffb77",
    16107 => x"b9a00800", 16108 => x"fbfffc09", 16109 => x"34010002",
    16110 => x"59610004", 16111 => x"e0000029", 16112 => x"b9a00800",
    16113 => x"fbfffc1a", 16114 => x"e0000012", 16115 => x"ba000800",
    16116 => x"fbfffd74", 16117 => x"34010004", 16118 => x"e3fffff8",
    16119 => x"29610064", 16120 => x"44200020", 16121 => x"29610068",
    16122 => x"4420001e", 16123 => x"29610000", 16124 => x"5c320009",
    16125 => x"34010005", 16126 => x"e3fffff0", 16127 => x"ba200800",
    16128 => x"fbfffdb5", 16129 => x"34010006", 16130 => x"e3ffffec",
    16131 => x"296100ec", 16132 => x"44200014", 16133 => x"b9600800",
    16134 => x"fbffff6f", 16135 => x"34010008", 16136 => x"e3ffffe6",
    16137 => x"29610000", 16138 => x"5c370004", 16139 => x"b9a00800",
    16140 => x"fbfffbff", 16141 => x"44200007", 16142 => x"29610064",
    16143 => x"44200005", 16144 => x"29610000", 16145 => x"5c320007",
    16146 => x"296100ec", 16147 => x"5c200005", 16148 => x"29610010",
    16149 => x"34210001", 16150 => x"59610010", 16151 => x"59730004",
    16152 => x"ba000800", 16153 => x"ba801000", 16154 => x"b9c01800",
    16155 => x"fbfffcf6", 16156 => x"29610064", 16157 => x"4420001c",
    16158 => x"ba801000", 16159 => x"ba200800", 16160 => x"b9c01800",
    16161 => x"fbfffdca", 16162 => x"29620004", 16163 => x"34010008",
    16164 => x"5c410015", 16165 => x"29610000", 16166 => x"34150000",
    16167 => x"5c32000c", 16168 => x"e0000008", 16169 => x"0aa10090",
    16170 => x"ba801000", 16171 => x"b9c01800", 16172 => x"b5610800",
    16173 => x"34210144", 16174 => x"fbfffdbd", 16175 => x"36b50001",
    16176 => x"29e10000", 16177 => x"3421ffff", 16178 => x"4835fff7",
    16179 => x"29810000", 16180 => x"49c10005", 16181 => x"bac00800",
    16182 => x"ba801000", 16183 => x"b9c01800", 16184 => x"fbfffe78",
    16185 => x"2b230000", 16186 => x"78020002", 16187 => x"28610080",
    16188 => x"a0220800", 16189 => x"4420ff82", 16190 => x"78010001",
    16191 => x"38216a74", 16192 => x"28220000", 16193 => x"34420001",
    16194 => x"58220000", 16195 => x"34010001", 16196 => x"d0410000",
    16197 => x"2b9d0004", 16198 => x"2b8b0044", 16199 => x"2b8c0040",
    16200 => x"2b8d003c", 16201 => x"2b8e0038", 16202 => x"2b8f0034",
    16203 => x"2b900030", 16204 => x"2b91002c", 16205 => x"2b920028",
    16206 => x"2b930024", 16207 => x"2b940020", 16208 => x"2b95001c",
    16209 => x"2b960018", 16210 => x"2b970014", 16211 => x"2b980010",
    16212 => x"2b99000c", 16213 => x"2b9b0008", 16214 => x"379c0048",
    16215 => x"c3a00000", 16216 => x"78010001", 16217 => x"38216d10",
    16218 => x"28220000", 16219 => x"78030001", 16220 => x"78010001",
    16221 => x"38216d0c", 16222 => x"38633d78", 16223 => x"58220000",
    16224 => x"28610000", 16225 => x"58410000", 16226 => x"c3a00000",
    16227 => x"379cffd4", 16228 => x"5b8b0028", 16229 => x"5b8c0024",
    16230 => x"5b8d0020", 16231 => x"5b8e001c", 16232 => x"5b8f0018",
    16233 => x"5b900014", 16234 => x"5b910010", 16235 => x"5b92000c",
    16236 => x"5b930008", 16237 => x"5b9d0004", 16238 => x"b8205800",
    16239 => x"b8408000", 16240 => x"b8609000", 16241 => x"fbffc101",
    16242 => x"78010001", 16243 => x"38216dd4", 16244 => x"28240000",
    16245 => x"78010001", 16246 => x"38216d08", 16247 => x"58240000",
    16248 => x"78010001", 16249 => x"28860000", 16250 => x"38216d10",
    16251 => x"28220000", 16252 => x"78010001", 16253 => x"38216d0c",
    16254 => x"00c50010", 16255 => x"58220000", 16256 => x"78010001",
    16257 => x"38216db0", 16258 => x"20a5003f", 16259 => x"00c60018",
    16260 => x"58250000", 16261 => x"78010001", 16262 => x"38216da8",
    16263 => x"20c60007", 16264 => x"58260000", 16265 => x"78010001",
    16266 => x"38216a78", 16267 => x"582b0000", 16268 => x"58200010",
    16269 => x"58800040", 16270 => x"58800044", 16271 => x"58800000",
    16272 => x"58800028", 16273 => x"58800024", 16274 => x"58800004",
    16275 => x"58800020", 16276 => x"340303e8", 16277 => x"58830048",
    16278 => x"78040001", 16279 => x"38843d3c", 16280 => x"28830000",
    16281 => x"5840001c", 16282 => x"58430000", 16283 => x"34020004",
    16284 => x"5d620004", 16285 => x"34020007", 16286 => x"58220004",
    16287 => x"e0000006", 16288 => x"34020009", 16289 => x"58220004",
    16290 => x"34010003", 16291 => x"5d610002", 16292 => x"ba002800",
    16293 => x"78010001", 16294 => x"b8a01000", 16295 => x"38216a90",
    16296 => x"780d0001", 16297 => x"fbfffc55", 16298 => x"39ad6db0",
    16299 => x"29a30000", 16300 => x"78010001", 16301 => x"38216b2c",
    16302 => x"ba001000", 16303 => x"780f0001", 16304 => x"780e0001",
    16305 => x"fbfffcd6", 16306 => x"340c0000", 16307 => x"39ef6da8",
    16308 => x"39ce6a78", 16309 => x"34130001", 16310 => x"e000000c",
    16311 => x"09910090", 16312 => x"29a40000", 16313 => x"ba001000",
    16314 => x"b5d10800", 16315 => x"34840001", 16316 => x"b48c1800",
    16317 => x"34210144", 16318 => x"b5d18800", 16319 => x"fbfffcc8",
    16320 => x"358c0001", 16321 => x"5a33013c", 16322 => x"29e10000",
    16323 => x"3421ffff", 16324 => x"482cfff3", 16325 => x"34010002",
    16326 => x"5d610006", 16327 => x"78010001", 16328 => x"38216d0c",
    16329 => x"28210000", 16330 => x"34020006", 16331 => x"5822001c",
    16332 => x"780e0001", 16333 => x"780d0001", 16334 => x"340c0000",
    16335 => x"39ce6db0", 16336 => x"39ad6a78", 16337 => x"e0000008",
    16338 => x"3d810005", 16339 => x"b9801000", 16340 => x"b5a10800",
    16341 => x"3421025c", 16342 => x"34030200", 16343 => x"fbfffdc0",
    16344 => x"358c0001", 16345 => x"29c20000", 16346 => x"484cfff8",
    16347 => x"34010001", 16348 => x"5d61001d", 16349 => x"78010001",
    16350 => x"38216d08", 16351 => x"28210000", 16352 => x"28210004",
    16353 => x"20210002", 16354 => x"44200012", 16355 => x"78010001",
    16356 => x"78040001", 16357 => x"38216a78", 16358 => x"38846a90",
    16359 => x"58240094", 16360 => x"78040001", 16361 => x"38846b2c",
    16362 => x"58240098", 16363 => x"78010001", 16364 => x"38216da8",
    16365 => x"28240000", 16366 => x"78010001", 16367 => x"38216b0c",
    16368 => x"b4441000", 16369 => x"ba401800", 16370 => x"fbfffae7",
    16371 => x"e0000006", 16372 => x"78020001", 16373 => x"34010000",
    16374 => x"3842399c", 16375 => x"fbffc08e", 16376 => x"e0000020",
    16377 => x"78010001", 16378 => x"3d6b0002", 16379 => x"382141b4",
    16380 => x"78040001", 16381 => x"78050001", 16382 => x"b42b5800",
    16383 => x"38846db0", 16384 => x"38a56da8", 16385 => x"29630000",
    16386 => x"28840000", 16387 => x"28a50000", 16388 => x"78020001",
    16389 => x"34010000", 16390 => x"384239d8", 16391 => x"fbffc07e",
    16392 => x"78010001", 16393 => x"38216d08", 16394 => x"28210000",
    16395 => x"78020002", 16396 => x"e0000003", 16397 => x"2823007c",
    16398 => x"5b83002c", 16399 => x"28230080", 16400 => x"a0621800",
    16401 => x"4460fffc", 16402 => x"34020001", 16403 => x"58220064",
    16404 => x"28220028", 16405 => x"38420001", 16406 => x"58220028",
    16407 => x"fbffc064", 16408 => x"2b9d0004", 16409 => x"2b8b0028",
    16410 => x"2b8c0024", 16411 => x"2b8d0020", 16412 => x"2b8e001c",
    16413 => x"2b8f0018", 16414 => x"2b900014", 16415 => x"2b910010",
    16416 => x"2b92000c", 16417 => x"2b930008", 16418 => x"379c002c",
    16419 => x"c3a00000", 16420 => x"379cfffc", 16421 => x"5b9d0004",
    16422 => x"78020001", 16423 => x"38426a78", 16424 => x"b8201800",
    16425 => x"28410004", 16426 => x"64640000", 16427 => x"7c210008",
    16428 => x"b8810800", 16429 => x"44200006", 16430 => x"78020001",
    16431 => x"34010000", 16432 => x"38423a0c", 16433 => x"fbffc054",
    16434 => x"e0000006", 16435 => x"3463ffff", 16436 => x"08630090",
    16437 => x"b4431000", 16438 => x"34410144", 16439 => x"fbfffc7e",
    16440 => x"2b9d0004", 16441 => x"379c0004", 16442 => x"c3a00000",
    16443 => x"379cfffc", 16444 => x"5b9d0004", 16445 => x"44200008",
    16446 => x"3421ffff", 16447 => x"08210090", 16448 => x"78020001",
    16449 => x"38426a78", 16450 => x"b4220800", 16451 => x"34210144",
    16452 => x"fbfffc9b", 16453 => x"2b9d0004", 16454 => x"379c0004",
    16455 => x"c3a00000", 16456 => x"78020001", 16457 => x"b8201800",
    16458 => x"38426a78", 16459 => x"5c200004", 16460 => x"28410004",
    16461 => x"64210008", 16462 => x"c3a00000", 16463 => x"28450004",
    16464 => x"34040008", 16465 => x"34010000", 16466 => x"5ca40006",
    16467 => x"3463ffff", 16468 => x"08630090", 16469 => x"b4431000",
    16470 => x"2841017c", 16471 => x"7c210000", 16472 => x"c3a00000",
    16473 => x"379cffe8", 16474 => x"5b8b0018", 16475 => x"5b8c0014",
    16476 => x"5b8d0010", 16477 => x"5b8e000c", 16478 => x"5b8f0008",
    16479 => x"5b9d0004", 16480 => x"3403ffff", 16481 => x"b8407800",
    16482 => x"5c230016", 16483 => x"34010000", 16484 => x"780c0001",
    16485 => x"780d0001", 16486 => x"fbfffff3", 16487 => x"340b0000",
    16488 => x"398c6da8", 16489 => x"39ad6a78", 16490 => x"340e0004",
    16491 => x"e0000009", 16492 => x"09610090", 16493 => x"b5a10800",
    16494 => x"2821013c", 16495 => x"5c2e0004", 16496 => x"35610001",
    16497 => x"b9e01000", 16498 => x"fbfffdec", 16499 => x"356b0001",
    16500 => x"29810000", 16501 => x"3421ffff", 16502 => x"482bfff6",
    16503 => x"e0000002", 16504 => x"fbfffde6", 16505 => x"2b9d0004",
    16506 => x"2b8b0018", 16507 => x"2b8c0014", 16508 => x"2b8d0010",
    16509 => x"2b8e000c", 16510 => x"2b8f0008", 16511 => x"379c0018",
    16512 => x"c3a00000", 16513 => x"379cfff0", 16514 => x"5b8b0010",
    16515 => x"5b8c000c", 16516 => x"5b8d0008", 16517 => x"5b9d0004",
    16518 => x"780b0001", 16519 => x"b8406800", 16520 => x"b8606000",
    16521 => x"396b6b2c", 16522 => x"44200007", 16523 => x"3421ffff",
    16524 => x"082b0090", 16525 => x"78010001", 16526 => x"38216a78",
    16527 => x"b5610800", 16528 => x"342b0144", 16529 => x"45a0000b",
    16530 => x"2962006c", 16531 => x"34041f40", 16532 => x"34030000",
    16533 => x"3c420001", 16534 => x"1441001f", 16535 => x"f80002e6",
    16536 => x"3c210012", 16537 => x"0044000e", 16538 => x"b8242000",
    16539 => x"59a40000", 16540 => x"4580000b", 16541 => x"29620068",
    16542 => x"34030000", 16543 => x"34041f40", 16544 => x"3c420001",
    16545 => x"1441001f", 16546 => x"f80002db", 16547 => x"3c210012",
    16548 => x"0042000e", 16549 => x"b8221000", 16550 => x"59820000",
    16551 => x"2b9d0004", 16552 => x"2b8b0010", 16553 => x"2b8c000c",
    16554 => x"2b8d0008", 16555 => x"379c0010", 16556 => x"c3a00000",
    16557 => x"379cfff0", 16558 => x"5b8b0010", 16559 => x"5b8c000c",
    16560 => x"5b8d0008", 16561 => x"5b9d0004", 16562 => x"b8205800",
    16563 => x"b8406800", 16564 => x"78010001", 16565 => x"3d620005",
    16566 => x"38216a78", 16567 => x"b4220800", 16568 => x"28240274",
    16569 => x"b8606000", 16570 => x"4c800003", 16571 => x"34844000",
    16572 => x"e0000004", 16573 => x"34013fff", 16574 => x"4c240002",
    16575 => x"3484c000", 16576 => x"3c840001", 16577 => x"34010000",
    16578 => x"20823ffe", 16579 => x"34030000", 16580 => x"34041f40",
    16581 => x"f80002b8", 16582 => x"3c210012", 16583 => x"0044000e",
    16584 => x"b8242000", 16585 => x"59a40000", 16586 => x"4580000c",
    16587 => x"78010001", 16588 => x"38216cf4", 16589 => x"28220000",
    16590 => x"3d630005", 16591 => x"78010001", 16592 => x"38216a78",
    16593 => x"b4230800", 16594 => x"28210260", 16595 => x"94410800",
    16596 => x"20210001", 16597 => x"59810000", 16598 => x"3d6b0005",
    16599 => x"78020001", 16600 => x"38426a78", 16601 => x"b44b1000",
    16602 => x"28410278", 16603 => x"2b9d0004", 16604 => x"2b8b0010",
    16605 => x"2b8c000c", 16606 => x"2b8d0008", 16607 => x"379c0010",
    16608 => x"c3a00000", 16609 => x"379cffec", 16610 => x"5b8b0014",
    16611 => x"5b8c0010", 16612 => x"5b9d000c", 16613 => x"780b0001",
    16614 => x"396b6a78", 16615 => x"29610000", 16616 => x"4c010016",
    16617 => x"78010001", 16618 => x"38216a74", 16619 => x"282c0000",
    16620 => x"29620004", 16621 => x"78010001", 16622 => x"3821415c",
    16623 => x"fbfff9cb", 16624 => x"29640000", 16625 => x"b8201800",
    16626 => x"296500a0", 16627 => x"29660064", 16628 => x"296700ec",
    16629 => x"29680050", 16630 => x"296200d8", 16631 => x"29610010",
    16632 => x"5b820004", 16633 => x"5b810008", 16634 => x"78010001",
    16635 => x"38213a3c", 16636 => x"b9801000", 16637 => x"fbffea74",
    16638 => x"2b9d000c", 16639 => x"2b8b0014", 16640 => x"2b8c0010",
    16641 => x"379c0014", 16642 => x"c3a00000", 16643 => x"379cfffc",
    16644 => x"5b9d0004", 16645 => x"5c200004", 16646 => x"78010001",
    16647 => x"38216b2c", 16648 => x"e0000007", 16649 => x"3421ffff",
    16650 => x"08210090", 16651 => x"78020001", 16652 => x"38426a78",
    16653 => x"b4220800", 16654 => x"34210144", 16655 => x"fbfffc84",
    16656 => x"2b9d0004", 16657 => x"379c0004", 16658 => x"c3a00000",
    16659 => x"379cfff0", 16660 => x"5b8b0010", 16661 => x"5b8c000c",
    16662 => x"5b8d0008", 16663 => x"5b9d0004", 16664 => x"780d0001",
    16665 => x"780c0001", 16666 => x"b8205800", 16667 => x"39ad6a78",
    16668 => x"398c6cf4", 16669 => x"44400010", 16670 => x"34020001",
    16671 => x"fbfff942", 16672 => x"3d610005", 16673 => x"b5a16800",
    16674 => x"35a1025c", 16675 => x"fbfffc7b", 16676 => x"29820000",
    16677 => x"34010001", 16678 => x"bc2b0800", 16679 => x"b8220800",
    16680 => x"78020001", 16681 => x"59810000", 16682 => x"38423a90",
    16683 => x"34010000", 16684 => x"e000000d", 16685 => x"34030001",
    16686 => x"29840000", 16687 => x"bc611800", 16688 => x"a4601800",
    16689 => x"a0641800", 16690 => x"59830000", 16691 => x"29a30124",
    16692 => x"44230002", 16693 => x"fbfff92c", 16694 => x"78020001",
    16695 => x"34010000", 16696 => x"38423ab0", 16697 => x"b9601800",
    16698 => x"fbffbf4b", 16699 => x"2b9d0004", 16700 => x"2b8b0010",
    16701 => x"2b8c000c", 16702 => x"2b8d0008", 16703 => x"379c0010",
    16704 => x"c3a00000", 16705 => x"08210090", 16706 => x"78020001",
    16707 => x"38426a78", 16708 => x"b4411000", 16709 => x"2841013c",
    16710 => x"2843013c", 16711 => x"34020004", 16712 => x"7c210001",
    16713 => x"5c620002", 16714 => x"38210002", 16715 => x"c3a00000",
    16716 => x"4c200005", 16717 => x"78010001", 16718 => x"38216a78",
    16719 => x"28210050", 16720 => x"c3a00000", 16721 => x"78020001",
    16722 => x"38426a78", 16723 => x"5c200003", 16724 => x"284100d8",
    16725 => x"c3a00000", 16726 => x"3421ffff", 16727 => x"08210090",
    16728 => x"b4411000", 16729 => x"28410168", 16730 => x"c3a00000",
    16731 => x"78030001", 16732 => x"38636d08", 16733 => x"4c200007",
    16734 => x"78010001", 16735 => x"38216a78", 16736 => x"58220050",
    16737 => x"28610000", 16738 => x"58220040", 16739 => x"c3a00000",
    16740 => x"2024000f", 16741 => x"28630000", 16742 => x"3c840010",
    16743 => x"2045ffff", 16744 => x"b8a42000", 16745 => x"58640044",
    16746 => x"78030001", 16747 => x"38636a78", 16748 => x"5c200003",
    16749 => x"586200d8", 16750 => x"c3a00000", 16751 => x"3421ffff",
    16752 => x"08210090", 16753 => x"b4611800", 16754 => x"58620168",
    16755 => x"c3a00000", 16756 => x"379cffc0", 16757 => x"5b8b0040",
    16758 => x"5b8c003c", 16759 => x"5b8d0038", 16760 => x"5b8e0034",
    16761 => x"5b8f0030", 16762 => x"5b90002c", 16763 => x"5b910028",
    16764 => x"5b920024", 16765 => x"5b930020", 16766 => x"5b94001c",
    16767 => x"5b950018", 16768 => x"5b960014", 16769 => x"5b970010",
    16770 => x"5b98000c", 16771 => x"5b990008", 16772 => x"5b9d0004",
    16773 => x"78010001", 16774 => x"38216a78", 16775 => x"28220000",
    16776 => x"34010001", 16777 => x"5c410004", 16778 => x"78010001",
    16779 => x"38216b0c", 16780 => x"fbfff99a", 16781 => x"78100001",
    16782 => x"780c0001", 16783 => x"780d0001", 16784 => x"78160001",
    16785 => x"78140001", 16786 => x"78130001", 16787 => x"78120001",
    16788 => x"78110001", 16789 => x"340b0001", 16790 => x"3a106da8",
    16791 => x"398c6a78", 16792 => x"340e0001", 16793 => x"39ad6d08",
    16794 => x"3ad63ae4", 16795 => x"34150002", 16796 => x"3a943b2c",
    16797 => x"34190003", 16798 => x"3a733b5c", 16799 => x"34180004",
    16800 => x"3a523b80", 16801 => x"3a313b08", 16802 => x"e0000058",
    16803 => x"3577ffff", 16804 => x"0aef0090", 16805 => x"b58f7800",
    16806 => x"29e1013c", 16807 => x"442e0011", 16808 => x"29a10000",
    16809 => x"bdcb1000", 16810 => x"28210020", 16811 => x"00210008",
    16812 => x"202100ff", 16813 => x"a0220800", 16814 => x"5c20000a",
    16815 => x"bac01000", 16816 => x"b9601800", 16817 => x"fbffbed4",
    16818 => x"b9600800", 16819 => x"fbfffe88", 16820 => x"b9600800",
    16821 => x"34020000", 16822 => x"fbfffc3f", 16823 => x"59ee013c",
    16824 => x"0ae10090", 16825 => x"b5817800", 16826 => x"29e3013c",
    16827 => x"44750018", 16828 => x"48750003", 16829 => x"5c6e003c",
    16830 => x"e0000004", 16831 => x"44790020", 16832 => x"5c780039",
    16833 => x"e000002a", 16834 => x"298100ec", 16835 => x"44200036",
    16836 => x"29a10000", 16837 => x"bdcb1000", 16838 => x"28210020",
    16839 => x"00210008", 16840 => x"202100ff", 16841 => x"a0220800",
    16842 => x"4420002f", 16843 => x"34010000", 16844 => x"ba201000",
    16845 => x"b9601800", 16846 => x"fbffbeb7", 16847 => x"b9600800",
    16848 => x"fbfffe54", 16849 => x"59f5013c", 16850 => x"e0000027",
    16851 => x"29e1017c", 16852 => x"44200025", 16853 => x"29840014",
    16854 => x"34010000", 16855 => x"ba801000", 16856 => x"b9601800",
    16857 => x"fbffbeac", 16858 => x"29820014", 16859 => x"b9600800",
    16860 => x"fbfffc82", 16861 => x"59f9013c", 16862 => x"e000001b",
    16863 => x"b5810800", 16864 => x"34210144", 16865 => x"fbfffbb2",
    16866 => x"5c200017", 16867 => x"ba601000", 16868 => x"b9601800",
    16869 => x"fbffbea0", 16870 => x"b9600800", 16871 => x"34020001",
    16872 => x"fbfffc0d", 16873 => x"59f8013c", 16874 => x"e000000f",
    16875 => x"298100ec", 16876 => x"44200003", 16877 => x"29e1017c",
    16878 => x"5c20000b", 16879 => x"0af70090", 16880 => x"34010000",
    16881 => x"ba401000", 16882 => x"b9601800", 16883 => x"fbffbe92",
    16884 => x"b9600800", 16885 => x"34020000", 16886 => x"b597b800",
    16887 => x"fbfffbfe", 16888 => x"5aee013c", 16889 => x"356b0001",
    16890 => x"2a010000", 16891 => x"482bffa8", 16892 => x"2b9d0004",
    16893 => x"2b8b0040", 16894 => x"2b8c003c", 16895 => x"2b8d0038",
    16896 => x"2b8e0034", 16897 => x"2b8f0030", 16898 => x"2b90002c",
    16899 => x"2b910028", 16900 => x"2b920024", 16901 => x"2b930020",
    16902 => x"2b94001c", 16903 => x"2b950018", 16904 => x"2b960014",
    16905 => x"2b970010", 16906 => x"2b98000c", 16907 => x"2b990008",
    16908 => x"379c0040", 16909 => x"c3a00000", 16910 => x"379cfff0",
    16911 => x"5b8b0010", 16912 => x"5b8c000c", 16913 => x"5b8d0008",
    16914 => x"5b9d0004", 16915 => x"fbffbe5f", 16916 => x"78020001",
    16917 => x"34010000", 16918 => x"38423bac", 16919 => x"fbffbe6e",
    16920 => x"34020000", 16921 => x"3401ffff", 16922 => x"fbffff41",
    16923 => x"34010001", 16924 => x"fbfffc1f", 16925 => x"380bffff",
    16926 => x"b8206800", 16927 => x"b9601000", 16928 => x"3401ffff",
    16929 => x"fbffff3a", 16930 => x"34010001", 16931 => x"fbfffc18",
    16932 => x"78040001", 16933 => x"38843d7c", 16934 => x"28830000",
    16935 => x"b8206000", 16936 => x"b9801000", 16937 => x"b9a00800",
    16938 => x"fbfffbe0", 16939 => x"78020001", 16940 => x"b8202800",
    16941 => x"b9a01800", 16942 => x"b9802000", 16943 => x"34010000",
    16944 => x"38423bd0", 16945 => x"fbffbe54", 16946 => x"34020000",
    16947 => x"34010000", 16948 => x"fbffff27", 16949 => x"34010000",
    16950 => x"fbfffc05", 16951 => x"b8206000", 16952 => x"b9601000",
    16953 => x"34010000", 16954 => x"fbffff21", 16955 => x"34010000",
    16956 => x"fbfffbff", 16957 => x"78040001", 16958 => x"38843d80",
    16959 => x"28830000", 16960 => x"b8205800", 16961 => x"b9601000",
    16962 => x"b9800800", 16963 => x"fbfffbc7", 16964 => x"78020001",
    16965 => x"b8202800", 16966 => x"b9801800", 16967 => x"b9602000",
    16968 => x"38423c00", 16969 => x"34010000", 16970 => x"fbffbe3b",
    16971 => x"34010002", 16972 => x"fbfffbef", 16973 => x"78020001",
    16974 => x"b8201800", 16975 => x"38423c30", 16976 => x"34010000",
    16977 => x"fbffbe34", 16978 => x"2b9d0004", 16979 => x"2b8b0010",
    16980 => x"2b8c000c", 16981 => x"2b8d0008", 16982 => x"379c0010",
    16983 => x"c3a00000", 16984 => x"379cfff0", 16985 => x"5b8b0010",
    16986 => x"5b8c000c", 16987 => x"5b8d0008", 16988 => x"5b9d0004",
    16989 => x"78010001", 16990 => x"780b0001", 16991 => x"38213cd8",
    16992 => x"780c0001", 16993 => x"396bf800", 16994 => x"282d0000",
    16995 => x"398c3cc4", 16996 => x"e0000005", 16997 => x"b9800800",
    16998 => x"fbffe90b", 16999 => x"340103e8", 17000 => x"fbffef40",
    17001 => x"29610000", 17002 => x"5c2dfffb", 17003 => x"2b9d0004",
    17004 => x"2b8b0010", 17005 => x"2b8c000c", 17006 => x"2b8d0008",
    17007 => x"379c0010", 17008 => x"c3a00000", 17009 => x"c3a00000",
    17010 => x"379cfff8", 17011 => x"5b8b0008", 17012 => x"5b9d0004",
    17013 => x"28240014", 17014 => x"b8201800", 17015 => x"b8403000",
    17016 => x"44800015", 17017 => x"28250010", 17018 => x"20a50002",
    17019 => x"5ca00007", 17020 => x"b4862000", 17021 => x"b8800800",
    17022 => x"2b9d0004", 17023 => x"2b8b0008", 17024 => x"379c0008",
    17025 => x"c3a00000", 17026 => x"346b0030", 17027 => x"b4861000",
    17028 => x"b9600800", 17029 => x"34030040", 17030 => x"f80001cc",
    17031 => x"b9602000", 17032 => x"b8800800", 17033 => x"2b9d0004",
    17034 => x"2b8b0008", 17035 => x"379c0008", 17036 => x"c3a00000",
    17037 => x"28250010", 17038 => x"20a70004", 17039 => x"5ce4ffeb",
    17040 => x"2825001c", 17041 => x"34040000", 17042 => x"44a7ffeb",
    17043 => x"342b0030", 17044 => x"34040040", 17045 => x"b9601800",
    17046 => x"d8a00000", 17047 => x"b9602000", 17048 => x"e3fffff0",
    17049 => x"379cfff4", 17050 => x"5b8b0008", 17051 => x"5b9d0004",
    17052 => x"28220014", 17053 => x"b8205800", 17054 => x"44400013",
    17055 => x"2961000c", 17056 => x"b4411000", 17057 => x"28430000",
    17058 => x"78040001", 17059 => x"38843d84", 17060 => x"28820000",
    17061 => x"3401ffec", 17062 => x"5c620007", 17063 => x"78020001",
    17064 => x"38426cf8", 17065 => x"28430000", 17066 => x"34010000",
    17067 => x"584b0000", 17068 => x"5963007c", 17069 => x"2b9d0004",
    17070 => x"2b8b0008", 17071 => x"379c000c", 17072 => x"c3a00000",
    17073 => x"28230010", 17074 => x"20630004", 17075 => x"5c62ffec",
    17076 => x"2825001c", 17077 => x"2822000c", 17078 => x"3783000c",
    17079 => x"34040004", 17080 => x"d8a00000", 17081 => x"2b83000c",
    17082 => x"e3ffffe8", 17083 => x"379cfff0", 17084 => x"5b8b0010",
    17085 => x"5b8c000c", 17086 => x"5b8d0008", 17087 => x"5b9d0004",
    17088 => x"b8205800", 17089 => x"44400047", 17090 => x"2822000c",
    17091 => x"58200080", 17092 => x"582000b0", 17093 => x"58220090",
    17094 => x"340c0000", 17095 => x"b9600800", 17096 => x"fbffffaa",
    17097 => x"59610028", 17098 => x"4022003f", 17099 => x"5c400006",
    17100 => x"78040001", 17101 => x"38843d84", 17102 => x"28230000",
    17103 => x"28820000", 17104 => x"4462005d", 17105 => x"34010000",
    17106 => x"45800030", 17107 => x"3583ffff", 17108 => x"346c0028",
    17109 => x"b58c0800", 17110 => x"b4210800", 17111 => x"b5610800",
    17112 => x"28220000", 17113 => x"5c40000f", 17114 => x"34010000",
    17115 => x"44620027", 17116 => x"34620027", 17117 => x"b4421000",
    17118 => x"b4421000", 17119 => x"b5621000", 17120 => x"e0000002",
    17121 => x"44610044", 17122 => x"28410000", 17123 => x"3463ffff",
    17124 => x"3442fffc", 17125 => x"4420fffc", 17126 => x"596300b0",
    17127 => x"346c0028", 17128 => x"346d0024", 17129 => x"b5ad6800",
    17130 => x"b5ad6800", 17131 => x"b56d6800", 17132 => x"29a20000",
    17133 => x"b9600800", 17134 => x"b58c6000", 17135 => x"fbffff83",
    17136 => x"b58c6000", 17137 => x"b56c1000", 17138 => x"29a40000",
    17139 => x"28430000", 17140 => x"296c00b0", 17141 => x"34840040",
    17142 => x"3463ffff", 17143 => x"59610028", 17144 => x"59a40000",
    17145 => x"58430000", 17146 => x"35830020", 17147 => x"b4631800",
    17148 => x"b4631800", 17149 => x"b5631800", 17150 => x"2824000c",
    17151 => x"28620000", 17152 => x"b4441000", 17153 => x"59620074",
    17154 => x"2b9d0004", 17155 => x"2b8b0010", 17156 => x"2b8c000c",
    17157 => x"2b8d0008", 17158 => x"379c0010", 17159 => x"c3a00000",
    17160 => x"28210028", 17161 => x"296300b0", 17162 => x"34050002",
    17163 => x"4024003f", 17164 => x"eca32800", 17165 => x"64840002",
    17166 => x"a0852000", 17167 => x"4482ffc5", 17168 => x"34620020",
    17169 => x"b4421000", 17170 => x"b4421000", 17171 => x"b5621000",
    17172 => x"28450000", 17173 => x"34640025", 17174 => x"28220004",
    17175 => x"b4842000", 17176 => x"b4842000", 17177 => x"b4a21000",
    17178 => x"b5642000", 17179 => x"58820000", 17180 => x"2824000c",
    17181 => x"34610021", 17182 => x"b4210800", 17183 => x"b4210800",
    17184 => x"b5610800", 17185 => x"b4852800", 17186 => x"346c0001",
    17187 => x"58250000", 17188 => x"e3ffffa3", 17189 => x"34010000",
    17190 => x"596000b0", 17191 => x"2b9d0004", 17192 => x"2b8b0010",
    17193 => x"2b8c000c", 17194 => x"2b8d0008", 17195 => x"379c0010",
    17196 => x"c3a00000", 17197 => x"35820024", 17198 => x"b4421000",
    17199 => x"b4421000", 17200 => x"b5621800", 17201 => x"2c250004",
    17202 => x"28640000", 17203 => x"35820028", 17204 => x"b4421000",
    17205 => x"b4421000", 17206 => x"b5621000", 17207 => x"34a5ffff",
    17208 => x"34840040", 17209 => x"58450000", 17210 => x"58640000",
    17211 => x"596c00b0", 17212 => x"e3ffffbe", 17213 => x"379cffec",
    17214 => x"5b8b0014", 17215 => x"5b8c0010", 17216 => x"5b8d000c",
    17217 => x"5b8e0008", 17218 => x"5b9d0004", 17219 => x"b8406000",
    17220 => x"34020001", 17221 => x"b8205800", 17222 => x"b8607000",
    17223 => x"b8806800", 17224 => x"fbffff73", 17225 => x"b9600800",
    17226 => x"34020000", 17227 => x"fbffff70", 17228 => x"b8202800",
    17229 => x"4420001e", 17230 => x"28a10018", 17231 => x"5c2cfffa",
    17232 => x"28a1001c", 17233 => x"5c2efff8", 17234 => x"28a10020",
    17235 => x"5c2dfff6", 17236 => x"296100b0", 17237 => x"59650028",
    17238 => x"28a2000c", 17239 => x"34210020", 17240 => x"b4210800",
    17241 => x"b4210800", 17242 => x"b5610800", 17243 => x"28230000",
    17244 => x"34010000", 17245 => x"b4431800", 17246 => x"59630074",
    17247 => x"28a30014", 17248 => x"59600078", 17249 => x"34630001",
    17250 => x"c8621000", 17251 => x"59620070", 17252 => x"2b9d0004",
    17253 => x"2b8b0014", 17254 => x"2b8c0010", 17255 => x"2b8d000c",
    17256 => x"2b8e0008", 17257 => x"379c0014", 17258 => x"c3a00000",
    17259 => x"3401fffe", 17260 => x"e3fffff8", 17261 => x"379cfff8",
    17262 => x"5b8b0008", 17263 => x"5b9d0004", 17264 => x"b8205800",
    17265 => x"fbffffcc", 17266 => x"4c200005", 17267 => x"2b9d0004",
    17268 => x"2b8b0008", 17269 => x"379c0008", 17270 => x"c3a00000",
    17271 => x"29610074", 17272 => x"59600028", 17273 => x"2b9d0004",
    17274 => x"2b8b0008", 17275 => x"379c0008", 17276 => x"c3a00000",
    17277 => x"2045ffff", 17278 => x"00460010", 17279 => x"2088ffff",
    17280 => x"00890010", 17281 => x"89053800", 17282 => x"89064000",
    17283 => x"89252800", 17284 => x"00ea0010", 17285 => x"89263000",
    17286 => x"b5052800", 17287 => x"b4aa2800", 17288 => x"50a80003",
    17289 => x"78080001", 17290 => x"b4c83000", 17291 => x"88431000",
    17292 => x"88812000", 17293 => x"00a10010", 17294 => x"3ca50010",
    17295 => x"b4c13000", 17296 => x"20e7ffff", 17297 => x"b4440800",
    17298 => x"b4260800", 17299 => x"b4a71000", 17300 => x"c3a00000",
    17301 => x"44600008", 17302 => x"34040020", 17303 => x"c8832000",
    17304 => x"48800006", 17305 => x"c8041000", 17306 => x"34030000",
    17307 => x"80221000", 17308 => x"b8600800", 17309 => x"c3a00000",
    17310 => x"bc242000", 17311 => x"80431000", 17312 => x"80231800",
    17313 => x"b8821000", 17314 => x"b8600800", 17315 => x"e3fffffa",
    17316 => x"379cfff8", 17317 => x"5b8b0008", 17318 => x"5b9d0004",
    17319 => x"44400022", 17320 => x"b8412000", 17321 => x"3403000f",
    17322 => x"5483000b", 17323 => x"78030001", 17324 => x"386341c8",
    17325 => x"3c210004", 17326 => x"b4621000", 17327 => x"b4410800",
    17328 => x"40210000", 17329 => x"2b9d0004", 17330 => x"2b8b0008",
    17331 => x"379c0008", 17332 => x"c3a00000", 17333 => x"340b0000",
    17334 => x"4c200003", 17335 => x"c8010800", 17336 => x"340b0001",
    17337 => x"4c400003", 17338 => x"c8021000", 17339 => x"196b0001",
    17340 => x"90c01800", 17341 => x"20630002", 17342 => x"44600008",
    17343 => x"8c220800", 17344 => x"45600002", 17345 => x"c8010800",
    17346 => x"2b9d0004", 17347 => x"2b8b0008", 17348 => x"379c0008",
    17349 => x"c3a00000", 17350 => x"34030000", 17351 => x"f800004a",
    17352 => x"e3fffff8", 17353 => x"90000800", 17354 => x"20210001",
    17355 => x"3c210001", 17356 => x"d0010000", 17357 => x"90e00800",
    17358 => x"bba0f000", 17359 => x"342100a0", 17360 => x"c0200000",
    17361 => x"379cfff8", 17362 => x"5b8b0008", 17363 => x"5b9d0004",
    17364 => x"44400015", 17365 => x"340b0000", 17366 => x"4c200003",
    17367 => x"c8010800", 17368 => x"340b0001", 17369 => x"1443001f",
    17370 => x"90c02000", 17371 => x"98621000", 17372 => x"20840002",
    17373 => x"c8431000", 17374 => x"44800008", 17375 => x"c4220800",
    17376 => x"45600002", 17377 => x"c8010800", 17378 => x"2b9d0004",
    17379 => x"2b8b0008", 17380 => x"379c0008", 17381 => x"c3a00000",
    17382 => x"34030001", 17383 => x"f800002a", 17384 => x"e3fffff8",
    17385 => x"90000800", 17386 => x"20210001", 17387 => x"3c210001",
    17388 => x"d0010000", 17389 => x"90e00800", 17390 => x"bba0f000",
    17391 => x"342100a0", 17392 => x"c0200000", 17393 => x"379cfffc",
    17394 => x"5b9d0004", 17395 => x"44400006", 17396 => x"34030000",
    17397 => x"f800001c", 17398 => x"2b9d0004", 17399 => x"379c0004",
    17400 => x"c3a00000", 17401 => x"90000800", 17402 => x"20210001",
    17403 => x"3c210001", 17404 => x"d0010000", 17405 => x"90e00800",
    17406 => x"bba0f000", 17407 => x"342100a0", 17408 => x"c0200000",
    17409 => x"379cfffc", 17410 => x"5b9d0004", 17411 => x"44400006",
    17412 => x"34030001", 17413 => x"f800000c", 17414 => x"2b9d0004",
    17415 => x"379c0004", 17416 => x"c3a00000", 17417 => x"90000800",
    17418 => x"20210001", 17419 => x"3c210001", 17420 => x"d0010000",
    17421 => x"90e00800", 17422 => x"bba0f000", 17423 => x"342100a0",
    17424 => x"c0200000", 17425 => x"f4222000", 17426 => x"44800018",
    17427 => x"34040001", 17428 => x"4c40000b", 17429 => x"34050000",
    17430 => x"54410003", 17431 => x"c8220800", 17432 => x"b8a42800",
    17433 => x"00840001", 17434 => x"00420001", 17435 => x"5c80fffb",
    17436 => x"5c600002", 17437 => x"b8a00800", 17438 => x"c3a00000",
    17439 => x"3c420001", 17440 => x"3c840001", 17441 => x"f4222800",
    17442 => x"7c860000", 17443 => x"a0c52800", 17444 => x"44a00002",
    17445 => x"4c40fffa", 17446 => x"34050000", 17447 => x"4480fff5",
    17448 => x"34050000", 17449 => x"e3ffffed", 17450 => x"34040001",
    17451 => x"34050000", 17452 => x"e3ffffea", 17453 => x"1422001f",
    17454 => x"98410800", 17455 => x"c8220800", 17456 => x"c3a00000",
    17457 => x"34060003", 17458 => x"b8202000", 17459 => x"b8402800",
    17460 => x"50c3000c", 17461 => x"b8413000", 17462 => x"20c60003",
    17463 => x"5cc0000b", 17464 => x"34010003", 17465 => x"28860000",
    17466 => x"28a20000", 17467 => x"5cc20005", 17468 => x"3463fffc",
    17469 => x"34840004", 17470 => x"34a50004", 17471 => x"5461fffa",
    17472 => x"34010000", 17473 => x"4460000e", 17474 => x"40860000",
    17475 => x"40a10000", 17476 => x"3462ffff", 17477 => x"44c10006",
    17478 => x"e000000a", 17479 => x"40860000", 17480 => x"40a10000",
    17481 => x"3442ffff", 17482 => x"5cc10006", 17483 => x"34840001",
    17484 => x"34a50001", 17485 => x"5c40fffa", 17486 => x"34010000",
    17487 => x"c3a00000", 17488 => x"c8c10800", 17489 => x"c3a00000",
    17490 => x"3404000f", 17491 => x"b8203800", 17492 => x"b8403000",
    17493 => x"5083002d", 17494 => x"b8412000", 17495 => x"20840003",
    17496 => x"5c80002b", 17497 => x"b8402000", 17498 => x"b8202800",
    17499 => x"b8603000", 17500 => x"3407000f", 17501 => x"28880000",
    17502 => x"34c6fff0", 17503 => x"58a80000", 17504 => x"28880004",
    17505 => x"58a80004", 17506 => x"28880008", 17507 => x"58a80008",
    17508 => x"2888000c", 17509 => x"34840010", 17510 => x"58a8000c",
    17511 => x"34a50010", 17512 => x"54c7fff5", 17513 => x"3463fff0",
    17514 => x"00660004", 17515 => x"2063000f", 17516 => x"34c60001",
    17517 => x"3cc60004", 17518 => x"b4263800", 17519 => x"b4463000",
    17520 => x"34020003", 17521 => x"50430011", 17522 => x"34020000",
    17523 => x"34080003", 17524 => x"b4c22000", 17525 => x"28850000",
    17526 => x"b4e22000", 17527 => x"34420004", 17528 => x"58850000",
    17529 => x"c8622000", 17530 => x"5488fffa", 17531 => x"3463fffc",
    17532 => x"00620002", 17533 => x"20630003", 17534 => x"34420001",
    17535 => x"3c420002", 17536 => x"b4e23800", 17537 => x"b4c23000",
    17538 => x"44600008", 17539 => x"34020000", 17540 => x"b4c22000",
    17541 => x"40850000", 17542 => x"b4e22000", 17543 => x"34420001",
    17544 => x"30850000", 17545 => x"5c43fffb", 17546 => x"c3a00000",
    17547 => x"b8203800", 17548 => x"b8403000", 17549 => x"5041000c",
    17550 => x"b4432000", 17551 => x"5024000a", 17552 => x"4460003f",
    17553 => x"b4231000", 17554 => x"3484ffff", 17555 => x"40850000",
    17556 => x"3442ffff", 17557 => x"3463ffff", 17558 => x"30450000",
    17559 => x"5c60fffb", 17560 => x"c3a00000", 17561 => x"3404000f",
    17562 => x"5083002d", 17563 => x"b8412000", 17564 => x"20840003",
    17565 => x"5c80002b", 17566 => x"b8402000", 17567 => x"b8202800",
    17568 => x"b8603000", 17569 => x"3407000f", 17570 => x"28880000",
    17571 => x"34c6fff0", 17572 => x"58a80000", 17573 => x"28880004",
    17574 => x"58a80004", 17575 => x"28880008", 17576 => x"58a80008",
    17577 => x"2888000c", 17578 => x"34840010", 17579 => x"58a8000c",
    17580 => x"34a50010", 17581 => x"54c7fff5", 17582 => x"3463fff0",
    17583 => x"00660004", 17584 => x"2063000f", 17585 => x"34c60001",
    17586 => x"3cc60004", 17587 => x"b4263800", 17588 => x"b4463000",
    17589 => x"34020003", 17590 => x"50430011", 17591 => x"34020000",
    17592 => x"34080003", 17593 => x"b4c22000", 17594 => x"28850000",
    17595 => x"b4e22000", 17596 => x"34420004", 17597 => x"58850000",
    17598 => x"c8622000", 17599 => x"5488fffa", 17600 => x"3463fffc",
    17601 => x"00620002", 17602 => x"20630003", 17603 => x"34420001",
    17604 => x"3c420002", 17605 => x"b4e23800", 17606 => x"b4c23000",
    17607 => x"44600008", 17608 => x"34020000", 17609 => x"b4c22000",
    17610 => x"40850000", 17611 => x"b4e22000", 17612 => x"34420001",
    17613 => x"30850000", 17614 => x"5c43fffb", 17615 => x"c3a00000",
    17616 => x"20250003", 17617 => x"b8202000", 17618 => x"44a0000b",
    17619 => x"4460002c", 17620 => x"3463ffff", 17621 => x"204600ff",
    17622 => x"e0000003", 17623 => x"44600028", 17624 => x"3463ffff",
    17625 => x"30860000", 17626 => x"34840001", 17627 => x"20850003",
    17628 => x"5ca0fffb", 17629 => x"34050003", 17630 => x"50a3001a",
    17631 => x"204500ff", 17632 => x"3ca60008", 17633 => x"340a000f",
    17634 => x"b8c52800", 17635 => x"3ca60010", 17636 => x"b8804000",
    17637 => x"b8c53000", 17638 => x"b8603800", 17639 => x"b8802800",
    17640 => x"3409000f", 17641 => x"546a0017", 17642 => x"34040000",
    17643 => x"34070003", 17644 => x"b5042800", 17645 => x"34840004",
    17646 => x"58a60000", 17647 => x"c8642800", 17648 => x"54a7fffc",
    17649 => x"3463fffc", 17650 => x"00640002", 17651 => x"20630003",
    17652 => x"34840001", 17653 => x"3c840002", 17654 => x"b5044000",
    17655 => x"b9002000", 17656 => x"44600007", 17657 => x"204200ff",
    17658 => x"34050000", 17659 => x"b4853000", 17660 => x"30c20000",
    17661 => x"34a50001", 17662 => x"5c65fffd", 17663 => x"c3a00000",
    17664 => x"58a60000", 17665 => x"58a60004", 17666 => x"58a60008",
    17667 => x"58a6000c", 17668 => x"34e7fff0", 17669 => x"34a50010",
    17670 => x"54e9fffa", 17671 => x"3463fff0", 17672 => x"00680004",
    17673 => x"2063000f", 17674 => x"35080001", 17675 => x"3d080004",
    17676 => x"b4884000", 17677 => x"34040003", 17678 => x"5464ffdc",
    17679 => x"b9002000", 17680 => x"e3ffffe8", 17681 => x"78030001",
    17682 => x"38634d50", 17683 => x"28670000", 17684 => x"b8204800",
    17685 => x"34030000", 17686 => x"34060001", 17687 => x"e0000009",
    17688 => x"40840000", 17689 => x"b4e44000", 17690 => x"41080001",
    17691 => x"21080003", 17692 => x"45060012", 17693 => x"c8a40800",
    17694 => x"5c200013", 17695 => x"44810012", 17696 => x"b5232800",
    17697 => x"40a50000", 17698 => x"b4432000", 17699 => x"34630001",
    17700 => x"b4e54000", 17701 => x"41080001", 17702 => x"21080003",
    17703 => x"5d06fff1", 17704 => x"40840000", 17705 => x"34a50020",
    17706 => x"b4e44000", 17707 => x"41080001", 17708 => x"21080003",
    17709 => x"5d06fff0", 17710 => x"34840020", 17711 => x"c8a40800",
    17712 => x"4420ffef", 17713 => x"c3a00000", 17714 => x"b8412800",
    17715 => x"20a50003", 17716 => x"b8403800", 17717 => x"b8202000",
    17718 => x"5ca00018", 17719 => x"78040001", 17720 => x"388442c8",
    17721 => x"28430000", 17722 => x"28880000", 17723 => x"78040001",
    17724 => x"388442cc", 17725 => x"28870000", 17726 => x"a4603000",
    17727 => x"b4682000", 17728 => x"a0c43000", 17729 => x"a0c73000",
    17730 => x"b8202000", 17731 => x"5cc5000a", 17732 => x"58830000",
    17733 => x"34420004", 17734 => x"28430000", 17735 => x"34840004",
    17736 => x"a4603000", 17737 => x"b4682800", 17738 => x"a0c52800",
    17739 => x"a0a72800", 17740 => x"44a0fff8", 17741 => x"b8403800",
    17742 => x"34030000", 17743 => x"b4e32800", 17744 => x"40a50000",
    17745 => x"b4833000", 17746 => x"34630001", 17747 => x"30c50000",
    17748 => x"5ca0fffb", 17749 => x"c3a00000", 17750 => x"20220003",
    17751 => x"4440002c", 17752 => x"40230000", 17753 => x"34020000",
    17754 => x"44600027", 17755 => x"b8201000", 17756 => x"e0000003",
    17757 => x"40430000", 17758 => x"44600022", 17759 => x"34420001",
    17760 => x"20430003", 17761 => x"5c60fffc", 17762 => x"78040001",
    17763 => x"388442c8", 17764 => x"28430000", 17765 => x"28860000",
    17766 => x"78040001", 17767 => x"388442cc", 17768 => x"28850000",
    17769 => x"a4602000", 17770 => x"b4661800", 17771 => x"a0641800",
    17772 => x"a0651800", 17773 => x"5c600011", 17774 => x"34420004",
    17775 => x"28430000", 17776 => x"b4662000", 17777 => x"a4601800",
    17778 => x"a0831800", 17779 => x"a0651800", 17780 => x"5c60000a",
    17781 => x"34420004", 17782 => x"28430000", 17783 => x"b4662000",
    17784 => x"a4601800", 17785 => x"a0831800", 17786 => x"a0651800",
    17787 => x"4460fff3", 17788 => x"e0000002", 17789 => x"34420001",
    17790 => x"40430000", 17791 => x"5c60fffe", 17792 => x"c8411000",
    17793 => x"b8400800", 17794 => x"c3a00000", 17795 => x"b8201000",
    17796 => x"e3ffffde", 17797 => x"34060000", 17798 => x"44600017",
    17799 => x"b8413800", 17800 => x"20e70003", 17801 => x"3464ffff",
    17802 => x"44e00015", 17803 => x"40230000", 17804 => x"40450000",
    17805 => x"5c65000f", 17806 => x"34060000", 17807 => x"4480000e",
    17808 => x"34210001", 17809 => x"34420001", 17810 => x"5c600004",
    17811 => x"e000000a", 17812 => x"44800033", 17813 => x"44600032",
    17814 => x"40230000", 17815 => x"40450000", 17816 => x"3484ffff",
    17817 => x"34210001", 17818 => x"34420001", 17819 => x"4465fff9",
    17820 => x"c8653000", 17821 => x"b8c00800", 17822 => x"c3a00000",
    17823 => x"b8202800", 17824 => x"34010003", 17825 => x"b8402000",
    17826 => x"50230028", 17827 => x"28a10000", 17828 => x"28420000",
    17829 => x"5c220025", 17830 => x"3463fffc", 17831 => x"b8e03000",
    17832 => x"4460fff5", 17833 => x"78020001", 17834 => x"384242c8",
    17835 => x"28490000", 17836 => x"78020001", 17837 => x"384242cc",
    17838 => x"28480000", 17839 => x"a4201000", 17840 => x"b4290800",
    17841 => x"a0220800", 17842 => x"a0280800", 17843 => x"34070003",
    17844 => x"5c20ffe9", 17845 => x"34a50004", 17846 => x"34840004",
    17847 => x"54670006", 17848 => x"b8a00800", 17849 => x"b8801000",
    17850 => x"44600014", 17851 => x"3464ffff", 17852 => x"e3ffffcf",
    17853 => x"28a10000", 17854 => x"288a0000", 17855 => x"b4293000",
    17856 => x"a4201000", 17857 => x"a0c21000", 17858 => x"a0481000",
    17859 => x"5c2a0007", 17860 => x"3463fffc", 17861 => x"44600002",
    17862 => x"4440ffef", 17863 => x"34060000", 17864 => x"b8c00800",
    17865 => x"c3a00000", 17866 => x"b8801000", 17867 => x"b8a00800",
    17868 => x"3464ffff", 17869 => x"e3ffffbe", 17870 => x"40a30000",
    17871 => x"40850000", 17872 => x"c8653000", 17873 => x"e3ffffcc",
    17874 => x"b8412000", 17875 => x"20840003", 17876 => x"74650003",
    17877 => x"64840000", 17878 => x"b8403000", 17879 => x"a0852000",
    17880 => x"b8202800", 17881 => x"44800015", 17882 => x"78040001",
    17883 => x"388442c8", 17884 => x"28890000", 17885 => x"78040001",
    17886 => x"388442cc", 17887 => x"28880000", 17888 => x"340a0003",
    17889 => x"e0000006", 17890 => x"58a40000", 17891 => x"3463fffc",
    17892 => x"34a50004", 17893 => x"34420004", 17894 => x"51430007",
    17895 => x"28440000", 17896 => x"a4803800", 17897 => x"b4893000",
    17898 => x"a0e63000", 17899 => x"a0c83000", 17900 => x"44c0fff6",
    17901 => x"b8403000", 17902 => x"44600014", 17903 => x"40c20000",
    17904 => x"3463ffff", 17905 => x"34a40001", 17906 => x"30a20000",
    17907 => x"44400009", 17908 => x"34c20001", 17909 => x"4460000e",
    17910 => x"40450000", 17911 => x"3463ffff", 17912 => x"34420001",
    17913 => x"30850000", 17914 => x"34840001", 17915 => x"5ca0fffa",
    17916 => x"34020000", 17917 => x"44600007", 17918 => x"b4822800",
    17919 => x"30a00000", 17920 => x"34420001", 17921 => x"5c62fffd",
    17922 => x"c3a00000", 17923 => x"c3a00000", 17924 => x"c3a00000",
    17925 => x"57522043", 17926 => x"6f72653a", 17927 => x"20737461",
    17928 => x"7274696e", 17929 => x"67207570", 17930 => x"2e2e2e0a",
    17931 => x"00000000", 17932 => x"556e6162", 17933 => x"6c652074",
    17934 => x"6f206465", 17935 => x"7465726d", 17936 => x"696e6520",
    17937 => x"4d414320", 17938 => x"61646472", 17939 => x"6573730a",
    17940 => x"00000000", 17941 => x"4c6f6361", 17942 => x"6c204d41",
    17943 => x"43206164", 17944 => x"64726573", 17945 => x"733a2025",
    17946 => x"3032783a", 17947 => x"25303278", 17948 => x"3a253032",
    17949 => x"783a2530", 17950 => x"32783a25", 17951 => x"3032783a",
    17952 => x"25303278", 17953 => x"0a000000", 17954 => x"4c696e6b",
    17955 => x"2075702e", 17956 => x"0a000000", 17957 => x"4c696e6b",
    17958 => x"20646f77", 17959 => x"6e2e0a00", 17960 => x"25750000",
    17961 => x"25752575", 17962 => x"00000000", 17963 => x"0a0a5054",
    17964 => x"50207374", 17965 => x"61747573", 17966 => x"3a200000",
    17967 => x"25730000", 17968 => x"0a0a5379", 17969 => x"6e632069",
    17970 => x"6e666f20", 17971 => x"6e6f7420", 17972 => x"76616c69",
    17973 => x"640a0a00", 17974 => x"0a0a5379", 17975 => x"6e636872",
    17976 => x"6f6e697a", 17977 => x"6174696f", 17978 => x"6e207374",
    17979 => x"61747573", 17980 => x"3a0a0a00", 17981 => x"57522050",
    17982 => x"54502043", 17983 => x"6f726520", 17984 => x"53796e63",
    17985 => x"204d6f6e", 17986 => x"69746f72", 17987 => x"20762031",
    17988 => x"2e300000", 17989 => x"45736320", 17990 => x"3d206578",
    17991 => x"69740000", 17992 => x"0a0a5441", 17993 => x"49205469",
    17994 => x"6d653a20", 17995 => x"20202020", 17996 => x"20202020",
    17997 => x"20202020", 17998 => x"20202020", 17999 => x"20000000",
    18000 => x"0a0a4c69", 18001 => x"6e6b2073", 18002 => x"74617475",
    18003 => x"733a0000", 18004 => x"25733a20", 18005 => x"00000000",
    18006 => x"77727531", 18007 => x"00000000", 18008 => x"4c696e6b",
    18009 => x"20757020", 18010 => x"20200000", 18011 => x"4c696e6b",
    18012 => x"20646f77", 18013 => x"6e200000", 18014 => x"2852583a",
    18015 => x"2025642c", 18016 => x"2054583a", 18017 => x"20256429",
    18018 => x"2c206d6f", 18019 => x"64653a20", 18020 => x"00000000",
    18021 => x"5752204f", 18022 => x"66660000", 18023 => x"436c6f63",
    18024 => x"6b206f66", 18025 => x"66736574", 18026 => x"3a202020",
    18027 => x"20202020", 18028 => x"20202020", 18029 => x"20202020",
    18030 => x"20200000", 18031 => x"2532692e", 18032 => x"25303969",
    18033 => x"20730000", 18034 => x"25396920", 18035 => x"6e730000",
    18036 => x"0a4f6e65", 18037 => x"2d776179", 18038 => x"2064656c",
    18039 => x"61792061", 18040 => x"76657261", 18041 => x"6765643a",
    18042 => x"20202020", 18043 => x"20202000", 18044 => x"0a4f6273",
    18045 => x"65727665", 18046 => x"64206472", 18047 => x"6966743a",
    18048 => x"20202020", 18049 => x"20202020", 18050 => x"20202020",
    18051 => x"20202000", 18052 => x"5752204d", 18053 => x"61737465",
    18054 => x"72202000", 18055 => x"57522053", 18056 => x"6c617665",
    18057 => x"20202000", 18058 => x"57522055", 18059 => x"6e6b6e6f",
    18060 => x"776e2020", 18061 => x"20000000", 18062 => x"4c6f636b",
    18063 => x"65642020", 18064 => x"00000000", 18065 => x"4e6f4c6f",
    18066 => x"636b2020", 18067 => x"00000000", 18068 => x"43616c69",
    18069 => x"62726174", 18070 => x"65642020", 18071 => x"00000000",
    18072 => x"556e6361", 18073 => x"6c696272", 18074 => x"61746564",
    18075 => x"20200000", 18076 => x"0a495076", 18077 => x"343a2000",
    18078 => x"424f4f54", 18079 => x"50207275", 18080 => x"6e6e696e",
    18081 => x"67000000", 18082 => x"25642e25", 18083 => x"642e2564",
    18084 => x"2e256400", 18085 => x"53657276", 18086 => x"6f207374",
    18087 => x"6174653a", 18088 => x"20202020", 18089 => x"20202020",
    18090 => x"20202020", 18091 => x"20202000", 18092 => x"50686173",
    18093 => x"65207472", 18094 => x"61636b69", 18095 => x"6e673a20",
    18096 => x"20202020", 18097 => x"20202020", 18098 => x"20202000",
    18099 => x"4f4e0a00", 18100 => x"4f46460a", 18101 => x"00000000",
    18102 => x"41757820", 18103 => x"636c6f63", 18104 => x"6b207374",
    18105 => x"61747573", 18106 => x"3a202020", 18107 => x"20202020",
    18108 => x"20202000", 18109 => x"656e6162", 18110 => x"6c656400",
    18111 => x"2c206c6f", 18112 => x"636b6564", 18113 => x"00000000",
    18114 => x"0a54696d", 18115 => x"696e6720", 18116 => x"70617261",
    18117 => x"6d657465", 18118 => x"72733a0a", 18119 => x"0a000000",
    18120 => x"526f756e", 18121 => x"642d7472", 18122 => x"69702074",
    18123 => x"696d6520", 18124 => x"286d7529", 18125 => x"3a202020",
    18126 => x"20000000", 18127 => x"25732070", 18128 => x"730a0000",
    18129 => x"4d617374", 18130 => x"65722d73", 18131 => x"6c617665",
    18132 => x"2064656c", 18133 => x"61793a20", 18134 => x"20202020",
    18135 => x"20000000", 18136 => x"4d617374", 18137 => x"65722050",
    18138 => x"48592064", 18139 => x"656c6179", 18140 => x"733a2020",
    18141 => x"20202020", 18142 => x"20000000", 18143 => x"54583a20",
    18144 => x"25642070", 18145 => x"732c2052", 18146 => x"583a2025",
    18147 => x"64207073", 18148 => x"0a000000", 18149 => x"536c6176",
    18150 => x"65205048", 18151 => x"59206465", 18152 => x"6c617973",
    18153 => x"3a202020", 18154 => x"20202020", 18155 => x"20000000",
    18156 => x"546f7461", 18157 => x"6c206c69", 18158 => x"6e6b2061",
    18159 => x"73796d6d", 18160 => x"65747279", 18161 => x"3a202020",
    18162 => x"20000000", 18163 => x"25396420", 18164 => x"70730a00",
    18165 => x"4361626c", 18166 => x"65207274", 18167 => x"74206465",
    18168 => x"6c61793a", 18169 => x"20202020", 18170 => x"20202020",
    18171 => x"20000000", 18172 => x"436c6f63", 18173 => x"6b206f66",
    18174 => x"66736574", 18175 => x"3a202020", 18176 => x"20202020",
    18177 => x"20202020", 18178 => x"20000000", 18179 => x"50686173",
    18180 => x"65207365", 18181 => x"74706f69", 18182 => x"6e743a20",
    18183 => x"20202020", 18184 => x"20202020", 18185 => x"20000000",
    18186 => x"536b6577", 18187 => x"3a202020", 18188 => x"20202020",
    18189 => x"20202020", 18190 => x"20202020", 18191 => x"20202020",
    18192 => x"20000000", 18193 => x"4d616e75", 18194 => x"616c2070",
    18195 => x"68617365", 18196 => x"2061646a", 18197 => x"7573746d",
    18198 => x"656e743a", 18199 => x"20000000", 18200 => x"55706461",
    18201 => x"74652063", 18202 => x"6f756e74", 18203 => x"65723a20",
    18204 => x"20202020", 18205 => x"20202020", 18206 => x"20000000",
    18207 => x"2539640a", 18208 => x"00000000", 18209 => x"2d2d0000",
    18210 => x"6c6e6b3a", 18211 => x"25642072", 18212 => x"783a2564",
    18213 => x"2074783a", 18214 => x"25642000", 18215 => x"6c6f636b",
    18216 => x"3a256420", 18217 => x"00000000", 18218 => x"7074703a",
    18219 => x"25732000", 18220 => x"73763a25", 18221 => x"64200000",
    18222 => x"73733a27", 18223 => x"25732720", 18224 => x"00000000",
    18225 => x"6175783a", 18226 => x"25782000", 18227 => x"7365633a",
    18228 => x"2564206e", 18229 => x"7365633a", 18230 => x"25642000",
    18231 => x"6d753a25", 18232 => x"73200000", 18233 => x"646d733a",
    18234 => x"25732000", 18235 => x"6474786d", 18236 => x"3a256420",
    18237 => x"6472786d", 18238 => x"3a256420", 18239 => x"00000000",
    18240 => x"64747873", 18241 => x"3a256420", 18242 => x"64727873",
    18243 => x"3a256420", 18244 => x"00000000", 18245 => x"6173796d",
    18246 => x"3a256420", 18247 => x"00000000", 18248 => x"63727474",
    18249 => x"3a257320", 18250 => x"00000000", 18251 => x"636b6f3a",
    18252 => x"25642000", 18253 => x"73657470", 18254 => x"3a256420",
    18255 => x"00000000", 18256 => x"75636e74", 18257 => x"3a256420",
    18258 => x"00000000", 18259 => x"68643a25", 18260 => x"64206d64",
    18261 => x"3a256420", 18262 => x"61643a25", 18263 => x"64200000",
    18264 => x"74656d70", 18265 => x"3a202564", 18266 => x"2e253034",
    18267 => x"64204300", 18268 => x"756e6b6e", 18269 => x"6f776e00",
    18270 => x"64696167", 18271 => x"2d66736d", 18272 => x"2d312d25",
    18273 => x"733a2025", 18274 => x"3039642e", 18275 => x"25303364",
    18276 => x"3a200000", 18277 => x"454e5445", 18278 => x"52202573",
    18279 => x"2c207061", 18280 => x"636b6574", 18281 => x"206c656e",
    18282 => x"2025690a", 18283 => x"00000000", 18284 => x"25733a20",
    18285 => x"7265656e", 18286 => x"74657220", 18287 => x"696e2025",
    18288 => x"69206d73", 18289 => x"0a000000", 18290 => x"4c454156",
    18291 => x"45202573", 18292 => x"20286e65", 18293 => x"78743a20",
    18294 => x"25336929", 18295 => x"0a0a0000", 18296 => x"52454356",
    18297 => x"20253032", 18298 => x"64206279", 18299 => x"74657320",
    18300 => x"61742025", 18301 => x"642e2530", 18302 => x"39642028",
    18303 => x"74797065", 18304 => x"2025782c", 18305 => x"20257329",
    18306 => x"0a000000", 18307 => x"66736d20", 18308 => x"666f7220",
    18309 => x"25733a20", 18310 => x"4572726f", 18311 => x"72202569",
    18312 => x"20696e20", 18313 => x"25730a00", 18314 => x"66736d3a",
    18315 => x"20556e6b", 18316 => x"6e6f776e", 18317 => x"20737461",
    18318 => x"74652066", 18319 => x"6f722070", 18320 => x"6f727420",
    18321 => x"25730a00", 18322 => x"70707369", 18323 => x"00000000",
    18324 => x"25732d25", 18325 => x"692d2573", 18326 => x"3a200000",
    18327 => x"25733a20", 18328 => x"6572726f", 18329 => x"72207061",
    18330 => x"7273696e", 18331 => x"67202225", 18332 => x"73220a00",
    18333 => x"64696167", 18334 => x"2d636f6e", 18335 => x"66696700",
    18336 => x"64696167", 18337 => x"2d657874", 18338 => x"656e7369",
    18339 => x"6f6e0000", 18340 => x"64696167", 18341 => x"2d626d63",
    18342 => x"00000000", 18343 => x"64696167", 18344 => x"2d736572",
    18345 => x"766f0000", 18346 => x"64696167", 18347 => x"2d667261",
    18348 => x"6d657300", 18349 => x"64696167", 18350 => x"2d74696d",
    18351 => x"65000000", 18352 => x"64696167", 18353 => x"2d66736d",
    18354 => x"00000000", 18355 => x"50505369", 18356 => x"20666f72",
    18357 => x"20575250", 18358 => x"432e2043", 18359 => x"6f6d6d69",
    18360 => x"74202573", 18361 => x"2c206275", 18362 => x"696c7420",
    18363 => x"6f6e2041", 18364 => x"75672032", 18365 => x"35203230",
    18366 => x"31360a00", 18367 => x"70707369", 18368 => x"2d763230",
    18369 => x"31342e30", 18370 => x"372d3137", 18371 => x"332d6762",
    18372 => x"32303363", 18373 => x"63390000", 18374 => x"4c6f636b",
    18375 => x"696e6720", 18376 => x"504c4c00", 18377 => x"0a4c6f63",
    18378 => x"6b207469", 18379 => x"6d656f75", 18380 => x"742e0000",
    18381 => x"2e000000", 18382 => x"4c696e6b", 18383 => x"20646f77",
    18384 => x"6e3a2050", 18385 => x"54502073", 18386 => x"746f700a",
    18387 => x"00000000", 18388 => x"4c696e6b", 18389 => x"2075703a",
    18390 => x"20505450", 18391 => x"20737461", 18392 => x"72740a00",
    18393 => x"77723100", 18394 => x"25732573", 18395 => x"25303278",
    18396 => x"2d253032", 18397 => x"782d2530", 18398 => x"32782d25",
    18399 => x"3032782d", 18400 => x"25303278", 18401 => x"2d253032",
    18402 => x"782d2530", 18403 => x"32782d25", 18404 => x"3032782d",
    18405 => x"25303278", 18406 => x"2d253032", 18407 => x"780a0000",
    18408 => x"25732573", 18409 => x"25732028", 18410 => x"73697a65",
    18411 => x"20256929", 18412 => x"0a000000", 18413 => x"25732573",
    18414 => x"00000000", 18415 => x"25303278", 18416 => x"00000000",
    18417 => x"25735645", 18418 => x"5253494f", 18419 => x"4e3a2075",
    18420 => x"6e737570", 18421 => x"706f7274", 18422 => x"65642028",
    18423 => x"2569290a", 18424 => x"00000000", 18425 => x"25735645",
    18426 => x"5253494f", 18427 => x"4e3a2025", 18428 => x"69202874",
    18429 => x"79706520", 18430 => x"25692c20", 18431 => x"6c656e20",
    18432 => x"25692c20", 18433 => x"646f6d61", 18434 => x"696e2025",
    18435 => x"69290a00", 18436 => x"2573464c", 18437 => x"4147533a",
    18438 => x"20307825", 18439 => x"30347820", 18440 => x"28636f72",
    18441 => x"72656374", 18442 => x"696f6e20", 18443 => x"2530386c",
    18444 => x"75290a00", 18445 => x"504f5254", 18446 => x"3a200000",
    18447 => x"25735245", 18448 => x"53543a20", 18449 => x"73657120",
    18450 => x"25692c20", 18451 => x"6374726c", 18452 => x"2025692c",
    18453 => x"206c6f67", 18454 => x"2d696e74", 18455 => x"65727661",
    18456 => x"6c202569", 18457 => x"0a000000", 18458 => x"25734d45",
    18459 => x"53534147", 18460 => x"453a2028", 18461 => x"45292053",
    18462 => x"594e430a", 18463 => x"00000000", 18464 => x"25732573",
    18465 => x"256c752e", 18466 => x"25303969", 18467 => x"0a000000",
    18468 => x"4d53472d", 18469 => x"53594e43", 18470 => x"3a200000",
    18471 => x"25734d45", 18472 => x"53534147", 18473 => x"453a2028",
    18474 => x"45292044", 18475 => x"454c4159", 18476 => x"5f524551",
    18477 => x"0a000000", 18478 => x"4d53472d", 18479 => x"44454c41",
    18480 => x"595f5245", 18481 => x"513a2000", 18482 => x"25734d45",
    18483 => x"53534147", 18484 => x"453a2028", 18485 => x"47292046",
    18486 => x"4f4c4c4f", 18487 => x"575f5550", 18488 => x"0a000000",
    18489 => x"4d53472d", 18490 => x"464f4c4c", 18491 => x"4f575f55",
    18492 => x"503a2000", 18493 => x"25734d45", 18494 => x"53534147",
    18495 => x"453a2028", 18496 => x"47292044", 18497 => x"454c4159",
    18498 => x"5f524553", 18499 => x"500a0000", 18500 => x"4d53472d",
    18501 => x"44454c41", 18502 => x"595f5245", 18503 => x"53503a20",
    18504 => x"00000000", 18505 => x"25734d45", 18506 => x"53534147",
    18507 => x"453a2028", 18508 => x"47292041", 18509 => x"4e4e4f55",
    18510 => x"4e43450a", 18511 => x"00000000", 18512 => x"4d53472d",
    18513 => x"414e4e4f", 18514 => x"554e4345", 18515 => x"3a207374",
    18516 => x"616d7020", 18517 => x"00000000", 18518 => x"25732573",
    18519 => x"25303278", 18520 => x"2d253032", 18521 => x"782d2530",
    18522 => x"34780a00", 18523 => x"4d53472d", 18524 => x"414e4e4f",
    18525 => x"554e4345", 18526 => x"3a206772", 18527 => x"616e646d",
    18528 => x"61737465", 18529 => x"722d7175", 18530 => x"616c6974",
    18531 => x"79200000", 18532 => x"25734d53", 18533 => x"472d414e",
    18534 => x"4e4f554e", 18535 => x"43453a20", 18536 => x"6772616e",
    18537 => x"646d6173", 18538 => x"7465722d", 18539 => x"7072696f",
    18540 => x"20256920", 18541 => x"25690a00", 18542 => x"25732573",
    18543 => x"25303278", 18544 => x"2d253032", 18545 => x"782d2530",
    18546 => x"32782d25", 18547 => x"3032782d", 18548 => x"25303278",
    18549 => x"2d253032", 18550 => x"782d2530", 18551 => x"32782d25",
    18552 => x"3032780a", 18553 => x"00000000", 18554 => x"4d53472d",
    18555 => x"414e4e4f", 18556 => x"554e4345", 18557 => x"3a206772",
    18558 => x"616e646d", 18559 => x"61737465", 18560 => x"722d6964",
    18561 => x"20000000", 18562 => x"25734d45", 18563 => x"53534147",
    18564 => x"453a2028", 18565 => x"47292053", 18566 => x"49474e41",
    18567 => x"4c494e47", 18568 => x"0a000000", 18569 => x"4d53472d",
    18570 => x"5349474e", 18571 => x"414c494e", 18572 => x"473a2074",
    18573 => x"61726765", 18574 => x"742d706f", 18575 => x"72742000",
    18576 => x"2573544c", 18577 => x"563a2074", 18578 => x"6f6f2073",
    18579 => x"686f7274", 18580 => x"20282569", 18581 => x"202d2025",
    18582 => x"69203d20", 18583 => x"2569290a", 18584 => x"00000000",
    18585 => x"2573544c", 18586 => x"563a2074", 18587 => x"79706520",
    18588 => x"25303478", 18589 => x"206c656e", 18590 => x"20256920",
    18591 => x"6f756920", 18592 => x"25303278", 18593 => x"3a253032",
    18594 => x"783a2530", 18595 => x"32782073", 18596 => x"75622025",
    18597 => x"3032783a", 18598 => x"25303278", 18599 => x"3a253032",
    18600 => x"780a0000", 18601 => x"2573544c", 18602 => x"563a2074",
    18603 => x"6f6f2073", 18604 => x"686f7274", 18605 => x"20286578",
    18606 => x"70656374", 18607 => x"65642025", 18608 => x"692c2074",
    18609 => x"6f74616c", 18610 => x"20256929", 18611 => x"0a000000",
    18612 => x"544c563a", 18613 => x"20000000", 18614 => x"746c762d",
    18615 => x"636f6e74", 18616 => x"656e7400", 18617 => x"44554d50",
    18618 => x"3a200000", 18619 => x"7061796c", 18620 => x"6f616400",
    18621 => x"20696e76", 18622 => x"616c6964", 18623 => x"00000000",
    18624 => x"25735449", 18625 => x"4d453a20", 18626 => x"28256c69",
    18627 => x"202d2030", 18628 => x"78256c78", 18629 => x"2920256c",
    18630 => x"692e2530", 18631 => x"366c6925", 18632 => x"730a0000",
    18633 => x"2573564c", 18634 => x"414e2025", 18635 => x"690a0000",
    18636 => x"25734554", 18637 => x"483a2025", 18638 => x"30347820",
    18639 => x"28253032", 18640 => x"783a2530", 18641 => x"32783a25",
    18642 => x"3032783a", 18643 => x"25303278", 18644 => x"3a253032",
    18645 => x"783a2530", 18646 => x"3278202d", 18647 => x"3e202530",
    18648 => x"32783a25", 18649 => x"3032783a", 18650 => x"25303278",
    18651 => x"3a253032", 18652 => x"783a2530", 18653 => x"32783a25",
    18654 => x"30327829", 18655 => x"0a000000", 18656 => x"25734950",
    18657 => x"3a202569", 18658 => x"20282569", 18659 => x"2e25692e",
    18660 => x"25692e25", 18661 => x"69202d3e", 18662 => x"2025692e",
    18663 => x"25692e25", 18664 => x"692e2569", 18665 => x"29206c65",
    18666 => x"6e202569", 18667 => x"0a000000", 18668 => x"25735544",
    18669 => x"503a2028", 18670 => x"2569202d", 18671 => x"3e202569",
    18672 => x"29206c65", 18673 => x"6e202569", 18674 => x"0a000000",
    18675 => x"25733a20", 18676 => x"256c690a", 18677 => x"00000000",
    18678 => x"5761726e", 18679 => x"696e673a", 18680 => x"2025733a",
    18681 => x"2063616e", 18682 => x"206e6f74", 18683 => x"2061646a",
    18684 => x"75737420", 18685 => x"66726571", 18686 => x"5f707062",
    18687 => x"20256c69", 18688 => x"0a000000", 18689 => x"25733a20",
    18690 => x"25396c75", 18691 => x"2e253039", 18692 => x"6c690a00",
    18693 => x"25733a20", 18694 => x"736e743d", 18695 => x"25642c20",
    18696 => x"7365633d", 18697 => x"25642c20", 18698 => x"6e736563",
    18699 => x"3d25640a", 18700 => x"00000000", 18701 => x"73656e64",
    18702 => x"3a200000", 18703 => x"72656376", 18704 => x"3a200000",
    18705 => x"696e6974", 18706 => x"69616c69", 18707 => x"7a696e67",
    18708 => x"00000000", 18709 => x"6661756c", 18710 => x"74790000",
    18711 => x"64697361", 18712 => x"626c6564", 18713 => x"00000000",
    18714 => x"6c697374", 18715 => x"656e696e", 18716 => x"67000000",
    18717 => x"756e6361", 18718 => x"6c696272", 18719 => x"61746564",
    18720 => x"00000000", 18721 => x"736c6176", 18722 => x"65000000",
    18723 => x"756e6361", 18724 => x"6c696272", 18725 => x"61746564",
    18726 => x"2f77722d", 18727 => x"70726573", 18728 => x"656e7400",
    18729 => x"6d617374", 18730 => x"65722f77", 18731 => x"722d6d2d",
    18732 => x"6c6f636b", 18733 => x"00000000", 18734 => x"756e6361",
    18735 => x"6c696272", 18736 => x"61746564", 18737 => x"2f77722d",
    18738 => x"732d6c6f", 18739 => x"636b0000", 18740 => x"756e6361",
    18741 => x"6c696272", 18742 => x"61746564", 18743 => x"2f77722d",
    18744 => x"6c6f636b", 18745 => x"65640000", 18746 => x"77722d63",
    18747 => x"616c6962", 18748 => x"72617469", 18749 => x"6f6e0000",
    18750 => x"77722d63", 18751 => x"616c6962", 18752 => x"72617465",
    18753 => x"64000000", 18754 => x"77722d72", 18755 => x"6573702d",
    18756 => x"63616c69", 18757 => x"622d7265", 18758 => x"71000000",
    18759 => x"77722d6c", 18760 => x"696e6b2d", 18761 => x"6f6e0000",
    18762 => x"686f6f6b", 18763 => x"3a202573", 18764 => x"0a000000",
    18765 => x"5432206f", 18766 => x"72205433", 18767 => x"20696e63",
    18768 => x"6f727265", 18769 => x"63742c20", 18770 => x"64697363",
    18771 => x"61726469", 18772 => x"6e672074", 18773 => x"75706c65",
    18774 => x"0a000000", 18775 => x"48616e64", 18776 => x"7368616b",
    18777 => x"65206661", 18778 => x"696c7572", 18779 => x"653a206e",
    18780 => x"6f77206e", 18781 => x"6f6e2d77", 18782 => x"72202573",
    18783 => x"0a000000", 18784 => x"52657472", 18785 => x"79206f6e",
    18786 => x"2074696d", 18787 => x"656f7574", 18788 => x"0a000000",
    18789 => x"25733a20", 18790 => x"73756273", 18791 => x"74617465",
    18792 => x"2025690a", 18793 => x"00000000", 18794 => x"54783d3e",
    18795 => x"3e736361", 18796 => x"6c656450", 18797 => x"69636f73",
    18798 => x"65636f6e", 18799 => x"64732e6d", 18800 => x"7362203d",
    18801 => x"20307825", 18802 => x"780a0000", 18803 => x"54783d3e",
    18804 => x"3e736361", 18805 => x"6c656450", 18806 => x"69636f73",
    18807 => x"65636f6e", 18808 => x"64732e6c", 18809 => x"7362203d",
    18810 => x"20307825", 18811 => x"780a0000", 18812 => x"52782066",
    18813 => x"69786564", 18814 => x"2064656c", 18815 => x"6179203d",
    18816 => x"2025640a", 18817 => x"00000000", 18818 => x"52783d3e",
    18819 => x"3e736361", 18820 => x"6c656450", 18821 => x"69636f73",
    18822 => x"65636f6e", 18823 => x"64732e6d", 18824 => x"7362203d",
    18825 => x"20307825", 18826 => x"780a0000", 18827 => x"52783d3e",
    18828 => x"3e736361", 18829 => x"6c656450", 18830 => x"69636f73",
    18831 => x"65636f6e", 18832 => x"64732e6c", 18833 => x"7362203d",
    18834 => x"20307825", 18835 => x"780a0000", 18836 => x"4552524f",
    18837 => x"523a204e", 18838 => x"65772063", 18839 => x"6c617373",
    18840 => x"2025690a", 18841 => x"00000000", 18842 => x"4255473a",
    18843 => x"20547279", 18844 => x"696e6720", 18845 => x"746f2073",
    18846 => x"656e6420", 18847 => x"696e7661", 18848 => x"6c696420",
    18849 => x"77725f6d", 18850 => x"7367206d", 18851 => x"6f64653d",
    18852 => x"25782069", 18853 => x"643d2578", 18854 => x"00000000",
    18855 => x"68616e64", 18856 => x"6c652053", 18857 => x"69676e61",
    18858 => x"6c696e67", 18859 => x"206d7367", 18860 => x"2c206661",
    18861 => x"696c6564", 18862 => x"2c205468", 18863 => x"69732069",
    18864 => x"73206e6f", 18865 => x"74206f72", 18866 => x"67616e69",
    18867 => x"7a617469", 18868 => x"6f6e2065", 18869 => x"7874656e",
    18870 => x"73696f6e", 18871 => x"20544c56", 18872 => x"203d2030",
    18873 => x"7825780a", 18874 => x"00000000", 18875 => x"68616e64",
    18876 => x"6c652053", 18877 => x"69676e61", 18878 => x"6c696e67",
    18879 => x"206d7367", 18880 => x"2c206661", 18881 => x"696c6564",
    18882 => x"2c206e6f", 18883 => x"74204345", 18884 => x"524e2773",
    18885 => x"204f5549", 18886 => x"203d2030", 18887 => x"7825780a",
    18888 => x"00000000", 18889 => x"68616e64", 18890 => x"6c652053",
    18891 => x"69676e61", 18892 => x"6c696e67", 18893 => x"206d7367",
    18894 => x"2c206661", 18895 => x"696c6564", 18896 => x"2c206e6f",
    18897 => x"74205768", 18898 => x"69746520", 18899 => x"52616262",
    18900 => x"6974206d", 18901 => x"61676963", 18902 => x"206e756d",
    18903 => x"62657220", 18904 => x"3d203078", 18905 => x"25780a00",
    18906 => x"68616e64", 18907 => x"6c652053", 18908 => x"69676e61",
    18909 => x"6c696e67", 18910 => x"206d7367", 18911 => x"2c206661",
    18912 => x"696c6564", 18913 => x"2c206e6f", 18914 => x"74207375",
    18915 => x"70706f72", 18916 => x"74656420", 18917 => x"76657273",
    18918 => x"696f6e20", 18919 => x"6e756d62", 18920 => x"6572203d",
    18921 => x"20307825", 18922 => x"780a0000", 18923 => x"25732825",
    18924 => x"6429204d", 18925 => x"65737361", 18926 => x"67652063",
    18927 => x"616e2774", 18928 => x"20626520", 18929 => x"73656e74",
    18930 => x"0a000000", 18931 => x"53454e54", 18932 => x"20253032",
    18933 => x"64206279", 18934 => x"74657320", 18935 => x"61742025",
    18936 => x"642e2530", 18937 => x"39642028", 18938 => x"2573290a",
    18939 => x"00000000", 18940 => x"556e696e", 18941 => x"69746961",
    18942 => x"6c697a65", 18943 => x"64000000", 18944 => x"20287761",
    18945 => x"69742066", 18946 => x"6f722068", 18947 => x"77290000",
    18948 => x"4552524f", 18949 => x"523a2025", 18950 => x"733a2054",
    18951 => x"696d6573", 18952 => x"74616d70", 18953 => x"73496e63",
    18954 => x"6f727265", 18955 => x"63743a20", 18956 => x"25642025",
    18957 => x"64202564", 18958 => x"2025640a", 18959 => x"00000000",
    18960 => x"2573203d", 18961 => x"2025643a", 18962 => x"25643a25",
    18963 => x"640a0000", 18964 => x"73657276", 18965 => x"6f3a7431",
    18966 => x"00000000", 18967 => x"73657276", 18968 => x"6f3a7432",
    18969 => x"00000000", 18970 => x"73657276", 18971 => x"6f3a7433",
    18972 => x"00000000", 18973 => x"73657276", 18974 => x"6f3a7434",
    18975 => x"00000000", 18976 => x"2d3e6d64", 18977 => x"656c6179",
    18978 => x"00000000", 18979 => x"504c4c20", 18980 => x"4f75744f",
    18981 => x"664c6f63", 18982 => x"6b2c2073", 18983 => x"686f756c",
    18984 => x"64207265", 18985 => x"73746172", 18986 => x"74207379",
    18987 => x"6e630a00", 18988 => x"73657276", 18989 => x"6f3a6275",
    18990 => x"73790a00", 18991 => x"6f666673", 18992 => x"65745f68",
    18993 => x"773a2025", 18994 => x"6c692e25", 18995 => x"30396c69",
    18996 => x"20282b25", 18997 => x"6c69290a", 18998 => x"00000000",
    18999 => x"77725f73", 19000 => x"6572766f", 19001 => x"20737461",
    19002 => x"74653a20", 19003 => x"25732573", 19004 => x"0a000000",
    19005 => x"6f6c6473", 19006 => x"65747020", 19007 => x"25692c20",
    19008 => x"6f666673", 19009 => x"65742025", 19010 => x"693a2530",
    19011 => x"34690a00", 19012 => x"61646a75", 19013 => x"73742070",
    19014 => x"68617365", 19015 => x"2025690a", 19016 => x"00000000",
    19017 => x"53594e43", 19018 => x"5f4e5345", 19019 => x"43000000",
    19020 => x"53594e43", 19021 => x"5f534543", 19022 => x"00000000",
    19023 => x"53594e43", 19024 => x"5f504841", 19025 => x"53450000",
    19026 => x"54524143", 19027 => x"4b5f5048", 19028 => x"41534500",
    19029 => x"57414954", 19030 => x"5f4f4646", 19031 => x"5345545f",
    19032 => x"53544142", 19033 => x"4c450000", 19034 => x"7072652d",
    19035 => x"6d617374", 19036 => x"65720000", 19037 => x"70617373",
    19038 => x"69766500", 19039 => x"25733a20", 19040 => x"63616e27",
    19041 => x"7420696e", 19042 => x"69742065", 19043 => x"7874656e",
    19044 => x"73696f6e", 19045 => x"0a000000", 19046 => x"636c6f63",
    19047 => x"6b20636c", 19048 => x"61737320", 19049 => x"3d202564",
    19050 => x"0a000000", 19051 => x"636c6f63", 19052 => x"6b206163",
    19053 => x"63757261", 19054 => x"6379203d", 19055 => x"2025640a",
    19056 => x"00000000", 19057 => x"70705f73", 19058 => x"6c617665",
    19059 => x"203a2044", 19060 => x"656c6179", 19061 => x"20526573",
    19062 => x"7020646f", 19063 => x"65736e27", 19064 => x"74206d61",
    19065 => x"74636820", 19066 => x"44656c61", 19067 => x"79205265",
    19068 => x"710a0000", 19069 => x"4e657720", 19070 => x"666f7265",
    19071 => x"69676e20", 19072 => x"4d617374", 19073 => x"65722025",
    19074 => x"69206164", 19075 => x"6465640a", 19076 => x"00000000",
    19077 => x"4552524f", 19078 => x"523a2025", 19079 => x"733a2046",
    19080 => x"6f6c6c6f", 19081 => x"77207570", 19082 => x"206d6573",
    19083 => x"73616765", 19084 => x"20697320", 19085 => x"6e6f7420",
    19086 => x"66726f6d", 19087 => x"20637572", 19088 => x"72656e74",
    19089 => x"20706172", 19090 => x"656e740a", 19091 => x"00000000",
    19092 => x"4552524f", 19093 => x"523a2025", 19094 => x"733a2053",
    19095 => x"6c617665", 19096 => x"20776173", 19097 => x"206e6f74",
    19098 => x"20776169", 19099 => x"74696e67", 19100 => x"20612066",
    19101 => x"6f6c6c6f", 19102 => x"77207570", 19103 => x"206d6573",
    19104 => x"73616765", 19105 => x"0a000000", 19106 => x"4552524f",
    19107 => x"523a2025", 19108 => x"733a2053", 19109 => x"65717565",
    19110 => x"6e636549", 19111 => x"44202564", 19112 => x"20646f65",
    19113 => x"736e2774", 19114 => x"206d6174", 19115 => x"6368206c",
    19116 => x"61737420", 19117 => x"53796e63", 19118 => x"206d6573",
    19119 => x"73616765", 19120 => x"2025640a", 19121 => x"00000000",
    19122 => x"416e6e6f", 19123 => x"756e6365", 19124 => x"206d6573",
    19125 => x"73616765", 19126 => x"2066726f", 19127 => x"6d20616e",
    19128 => x"6f746865", 19129 => x"7220666f", 19130 => x"72656967",
    19131 => x"6e206d61", 19132 => x"73746572", 19133 => x"0a000000",
    19134 => x"25733a25", 19135 => x"693a2045", 19136 => x"72726f72",
    19137 => x"20310a00", 19138 => x"25733a25", 19139 => x"693a2045",
    19140 => x"72726f72", 19141 => x"20320a00", 19142 => x"42657374",
    19143 => x"20666f72", 19144 => x"6569676e", 19145 => x"206d6173",
    19146 => x"74657220", 19147 => x"69732025", 19148 => x"692f2569",
    19149 => x"0a000000", 19150 => x"25733a20", 19151 => x"6572726f",
    19152 => x"720a0000", 19153 => x"25733a20", 19154 => x"70617373",
    19155 => x"6976650a", 19156 => x"00000000", 19157 => x"25733a20",
    19158 => x"6d617374", 19159 => x"65720a00", 19160 => x"4e657720",
    19161 => x"55544320", 19162 => x"6f666673", 19163 => x"65743a20",
    19164 => x"25690a00", 19165 => x"25733a20", 19166 => x"736c6176",
    19167 => x"650a0000", 19168 => x"73796e63", 19169 => x"00000000",
    19170 => x"64656c61", 19171 => x"795f7265", 19172 => x"71000000",
    19173 => x"7064656c", 19174 => x"61795f72", 19175 => x"65710000",
    19176 => x"7064656c", 19177 => x"61795f72", 19178 => x"65737000",
    19179 => x"64656c61", 19180 => x"795f7265", 19181 => x"73700000",
    19182 => x"7064656c", 19183 => x"61795f72", 19184 => x"6573705f",
    19185 => x"666f6c6c", 19186 => x"6f775f75", 19187 => x"70000000",
    19188 => x"616e6e6f", 19189 => x"756e6365", 19190 => x"00000000",
    19191 => x"7369676e", 19192 => x"616c696e", 19193 => x"67000000",
    19194 => x"6d616e61", 19195 => x"67656d65", 19196 => x"6e740000",
    19197 => x"4552524f", 19198 => x"523a2042", 19199 => x"55473a20",
    19200 => x"25732064", 19201 => x"6f65736e", 19202 => x"27742073",
    19203 => x"7570706f", 19204 => x"7274206e", 19205 => x"65676174",
    19206 => x"69766573", 19207 => x"0a000000", 19208 => x"4552524f",
    19209 => x"523a204e", 19210 => x"65676174", 19211 => x"69766520",
    19212 => x"76616c75", 19213 => x"65206361", 19214 => x"6e6e6f74",
    19215 => x"20626520", 19216 => x"636f6e76", 19217 => x"65727465",
    19218 => x"6420696e", 19219 => x"746f2074", 19220 => x"696d6573",
    19221 => x"74616d70", 19222 => x"0a000000", 19223 => x"4552524f",
    19224 => x"523a2074", 19225 => x"6f5f5469", 19226 => x"6d65496e",
    19227 => x"7465726e", 19228 => x"616c3a20", 19229 => x"7365636f",
    19230 => x"6e647320", 19231 => x"6669656c", 19232 => x"64206973",
    19233 => x"20686967", 19234 => x"68657220", 19235 => x"7468616e",
    19236 => x"20736967", 19237 => x"6e656420", 19238 => x"696e7465",
    19239 => x"67657220", 19240 => x"28333262", 19241 => x"69747329",
    19242 => x"0a000000", 19243 => x"2d000000", 19244 => x"25732564",
    19245 => x"2e253039", 19246 => x"64000000", 19247 => x"6572726f",
    19248 => x"7220696e", 19249 => x"20745f6f", 19250 => x"70732d3e",
    19251 => x"73657276", 19252 => x"6f5f696e", 19253 => x"69740000",
    19254 => x"496e6974", 19255 => x"69616c69", 19256 => x"7a65643a",
    19257 => x"206f6273", 19258 => x"5f647269", 19259 => x"66742025",
    19260 => x"6c6c690a", 19261 => x"00000000", 19262 => x"636f7272",
    19263 => x"65637469", 19264 => x"6f6e2066", 19265 => x"69656c64",
    19266 => x"20313a20", 19267 => x"25730a00", 19268 => x"64697363",
    19269 => x"61726420", 19270 => x"54332f54", 19271 => x"343a2077",
    19272 => x"65206d69", 19273 => x"73732054", 19274 => x"312f5432",
    19275 => x"0a000000", 19276 => x"636f7272", 19277 => x"65637469",
    19278 => x"6f6e2066", 19279 => x"69656c64", 19280 => x"20323a20",
    19281 => x"25730a00", 19282 => x"54313a20", 19283 => x"25730a00",
    19284 => x"54323a20", 19285 => x"25730a00", 19286 => x"54333a20",
    19287 => x"25730a00", 19288 => x"54343a20", 19289 => x"25730a00",
    19290 => x"4d617374", 19291 => x"65722074", 19292 => x"6f20736c",
    19293 => x"6176653a", 19294 => x"2025730a", 19295 => x"00000000",
    19296 => x"536c6176", 19297 => x"6520746f", 19298 => x"206d6173",
    19299 => x"7465723a", 19300 => x"2025730a", 19301 => x"00000000",
    19302 => x"6d65616e", 19303 => x"50617468", 19304 => x"44656c61",
    19305 => x"793a2025", 19306 => x"730a0000", 19307 => x"73657276",
    19308 => x"6f206162", 19309 => x"6f727465", 19310 => x"642c2064",
    19311 => x"656c6179", 19312 => x"20677265", 19313 => x"61746572",
    19314 => x"20746861", 19315 => x"6e203120", 19316 => x"7365636f",
    19317 => x"6e640a00", 19318 => x"73657276", 19319 => x"6f206162",
    19320 => x"6f727465", 19321 => x"642c2064", 19322 => x"656c6179",
    19323 => x"20256420", 19324 => x"6f722025", 19325 => x"64206772",
    19326 => x"65617465", 19327 => x"72207468", 19328 => x"616e2063",
    19329 => x"6f6e6669", 19330 => x"67757265", 19331 => x"64206d61",
    19332 => x"78696d75", 19333 => x"6d202564", 19334 => x"0a000000",
    19335 => x"5472696d", 19336 => x"20746f6f", 19337 => x"2d6c6f6e",
    19338 => x"67206d70", 19339 => x"643a2025", 19340 => x"690a0000",
    19341 => x"41667465", 19342 => x"72206176", 19343 => x"67282569",
    19344 => x"292c206d", 19345 => x"65616e50", 19346 => x"61746844",
    19347 => x"656c6179", 19348 => x"3a202569", 19349 => x"0a000000",
    19350 => x"4f666673", 19351 => x"65742066", 19352 => x"726f6d20",
    19353 => x"6d617374", 19354 => x"65723a20", 19355 => x"20202020",
    19356 => x"25730a00", 19357 => x"73657276", 19358 => x"6f206162",
    19359 => x"6f727465", 19360 => x"642c206f", 19361 => x"66667365",
    19362 => x"74206772", 19363 => x"65617465", 19364 => x"72207468",
    19365 => x"616e2031", 19366 => x"20736563", 19367 => x"6f6e640a",
    19368 => x"00000000", 19369 => x"73657276", 19370 => x"6f206162",
    19371 => x"6f727465", 19372 => x"642c206f", 19373 => x"66667365",
    19374 => x"74206772", 19375 => x"65617465", 19376 => x"72207468",
    19377 => x"616e2063", 19378 => x"6f6e6669", 19379 => x"67757265",
    19380 => x"64206d61", 19381 => x"78696d75", 19382 => x"6d202564",
    19383 => x"0a000000", 19384 => x"4f627365", 19385 => x"72766564",
    19386 => x"20647269", 19387 => x"66743a20", 19388 => x"2539690a",
    19389 => x"00000000", 19390 => x"74696d65", 19391 => x"6f757420",
    19392 => x"65787069", 19393 => x"7265643a", 19394 => x"2025730a",
    19395 => x"00000000", 19396 => x"50505f54", 19397 => x"4f5f4445",
    19398 => x"4c415952", 19399 => x"45510000", 19400 => x"50505f54",
    19401 => x"4f5f5359", 19402 => x"4e430000", 19403 => x"50505f54",
    19404 => x"4f5f414e", 19405 => x"4e5f5245", 19406 => x"43454950",
    19407 => x"54000000", 19408 => x"50505f54", 19409 => x"4f5f414e",
    19410 => x"4e5f494e", 19411 => x"54455256", 19412 => x"414c0000",
    19413 => x"50505f54", 19414 => x"4f5f4641", 19415 => x"554c5459",
    19416 => x"00000000", 19417 => x"50505f54", 19418 => x"4f5f4558",
    19419 => x"545f3000", 19420 => x"50505f54", 19421 => x"4f5f4558",
    19422 => x"545f3100", 19423 => x"50505f54", 19424 => x"4f5f4558",
    19425 => x"545f3200", 19426 => x"536c6176", 19427 => x"65204f6e",
    19428 => x"6c792c20", 19429 => x"636c6f63", 19430 => x"6b20636c",
    19431 => x"61737320", 19432 => x"73657420", 19433 => x"746f2032",
    19434 => x"35350a00", 19435 => x"1b5b3125", 19436 => x"63000000",
    19437 => x"436f6d6d", 19438 => x"616e6420", 19439 => x"22257322",
    19440 => x"3a206572", 19441 => x"726f7220", 19442 => x"25640a00",
    19443 => x"556e7265", 19444 => x"636f676e", 19445 => x"697a6564",
    19446 => x"20636f6d", 19447 => x"6d616e64", 19448 => x"20222573",
    19449 => x"222e0a00", 19450 => x"77726323", 19451 => x"20000000",
    19452 => x"25630000", 19453 => x"456d7074", 19454 => x"7920696e",
    19455 => x"69742073", 19456 => x"63726970", 19457 => x"742e2e2e",
    19458 => x"0a000000", 19459 => x"65786563", 19460 => x"7574696e",
    19461 => x"673a2025", 19462 => x"730a0000", 19463 => x"57522043",
    19464 => x"6f726520", 19465 => x"6275696c", 19466 => x"643a2025",
    19467 => x"7325730a", 19468 => x"00000000", 19469 => x"2028756e",
    19470 => x"73757070", 19471 => x"6f727465", 19472 => x"64206465",
    19473 => x"76656c6f", 19474 => x"70657220", 19475 => x"6275696c",
    19476 => x"64290000", 19477 => x"4275696c", 19478 => x"743a2025",
    19479 => x"73202573", 19480 => x"0a000000", 19481 => x"4275696c",
    19482 => x"7420666f", 19483 => x"72202564", 19484 => x"206b4220",
    19485 => x"52414d2c", 19486 => x"20737461", 19487 => x"636b2069",
    19488 => x"73202564", 19489 => x"20627974", 19490 => x"65730a00",
    19491 => x"5741524e", 19492 => x"494e473a", 19493 => x"20686172",
    19494 => x"64776172", 19495 => x"65207361", 19496 => x"79732025",
    19497 => x"696b4220", 19498 => x"3c3d2052", 19499 => x"414d203c",
    19500 => x"2025696b", 19501 => x"420a0000", 19502 => x"76657200",
    19503 => x"696e6974", 19504 => x"00000000", 19505 => x"636c0000",
    19506 => x"73746174", 19507 => x"00000000", 19508 => x"73707300",
    19509 => x"67707300", 19510 => x"25642025", 19511 => x"640a0000",
    19512 => x"73746172", 19513 => x"74000000", 19514 => x"73746f70",
    19515 => x"00000000", 19516 => x"73646163", 19517 => x"00000000",
    19518 => x"67646163", 19519 => x"00000000", 19520 => x"63686563",
    19521 => x"6b76636f", 19522 => x"00000000", 19523 => x"706c6c00",
    19524 => x"64657465", 19525 => x"63740000", 19526 => x"4e6f2053",
    19527 => x"46502e0a", 19528 => x"00000000", 19529 => x"65726173",
    19530 => x"65000000", 19531 => x"436f756c", 19532 => x"64206e6f",
    19533 => x"74206572", 19534 => x"61736520", 19535 => x"44420a00",
    19536 => x"61646400", 19537 => x"53465020", 19538 => x"44422069",
    19539 => x"73206675", 19540 => x"6c6c0a00", 19541 => x"49324320",
    19542 => x"6572726f", 19543 => x"720a0000", 19544 => x"25642053",
    19545 => x"46507320", 19546 => x"696e2044", 19547 => x"420a0000",
    19548 => x"73686f77", 19549 => x"00000000", 19550 => x"53465020",
    19551 => x"64617461", 19552 => x"62617365", 19553 => x"20656d70",
    19554 => x"74792e2e", 19555 => x"2e0a0000", 19556 => x"53465020",
    19557 => x"64617461", 19558 => x"62617365", 19559 => x"20636f72",
    19560 => x"72757074", 19561 => x"65642e2e", 19562 => x"2e0a0000",
    19563 => x"25643a20", 19564 => x"504e3a00", 19565 => x"20645478",
    19566 => x"3a202564", 19567 => x"2c206452", 19568 => x"783a2025",
    19569 => x"642c2061", 19570 => x"6c706861", 19571 => x"3a202564",
    19572 => x"0a000000", 19573 => x"6d617463", 19574 => x"68000000",
    19575 => x"52756e20", 19576 => x"73667020", 19577 => x"64657465",
    19578 => x"63742066", 19579 => x"69727374", 19580 => x"0a000000",
    19581 => x"53465020", 19582 => x"6d617463", 19583 => x"6865642c",
    19584 => x"20645478", 19585 => x"3d25642c", 19586 => x"20645278",
    19587 => x"3d25642c", 19588 => x"20616c70", 19589 => x"68613d25",
    19590 => x"640a0000", 19591 => x"436f756c", 19592 => x"64206e6f",
    19593 => x"74206d61", 19594 => x"74636820", 19595 => x"746f2044",
    19596 => x"420a0000", 19597 => x"656e6100", 19598 => x"73667000",
    19599 => x"73746174", 19600 => x"69737469", 19601 => x"6373206e",
    19602 => x"6f77206f", 19603 => x"66660a00", 19604 => x"62747300",
    19605 => x"6f666600", 19606 => x"70747000", 19607 => x"676d0000",
    19608 => x"6d6f6465", 19609 => x"00000000", 19610 => x"6772616e",
    19611 => x"646d6173", 19612 => x"74657200", 19613 => x"666f7263",
    19614 => x"65000000", 19615 => x"466f756e", 19616 => x"64207068",
    19617 => x"61736520", 19618 => x"7472616e", 19619 => x"73697469",
    19620 => x"6f6e2069", 19621 => x"6e204545", 19622 => x"50524f4d",
    19623 => x"3a202564", 19624 => x"70730a00", 19625 => x"4d656173",
    19626 => x"7572696e", 19627 => x"67207432", 19628 => x"2f743420",
    19629 => x"70686173", 19630 => x"65207472", 19631 => x"616e7369",
    19632 => x"74696f6e", 19633 => x"2e2e2e0a", 19634 => x"00000000",
    19635 => x"63616c69", 19636 => x"62726174", 19637 => x"696f6e00",
    19638 => x"73657400", 19639 => x"73657473", 19640 => x"65630000",
    19641 => x"7365746e", 19642 => x"73656300", 19643 => x"72617700",
    19644 => x"2573202b", 19645 => x"2564206e", 19646 => x"616e6f73",
    19647 => x"65636f6e", 19648 => x"64732e0a", 19649 => x"00000000",
    19650 => x"74696d65", 19651 => x"00000000", 19652 => x"67756900",
    19653 => x"73646200", 19654 => x"67657400", 19655 => x"67657470",
    19656 => x"00000000", 19657 => x"73657470", 19658 => x"00000000",
    19659 => x"4d41432d", 19660 => x"61646472", 19661 => x"6573733a",
    19662 => x"20253032", 19663 => x"783a2530", 19664 => x"32783a25",
    19665 => x"3032783a", 19666 => x"25303278", 19667 => x"3a253032",
    19668 => x"783a2530", 19669 => x"32780a00", 19670 => x"6d616300",
    19671 => x"45455052", 19672 => x"4f4d206e", 19673 => x"6f742066",
    19674 => x"6f756e64", 19675 => x"2e2e0a00", 19676 => x"436f756c",
    19677 => x"64206e6f", 19678 => x"74206572", 19679 => x"61736520",
    19680 => x"696e6974", 19681 => x"20736372", 19682 => x"6970740a",
    19683 => x"00000000", 19684 => x"436f756c", 19685 => x"64206e6f",
    19686 => x"74206164", 19687 => x"64207468", 19688 => x"6520636f",
    19689 => x"6d6d616e", 19690 => x"640a0000", 19691 => x"4f4b2e0a",
    19692 => x"00000000", 19693 => x"626f6f74", 19694 => x"00000000",
    19695 => x"4f4e0000", 19696 => x"4f464600", 19697 => x"656e6162",
    19698 => x"6c650000", 19699 => x"64697361", 19700 => x"626c6500",
    19701 => x"70686173", 19702 => x"65207472", 19703 => x"61636b69",
    19704 => x"6e672025", 19705 => x"730a0000", 19706 => x"70747261",
    19707 => x"636b0000", 19708 => x"41766169", 19709 => x"6c61626c",
    19710 => x"6520636f", 19711 => x"6d6d616e", 19712 => x"64733a0a",
    19713 => x"00000000", 19714 => x"20202573", 19715 => x"0a000000",
    19716 => x"68656c70", 19717 => x"00000000", 19718 => x"55736167",
    19719 => x"653a2072", 19720 => x"65667265", 19721 => x"7368203c",
    19722 => x"7365636f", 19723 => x"6e64733e", 19724 => x"0a000000",
    19725 => x"72656672", 19726 => x"65736800", 19727 => x"49502d61",
    19728 => x"64647265", 19729 => x"73733a20", 19730 => x"696e2074",
    19731 => x"7261696e", 19732 => x"696e670a", 19733 => x"00000000",
    19734 => x"49502d61", 19735 => x"64647265", 19736 => x"73733a20",
    19737 => x"25642e25", 19738 => x"642e2564", 19739 => x"2e25640a",
    19740 => x"00000000", 19741 => x"69700000", 19742 => x"50505349",
    19743 => x"20766572", 19744 => x"626f7369", 19745 => x"74793a20",
    19746 => x"2530386c", 19747 => x"780a0000", 19748 => x"76657262",
    19749 => x"6f736500", 19750 => x"25732c20", 19751 => x"25732025",
    19752 => x"642c2025", 19753 => x"642c2025", 19754 => x"3032643a",
    19755 => x"25303264", 19756 => x"3a253032", 19757 => x"64000000",
    19758 => x"1b5b3025", 19759 => x"643b3325", 19760 => x"646d0000",
    19761 => x"1b5b6d00", 19762 => x"1b5b2564", 19763 => x"3b256466",
    19764 => x"00000000", 19765 => x"1b5b324a", 19766 => x"1b5b313b",
    19767 => x"31480000", 19768 => x"53756e00", 19769 => x"4d6f6e00",
    19770 => x"54756500", 19771 => x"57656400", 19772 => x"54687500",
    19773 => x"46726900", 19774 => x"53617400", 19775 => x"4a616e00",
    19776 => x"46656200", 19777 => x"4d617200", 19778 => x"41707200",
    19779 => x"4d617900", 19780 => x"4a756e00", 19781 => x"4a756c00",
    19782 => x"41756700", 19783 => x"53657000", 19784 => x"4f637400",
    19785 => x"4e6f7600", 19786 => x"44656300", 19787 => x"4c6f6f70",
    19788 => x"73207065", 19789 => x"72206a69", 19790 => x"6666793a",
    19791 => x"2025690a", 19792 => x"00000000", 19793 => x"77723000",
    19794 => x"44697363", 19795 => x"6f766572", 19796 => x"65642049",
    19797 => x"50206164", 19798 => x"64726573", 19799 => x"73202825",
    19800 => x"642e2564", 19801 => x"2e25642e", 19802 => x"25642921",
    19803 => x"0a000000", 19804 => x"30313233", 19805 => x"34353637",
    19806 => x"38396162", 19807 => x"63646566", 19808 => x"00000000",
    19809 => x"49443a20", 19810 => x"25780a00", 19811 => x"7066696c",
    19812 => x"7465723a", 19813 => x"2077726f", 19814 => x"6e67206d",
    19815 => x"61676963", 19816 => x"206e756d", 19817 => x"62657220",
    19818 => x"28676f74", 19819 => x"20307825", 19820 => x"78290a00",
    19821 => x"7066696c", 19822 => x"7465723a", 19823 => x"2077726f",
    19824 => x"6e672072", 19825 => x"756c652d", 19826 => x"7365742c",
    19827 => x"2063616e", 19828 => x"27742061", 19829 => x"70706c79",
    19830 => x"0a000000", 19831 => x"696e7661", 19832 => x"6c696420",
    19833 => x"64657363", 19834 => x"72697074", 19835 => x"6f722040",
    19836 => x"2578203d", 19837 => x"2025780a", 19838 => x"00000000",
    19839 => x"5761726e", 19840 => x"696e673a", 19841 => x"20747820",
    19842 => x"6e6f7420", 19843 => x"7465726d", 19844 => x"696e6174",
    19845 => x"65642069", 19846 => x"6e66696e", 19847 => x"69746520",
    19848 => x"6d63723d", 19849 => x"30782578", 19850 => x"0a000000",
    19851 => x"5761726e", 19852 => x"696e673a", 19853 => x"20747820",
    19854 => x"74696d65", 19855 => x"7374616d", 19856 => x"70206e65",
    19857 => x"76657220", 19858 => x"62656361", 19859 => x"6d652061",
    19860 => x"7661696c", 19861 => x"61626c65", 19862 => x"0a000000",
    19863 => x"6d696e69", 19864 => x"635f7478", 19865 => x"5f667261",
    19866 => x"6d653a20", 19867 => x"756e6d61", 19868 => x"74636865",
    19869 => x"64206669", 19870 => x"64202564", 19871 => x"20767320",
    19872 => x"25640a00", 19873 => x"6e616e6f", 19874 => x"7365636f",
    19875 => x"6e647300", 19876 => x"41646a75", 19877 => x"73743a20",
    19878 => x"636f756e", 19879 => x"74657220", 19880 => x"3d202573",
    19881 => x"205b2563", 19882 => x"25645d0a", 19883 => x"00000000",
    19884 => x"64657620", 19885 => x"20307825", 19886 => x"30386c78",
    19887 => x"20402025", 19888 => x"30366c78", 19889 => x"2c202573",
    19890 => x"0a000000", 19891 => x"66706761", 19892 => x"2d617265",
    19893 => x"61000000", 19894 => x"4572726f", 19895 => x"72202564",
    19896 => x"20776869", 19897 => x"6c652072", 19898 => x"65616469",
    19899 => x"6e672074", 19900 => x"32347020", 19901 => x"66726f6d",
    19902 => x"2073746f", 19903 => x"72616765", 19904 => x"0a000000",
    19905 => x"74323470", 19906 => x"20726561", 19907 => x"64206672",
    19908 => x"6f6d2073", 19909 => x"746f7261", 19910 => x"67653a20",
    19911 => x"25642070", 19912 => x"730a0000", 19913 => x"52585453",
    19914 => x"2063616c", 19915 => x"69627261", 19916 => x"74696f6e",
    19917 => x"20657272", 19918 => x"6f722e0a", 19919 => x"00000000",
    19920 => x"52585453", 19921 => x"2063616c", 19922 => x"69627261",
    19923 => x"74696f6e", 19924 => x"3a205240", 19925 => x"25647073",
    19926 => x"2c204640", 19927 => x"25647073", 19928 => x"2c207472",
    19929 => x"616e7369", 19930 => x"74696f6e", 19931 => x"40256470",
    19932 => x"730a0000", 19933 => x"57616974", 19934 => x"696e6720",
    19935 => x"666f7220", 19936 => x"6c696e6b", 19937 => x"2e2e2e0a",
    19938 => x"00000000", 19939 => x"4c6f636b", 19940 => x"696e6720",
    19941 => x"504c4c2e", 19942 => x"2e2e0a00", 19943 => x"43616c69",
    19944 => x"62726174", 19945 => x"696e6720", 19946 => x"52582074",
    19947 => x"696d6573", 19948 => x"74616d70", 19949 => x"65722e2e",
    19950 => x"2e0a0000", 19951 => x"4661696c", 19952 => x"65640000",
    19953 => x"53756363", 19954 => x"65737300", 19955 => x"57726f74",
    19956 => x"65206e65", 19957 => x"77207432", 19958 => x"34702076",
    19959 => x"616c7565", 19960 => x"3a202564", 19961 => x"20707320",
    19962 => x"28257329", 19963 => x"0a000000", 19964 => x"43616e27",
    19965 => x"74207361", 19966 => x"76652070", 19967 => x"65727369",
    19968 => x"7374656e", 19969 => x"74204d41", 19970 => x"43206164",
    19971 => x"64726573", 19972 => x"730a0000", 19973 => x"25733a20",
    19974 => x"5573696e", 19975 => x"67205731", 19976 => x"20736572",
    19977 => x"69616c20", 19978 => x"6e756d62", 19979 => x"65720a00",
    19980 => x"6f666673", 19981 => x"65742025", 19982 => x"34692028",
    19983 => x"30782530", 19984 => x"3378293a", 19985 => x"20253369",
    19986 => x"20283078", 19987 => x"25303278", 19988 => x"290a0000",
    19989 => x"77726974", 19990 => x"65283078", 19991 => x"25782c20",
    19992 => x"2569293a", 19993 => x"20726573", 19994 => x"756c7420",
    19995 => x"3d202569", 19996 => x"0a000000", 19997 => x"72656164",
    19998 => x"28307825", 19999 => x"782c2025", 20000 => x"69293a20",
    20001 => x"72657375", 20002 => x"6c74203d", 20003 => x"2025690a",
    20004 => x"00000000", 20005 => x"64657669", 20006 => x"63652025",
    20007 => x"693a2025", 20008 => x"30387825", 20009 => x"3038780a",
    20010 => x"00000000", 20011 => x"74656d70", 20012 => x"3a202564",
    20013 => x"2e253034", 20014 => x"640a0000", 20015 => x"77310000",
    20016 => x"77317200", 20017 => x"77317700", 20018 => x"456e6162",
    20019 => x"6c655461", 20020 => x"67676572", 20021 => x"20256420",
    20022 => x"25640a00", 20023 => x"25733a20", 20024 => x"63682025",
    20025 => x"642c204f", 20026 => x"43455220", 20027 => x"30782578",
    20028 => x"2c205243", 20029 => x"45522030", 20030 => x"7825780a",
    20031 => x"00000000", 20032 => x"3c756e6b", 20033 => x"6e6f776e",
    20034 => x"3e000000", 20035 => x"4558543a", 20036 => x"20444d54",
    20037 => x"44206c6f", 20038 => x"636b6564", 20039 => x"2e0a0000",
    20040 => x"4558543a", 20041 => x"20435379", 20042 => x"6e632063",
    20043 => x"6f6d706c", 20044 => x"6574652e", 20045 => x"0a000000",
    20046 => x"4558543a", 20047 => x"20416c69", 20048 => x"676e2074",
    20049 => x"61726765", 20050 => x"74202564", 20051 => x"2c207374",
    20052 => x"65702025", 20053 => x"642e0a00", 20054 => x"4558543a",
    20055 => x"20416c69", 20056 => x"676e2064", 20057 => x"6f6e652e",
    20058 => x"0a000000", 20059 => x"72656620", 20060 => x"2564206f",
    20061 => x"75742025", 20062 => x"64206964", 20063 => x"78202578",
    20064 => x"200a0000", 20065 => x"4d504c4c", 20066 => x"5f537461",
    20067 => x"7274205b", 20068 => x"64616320", 20069 => x"25645d0a",
    20070 => x"00000000", 20071 => x"736f6674", 20072 => x"706c6c3a",
    20073 => x"20617474", 20074 => x"656d7074", 20075 => x"696e6720",
    20076 => x"746f2065", 20077 => x"6e61626c", 20078 => x"6520474d",
    20079 => x"206d6f64", 20080 => x"65206f6e", 20081 => x"206e6f6e",
    20082 => x"2d474d20", 20083 => x"68617264", 20084 => x"77617265",
    20085 => x"2e0a0000", 20086 => x"736f6674", 20087 => x"706c6c3a",
    20088 => x"206d6f64", 20089 => x"65202573", 20090 => x"2c202564",
    20091 => x"20726566", 20092 => x"20636861", 20093 => x"6e6e656c",
    20094 => x"732c2025", 20095 => x"64206f75", 20096 => x"74206368",
    20097 => x"616e6e65", 20098 => x"6c730a00", 20099 => x"43616e27",
    20100 => x"74207374", 20101 => x"61727420", 20102 => x"6368616e",
    20103 => x"6e656c20", 20104 => x"25642c20", 20105 => x"74686520",
    20106 => x"504c4c20", 20107 => x"6973206e", 20108 => x"6f742072",
    20109 => x"65616479", 20110 => x"0a000000", 20111 => x"736f6674",
    20112 => x"706c6c3a", 20113 => x"20697271", 20114 => x"73202564",
    20115 => x"20736571", 20116 => x"20257320", 20117 => x"6d6f6465",
    20118 => x"20256420", 20119 => x"616c6967", 20120 => x"6e6d656e",
    20121 => x"745f7374", 20122 => x"61746520", 20123 => x"25642048",
    20124 => x"4c256420", 20125 => x"4d4c2564", 20126 => x"2048593d",
    20127 => x"2564204d", 20128 => x"593d2564", 20129 => x"2044656c",
    20130 => x"436e743d", 20131 => x"25640a00", 20132 => x"456e6162",
    20133 => x"6c696e67", 20134 => x"20707472", 20135 => x"61636b65",
    20136 => x"72206368", 20137 => x"616e6e65", 20138 => x"6c3a2025",
    20139 => x"640a0000", 20140 => x"44697361", 20141 => x"626c696e",
    20142 => x"67207074", 20143 => x"7261636b", 20144 => x"65722074",
    20145 => x"61676765", 20146 => x"723a2025", 20147 => x"640a0000",
    20148 => x"6c6f636b", 20149 => x"696e6700", 20150 => x"616c6967",
    20151 => x"6e696e67", 20152 => x"00000000", 20153 => x"736f6674",
    20154 => x"706c6c3a", 20155 => x"20646973", 20156 => x"61626c65",
    20157 => x"64206175", 20158 => x"78206368", 20159 => x"616e6e65",
    20160 => x"6c202564", 20161 => x"0a000000", 20162 => x"736f6674",
    20163 => x"706c6c3a", 20164 => x"20656e61", 20165 => x"626c6564",
    20166 => x"20617578", 20167 => x"20636861", 20168 => x"6e6e656c",
    20169 => x"2025640a", 20170 => x"00000000", 20171 => x"736f6674",
    20172 => x"706c6c3a", 20173 => x"20636861", 20174 => x"6e6e656c",
    20175 => x"20256420", 20176 => x"6c6f636b", 20177 => x"6564205b",
    20178 => x"616c6967", 20179 => x"6e696e67", 20180 => x"20402025",
    20181 => x"64207073", 20182 => x"5d0a0000", 20183 => x"736f6674",
    20184 => x"706c6c3a", 20185 => x"20636861", 20186 => x"6e6e656c",
    20187 => x"20256420", 20188 => x"70686173", 20189 => x"6520616c",
    20190 => x"69676e65", 20191 => x"640a0000", 20192 => x"736f6674",
    20193 => x"706c6c3a", 20194 => x"20617578", 20195 => x"20636861",
    20196 => x"6e6e656c", 20197 => x"20256420", 20198 => x"6f72206d",
    20199 => x"706c6c20", 20200 => x"6c6f7374", 20201 => x"206c6f63",
    20202 => x"6b0a0000", 20203 => x"536f6674", 20204 => x"504c4c20",
    20205 => x"56434f20", 20206 => x"46726571", 20207 => x"75656e63",
    20208 => x"792f4150", 20209 => x"52207465", 20210 => x"73743a0a",
    20211 => x"00000000", 20212 => x"444d5444", 20213 => x"2056434f",
    20214 => x"3a20204c", 20215 => x"6f773d25", 20216 => x"6420487a",
    20217 => x"2048693d", 20218 => x"25642048", 20219 => x"7a2c2041",
    20220 => x"5052203d", 20221 => x"20256420", 20222 => x"70706d2e",
    20223 => x"0a000000", 20224 => x"52454620", 20225 => x"56434f3a",
    20226 => x"2020204c", 20227 => x"6f773d25", 20228 => x"6420487a",
    20229 => x"2048693d", 20230 => x"25642048", 20231 => x"7a2c2041",
    20232 => x"5052203d", 20233 => x"20256420", 20234 => x"70706d2e",
    20235 => x"0a000000", 20236 => x"45585420", 20237 => x"636c6f63",
    20238 => x"6b3a2046", 20239 => x"7265713d", 20240 => x"25642048",
    20241 => x"7a0a0000", 20242 => x"73746172", 20243 => x"742d6578",
    20244 => x"74000000", 20245 => x"77616974", 20246 => x"2d657874",
    20247 => x"00000000", 20248 => x"73746172", 20249 => x"742d6865",
    20250 => x"6c706572", 20251 => x"00000000", 20252 => x"77616974",
    20253 => x"2d68656c", 20254 => x"70657200", 20255 => x"73746172",
    20256 => x"742d6d61", 20257 => x"696e0000", 20258 => x"77616974",
    20259 => x"2d6d6169", 20260 => x"6e000000", 20261 => x"72656164",
    20262 => x"79000000", 20263 => x"636c6561", 20264 => x"722d6461",
    20265 => x"63730000", 20266 => x"77616974", 20267 => x"2d636c65",
    20268 => x"61722d64", 20269 => x"61637300", 20270 => x"66726565",
    20271 => x"6d617374", 20272 => x"65720000", 20273 => x"53746163",
    20274 => x"6b206f76", 20275 => x"6572666c", 20276 => x"6f77210a",
    20277 => x"00000000", 20278 => x"badc0ffe", 20279 => x"3b9ac9ff",
    20280 => x"3b9aca00", 20281 => x"000f4240", 20282 => x"00080030",
    20283 => x"d4a51000", 20284 => x"c4653600", 20285 => x"7ffffffe",
    20286 => x"80000001", 20287 => x"fff06000", 20288 => x"0007d000",
    20289 => x"41c64e6d", 20290 => x"00010043", 20291 => x"00010044",
    20292 => x"00015180", 20293 => x"000186a0", 20294 => x"00062000",
    20295 => x"005ee000", 20296 => x"01000001", 20297 => x"11223344",
    20298 => x"e0001fff", 20299 => x"0fffffff", 20300 => x"059682f0",
    20301 => x"0ee6b27f", 20302 => x"7fffffff", 20303 => x"01312d02",
    20304 => x"01312d0a", 20305 => x"c0a80001", 20306 => x"4b002f40",
    20307 => x"003d0137", 20308 => x"8000001f", 20309 => x"009895b6",
    20310 => x"c4000001", 20311 => x"00ffffff", 20312 => x"fffdb610",
    20313 => x"000249f0", 20314 => x"05f5e100", 20315 => x"0bebc200",
    20316 => x"fa0a1f00", 20317 => x"fff0bdc0", 20318 => x"01312d03",
    20319 => x"03b9aca0", 20320 => x"07735940", 20321 => x"5344422d",
    20322 => x"011b1900", 20323 => x"00000000", 20324 => x"70705f64",
    20325 => x"6961675f", 20326 => x"70617273", 20327 => x"65000000",
    20328 => x"00000000", 20329 => x"00011e74", 20330 => x"00011e80",
    20331 => x"00011e90", 20332 => x"00011e9c", 20333 => x"00011ea8",
    20334 => x"00011eb4", 20335 => x"00011ec0", 20336 => x"00002094",
    20337 => x"00002104", 20338 => x"000023bc", 20339 => x"000023bc",
    20340 => x"000023bc", 20341 => x"000023bc", 20342 => x"000023bc",
    20343 => x"000023bc", 20344 => x"00002180", 20345 => x"000021f0",
    20346 => x"000023bc", 20347 => x"00002284", 20348 => x"00002390",
    20349 => x"77727063", 20350 => x"5f74696d", 20351 => x"655f6164",
    20352 => x"6a757374", 20353 => x"5f6f6666", 20354 => x"73657400",
    20355 => x"77727063", 20356 => x"5f74696d", 20357 => x"655f6164",
    20358 => x"6a757374", 20359 => x"00000000", 20360 => x"77727063",
    20361 => x"5f74696d", 20362 => x"655f7365", 20363 => x"74000000",
    20364 => x"77727063", 20365 => x"5f74696d", 20366 => x"655f6765",
    20367 => x"74000000", 20368 => x"77727063", 20369 => x"5f6e6574",
    20370 => x"5f73656e", 20371 => x"64000000", 20372 => x"77725f75",
    20373 => x"6e706163", 20374 => x"6b5f616e", 20375 => x"6e6f756e",
    20376 => x"63650000", 20377 => x"77725f70", 20378 => x"61636b5f",
    20379 => x"616e6e6f", 20380 => x"756e6365", 20381 => x"00000000",
    20382 => x"77725f68", 20383 => x"616e646c", 20384 => x"655f666f",
    20385 => x"6c6c6f77", 20386 => x"75700000", 20387 => x"77725f68",
    20388 => x"616e646c", 20389 => x"655f616e", 20390 => x"6e6f756e",
    20391 => x"63650000", 20392 => x"77725f65", 20393 => x"78656375",
    20394 => x"74655f73", 20395 => x"6c617665", 20396 => x"00000000",
    20397 => x"77725f73", 20398 => x"31000000", 20399 => x"77725f68",
    20400 => x"616e646c", 20401 => x"655f7265", 20402 => x"73700000",
    20403 => x"77725f6e", 20404 => x"65775f73", 20405 => x"6c617665",
    20406 => x"00000000", 20407 => x"77725f6d", 20408 => x"61737465",
    20409 => x"725f6d73", 20410 => x"67000000", 20411 => x"77725f6c",
    20412 => x"69737465", 20413 => x"6e696e67", 20414 => x"00000000",
    20415 => x"77725f6f", 20416 => x"70656e00", 20417 => x"77725f69",
    20418 => x"6e697400", 20419 => x"0000398c", 20420 => x"000039b4",
    20421 => x"000039d4", 20422 => x"00003a44", 20423 => x"00003a64",
    20424 => x"00003a80", 20425 => x"00003aa0", 20426 => x"00003b2c",
    20427 => x"00003b4c", 20428 => x"77725f63", 20429 => x"616c6962",
    20430 => x"72617469", 20431 => x"6f6e0000", 20432 => x"00004f30",
    20433 => x"00004f18", 20434 => x"00004f58", 20435 => x"00005068",
    20436 => x"00004fac", 20437 => x"000127f0", 20438 => x"00012924",
    20439 => x"00012930", 20440 => x"0001293c", 20441 => x"00012948",
    20442 => x"00012954", 20443 => x"77725f73", 20444 => x"6572766f",
    20445 => x"5f757064", 20446 => x"61746500", 20447 => x"70705f69",
    20448 => x"6e697469", 20449 => x"616c697a", 20450 => x"696e6700",
    20451 => x"73745f63", 20452 => x"6f6d5f73", 20453 => x"6c617665",
    20454 => x"5f68616e", 20455 => x"646c655f", 20456 => x"666f6c6c",
    20457 => x"6f777570", 20458 => x"00000000", 20459 => x"626d635f",
    20460 => x"64617461", 20461 => x"7365745f", 20462 => x"636d7000",
    20463 => x"626d635f", 20464 => x"73746174", 20465 => x"655f6465",
    20466 => x"63697369", 20467 => x"6f6e0000", 20468 => x"63466965",
    20469 => x"6c645f74", 20470 => x"6f5f5469", 20471 => x"6d65496e",
    20472 => x"7465726e", 20473 => x"616c0000", 20474 => x"00011d70",
    20475 => x"00013268", 20476 => x"0001296c", 20477 => x"00012484",
    20478 => x"0000001f", 20479 => x"0000001c", 20480 => x"0000001f",
    20481 => x"0000001e", 20482 => x"0000001f", 20483 => x"0000001e",
    20484 => x"0000001f", 20485 => x"0000001f", 20486 => x"0000001e",
    20487 => x"0000001f", 20488 => x"0000001e", 20489 => x"0000001f",
    20490 => x"0000001f", 20491 => x"0000001d", 20492 => x"0000001f",
    20493 => x"0000001e", 20494 => x"0000001f", 20495 => x"0000001e",
    20496 => x"0000001f", 20497 => x"0000001f", 20498 => x"0000001e",
    20499 => x"0000001f", 20500 => x"0000001e", 20501 => x"0000001f",
    20502 => x"000134e0", 20503 => x"000134e4", 20504 => x"000134e8",
    20505 => x"000134ec", 20506 => x"000134f0", 20507 => x"000134f4",
    20508 => x"000134f8", 20509 => x"000134fc", 20510 => x"00013500",
    20511 => x"00013504", 20512 => x"00013508", 20513 => x"0001350c",
    20514 => x"00013510", 20515 => x"00013514", 20516 => x"00013518",
    20517 => x"0001351c", 20518 => x"00013520", 20519 => x"00013524",
    20520 => x"00013528", 20521 => x"6765745f", 20522 => x"70657273",
    20523 => x"69737465", 20524 => x"6e745f6d", 20525 => x"61630000",
    20526 => x"73706c6c", 20527 => x"5f656e61", 20528 => x"626c655f",
    20529 => x"74616767", 20530 => x"65720000", 20531 => x"0000ed48",
    20532 => x"0000edd0", 20533 => x"0000ee04", 20534 => x"0000eea4",
    20535 => x"0000ef28", 20536 => x"0000ef48", 20537 => x"0000ee30",
    20538 => x"0000ed6c", 20539 => x"0000ecd4", 20540 => x"0000ed04",
    20541 => x"00000000", 20542 => x"00000000", 20543 => x"00000000",
    20544 => x"00000000", 20545 => x"00000001", 20546 => x"00000001",
    20547 => x"00000001", 20548 => x"00000001", 20549 => x"00000000",
    20550 => x"00000000", 20551 => x"00000000", 20552 => x"0000ece8",
    20553 => x"0000ece8", 20554 => x"00000000", 20555 => x"0000d9d0",
    20556 => x"00000000", 20557 => x"0000fba0", 20558 => x"0000fbc0",
    20559 => x"0000fbcc", 20560 => x"0000fbdc", 20561 => x"0000fbfc",
    20562 => x"0000fc0c", 20563 => x"0000fc60", 20564 => x"0000fc24",
    20565 => x"0000fb34", 20566 => x"0000fb78", 20567 => x"00000001",
    20568 => x"00013c48", 20569 => x"00000002", 20570 => x"00013c54",
    20571 => x"00000003", 20572 => x"00013c60", 20573 => x"00000004",
    20574 => x"00013c70", 20575 => x"00000005", 20576 => x"00013c7c",
    20577 => x"00000006", 20578 => x"00013c88", 20579 => x"00000007",
    20580 => x"0001245c", 20581 => x"00000008", 20582 => x"00013c94",
    20583 => x"00000009", 20584 => x"00013c9c", 20585 => x"0000000a",
    20586 => x"00013ca8", 20587 => x"00000000", 20588 => x"00000000",
    20589 => x"00013cd4", 20590 => x"00013268", 20591 => x"00013cb8",
    20592 => x"00012484", 20593 => x"0001245c", 20594 => x"00000000",
    20595 => x"00000000", 20596 => x"00000000", 20597 => x"00000000",
    20598 => x"00010000", 20599 => x"00000000", 20600 => x"00000000",
    20601 => x"00000000", 20602 => x"00020100", 20603 => x"00000000",
    20604 => x"00000000", 20605 => x"00000000", 20606 => x"00030101",
    20607 => x"00000000", 20608 => x"00000000", 20609 => x"00000000",
    20610 => x"00040201", 20611 => x"01000000", 20612 => x"00000000",
    20613 => x"00000000", 20614 => x"00050201", 20615 => x"01010000",
    20616 => x"00000000", 20617 => x"00000000", 20618 => x"00060302",
    20619 => x"01010100", 20620 => x"00000000", 20621 => x"00000000",
    20622 => x"00070302", 20623 => x"01010101", 20624 => x"00000000",
    20625 => x"00000000", 20626 => x"00080402", 20627 => x"02010101",
    20628 => x"01000000", 20629 => x"00000000", 20630 => x"00090403",
    20631 => x"02010101", 20632 => x"01010000", 20633 => x"00000000",
    20634 => x"000a0503", 20635 => x"02020101", 20636 => x"01010100",
    20637 => x"00000000", 20638 => x"000b0503", 20639 => x"02020101",
    20640 => x"01010101", 20641 => x"00000000", 20642 => x"000c0604",
    20643 => x"03020201", 20644 => x"01010101", 20645 => x"01000000",
    20646 => x"000d0604", 20647 => x"03020201", 20648 => x"01010101",
    20649 => x"01010000", 20650 => x"000e0704", 20651 => x"03020202",
    20652 => x"01010101", 20653 => x"01010100", 20654 => x"000f0705",
    20655 => x"03030202", 20656 => x"01010101", 20657 => x"01010101",
    20658 => x"fefefeff", 20659 => x"80808080", 20660 => x"00202020",
    20661 => x"20202020", 20662 => x"20202828", 20663 => x"28282820",
    20664 => x"20202020", 20665 => x"20202020", 20666 => x"20202020",
    20667 => x"20202020", 20668 => x"20881010", 20669 => x"10101010",
    20670 => x"10101010", 20671 => x"10101010", 20672 => x"10040404",
    20673 => x"04040404", 20674 => x"04040410", 20675 => x"10101010",
    20676 => x"10104141", 20677 => x"41414141", 20678 => x"01010101",
    20679 => x"01010101", 20680 => x"01010101", 20681 => x"01010101",
    20682 => x"01010101", 20683 => x"10101010", 20684 => x"10104242",
    20685 => x"42424242", 20686 => x"02020202", 20687 => x"02020202",
    20688 => x"02020202", 20689 => x"02020202", 20690 => x"02020202",
    20691 => x"10101010", 20692 => x"20000000", 20693 => x"00000000",
    20694 => x"00000000", 20695 => x"00000000", 20696 => x"00000000",
    20697 => x"00000000", 20698 => x"00000000", 20699 => x"00000000",
    20700 => x"00000000", 20701 => x"00000000", 20702 => x"00000000",
    20703 => x"00000000", 20704 => x"00000000", 20705 => x"00000000",
    20706 => x"00000000", 20707 => x"00000000", 20708 => x"00000000",
    20709 => x"00000000", 20710 => x"00000000", 20711 => x"00000000",
    20712 => x"00000000", 20713 => x"00000000", 20714 => x"00000000",
    20715 => x"00000000", 20716 => x"00000000", 20717 => x"00000000",
    20718 => x"00000000", 20719 => x"00000000", 20720 => x"00000000",
    20721 => x"00000000", 20722 => x"00000000", 20723 => x"00000000",
    20724 => x"00000000", 20725 => x"00000000", 20726 => x"00014d88",
    20727 => x"00014da8", 20728 => x"00014db8", 20729 => x"000003e8",
    20730 => x"00000001", 20731 => x"046362a0", 20732 => x"00000955",
    20733 => x"ffffffff", 20734 => x"000143fc", 20735 => x"00000000",
    20736 => x"00000000", 20737 => x"00000000", 20738 => x"00000000",
    20739 => x"00000000", 20740 => x"00000000", 20741 => x"00000000",
    20742 => x"00000000", 20743 => x"00014770", 20744 => x"00014890",
    20745 => x"00014874", 20746 => x"00014f34", 20747 => x"00014fb4",
    20748 => x"00000000", 20749 => x"00000000", 20750 => x"00000000",
    20751 => x"00000000", 20752 => x"00000000", 20753 => x"00000000",
    20754 => x"00000000", 20755 => x"00000000", 20756 => x"00000000",
    20757 => x"00000000", 20758 => x"00000000", 20759 => x"00000000",
    20760 => x"00000000", 20761 => x"00000000", 20762 => x"00000000",
    20763 => x"00000000", 20764 => x"00000000", 20765 => x"00000000",
    20766 => x"00000000", 20767 => x"00000000", 20768 => x"00000000",
    20769 => x"00000000", 20770 => x"00000000", 20771 => x"00000000",
    20772 => x"00000000", 20773 => x"00000000", 20774 => x"00000000",
    20775 => x"00000000", 20776 => x"00000000", 20777 => x"00000000",
    20778 => x"00000000", 20779 => x"00000000", 20780 => x"00000000",
    20781 => x"00000000", 20782 => x"00000000", 20783 => x"00000000",
    20784 => x"00000000", 20785 => x"00000000", 20786 => x"00000000",
    20787 => x"00000000", 20788 => x"00000000", 20789 => x"00000000",
    20790 => x"00000000", 20791 => x"00000000", 20792 => x"00000000",
    20793 => x"00000000", 20794 => x"00000000", 20795 => x"00000000",
    20796 => x"00000000", 20797 => x"00000000", 20798 => x"00000000",
    20799 => x"00000000", 20800 => x"00000000", 20801 => x"00000000",
    20802 => x"00000000", 20803 => x"00000000", 20804 => x"00000000",
    20805 => x"00000000", 20806 => x"00000000", 20807 => x"00000000",
    20808 => x"00000000", 20809 => x"00000000", 20810 => x"00000000",
    20811 => x"00000000", 20812 => x"00000000", 20813 => x"00000000",
    20814 => x"00000000", 20815 => x"00000000", 20816 => x"00000000",
    20817 => x"00000000", 20818 => x"00000000", 20819 => x"00000000",
    20820 => x"00000000", 20821 => x"00000000", 20822 => x"00000000",
    20823 => x"00000000", 20824 => x"00000000", 20825 => x"00000000",
    20826 => x"00000000", 20827 => x"00000000", 20828 => x"00000000",
    20829 => x"00000000", 20830 => x"00000000", 20831 => x"00000000",
    20832 => x"00000000", 20833 => x"00000000", 20834 => x"00000000",
    20835 => x"00000000", 20836 => x"00000000", 20837 => x"00000000",
    20838 => x"00000000", 20839 => x"00000000", 20840 => x"00000000",
    20841 => x"00000000", 20842 => x"00000000", 20843 => x"00000000",
    20844 => x"00000000", 20845 => x"00000000", 20846 => x"00000000",
    20847 => x"00000000", 20848 => x"00000000", 20849 => x"00000000",
    20850 => x"00000000", 20851 => x"00000000", 20852 => x"00000000",
    20853 => x"00000000", 20854 => x"00000000", 20855 => x"00000000",
    20856 => x"00000000", 20857 => x"00000000", 20858 => x"00000000",
    20859 => x"00000000", 20860 => x"00000000", 20861 => x"00000000",
    20862 => x"00000000", 20863 => x"00000000", 20864 => x"00000000",
    20865 => x"00000000", 20866 => x"00000000", 20867 => x"00000000",
    20868 => x"00000000", 20869 => x"00000000", 20870 => x"00000000",
    20871 => x"00000000", 20872 => x"00000000", 20873 => x"00000000",
    20874 => x"00000000", 20875 => x"00000000", 20876 => x"00000000",
    20877 => x"00000000", 20878 => x"00000000", 20879 => x"00000000",
    20880 => x"00000000", 20881 => x"00000000", 20882 => x"00000000",
    20883 => x"00000000", 20884 => x"00000000", 20885 => x"00000000",
    20886 => x"00000000", 20887 => x"00000000", 20888 => x"00000000",
    20889 => x"00000000", 20890 => x"00000000", 20891 => x"00000000",
    20892 => x"00000000", 20893 => x"00000000", 20894 => x"00000000",
    20895 => x"00000000", 20896 => x"00000000", 20897 => x"00000000",
    20898 => x"00000000", 20899 => x"00000000", 20900 => x"00000000",
    20901 => x"00000000", 20902 => x"00000000", 20903 => x"00000000",
    20904 => x"00000000", 20905 => x"00000000", 20906 => x"00000000",
    20907 => x"00000000", 20908 => x"00000000", 20909 => x"00000000",
    20910 => x"00000000", 20911 => x"00000000", 20912 => x"00000000",
    20913 => x"000147b8", 20914 => x"00000000", 20915 => x"00000000",
    20916 => x"00000000", 20917 => x"00000000", 20918 => x"00000000",
    20919 => x"00000000", 20920 => x"00000000", 20921 => x"00000000",
    20922 => x"00000000", 20923 => x"00000000", 20924 => x"00000000",
    20925 => x"00000000", 20926 => x"00000000", 20927 => x"00000000",
    20928 => x"00000000", 20929 => x"00000000", 20930 => x"00000000",
    20931 => x"00000000", 20932 => x"00000000", 20933 => x"00000000",
    20934 => x"00000000", 20935 => x"00000000", 20936 => x"00000000",
    20937 => x"00000000", 20938 => x"00000000", 20939 => x"00011f64",
    20940 => x"00011f64", 20941 => x"00000000", 20942 => x"00000001",
    20943 => x"00000000", 20944 => x"00000000", 20945 => x"00000000",
    20946 => x"00000000", 20947 => x"00000000", 20948 => x"00000000",
    20949 => x"00000000", 20950 => x"00000000", 20951 => x"00000000",
    20952 => x"00000000", 20953 => x"00000000", 20954 => x"00000000",
    20955 => x"00000000", 20956 => x"000143fc", 20957 => x"00015038",
    20958 => x"00000000", 20959 => x"00015078", 20960 => x"00015094",
    20961 => x"000150c4", 20962 => x"000150e4", 20963 => x"00000000",
    20964 => x"00000000", 20965 => x"00000000", 20966 => x"00000000",
    20967 => x"00000000", 20968 => x"00000000", 20969 => x"00000000",
    20970 => x"00000000", 20971 => x"00000000", 20972 => x"00015108",
    20973 => x"000003e8", 20974 => x"00000000", 20975 => x"00000000",
    20976 => x"00000000", 20977 => x"00000000", 20978 => x"000147cc",
    20979 => x"00014838", 20980 => x"00000000", 20981 => x"00000000",
    20982 => x"00000000", 20983 => x"00000000", 20984 => x"00000000",
    20985 => x"00000000", 20986 => x"00000000", 20987 => x"00000000",
    20988 => x"00000000", 20989 => x"00000000", 20990 => x"00000000",
    20991 => x"00000000", 20992 => x"00000000", 20993 => x"00000000",
    20994 => x"00000000", 20995 => x"00000000", 20996 => x"00000000",
    20997 => x"00000000", 20998 => x"00000000", 20999 => x"00000000",
    21000 => x"00000000", 21001 => x"00000000", 21002 => x"00000000",
    21003 => x"00000000", 21004 => x"00000000", 21005 => x"00000000",
    21006 => x"000015cc", 21007 => x"00001600", 21008 => x"00001680",
    21009 => x"00001688", 21010 => x"000016e0", 21011 => x"0000170c",
    21012 => x"00001764", 21013 => x"00001788", 21014 => x"0000184c",
    21015 => x"00001854", 21016 => x"0000185c", 21017 => x"000018c0",
    21018 => x"000018dc", 21019 => x"000016ac", 21020 => x"00000000",
    21021 => x"00002844", 21022 => x"000027c8", 21023 => x"0000276c",
    21024 => x"00002714", 21025 => x"00000000", 21026 => x"00000000",
    21027 => x"000026e4", 21028 => x"00002ad0", 21029 => x"00002ab0",
    21030 => x"000029e0", 21031 => x"000028c4", 21032 => x"00000000",
    21033 => x"00000001", 21034 => x"00012444", 21035 => x"00005244",
    21036 => x"00000002", 21037 => x"00012454", 21038 => x"00005410",
    21039 => x"00000003", 21040 => x"0001245c", 21041 => x"000054cc",
    21042 => x"00000004", 21043 => x"00012468", 21044 => x"000054dc",
    21045 => x"00000006", 21046 => x"0001296c", 21047 => x"00005688",
    21048 => x"00000008", 21049 => x"00012474", 21050 => x"000059c8",
    21051 => x"00000009", 21052 => x"00012484", 21053 => x"00005a3c",
    21054 => x"00000064", 21055 => x"0001248c", 21056 => x"000033c4",
    21057 => x"00000066", 21058 => x"000124a4", 21059 => x"0000353c",
    21060 => x"00000065", 21061 => x"000124b8", 21062 => x"00003668",
    21063 => x"00000067", 21064 => x"000124d0", 21065 => x"0000376c",
    21066 => x"00000068", 21067 => x"000124e8", 21068 => x"00003898",
    21069 => x"00000069", 21070 => x"000124f8", 21071 => x"00003bb4",
    21072 => x"0000006a", 21073 => x"00012508", 21074 => x"00003cc8",
    21075 => x"0000006b", 21076 => x"0001251c", 21077 => x"00003e4c",
    21078 => x"00000000", 21079 => x"00000000", 21080 => x"00000000",
    21081 => x"00000001", 21082 => x"00012444", 21083 => x"00005244",
    21084 => x"00000002", 21085 => x"00012454", 21086 => x"00005410",
    21087 => x"00000003", 21088 => x"0001245c", 21089 => x"000054cc",
    21090 => x"00000004", 21091 => x"00012468", 21092 => x"000054dc",
    21093 => x"00000005", 21094 => x"00012968", 21095 => x"000055f4",
    21096 => x"00000006", 21097 => x"0001296c", 21098 => x"00005688",
    21099 => x"00000007", 21100 => x"00012974", 21101 => x"00005904",
    21102 => x"00000008", 21103 => x"00012474", 21104 => x"000059c8",
    21105 => x"00000009", 21106 => x"00012484", 21107 => x"00005a3c",
    21108 => x"00000000", 21109 => x"00000000", 21110 => x"00000000",
    21111 => x"00002dc8", 21112 => x"00002ce8", 21113 => x"00000000",
    21114 => x"00002ca0", 21115 => x"00003160", 21116 => x"00003118",
    21117 => x"0000302c", 21118 => x"00002c10", 21119 => x"00002b84",
    21120 => x"00002fb4", 21121 => x"00002f3c", 21122 => x"00002ed4",
    21123 => x"00002e68", 21124 => x"00000001", 21125 => x"00012b80",
    21126 => x"00012b88", 21127 => x"00012b94", 21128 => x"00012ba0",
    21129 => x"00000000", 21130 => x"00000000", 21131 => x"00000000",
    21132 => x"00000000", 21133 => x"00012bc4", 21134 => x"00012bac",
    21135 => x"00012bb8", 21136 => x"00012bd0", 21137 => x"00012bdc",
    21138 => x"00012be8", 21139 => x"00000000", 21140 => x"00000000",
    21141 => x"00012f10", 21142 => x"00012f20", 21143 => x"00012f2c",
    21144 => x"00012f40", 21145 => x"00012f54", 21146 => x"00012f64",
    21147 => x"00012f70", 21148 => x"00012f7c", 21149 => x"bbfef060",
    21150 => x"00000000", 21151 => x"00000000", 21152 => x"00000000",
    21153 => x"00000000", 21154 => x"00000000", 21155 => x"00000000",
    21156 => x"00000000", 21157 => x"00000000", 21158 => x"00000000",
    21159 => x"00000000", 21160 => x"00000000", 21161 => x"00000000",
    21162 => x"00000001", 21163 => x"00000000", 21164 => x"000a03e8",
    21165 => x"00060100", 21166 => x"80800000", 21167 => x"00000000",
    21168 => x"00000000", 21169 => x"00000000", 21170 => x"00000000",
    21171 => x"00000000", 21172 => x"00000000", 21173 => x"44332211",
    21174 => x"00000000", 21175 => x"04000000", 21176 => x"1b8046e2",
    21177 => x"01000000", 21178 => x"9800cfea", 21179 => x"01000000",
    21180 => x"188157f3", 21181 => x"01000000", 21182 => x"0be0ffff",
    21183 => x"01000000", 21184 => x"88e0ffff", 21185 => x"01000000",
    21186 => x"08e1ffff", 21187 => x"01000000", 21188 => x"136023e0",
    21189 => x"01000000", 21190 => x"900020e3", 21191 => x"01000000",
    21192 => x"100100e0", 21193 => x"01000000", 21194 => x"230300e1",
    21195 => x"01000000", 21196 => x"2be31ef1", 21197 => x"01000000",
    21198 => x"33c300e1", 21199 => x"01000000", 21200 => x"4be37ffb",
    21201 => x"01000000", 21202 => x"bb250060", 21203 => x"00000000",
    21204 => x"c3250260", 21205 => x"00000000", 21206 => x"59031000",
    21207 => x"04000000", 21208 => x"61611000", 21209 => x"04000000",
    21210 => x"78c19400", 21211 => x"04000000", 21212 => x"80ebbc00",
    21213 => x"04000000", 21214 => x"53097afd", 21215 => x"01000000",
    21216 => x"c3108001", 21217 => x"04000000", 21218 => x"e90a8001",
    21219 => x"04000000", 21220 => x"f9508103", 21221 => x"04000000",
    21222 => x"00000000", 21223 => x"08000000", 21224 => x"00000004",
    21225 => x"00000008", 21226 => x"00000100", 21227 => x"00000200",
    21228 => x"00016dcc", 21229 => x"00000000", 21230 => x"00000000",
    21231 => x"0000ce42", 21232 => x"ab28633a", 21233 => x"00000000",
    21234 => x"00016d00", 21235 => x"00000000", 21236 => x"00000000",
    21237 => x"0000ce42", 21238 => x"650c2d4f", 21239 => x"00000000",
    21240 => x"00016dd4", 21241 => x"00000000", 21242 => x"00000000",
    21243 => x"0000ce42", 21244 => x"65158dc0", 21245 => x"00000000",
    21246 => x"00016d10", 21247 => x"00000000", 21248 => x"00000000",
    21249 => x"0000ce42", 21250 => x"de0d8ced", 21251 => x"00000000",
    21252 => x"00016dd0", 21253 => x"00000000", 21254 => x"00000000",
    21255 => x"0000ce42", 21256 => x"ff07fc47", 21257 => x"00000000",
    21258 => x"00016da4", 21259 => x"00000000", 21260 => x"00000000",
    21261 => x"0000ce42", 21262 => x"e2d13d04", 21263 => x"00000000",
    21264 => x"00016da0", 21265 => x"00000000", 21266 => x"00000000",
    21267 => x"0000ce42", 21268 => x"779c5443", 21269 => x"00000000",
    21270 => x"00016dc8", 21271 => x"00000000", 21272 => x"00000000",
    21273 => x"00000651", 21274 => x"68202b22", 21275 => x"00000000",
    21276 => x"00016dc0", 21277 => x"00000000", 21278 => x"00000000",
    21279 => x"00001103", 21280 => x"c0413599", 21281 => x"00000000",
    21282 => x"000136cc", 21283 => x"00000000", 21284 => x"00000001",
    21285 => x"00030000", 21286 => x"00000004", 21287 => x"00000000",
    21288 => x"00000000", 21289 => x"00000000", 21290 => x"00000000",
    21291 => x"00000000", 21292 => x"00000000", 21293 => x"00000000",
    21294 => x"00000000", 21295 => x"00000000", 21296 => x"00000000",
    21297 => x"00000000", 21298 => x"00000000", 21299 => x"00000000",
    21300 => x"00000000", 21301 => x"00000000", 21302 => x"00000000",
    21303 => x"00000000", 21304 => x"00000000", 21305 => x"00000000",
    21306 => x"00000000", 21307 => x"00000000", 21308 => x"00000000",
    21309 => x"00000000", 21310 => x"00000000", 21311 => x"00000000",
    21312 => x"00000000", 21313 => x"00000000", 21314 => x"00000000",
    21315 => x"00000000", 21316 => x"00000000", 21317 => x"00000000",
    21318 => x"00000000", 21319 => x"00000000", 21320 => x"00000000",
    21321 => x"00000000", 21322 => x"00000000", 21323 => x"00000000",
    21324 => x"00000000", 21325 => x"00000000", 21326 => x"00000000",
    21327 => x"00000000", 21328 => x"0000de94", 21329 => x"0000dec8",
    21330 => x"0000def8", 21331 => x"ffffffff", 21332 => x"000142d0",
    21333 => x"5b1157a7", 21334 => x"00000002", 21335 => x"00000000",
    21336 => x"00000000", 21337 => x"00000000", 21338 => x"00000000",
    21339 => x"00000000", 21340 => x"00000000", 21341 => x"00000000",
    21342 => x"00000000", 21343 => x"00000000", 21344 => x"00000000",
    21345 => x"00000000", 21346 => x"77727063", 21347 => x"2d76332e",
    21348 => x"302d3130", 21349 => x"2d673138", 21350 => x"39653666",
    21351 => x"62000000", 21352 => x"00000000", 21353 => x"00000000",
    21354 => x"41756720", 21355 => x"32352032", 21356 => x"30313600",
    21357 => x"00000000", 21358 => x"31323a30", 21359 => x"303a3334",
    21360 => x"00000000", 21361 => x"00000000", 21362 => x"000130b8",
    21363 => x"000086c0", 21364 => x"0001310c", 21365 => x"00008774",
    21366 => x"00013238", 21367 => x"000089dc", 21368 => x"000130c8",
    21369 => x"00008d8c", 21370 => x"00013258", 21371 => x"00008e90",
    21372 => x"00013260", 21373 => x"00008ef0", 21374 => x"000132cc",
    21375 => x"00008f8c", 21376 => x"00013308", 21377 => x"00009064",
    21378 => x"00013310", 21379 => x"000091c0", 21380 => x"00013314",
    21381 => x"000091d8", 21382 => x"00013358", 21383 => x"00009254",
    21384 => x"000130bc", 21385 => x"0000936c", 21386 => x"000133e8",
    21387 => x"0000947c", 21388 => x"00013410", 21389 => x"00009528",
    21390 => x"00013434", 21391 => x"00009594", 21392 => x"00013474",
    21393 => x"000095f4", 21394 => x"00013490", 21395 => x"000096e8",
    21396 => x"000138bc", 21397 => x"0000e144", 21398 => x"000138c0",
    21399 => x"0000e048", 21400 => x"000138c4", 21401 => x"0000df4c",
    21402 => x"00000000", 21403 => x"00000000", 21404 => x"00000000",
    21405 => x"00000000", 21406 => x"00000000", 21407 => x"00000000",
    21408 => x"00000000", 21409 => x"00000000", 21410 => x"00000000",
    21411 => x"00000000", 21412 => x"00000000", 21413 => x"00000000",
    21414 => x"00000000", 21415 => x"00000000", 21416 => x"00000000",
    21417 => x"00000000", 21418 => x"00000000", 21419 => x"00000000",
    21420 => x"00000000", 21421 => x"00000000", 21422 => x"00000000",
    21423 => x"00000000", 21424 => x"00000000", 21425 => x"00000000",
    21426 => x"00000000", 21427 => x"00000000", 21428 => x"00000000",
    21429 => x"00000000", 21430 => x"00000000", 21431 => x"00000000",
    21432 => x"00000000", 21433 => x"00000000", 21434 => x"00000000",
    21435 => x"00000000", 21436 => x"00000000", 21437 => x"00000000",
    21438 => x"00000000", 21439 => x"00000000", 21440 => x"00000000",
    21441 => x"00000000", 21442 => x"00000000", 21443 => x"00000000",
    21444 => x"00000000", 21445 => x"00000000", 21446 => x"00000000",
    21447 => x"00000000", 21448 => x"00000000", 21449 => x"00000000",
    21450 => x"00000000", 21451 => x"00000000", 21452 => x"00000000",
    21453 => x"00000000", 21454 => x"00000000", 21455 => x"00000000",
    21456 => x"00000000", 21457 => x"00000000", 21458 => x"00000000",
    21459 => x"00000000", 21460 => x"00000000", 21461 => x"00000000",
    21462 => x"00000000", 21463 => x"00000000", 21464 => x"00000000",
    21465 => x"00000000", 21466 => x"00000000", 21467 => x"00000000",
    21468 => x"00000000", 21469 => x"00000000", 21470 => x"00000000",
    21471 => x"00000000", 21472 => x"00000000", 21473 => x"00000000",
    21474 => x"00000000", 21475 => x"00000000", 21476 => x"00000000",
    21477 => x"00000000", 21478 => x"00000000", 21479 => x"00000000",
    21480 => x"00000000", 21481 => x"00000000", 21482 => x"00000000",
    21483 => x"00000000", 21484 => x"00000000", 21485 => x"00000000",
    21486 => x"00000000", 21487 => x"00000000", 21488 => x"00000000",
    21489 => x"00000000", 21490 => x"00000000", 21491 => x"00000000",
    21492 => x"00000000", 21493 => x"00000000", 21494 => x"00000000",
    21495 => x"00000000", 21496 => x"00000000", 21497 => x"00000000",
    21498 => x"00000000", 21499 => x"00000000", 21500 => x"00000000",
    21501 => x"00000000", 21502 => x"00000000", 21503 => x"00000000",
    21504 => x"00000000", 21505 => x"00000000", 21506 => x"00000000",
    21507 => x"00000000", 21508 => x"00000000", 21509 => x"00000000",
    21510 => x"00000000", 21511 => x"00000000", 21512 => x"00000000",
    21513 => x"00000000", 21514 => x"00000000", 21515 => x"00000000",
    21516 => x"00000000", 21517 => x"00000000", 21518 => x"00000000",
    21519 => x"00000000", 21520 => x"00000000", 21521 => x"00000000",
    21522 => x"00000000", 21523 => x"00000000", 21524 => x"00000000",
    21525 => x"00000000", 21526 => x"00000000", 21527 => x"00000000",
    21528 => x"00000000", 21529 => x"00000000", 21530 => x"00000000",
    21531 => x"00000000", 21532 => x"00000000", 21533 => x"00000000",
    21534 => x"00000000", 21535 => x"00000000", 21536 => x"00000000",
    21537 => x"00000000", 21538 => x"00000000", 21539 => x"00000000",
    21540 => x"00000000", 21541 => x"00000000", 21542 => x"00000000",
    21543 => x"00000000", 21544 => x"00000000", 21545 => x"00000000",
    21546 => x"00000000", 21547 => x"00000000", 21548 => x"00000000",
    21549 => x"00000000", 21550 => x"00000000", 21551 => x"00000000",
    21552 => x"00000000", 21553 => x"00000000", 21554 => x"00000000",
    21555 => x"00000000", 21556 => x"00000000", 21557 => x"00000000",
    21558 => x"00000000", 21559 => x"00000000", 21560 => x"00000000",
    21561 => x"00000000", 21562 => x"00000000", 21563 => x"00000000",
    21564 => x"00000000", 21565 => x"00000000", 21566 => x"00000000",
    21567 => x"00000000", 21568 => x"00000000", 21569 => x"00000000",
    21570 => x"00000000", 21571 => x"00000000", 21572 => x"00000000",
    21573 => x"00000000", 21574 => x"00000000", 21575 => x"00000000",
    21576 => x"00000000", 21577 => x"00000000", 21578 => x"00000000",
    21579 => x"00000000", 21580 => x"00000000", 21581 => x"00000000",
    21582 => x"00000000", 21583 => x"00000000", 21584 => x"00000000",
    21585 => x"00000000", 21586 => x"00000000", 21587 => x"00000000",
    21588 => x"00000000", 21589 => x"00000000", 21590 => x"00000000",
    21591 => x"00000000", 21592 => x"00000000", 21593 => x"00000000",
    21594 => x"00000000", 21595 => x"00000000", 21596 => x"00000000",
    21597 => x"00000000", 21598 => x"00000000", 21599 => x"00000000",
    21600 => x"00000000", 21601 => x"00000000", 21602 => x"00000000",
    21603 => x"00000000", 21604 => x"00000000", 21605 => x"00000000",
    21606 => x"00000000", 21607 => x"00000000", 21608 => x"00000000",
    21609 => x"00000000", 21610 => x"00000000", 21611 => x"00000000",
    21612 => x"00000000", 21613 => x"00000000", 21614 => x"00000000",
    21615 => x"00000000", 21616 => x"00000000", 21617 => x"00000000",
    21618 => x"00000000", 21619 => x"00000000", 21620 => x"00000000",
    21621 => x"00000000", 21622 => x"00000000", 21623 => x"00000000",
    21624 => x"00000000", 21625 => x"00000000", 21626 => x"00000000",
    21627 => x"00000000", 21628 => x"00000000", 21629 => x"00000000",
    21630 => x"00000000", 21631 => x"00000000", 21632 => x"00000000",
    21633 => x"00000000", 21634 => x"00000000", 21635 => x"00000000",
    21636 => x"00000000", 21637 => x"00000000", 21638 => x"00000000",
    21639 => x"00000000", 21640 => x"00000000", 21641 => x"00000000",
    21642 => x"00000000", 21643 => x"00000000", 21644 => x"00000000",
    21645 => x"00000000", 21646 => x"00000000", 21647 => x"00000000",
    21648 => x"00000000", 21649 => x"00000000", 21650 => x"00000000",
    21651 => x"00000000", 21652 => x"00000000", 21653 => x"00000000",
    21654 => x"00000000", 21655 => x"00000000", 21656 => x"00000000",
    21657 => x"00000000", 21658 => x"00000000", 21659 => x"00000000",
    21660 => x"00000000", 21661 => x"00000000", 21662 => x"00000000",
    21663 => x"00000000", 21664 => x"00000000", 21665 => x"00000000",
    21666 => x"00000000", 21667 => x"00000000", 21668 => x"00000000",
    21669 => x"00000000", 21670 => x"00000000", 21671 => x"00000000",
    21672 => x"00000000", 21673 => x"00000000", 21674 => x"00000000",
    21675 => x"00000000", 21676 => x"00000000", 21677 => x"00000000",
    21678 => x"00000000", 21679 => x"00000000", 21680 => x"00000000",
    21681 => x"00000000", 21682 => x"00000000", 21683 => x"00000000",
    21684 => x"00000000", 21685 => x"00000000", 21686 => x"00000000",
    21687 => x"00000000", 21688 => x"00000000", 21689 => x"00000000",
    21690 => x"00000000", 21691 => x"00000000", 21692 => x"00000000",
    21693 => x"00000000", 21694 => x"00000000", 21695 => x"00000000",
    21696 => x"00000000", 21697 => x"00000000", 21698 => x"00000000",
    21699 => x"00000000", 21700 => x"00000000", 21701 => x"00000000",
    21702 => x"00000000", 21703 => x"00000000", 21704 => x"00000000",
    21705 => x"00000000", 21706 => x"00000000", 21707 => x"00000000",
    21708 => x"00000000", 21709 => x"00000000", 21710 => x"00000000",
    21711 => x"00000000", 21712 => x"00000000", 21713 => x"00000000",
    21714 => x"00000000", 21715 => x"00000000", 21716 => x"00000000",
    21717 => x"00000000", 21718 => x"00000000", 21719 => x"00000000",
    21720 => x"00000000", 21721 => x"00000000", 21722 => x"00000000",
    21723 => x"00000000", 21724 => x"00000000", 21725 => x"00000000",
    21726 => x"00000000", 21727 => x"00000000", 21728 => x"00000000",
    21729 => x"00000000", 21730 => x"00000000", 21731 => x"00000000",
    21732 => x"00000000", 21733 => x"00000000", 21734 => x"00000000",
    21735 => x"00000000", 21736 => x"00000000", 21737 => x"00000000",
    21738 => x"00000000", 21739 => x"00000000", 21740 => x"00000000",
    21741 => x"00000000", 21742 => x"00000000", 21743 => x"00000000",
    21744 => x"00000000", 21745 => x"00000000", 21746 => x"00000000",
    21747 => x"00000000", 21748 => x"00000000", 21749 => x"00000000",
    21750 => x"00000000", 21751 => x"00000000", 21752 => x"00000000",
    21753 => x"00000000", 21754 => x"00000000", 21755 => x"00000000",
    21756 => x"00000000", 21757 => x"00000000", 21758 => x"00000000",
    21759 => x"00000000", 21760 => x"00000000", 21761 => x"00000000",
    21762 => x"00000000", 21763 => x"00000000", 21764 => x"00000000",
    21765 => x"00000000", 21766 => x"00000000", 21767 => x"00000000",
    21768 => x"00000000", 21769 => x"00000000", 21770 => x"00000000",
    21771 => x"00000000", 21772 => x"00000000", 21773 => x"00000000",
    21774 => x"00000000", 21775 => x"00000000", 21776 => x"00000000",
    21777 => x"00000000", 21778 => x"00000000", 21779 => x"00000000",
    21780 => x"00000000", 21781 => x"00000000", 21782 => x"00000000",
    21783 => x"00000000", 21784 => x"00000000", 21785 => x"00000000",
    21786 => x"00000000", 21787 => x"00000000", 21788 => x"00000000",
    21789 => x"00000000", 21790 => x"00000000", 21791 => x"00000000",
    21792 => x"00000000", 21793 => x"00000000", 21794 => x"00000000",
    21795 => x"00000000", 21796 => x"00000000", 21797 => x"00000000",
    21798 => x"00000000", 21799 => x"00000000", 21800 => x"00000000",
    21801 => x"00000000", 21802 => x"00000000", 21803 => x"00000000",
    21804 => x"00000000", 21805 => x"00000000", 21806 => x"00000000",
    21807 => x"00000000", 21808 => x"00000000", 21809 => x"00000000",
    21810 => x"00000000", 21811 => x"00000000", 21812 => x"00000000",
    21813 => x"00000000", 21814 => x"00000000", 21815 => x"00000000",
    21816 => x"00000000", 21817 => x"00000000", 21818 => x"00000000",
    21819 => x"00000000", 21820 => x"00000000", 21821 => x"00000000",
    21822 => x"00000000", 21823 => x"00000000", 21824 => x"00000000",
    21825 => x"00000000", 21826 => x"00000000", 21827 => x"00000000",
    21828 => x"00000000", 21829 => x"00000000", 21830 => x"00000000",
    21831 => x"00000000", 21832 => x"00000000", 21833 => x"00000000",
    21834 => x"00000000", 21835 => x"00000000", 21836 => x"00000000",
    21837 => x"00000000", 21838 => x"00000000", 21839 => x"00000000",
    21840 => x"00000000", 21841 => x"00000000", 21842 => x"00000000",
    21843 => x"00000000", 21844 => x"00000000", 21845 => x"00000000",
    21846 => x"00000000", 21847 => x"00000000", 21848 => x"00000000",
    21849 => x"00000000", 21850 => x"00000000", 21851 => x"00000000",
    21852 => x"00000000", 21853 => x"00000000", 21854 => x"00000000",
    21855 => x"00000000", 21856 => x"00000000", 21857 => x"00000000",
    21858 => x"00000000", 21859 => x"00000000", 21860 => x"00000000",
    21861 => x"00000000", 21862 => x"00000000", 21863 => x"00000000",
    21864 => x"00000000", 21865 => x"00000000", 21866 => x"00000000",
    21867 => x"00000000", 21868 => x"00000000", 21869 => x"00000000",
    21870 => x"00000000", 21871 => x"00000000", 21872 => x"00000000",
    21873 => x"00000000", 21874 => x"00000000", 21875 => x"00000000",
    21876 => x"00000000", 21877 => x"00000000", 21878 => x"00000000",
    21879 => x"00000000", 21880 => x"00000000", 21881 => x"00000000",
    21882 => x"00000000", 21883 => x"00000000", 21884 => x"00000000",
    21885 => x"00000000", 21886 => x"00000000", 21887 => x"00000000",
    21888 => x"00000000", 21889 => x"00000000", 21890 => x"00000000",
    21891 => x"00000000", 21892 => x"00000000", 21893 => x"00000000",
    21894 => x"00000000", 21895 => x"00000000", 21896 => x"00000000",
    21897 => x"00000000", 21898 => x"00000000", 21899 => x"00000000",
    21900 => x"00000000", 21901 => x"00000000", 21902 => x"00000000",
    21903 => x"00000000", 21904 => x"00000000", 21905 => x"00000000",
    21906 => x"00000000", 21907 => x"00000000", 21908 => x"00000000",
    21909 => x"00000000", 21910 => x"00000000", 21911 => x"00000000",
    21912 => x"00000000", 21913 => x"00000000", 21914 => x"00000000",
    21915 => x"00000000", 21916 => x"00000000", 21917 => x"00000000",
    21918 => x"00000000", 21919 => x"00000000", 21920 => x"00000000",
    21921 => x"00000000", 21922 => x"00000000", 21923 => x"00000000",
    21924 => x"00000000", 21925 => x"00000000", 21926 => x"00000000",
    21927 => x"00000000", 21928 => x"00000000", 21929 => x"00000000",
    21930 => x"00000000", 21931 => x"00000000", 21932 => x"00000000",
    21933 => x"00000000", 21934 => x"00000000", 21935 => x"00000000",
    21936 => x"00000000", 21937 => x"00000000", 21938 => x"00000000",
    21939 => x"00000000", 21940 => x"00000000", 21941 => x"00000000",
    21942 => x"00000000", 21943 => x"00000000", 21944 => x"00000000",
    21945 => x"00000000", 21946 => x"00000000", 21947 => x"00000000",
    21948 => x"00000000", 21949 => x"00000000", 21950 => x"00000000",
    21951 => x"00000000", 21952 => x"00000000", 21953 => x"00000000",
    21954 => x"00000000", 21955 => x"00000000", 21956 => x"00000000",
    21957 => x"00000000", 21958 => x"00000000", 21959 => x"00000000",
    21960 => x"00000000", 21961 => x"00000000", 21962 => x"00000000",
    21963 => x"00000000", 21964 => x"00000000", 21965 => x"00000000",
    21966 => x"00000000", 21967 => x"00000000", 21968 => x"00000000",
    21969 => x"00000000", 21970 => x"00000000", 21971 => x"00000000",
    21972 => x"00000000", 21973 => x"00000000", 21974 => x"00000000",
    21975 => x"00000000", 21976 => x"00000000", 21977 => x"00000000",
    21978 => x"00000000", 21979 => x"00000000", 21980 => x"00000000",
    21981 => x"00000000", 21982 => x"00000000", 21983 => x"00000000",
    21984 => x"00000000", 21985 => x"00000000", 21986 => x"00000000",
    21987 => x"00000000", 21988 => x"00000000", 21989 => x"00000000",
    21990 => x"00000000", 21991 => x"00000000", 21992 => x"00000000",
    21993 => x"00000000", 21994 => x"00000000", 21995 => x"00000000",
    21996 => x"00000000", 21997 => x"00000000", 21998 => x"00000000",
    21999 => x"00000000", 22000 => x"00000000", 22001 => x"00000000",
    22002 => x"00000000", 22003 => x"00000000", 22004 => x"00000000",
    22005 => x"00000000", 22006 => x"00000000", 22007 => x"00000000",
    22008 => x"00000000", 22009 => x"00000000", 22010 => x"00000000",
    22011 => x"00000000", 22012 => x"00000000", 22013 => x"00000000",
    22014 => x"00000000", 22015 => x"00000000", 22016 => x"00000000",
    22017 => x"00000000", 22018 => x"00000000", 22019 => x"00000000",
    22020 => x"00000000", 22021 => x"00000000", 22022 => x"00000000",
    22023 => x"00000000", 22024 => x"00000000", 22025 => x"00000000",
    22026 => x"00000000", 22027 => x"00000000", 22028 => x"00000000",
    22029 => x"00000000", 22030 => x"00000000", 22031 => x"00000000",
    22032 => x"00000000", 22033 => x"00000000", 22034 => x"00000000",
    22035 => x"00000000", 22036 => x"00000000", 22037 => x"00000000",
    22038 => x"00000000", 22039 => x"00000000", 22040 => x"00000000",
    22041 => x"00000000", 22042 => x"00000000", 22043 => x"00000000",
    22044 => x"00000000", 22045 => x"00000000", 22046 => x"00000000",
    22047 => x"00000000", 22048 => x"00000000", 22049 => x"00000000",
    22050 => x"00000000", 22051 => x"00000000", 22052 => x"00000000",
    22053 => x"00000000", 22054 => x"00000000", 22055 => x"00000000",
    22056 => x"00000000", 22057 => x"00000000", 22058 => x"00000000",
    22059 => x"00000000", 22060 => x"00000000", 22061 => x"00000000",
    22062 => x"00000000", 22063 => x"00000000", 22064 => x"00000000",
    22065 => x"00000000", 22066 => x"00000000", 22067 => x"00000000",
    22068 => x"00000000", 22069 => x"00000000", 22070 => x"00000000",
    22071 => x"00000000", 22072 => x"00000000", 22073 => x"00000000",
    22074 => x"00000000", 22075 => x"00000000", 22076 => x"00000000",
    22077 => x"00000000", 22078 => x"00000000", 22079 => x"00000000",
    22080 => x"00000000", 22081 => x"00000000", 22082 => x"00000000",
    22083 => x"00000000", 22084 => x"00000000", 22085 => x"00000000",
    22086 => x"00000000", 22087 => x"00000000", 22088 => x"00000000",
    22089 => x"00000000", 22090 => x"00000000", 22091 => x"00000000",
    22092 => x"00000000", 22093 => x"00000000", 22094 => x"00000000",
    22095 => x"00000000", 22096 => x"00000000", 22097 => x"00000000",
    22098 => x"00000000", 22099 => x"00000000", 22100 => x"00000000",
    22101 => x"00000000", 22102 => x"00000000", 22103 => x"00000000",
    22104 => x"00000000", 22105 => x"00000000", 22106 => x"00000000",
    22107 => x"00000000", 22108 => x"00000000", 22109 => x"00000000",
    22110 => x"00000000", 22111 => x"00000000", 22112 => x"00000000",
    22113 => x"00000000", 22114 => x"00000000", 22115 => x"00000000",
    22116 => x"00000000", 22117 => x"00000000", 22118 => x"00000000",
    22119 => x"00000000", 22120 => x"00000000", 22121 => x"00000000",
    22122 => x"00000000", 22123 => x"00000000", 22124 => x"00000000",
    22125 => x"00000000", 22126 => x"00000000", 22127 => x"00000000",
    22128 => x"00000000", 22129 => x"00000000", 22130 => x"00000000",
    22131 => x"00000000", 22132 => x"00000000", 22133 => x"00000000",
    22134 => x"00000000", 22135 => x"00000000", 22136 => x"00000000",
    22137 => x"00000000", 22138 => x"00000000", 22139 => x"00000000",
    22140 => x"00000000", 22141 => x"00000000", 22142 => x"00000000",
    22143 => x"00000000", 22144 => x"00000000", 22145 => x"00000000",
    22146 => x"00000000", 22147 => x"00000000", 22148 => x"00000000",
    22149 => x"00000000", 22150 => x"00000000", 22151 => x"00000000",
    22152 => x"00000000", 22153 => x"00000000", 22154 => x"00000000",
    22155 => x"00000000", 22156 => x"00000000", 22157 => x"00000000",
    22158 => x"00000000", 22159 => x"00000000", 22160 => x"00000000",
    22161 => x"00000000", 22162 => x"00000000", 22163 => x"00000000",
    22164 => x"00000000", 22165 => x"00000000", 22166 => x"00000000",
    22167 => x"00000000", 22168 => x"00000000", 22169 => x"00000000",
    22170 => x"00000000", 22171 => x"00000000", 22172 => x"00000000",
    22173 => x"00000000", 22174 => x"00000000", 22175 => x"00000000",
    22176 => x"00000000", 22177 => x"00000000", 22178 => x"00000000",
    22179 => x"00000000", 22180 => x"00000000", 22181 => x"00000000",
    22182 => x"00000000", 22183 => x"00000000", 22184 => x"00000000",
    22185 => x"00000000", 22186 => x"00000000", 22187 => x"00000000",
    22188 => x"00000000", 22189 => x"00000000", 22190 => x"00000000",
    22191 => x"00000000", 22192 => x"00000000", 22193 => x"00000000",
    22194 => x"00000000", 22195 => x"00000000", 22196 => x"00000000",
    22197 => x"00000000", 22198 => x"00000000", 22199 => x"00000000",
    22200 => x"00000000", 22201 => x"00000000", 22202 => x"00000000",
    22203 => x"00000000", 22204 => x"00000000", 22205 => x"00000000",
    22206 => x"00000000", 22207 => x"00000000", 22208 => x"00000000",
    22209 => x"00000000", 22210 => x"00000000", 22211 => x"00000000",
    22212 => x"00000000", 22213 => x"00000000", 22214 => x"00000000",
    22215 => x"00000000", 22216 => x"00000000", 22217 => x"00000000",
    22218 => x"00000000", 22219 => x"00000000", 22220 => x"00000000",
    22221 => x"00000000", 22222 => x"00000000", 22223 => x"00000000",
    22224 => x"00000000", 22225 => x"00000000", 22226 => x"00000000",
    22227 => x"00000000", 22228 => x"00000000", 22229 => x"00000000",
    22230 => x"00000000", 22231 => x"00000000", 22232 => x"00000000",
    22233 => x"00000000", 22234 => x"00000000", 22235 => x"00000000",
    22236 => x"00000000", 22237 => x"00000000", 22238 => x"00000000",
    22239 => x"00000000", 22240 => x"00000000", 22241 => x"00000000",
    22242 => x"00000000", 22243 => x"00000000", 22244 => x"00000000",
    22245 => x"00000000", 22246 => x"00000000", 22247 => x"00000000",
    22248 => x"00000000", 22249 => x"00000000", 22250 => x"00000000",
    22251 => x"00000000", 22252 => x"00000000", 22253 => x"00000000",
    22254 => x"00000000", 22255 => x"00000000", 22256 => x"00000000",
    22257 => x"00000000", 22258 => x"00000000", 22259 => x"00000000",
    22260 => x"00000000", 22261 => x"00000000", 22262 => x"00000000",
    22263 => x"00000000", 22264 => x"00000000", 22265 => x"00000000",
    22266 => x"00000000", 22267 => x"00000000", 22268 => x"00000000",
    22269 => x"00000000", 22270 => x"00000000", 22271 => x"00000000",
    22272 => x"00000000", 22273 => x"00000000", 22274 => x"00000000",
    22275 => x"00000000", 22276 => x"00000000", 22277 => x"00000000",
    22278 => x"00000000", 22279 => x"00000000", 22280 => x"00000000",
    22281 => x"00000000", 22282 => x"00000000", 22283 => x"00000000",
    22284 => x"00000000", 22285 => x"00000000", 22286 => x"00000000",
    22287 => x"00000000", 22288 => x"00000000", 22289 => x"00000000",
    22290 => x"00000000", 22291 => x"00000000", 22292 => x"00000000",
    22293 => x"00000000", 22294 => x"00000000", 22295 => x"00000000",
    22296 => x"00000000", 22297 => x"00000000", 22298 => x"00000000",
    22299 => x"00000000", 22300 => x"00000000", 22301 => x"00000000",
    22302 => x"00000000", 22303 => x"00000000", 22304 => x"00000000",
    22305 => x"00000000", 22306 => x"00000000", 22307 => x"00000000",
    22308 => x"00000000", 22309 => x"00000000", 22310 => x"00000000",
    22311 => x"00000000", 22312 => x"00000000", 22313 => x"00000000",
    22314 => x"00000000", 22315 => x"00000000", 22316 => x"00000000",
    22317 => x"00000000", 22318 => x"00000000", 22319 => x"00000000",
    22320 => x"00000000", 22321 => x"00000000", 22322 => x"00000000",
    22323 => x"00000000", 22324 => x"00000000", 22325 => x"00000000",
    22326 => x"00000000", 22327 => x"00000000", 22328 => x"00000000",
    22329 => x"00000000", 22330 => x"00000000", 22331 => x"00000000",
    22332 => x"00000000", 22333 => x"00000000", 22334 => x"00000000",
    22335 => x"00000000", 22336 => x"00000000", 22337 => x"00000000",
    22338 => x"00000000", 22339 => x"00000000", 22340 => x"00000000",
    22341 => x"00000000", 22342 => x"00000000", 22343 => x"00000000",
    22344 => x"00000000", 22345 => x"00000000", 22346 => x"00000000",
    22347 => x"00000000", 22348 => x"00000000", 22349 => x"00000000",
    22350 => x"00000000", 22351 => x"00000000", 22352 => x"00000000",
    22353 => x"00000000", 22354 => x"00000000", 22355 => x"00000000",
    22356 => x"00000000", 22357 => x"00000000", 22358 => x"00000000",
    22359 => x"00000000", 22360 => x"00000000", 22361 => x"00000000",
    22362 => x"00000000", 22363 => x"00000000", 22364 => x"00000000",
    22365 => x"00000000", 22366 => x"00000000", 22367 => x"00000000",
    22368 => x"00000000", 22369 => x"00000000", 22370 => x"00000000",
    22371 => x"00000000", 22372 => x"00000000", 22373 => x"00000000",
    22374 => x"00000000", 22375 => x"00000000", 22376 => x"00000000",
    22377 => x"00000000", 22378 => x"00000000", 22379 => x"00000000",
    22380 => x"00000000", 22381 => x"00000000", 22382 => x"00000000",
    22383 => x"00000000", 22384 => x"00000000", 22385 => x"00000000",
    22386 => x"00000000", 22387 => x"00000000", 22388 => x"00000000",
    22389 => x"00000000", 22390 => x"00000000", 22391 => x"00000000",
    22392 => x"00000000", 22393 => x"00000000", 22394 => x"00000000",
    22395 => x"00000000", 22396 => x"00000000", 22397 => x"00000000",
    22398 => x"00000000", 22399 => x"00000000", 22400 => x"00000000",
    22401 => x"00000000", 22402 => x"00000000", 22403 => x"00000000",
    22404 => x"00000000", 22405 => x"00000000", 22406 => x"00000000",
    22407 => x"00000000", 22408 => x"00000000", 22409 => x"00000000",
    22410 => x"00000000", 22411 => x"00000000", 22412 => x"00000000",
    22413 => x"00000000", 22414 => x"00000000", 22415 => x"00000000",
    22416 => x"00000000", 22417 => x"00000000", 22418 => x"00000000",
    22419 => x"00000000", 22420 => x"00000000", 22421 => x"00000000",
    22422 => x"00000000", 22423 => x"00000000", 22424 => x"00000000",
    22425 => x"00000000", 22426 => x"00000000", 22427 => x"00000000",
    22428 => x"00000000", 22429 => x"00000000", 22430 => x"00000000",
    22431 => x"00000000", 22432 => x"00000000", 22433 => x"00000000",
    22434 => x"00000000", 22435 => x"00000000", 22436 => x"00000000",
    22437 => x"00000000", 22438 => x"00000000", 22439 => x"00000000",
    22440 => x"00000000", 22441 => x"00000000", 22442 => x"00000000",
    22443 => x"00000000", 22444 => x"00000000", 22445 => x"00000000",
    22446 => x"00000000", 22447 => x"00000000", 22448 => x"00000000",
    22449 => x"00000000", 22450 => x"00000000", 22451 => x"00000000",
    22452 => x"00000000", 22453 => x"00000000", 22454 => x"00000000",
    22455 => x"00000000", 22456 => x"00000000", 22457 => x"00000000",
    22458 => x"00000000", 22459 => x"00000000", 22460 => x"00000000",
    22461 => x"00000000", 22462 => x"00000000", 22463 => x"00000000",
    22464 => x"00000000", 22465 => x"00000000", 22466 => x"00000000",
    22467 => x"00000000", 22468 => x"00000000", 22469 => x"00000000",
    22470 => x"00000000", 22471 => x"00000000", 22472 => x"00000000",
    22473 => x"00000000", 22474 => x"00000000", 22475 => x"00000000",
    22476 => x"00000000", 22477 => x"00000000", 22478 => x"00000000",
    22479 => x"00000000", 22480 => x"00000000", 22481 => x"00000000",
    22482 => x"00000000", 22483 => x"00000000", 22484 => x"00000000",
    22485 => x"00000000", 22486 => x"00000000", 22487 => x"00000000",
    22488 => x"00000000", 22489 => x"00000000", 22490 => x"00000000",
    22491 => x"00000000", 22492 => x"00000000", 22493 => x"00000000",
    22494 => x"00000000", 22495 => x"00000000", 22496 => x"00000000",
    22497 => x"00000000", 22498 => x"00000000", 22499 => x"00000000",
    22500 => x"00000000", 22501 => x"00000000", 22502 => x"00000000",
    22503 => x"00000000", 22504 => x"00000000", 22505 => x"00000000",
    22506 => x"00000000", 22507 => x"00000000", 22508 => x"00000000",
    22509 => x"00000000", 22510 => x"00000000", 22511 => x"00000000",
    22512 => x"00000000", 22513 => x"00000000", 22514 => x"00000000",
    22515 => x"00000000", 22516 => x"00000000", 22517 => x"00000000",
    22518 => x"00000000", 22519 => x"00000000", 22520 => x"00000000",
    22521 => x"00000000", 22522 => x"00000000", 22523 => x"00000000",
    22524 => x"00000000", 22525 => x"00000000", 22526 => x"00000000",
    22527 => x"00000000", 22528 => x"00000000", 22529 => x"00000000",
    22530 => x"00000000", 22531 => x"00000000", 22532 => x"00000000",
    22533 => x"00000000", 22534 => x"00000000", 22535 => x"00000000",
    22536 => x"00000000", 22537 => x"00000000", 22538 => x"00000000",
    22539 => x"00000000", 22540 => x"00000000", 22541 => x"00000000",
    22542 => x"00000000", 22543 => x"00000000", 22544 => x"00000000",
    22545 => x"00000000", 22546 => x"00000000", 22547 => x"00000000",
    22548 => x"00000000", 22549 => x"00000000", 22550 => x"00000000",
    22551 => x"00000000", 22552 => x"00000000", 22553 => x"00000000",
    22554 => x"00000000", 22555 => x"00000000", 22556 => x"00000000",
    22557 => x"00000000", 22558 => x"00000000", 22559 => x"00000000",
    22560 => x"00000000", 22561 => x"00000000", 22562 => x"00000000",
    22563 => x"00000000", 22564 => x"00000000", 22565 => x"00000000",
    22566 => x"00000000", 22567 => x"00000000", 22568 => x"00000000",
    22569 => x"00000000", 22570 => x"00000000", 22571 => x"00000000",
    22572 => x"00000000", 22573 => x"00000000", 22574 => x"00000000",
    22575 => x"00000000", 22576 => x"00000000", 22577 => x"00000000",
    22578 => x"00000000", 22579 => x"00000000", 22580 => x"00000000",
    22581 => x"00000000", 22582 => x"00000000", 22583 => x"00000000",
    22584 => x"00000000", 22585 => x"00000000", 22586 => x"00000000",
    22587 => x"00000000", 22588 => x"00000000", 22589 => x"00000000",
    22590 => x"00000000", 22591 => x"00000000", 22592 => x"00000000",
    22593 => x"00000000", 22594 => x"00000000", 22595 => x"00000000",
    22596 => x"00000000", 22597 => x"00000000", 22598 => x"00000000",
    22599 => x"00000000", 22600 => x"00000000", 22601 => x"00000000",
    22602 => x"00000000", 22603 => x"00000000", 22604 => x"00000000",
    22605 => x"00000000", 22606 => x"00000000", 22607 => x"00000000",
    22608 => x"00000000", 22609 => x"00000000", 22610 => x"00000000",
    22611 => x"00000000", 22612 => x"00000000", 22613 => x"00000000",
    22614 => x"00000000", 22615 => x"00000000", 22616 => x"00000000",
    22617 => x"00000000", 22618 => x"00000000", 22619 => x"00000000",
    22620 => x"00000000", 22621 => x"00000000", 22622 => x"00000000",
    22623 => x"00000000", 22624 => x"00000000", 22625 => x"00000000",
    22626 => x"00000000", 22627 => x"00000000", 22628 => x"00000000",
    22629 => x"00000000", 22630 => x"00000000", 22631 => x"00000000",
    22632 => x"00000000", 22633 => x"00000000", 22634 => x"00000000",
    22635 => x"00000000", 22636 => x"00000000", 22637 => x"00000000",
    22638 => x"00000000", 22639 => x"00000000", 22640 => x"00000000",
    22641 => x"00000000", 22642 => x"00000000", 22643 => x"00000000",
    22644 => x"00000000", 22645 => x"00000000", 22646 => x"00000000",
    22647 => x"00000000", 22648 => x"00000000", 22649 => x"00000000",
    22650 => x"00000000", 22651 => x"00000000", 22652 => x"00000000",
    22653 => x"00000000", 22654 => x"00000000", 22655 => x"00000000",
    22656 => x"00000000", 22657 => x"00000000", 22658 => x"00000000",
    22659 => x"00000000", 22660 => x"00000000", 22661 => x"00000000",
    22662 => x"00000000", 22663 => x"00000000", 22664 => x"00000000",
    22665 => x"00000000", 22666 => x"00000000", 22667 => x"00000000",
    22668 => x"00000000", 22669 => x"00000000", 22670 => x"00000000",
    22671 => x"00000000", 22672 => x"00000000", 22673 => x"00000000",
    22674 => x"00000000", 22675 => x"00000000", 22676 => x"00000000",
    22677 => x"00000000", 22678 => x"00000000", 22679 => x"00000000",
    22680 => x"00000000", 22681 => x"00000000", 22682 => x"00000000",
    22683 => x"00000000", 22684 => x"00000000", 22685 => x"00000000",
    22686 => x"00000000", 22687 => x"00000000", 22688 => x"00000000",
    22689 => x"00000000", 22690 => x"00000000", 22691 => x"00000000",
    22692 => x"00000000", 22693 => x"00000000", 22694 => x"00000000",
    22695 => x"00000000", 22696 => x"00000000", 22697 => x"00000000",
    22698 => x"00000000", 22699 => x"00000000", 22700 => x"00000000",
    22701 => x"00000000", 22702 => x"00000000", 22703 => x"00000000",
    22704 => x"00000000", 22705 => x"00000000", 22706 => x"00000000",
    22707 => x"00000000", 22708 => x"00000000", 22709 => x"00000000",
    22710 => x"00000000", 22711 => x"00000000", 22712 => x"00000000",
    22713 => x"00000000", 22714 => x"00000000", 22715 => x"00000000",
    22716 => x"00000000", 22717 => x"00000000", 22718 => x"00000000",
    22719 => x"00000000", 22720 => x"00000000", 22721 => x"00000000",
    22722 => x"00000000", 22723 => x"00000000", 22724 => x"00000000",
    22725 => x"00000000", 22726 => x"00000000", 22727 => x"00000000",
    22728 => x"00000000", 22729 => x"00000000", 22730 => x"00000000",
    22731 => x"00000000", 22732 => x"00000000", 22733 => x"00000000",
    22734 => x"00000000", 22735 => x"00000000", 22736 => x"00000000",
    22737 => x"00000000", 22738 => x"00000000", 22739 => x"00000000",
    22740 => x"00000000", 22741 => x"00000000", 22742 => x"00000000",
    22743 => x"00000000", 22744 => x"00000000", 22745 => x"00000000",
    22746 => x"00000000", 22747 => x"00000000", 22748 => x"00000000",
    22749 => x"00000000", 22750 => x"00000000", 22751 => x"00000000",
    22752 => x"00000000", 22753 => x"00000000", 22754 => x"00000000",
    22755 => x"00000000", 22756 => x"00000000", 22757 => x"00000000",
    22758 => x"00000000", 22759 => x"00000000", 22760 => x"00000000",
    22761 => x"00000000", 22762 => x"00000000", 22763 => x"00000000",
    22764 => x"00000000", 22765 => x"00000000", 22766 => x"00000000",
    22767 => x"00000000", 22768 => x"00000000", 22769 => x"00000000",
    22770 => x"00000000", 22771 => x"00000000", 22772 => x"00000000",
    22773 => x"00000000", 22774 => x"00000000", 22775 => x"00000000",
    22776 => x"00000000", 22777 => x"00000000", 22778 => x"00000000",
    22779 => x"00000000", 22780 => x"00000000", 22781 => x"00000000",
    22782 => x"00000000", 22783 => x"00000000", 22784 => x"00000000",
    22785 => x"00000000", 22786 => x"00000000", 22787 => x"00000000",
    22788 => x"00000000", 22789 => x"00000000", 22790 => x"00000000",
    22791 => x"00000000", 22792 => x"00000000", 22793 => x"00000000",
    22794 => x"00000000", 22795 => x"00000000", 22796 => x"00000000",
    22797 => x"00000000", 22798 => x"00000000", 22799 => x"00000000",
    22800 => x"00000000", 22801 => x"00000000", 22802 => x"00000000",
    22803 => x"00000000", 22804 => x"00000000", 22805 => x"00000000",
    22806 => x"00000000", 22807 => x"00000000", 22808 => x"00000000",
    22809 => x"00000000", 22810 => x"00000000", 22811 => x"00000000",
    22812 => x"00000000", 22813 => x"00000000", 22814 => x"00000000",
    22815 => x"00000000", 22816 => x"00000000", 22817 => x"00000000",
    22818 => x"00000000", 22819 => x"00000000", 22820 => x"00000000",
    22821 => x"00000000", 22822 => x"00000000", 22823 => x"00000000",
    22824 => x"00000000", 22825 => x"00000000", 22826 => x"00000000",
    22827 => x"00000000", 22828 => x"00000000", 22829 => x"00000000",
    22830 => x"00000000", 22831 => x"00000000", 22832 => x"00000000",
    22833 => x"00000000", 22834 => x"00000000", 22835 => x"00000000",
    22836 => x"00000000", 22837 => x"00000000", 22838 => x"00000000",
    22839 => x"00000000", 22840 => x"00000000", 22841 => x"00000000",
    22842 => x"00000000", 22843 => x"00000000", 22844 => x"00000000",
    22845 => x"00000000", 22846 => x"00000000", 22847 => x"00000000",
    22848 => x"00000000", 22849 => x"00000000", 22850 => x"00000000",
    22851 => x"00000000", 22852 => x"00000000", 22853 => x"00000000",
    22854 => x"00000000", 22855 => x"00000000", 22856 => x"00000000",
    22857 => x"00000000", 22858 => x"00000000", 22859 => x"00000000",
    22860 => x"00000000", 22861 => x"00000000", 22862 => x"00000000",
    22863 => x"00000000", 22864 => x"00000000", 22865 => x"00000000",
    22866 => x"00000000", 22867 => x"00000000", 22868 => x"00000000",
    22869 => x"00000000", 22870 => x"00000000", 22871 => x"00000000",
    22872 => x"00000000", 22873 => x"00000000", 22874 => x"00000000",
    22875 => x"00000000", 22876 => x"00000000", 22877 => x"00000000",
    22878 => x"00000000", 22879 => x"00000000", 22880 => x"00000000",
    22881 => x"00000000", 22882 => x"00000000", 22883 => x"00000000",
    22884 => x"00000000", 22885 => x"00000000", 22886 => x"00000000",
    22887 => x"00000000", 22888 => x"00000000", 22889 => x"00000000",
    22890 => x"00000000", 22891 => x"00000000", 22892 => x"00000000",
    22893 => x"00000000", 22894 => x"00000000", 22895 => x"00000000",
    22896 => x"00000000", 22897 => x"00000000", 22898 => x"00000000",
    22899 => x"00000000", 22900 => x"00000000", 22901 => x"00000000",
    22902 => x"00000000", 22903 => x"00000000", 22904 => x"00000000",
    22905 => x"00000000", 22906 => x"00000000", 22907 => x"00000000",
    22908 => x"00000000", 22909 => x"00000000", 22910 => x"00000000",
    22911 => x"00000000", 22912 => x"00000000", 22913 => x"00000000",
    22914 => x"00000000", 22915 => x"00000000", 22916 => x"00000000",
    22917 => x"00000000", 22918 => x"00000000", 22919 => x"00000000",
    22920 => x"00000000", 22921 => x"00000000", 22922 => x"00000000",
    22923 => x"00000000", 22924 => x"00000000", 22925 => x"00000000",
    22926 => x"00000000", 22927 => x"00000000", 22928 => x"00000000",
    22929 => x"00000000", 22930 => x"00000000", 22931 => x"00000000",
    22932 => x"00000000", 22933 => x"00000000", 22934 => x"00000000",
    22935 => x"00000000", 22936 => x"00000000", 22937 => x"00000000",
    22938 => x"00000000", 22939 => x"00000000", 22940 => x"00000000",
    22941 => x"00000000", 22942 => x"00000000", 22943 => x"00000000",
    22944 => x"00000000", 22945 => x"00000000", 22946 => x"00000000",
    22947 => x"00000000", 22948 => x"00000000", 22949 => x"00000000",
    22950 => x"00000000", 22951 => x"00000000", 22952 => x"00000000",
    22953 => x"00000000", 22954 => x"00000000", 22955 => x"00000000",
    22956 => x"00000000", 22957 => x"00000000", 22958 => x"00000000",
    22959 => x"00000000", 22960 => x"00000000", 22961 => x"00000000",
    22962 => x"00000000", 22963 => x"00000000", 22964 => x"00000000",
    22965 => x"00000000", 22966 => x"00000000", 22967 => x"00000000",
    22968 => x"00000000", 22969 => x"00000000", 22970 => x"00000000",
    22971 => x"00000000", 22972 => x"00000000", 22973 => x"00000000",
    22974 => x"00000000", 22975 => x"00000000", 22976 => x"00000000",
    22977 => x"00000000", 22978 => x"00000000", 22979 => x"00000000",
    22980 => x"00000000", 22981 => x"00000000", 22982 => x"00000000",
    22983 => x"00000000", 22984 => x"00000000", 22985 => x"00000000",
    22986 => x"00000000", 22987 => x"00000000", 22988 => x"00000000",
    22989 => x"00000000", 22990 => x"00000000", 22991 => x"00000000",
    22992 => x"00000000", 22993 => x"00000000", 22994 => x"00000000",
    22995 => x"00000000", 22996 => x"00000000", 22997 => x"00000000",
    22998 => x"00000000", 22999 => x"00000000", 23000 => x"00000000",
    23001 => x"00000000", 23002 => x"00000000", 23003 => x"00000000",
    23004 => x"00000000", 23005 => x"00000000", 23006 => x"00000000",
    23007 => x"00000000", 23008 => x"00000000", 23009 => x"00000000",
    23010 => x"00000000", 23011 => x"00000000", 23012 => x"00000000",
    23013 => x"00000000", 23014 => x"00000000", 23015 => x"00000000",
    23016 => x"00000000", 23017 => x"00000000", 23018 => x"00000000",
    23019 => x"00000000", 23020 => x"00000000", 23021 => x"00000000",
    23022 => x"00000000", 23023 => x"00000000", 23024 => x"00000000",
    23025 => x"00000000", 23026 => x"00000000", 23027 => x"00000000",
    23028 => x"00000000", 23029 => x"00000000", 23030 => x"00000000",
    23031 => x"00000000", 23032 => x"00000000", 23033 => x"00000000",
    23034 => x"00000000", 23035 => x"00000000", 23036 => x"00000000",
    23037 => x"00000000", 23038 => x"00000000", 23039 => x"00000000",
    23040 => x"00000000", 23041 => x"00000000", 23042 => x"00000000",
    23043 => x"00000000", 23044 => x"00000000", 23045 => x"00000000",
    23046 => x"00000000", 23047 => x"00000000", 23048 => x"00000000",
    23049 => x"00000000", 23050 => x"00000000", 23051 => x"00000000",
    23052 => x"00000000", 23053 => x"00000000", 23054 => x"00000000",
    23055 => x"00000000", 23056 => x"00000000", 23057 => x"00000000",
    23058 => x"00000000", 23059 => x"00000000", 23060 => x"00000000",
    23061 => x"00000000", 23062 => x"00000000", 23063 => x"00000000",
    23064 => x"00000000", 23065 => x"00000000", 23066 => x"00000000",
    23067 => x"00000000", 23068 => x"00000000", 23069 => x"00000000",
    23070 => x"00000000", 23071 => x"00000000", 23072 => x"00000000",
    23073 => x"00000000", 23074 => x"00000000", 23075 => x"00000000",
    23076 => x"00000000", 23077 => x"00000000", 23078 => x"00000000",
    23079 => x"00000000", 23080 => x"00000000", 23081 => x"00000000",
    23082 => x"00000000", 23083 => x"00000000", 23084 => x"00000000",
    23085 => x"00000000", 23086 => x"00000000", 23087 => x"00000000",
    23088 => x"00000000", 23089 => x"00000000", 23090 => x"00000000",
    23091 => x"00000000", 23092 => x"00000000", 23093 => x"00000000",
    23094 => x"00000000", 23095 => x"00000000", 23096 => x"00000000",
    23097 => x"00000000", 23098 => x"00000000", 23099 => x"00000000",
    23100 => x"00000000", 23101 => x"00000000", 23102 => x"00000000",
    23103 => x"00000000", 23104 => x"00000000", 23105 => x"00000000",
    23106 => x"00000000", 23107 => x"00000000", 23108 => x"00000000",
    23109 => x"00000000", 23110 => x"00000000", 23111 => x"00000000",
    23112 => x"00000000", 23113 => x"00000000", 23114 => x"00000000",
    23115 => x"00000000", 23116 => x"00000000", 23117 => x"00000000",
    23118 => x"00000000", 23119 => x"00000000", 23120 => x"00000000",
    23121 => x"00000000", 23122 => x"00000000", 23123 => x"00000000",
    23124 => x"00000000", 23125 => x"00000000", 23126 => x"00000000",
    23127 => x"00000000", 23128 => x"00000000", 23129 => x"00000000",
    23130 => x"00000000", 23131 => x"00000000", 23132 => x"00000000",
    23133 => x"00000000", 23134 => x"00000000", 23135 => x"00000000",
    23136 => x"00000000", 23137 => x"00000000", 23138 => x"00000000",
    23139 => x"00000000", 23140 => x"00000000", 23141 => x"00000000",
    23142 => x"00000000", 23143 => x"00000000", 23144 => x"00000000",
    23145 => x"00000000", 23146 => x"00000000", 23147 => x"00000000",
    23148 => x"00000000", 23149 => x"00000000", 23150 => x"00000000",
    23151 => x"00000000", 23152 => x"00000000", 23153 => x"00000000",
    23154 => x"00000000", 23155 => x"00000000", 23156 => x"00000000",
    23157 => x"00000000", 23158 => x"00000000", 23159 => x"00000000",
    23160 => x"00000000", 23161 => x"00000000", 23162 => x"00000000",
    23163 => x"00000000", 23164 => x"00000000", 23165 => x"00000000",
    23166 => x"00000000", 23167 => x"00000000", 23168 => x"00000000",
    23169 => x"00000000", 23170 => x"00000000", 23171 => x"00000000",
    23172 => x"00000000", 23173 => x"00000000", 23174 => x"00000000",
    23175 => x"00000000", 23176 => x"00000000", 23177 => x"00000000",
    23178 => x"00000000", 23179 => x"00000000", 23180 => x"00000000",
    23181 => x"00000000", 23182 => x"00000000", 23183 => x"00000000",
    23184 => x"00000000", 23185 => x"00000000", 23186 => x"00000000",
    23187 => x"00000000", 23188 => x"00000000", 23189 => x"00000000",
    23190 => x"00000000", 23191 => x"00000000", 23192 => x"00000000",
    23193 => x"00000000", 23194 => x"00000000", 23195 => x"00000000",
    23196 => x"00000000", 23197 => x"00000000", 23198 => x"00000000",
    23199 => x"00000000", 23200 => x"00000000", 23201 => x"00000000",
    23202 => x"00000000", 23203 => x"00000000", 23204 => x"00000000",
    23205 => x"00000000", 23206 => x"00000000", 23207 => x"00000000",
    23208 => x"00000000", 23209 => x"00000000", 23210 => x"00000000",
    23211 => x"00000000", 23212 => x"00000000", 23213 => x"00000000",
    23214 => x"00000000", 23215 => x"00000000", 23216 => x"00000000",
    23217 => x"00000000", 23218 => x"00000000", 23219 => x"00000000",
    23220 => x"00000000", 23221 => x"00000000", 23222 => x"00000000",
    23223 => x"00000000", 23224 => x"00000000", 23225 => x"00000000",
    23226 => x"00000000", 23227 => x"00000000", 23228 => x"00000000",
    23229 => x"00000000", 23230 => x"00000000", 23231 => x"00000000",
    23232 => x"00000000", 23233 => x"00000000", 23234 => x"00000000",
    23235 => x"00000000", 23236 => x"00000000", 23237 => x"00000000",
    23238 => x"00000000", 23239 => x"00000000", 23240 => x"00000000",
    23241 => x"00000000", 23242 => x"00000000", 23243 => x"00000000",
    23244 => x"00000000", 23245 => x"00000000", 23246 => x"00000000",
    23247 => x"00000000", 23248 => x"00000000", 23249 => x"00000000",
    23250 => x"00000000", 23251 => x"00000000", 23252 => x"00000000",
    23253 => x"00000000", 23254 => x"00000000", 23255 => x"00000000",
    23256 => x"00000000", 23257 => x"00000000", 23258 => x"00000000",
    23259 => x"00000000", 23260 => x"00000000", 23261 => x"00000000",
    23262 => x"00000000", 23263 => x"00000000", 23264 => x"00000000",
    23265 => x"00000000", 23266 => x"00000000", 23267 => x"00000000",
    23268 => x"00000000", 23269 => x"00000000", 23270 => x"00000000",
    23271 => x"00000000", 23272 => x"00000000", 23273 => x"00000000",
    23274 => x"00000000", 23275 => x"00000000", 23276 => x"00000000",
    23277 => x"00000000", 23278 => x"00000000", 23279 => x"00000000",
    23280 => x"00000000", 23281 => x"00000000", 23282 => x"00000000",
    23283 => x"00000000", 23284 => x"00000000", 23285 => x"00000000",
    23286 => x"00000000", 23287 => x"00000000", 23288 => x"00000000",
    23289 => x"00000000", 23290 => x"00000000", 23291 => x"00000000",
    23292 => x"00000000", 23293 => x"00000000", 23294 => x"00000000",
    23295 => x"00000000", 23296 => x"00000000", 23297 => x"00000000",
    23298 => x"00000000", 23299 => x"00000000", 23300 => x"00000000",
    23301 => x"00000000", 23302 => x"00000000", 23303 => x"00000000",
    23304 => x"00000000", 23305 => x"00000000", 23306 => x"00000000",
    23307 => x"00000000", 23308 => x"00000000", 23309 => x"00000000",
    23310 => x"00000000", 23311 => x"00000000", 23312 => x"00000000",
    23313 => x"00000000", 23314 => x"00000000", 23315 => x"00000000",
    23316 => x"00000000", 23317 => x"00000000", 23318 => x"00000000",
    23319 => x"00000000", 23320 => x"00000000", 23321 => x"00000000",
    23322 => x"00000000", 23323 => x"00000000", 23324 => x"00000000",
    23325 => x"00000000", 23326 => x"00000000", 23327 => x"00000000",
    23328 => x"00000000", 23329 => x"00000000", 23330 => x"00000000",
    23331 => x"00000000", 23332 => x"00000000", 23333 => x"00000000",
    23334 => x"00000000", 23335 => x"00000000", 23336 => x"00000000",
    23337 => x"00000000", 23338 => x"00000000", 23339 => x"00000000",
    23340 => x"00000000", 23341 => x"00000000", 23342 => x"00000000",
    23343 => x"00000000", 23344 => x"00000000", 23345 => x"00000000",
    23346 => x"00000000", 23347 => x"00000000", 23348 => x"00000000",
    23349 => x"00000000", 23350 => x"00000000", 23351 => x"00000000",
    23352 => x"00000000", 23353 => x"00000000", 23354 => x"00000000",
    23355 => x"00000000", 23356 => x"00000000", 23357 => x"00000000",
    23358 => x"00000000", 23359 => x"00000000", 23360 => x"00000000",
    23361 => x"00000000", 23362 => x"00000000", 23363 => x"00000000",
    23364 => x"00000000", 23365 => x"00000000", 23366 => x"00000000",
    23367 => x"00000000", 23368 => x"00000000", 23369 => x"00000000",
    23370 => x"00000000", 23371 => x"00000000", 23372 => x"00000000",
    23373 => x"00000000", 23374 => x"00000000", 23375 => x"00000000",
    23376 => x"00000000", 23377 => x"00000000", 23378 => x"00000000",
    23379 => x"00000000", 23380 => x"00000000", 23381 => x"00000000",
    23382 => x"00000000", 23383 => x"00000000", 23384 => x"00000000",
    23385 => x"00000000", 23386 => x"00000000", 23387 => x"00000000",
    23388 => x"00000000", 23389 => x"00000000", 23390 => x"00000000",
    23391 => x"00000000", 23392 => x"00000000", 23393 => x"00000000",
    23394 => x"00000000", 23395 => x"00000000", 23396 => x"00000000",
    23397 => x"00000000", 23398 => x"00000000", 23399 => x"00000000",
    23400 => x"00000000", 23401 => x"00000000", 23402 => x"00000000",
    23403 => x"00000000", 23404 => x"00000000", 23405 => x"00000000",
    23406 => x"00000000", 23407 => x"00000000", 23408 => x"00000000",
    23409 => x"00000000", 23410 => x"00000000", 23411 => x"00000000",
    23412 => x"00000000", 23413 => x"00000000", 23414 => x"00000000",
    23415 => x"00000000", 23416 => x"00000000", 23417 => x"00000000",
    23418 => x"00000000", 23419 => x"00000000", 23420 => x"00000000",
    23421 => x"00000000", 23422 => x"00000000", 23423 => x"00000000",
    23424 => x"00000000", 23425 => x"00000000", 23426 => x"00000000",
    23427 => x"00000000", 23428 => x"00000000", 23429 => x"00000000",
    23430 => x"00000000", 23431 => x"00000000", 23432 => x"00000000",
    23433 => x"00000000", 23434 => x"00000000", 23435 => x"00000000",
    23436 => x"00000000", 23437 => x"00000000", 23438 => x"00000000",
    23439 => x"00000000", 23440 => x"00000000", 23441 => x"00000000",
    23442 => x"00000000", 23443 => x"00000000", 23444 => x"00000000",
    23445 => x"00000000", 23446 => x"00000000", 23447 => x"00000000",
    23448 => x"00000000", 23449 => x"00000000", 23450 => x"00000000",
    23451 => x"00000000", 23452 => x"00000000", 23453 => x"00000000",
    23454 => x"00000000", 23455 => x"00000000", 23456 => x"00000000",
    23457 => x"00000000", 23458 => x"00000000", 23459 => x"00000000",
    23460 => x"00000000", 23461 => x"00000000", 23462 => x"00000000",
    23463 => x"00000000", 23464 => x"00000000", 23465 => x"00000000",
    23466 => x"00000000", 23467 => x"00000000", 23468 => x"00000000",
    23469 => x"00000000", 23470 => x"00000000", 23471 => x"00000000",
    23472 => x"00000000", 23473 => x"00000000", 23474 => x"00000000",
    23475 => x"00000000", 23476 => x"00000000", 23477 => x"00000000",
    23478 => x"00000000", 23479 => x"00000000", 23480 => x"00000000",
    23481 => x"00000000", 23482 => x"00000000", 23483 => x"00000000",
    23484 => x"00000000", 23485 => x"00000000", 23486 => x"00000000",
    23487 => x"00000000", 23488 => x"00000000", 23489 => x"00000000",
    23490 => x"00000000", 23491 => x"00000000", 23492 => x"00000000",
    23493 => x"00000000", 23494 => x"00000000", 23495 => x"00000000",
    23496 => x"00000000", 23497 => x"00000000", 23498 => x"00000000",
    23499 => x"00000000", 23500 => x"00000000", 23501 => x"00000000",
    23502 => x"00000000", 23503 => x"00000000", 23504 => x"00000000",
    23505 => x"00000000", 23506 => x"00000000", 23507 => x"00000000",
    23508 => x"00000000", 23509 => x"00000000", 23510 => x"00000000",
    23511 => x"00000000", 23512 => x"00000000", 23513 => x"00000000",
    23514 => x"00000000", 23515 => x"00000000", 23516 => x"00000000",
    23517 => x"00000000", 23518 => x"00000000", 23519 => x"00000000",
    23520 => x"00000000", 23521 => x"00000000", 23522 => x"00000000",
    23523 => x"00000000", 23524 => x"00000000", 23525 => x"00000000",
    23526 => x"00000000", 23527 => x"00000000", 23528 => x"00000000",
    23529 => x"00000000", 23530 => x"00000000", 23531 => x"00000000",
    23532 => x"00000000", 23533 => x"00000000", 23534 => x"00000000",
    23535 => x"00000000", 23536 => x"00000000", 23537 => x"00000000",
    23538 => x"00000000", 23539 => x"00000000", 23540 => x"00000000",
    23541 => x"00000000", 23542 => x"00000000", 23543 => x"00000000",
    23544 => x"00000000", 23545 => x"00000000", 23546 => x"00000000",
    23547 => x"00000000", 23548 => x"00000000", 23549 => x"00000000",
    23550 => x"00000000", 23551 => x"00000000", 23552 => x"00000000",
    23553 => x"00000000", 23554 => x"00000000", 23555 => x"00000000",
    23556 => x"00000000", 23557 => x"00000000", 23558 => x"00000000",
    23559 => x"00000000", 23560 => x"00000000", 23561 => x"00000000",
    23562 => x"00000000", 23563 => x"00000000", 23564 => x"00000000",
    23565 => x"00000000", 23566 => x"00000000", 23567 => x"00000000",
    23568 => x"00000000", 23569 => x"00000000", 23570 => x"00000000",
    23571 => x"00000000", 23572 => x"00000000", 23573 => x"00000000",
    23574 => x"00000000", 23575 => x"00000000", 23576 => x"00000000",
    23577 => x"00000000", 23578 => x"00000000", 23579 => x"00000000",
    23580 => x"00000000", 23581 => x"00000000", 23582 => x"00000000",
    23583 => x"00000000", 23584 => x"00000000", 23585 => x"00000000",
    23586 => x"00000000", 23587 => x"00000000", 23588 => x"00000000",
    23589 => x"00000000", 23590 => x"00000000", 23591 => x"00000000",
    23592 => x"00000000", 23593 => x"00000000", 23594 => x"00000000",
    23595 => x"00000000", 23596 => x"00000000", 23597 => x"00000000",
    23598 => x"00000000", 23599 => x"00000000", 23600 => x"00000000",
    23601 => x"00000000", 23602 => x"00000000", 23603 => x"00000000",
    23604 => x"00000000", 23605 => x"00000000", 23606 => x"00000000",
    23607 => x"00000000", 23608 => x"00000000", 23609 => x"00000000",
    23610 => x"00000000", 23611 => x"00000000", 23612 => x"00000000",
    23613 => x"00000000", 23614 => x"00000000", 23615 => x"00000000",
    23616 => x"00000000", 23617 => x"00000000", 23618 => x"00000000",
    23619 => x"00000000", 23620 => x"00000000", 23621 => x"00000000",
    23622 => x"00000000", 23623 => x"00000000", 23624 => x"00000000",
    23625 => x"00000000", 23626 => x"00000000", 23627 => x"00000000",
    23628 => x"00000000", 23629 => x"00000000", 23630 => x"00000000",
    23631 => x"00000000", 23632 => x"00000000", 23633 => x"00000000",
    23634 => x"00000000", 23635 => x"00000000", 23636 => x"00000000",
    23637 => x"00000000", 23638 => x"00000000", 23639 => x"00000000",
    23640 => x"00000000", 23641 => x"00000000", 23642 => x"00000000",
    23643 => x"00000000", 23644 => x"00000000", 23645 => x"00000000",
    23646 => x"00000000", 23647 => x"00000000", 23648 => x"00000000",
    23649 => x"00000000", 23650 => x"00000000", 23651 => x"00000000",
    23652 => x"00000000", 23653 => x"00000000", 23654 => x"00000000",
    23655 => x"00000000", 23656 => x"00000000", 23657 => x"00000000",
    23658 => x"00000000", 23659 => x"00000000", 23660 => x"00000000",
    23661 => x"00000000", 23662 => x"00000000", 23663 => x"00000000",
    23664 => x"00000000", 23665 => x"00000000", 23666 => x"00000000",
    23667 => x"00000000", 23668 => x"00000000", 23669 => x"00000000",
    23670 => x"00000000", 23671 => x"00000000", 23672 => x"00000000",
    23673 => x"00000000", 23674 => x"00000000", 23675 => x"00000000",
    23676 => x"00000000", 23677 => x"00000000", 23678 => x"00000000",
    23679 => x"00000000", 23680 => x"00000000", 23681 => x"00000000",
    23682 => x"00000000", 23683 => x"00000000", 23684 => x"00000000",
    23685 => x"00000000", 23686 => x"00000000", 23687 => x"00000000",
    23688 => x"00000000", 23689 => x"00000000", 23690 => x"00000000",
    23691 => x"00000000", 23692 => x"00000000", 23693 => x"00000000",
    23694 => x"00000000", 23695 => x"00000000", 23696 => x"00000000",
    23697 => x"00000000", 23698 => x"00000000", 23699 => x"00000000",
    23700 => x"00000000", 23701 => x"00000000", 23702 => x"00000000",
    23703 => x"00000000", 23704 => x"00000000", 23705 => x"00000000",
    23706 => x"00000000", 23707 => x"00000000", 23708 => x"00000000",
    23709 => x"00000000", 23710 => x"00000000", 23711 => x"00000000",
    23712 => x"00000000", 23713 => x"00000000", 23714 => x"00000000",
    23715 => x"00000000", 23716 => x"00000000", 23717 => x"00000000",
    23718 => x"00000000", 23719 => x"00000000", 23720 => x"00000000",
    23721 => x"00000000", 23722 => x"00000000", 23723 => x"00000000",
    23724 => x"00000000", 23725 => x"00000000", 23726 => x"00000000",
    23727 => x"00000000", 23728 => x"00000000", 23729 => x"00000000",
    23730 => x"00000000", 23731 => x"00000000", 23732 => x"00000000",
    23733 => x"00000000", 23734 => x"00000000", 23735 => x"00000000",
    23736 => x"00000000", 23737 => x"00000000", 23738 => x"00000000",
    23739 => x"00000000", 23740 => x"00000000", 23741 => x"00000000",
    23742 => x"00000000", 23743 => x"00000000", 23744 => x"00000000",
    23745 => x"00000000", 23746 => x"00000000", 23747 => x"00000000",
    23748 => x"00000000", 23749 => x"00000000", 23750 => x"00000000",
    23751 => x"00000000", 23752 => x"00000000", 23753 => x"00000000",
    23754 => x"00000000", 23755 => x"00000000", 23756 => x"00000000",
    23757 => x"00000000", 23758 => x"00000000", 23759 => x"00000000",
    23760 => x"00000000", 23761 => x"00000000", 23762 => x"00000000",
    23763 => x"00000000", 23764 => x"00000000", 23765 => x"00000000",
    23766 => x"00000000", 23767 => x"00000000", 23768 => x"00000000",
    23769 => x"00000000", 23770 => x"00000000", 23771 => x"00000000",
    23772 => x"00000000", 23773 => x"00000000", 23774 => x"00000000",
    23775 => x"00000000", 23776 => x"00000000", 23777 => x"00000000",
    23778 => x"00000000", 23779 => x"00000000", 23780 => x"00000000",
    23781 => x"00000000", 23782 => x"00000000", 23783 => x"00000000",
    23784 => x"00000000", 23785 => x"00000000", 23786 => x"00000000",
    23787 => x"00000000", 23788 => x"00000000", 23789 => x"00000000",
    23790 => x"00000000", 23791 => x"00000000", 23792 => x"00000000",
    23793 => x"00000000", 23794 => x"00000000", 23795 => x"00000000",
    23796 => x"00000000", 23797 => x"00000000", 23798 => x"00000000",
    23799 => x"00000000", 23800 => x"00000000", 23801 => x"00000000",
    23802 => x"00000000", 23803 => x"00000000", 23804 => x"00000000",
    23805 => x"00000000", 23806 => x"00000000", 23807 => x"00000000",
    23808 => x"00000000", 23809 => x"00000000", 23810 => x"00000000",
    23811 => x"00000000", 23812 => x"00000000", 23813 => x"00000000",
    23814 => x"00000000", 23815 => x"00000000", 23816 => x"00000000",
    23817 => x"00000000", 23818 => x"00000000", 23819 => x"00000000",
    23820 => x"00000000", 23821 => x"00000000", 23822 => x"00000000",
    23823 => x"00000000", 23824 => x"00000000", 23825 => x"00000000",
    23826 => x"00000000", 23827 => x"00000000", 23828 => x"00000000",
    23829 => x"00000000", 23830 => x"00000000", 23831 => x"00000000",
    23832 => x"00000000", 23833 => x"00000000", 23834 => x"00000000",
    23835 => x"00000000", 23836 => x"00000000", 23837 => x"00000000",
    23838 => x"00000000", 23839 => x"00000000", 23840 => x"00000000",
    23841 => x"00000000", 23842 => x"00000000", 23843 => x"00000000",
    23844 => x"00000000", 23845 => x"00000000", 23846 => x"00000000",
    23847 => x"00000000", 23848 => x"00000000", 23849 => x"00000000",
    23850 => x"00000000", 23851 => x"00000000", 23852 => x"00000000",
    23853 => x"00000000", 23854 => x"00000000", 23855 => x"00000000",
    23856 => x"00000000", 23857 => x"00000000", 23858 => x"00000000",
    23859 => x"00000000", 23860 => x"00000000", 23861 => x"00000000",
    23862 => x"00000000", 23863 => x"00000000", 23864 => x"00000000",
    23865 => x"00000000", 23866 => x"00000000", 23867 => x"00000000",
    23868 => x"00000000", 23869 => x"00000000", 23870 => x"00000000",
    23871 => x"00000000", 23872 => x"00000000", 23873 => x"00000000",
    23874 => x"00000000", 23875 => x"00000000", 23876 => x"00000000",
    23877 => x"00000000", 23878 => x"00000000", 23879 => x"00000000",
    23880 => x"00000000", 23881 => x"00000000", 23882 => x"00000000",
    23883 => x"00000000", 23884 => x"00000000", 23885 => x"00000000",
    23886 => x"00000000", 23887 => x"00000000", 23888 => x"00000000",
    23889 => x"00000000", 23890 => x"00000000", 23891 => x"00000000",
    23892 => x"00000000", 23893 => x"00000000", 23894 => x"00000000",
    23895 => x"00000000", 23896 => x"00000000", 23897 => x"00000000",
    23898 => x"00000000", 23899 => x"00000000", 23900 => x"00000000",
    23901 => x"00000000", 23902 => x"00000000", 23903 => x"00000000",
    23904 => x"00000000", 23905 => x"00000000", 23906 => x"00000000",
    23907 => x"00000000", 23908 => x"00000000", 23909 => x"00000000",
    23910 => x"00000000", 23911 => x"00000000", 23912 => x"00000000",
    23913 => x"00000000", 23914 => x"00000000", 23915 => x"00000000",
    23916 => x"00000000", 23917 => x"00000000", 23918 => x"00000000",
    23919 => x"00000000", 23920 => x"00000000", 23921 => x"00000000",
    23922 => x"00000000", 23923 => x"00000000", 23924 => x"00000000",
    23925 => x"00000000", 23926 => x"00000000", 23927 => x"00000000",
    23928 => x"00000000", 23929 => x"00000000", 23930 => x"00000000",
    23931 => x"00000000", 23932 => x"00000000", 23933 => x"00000000",
    23934 => x"00000000", 23935 => x"00000000", 23936 => x"00000000",
    23937 => x"00000000", 23938 => x"00000000", 23939 => x"00000000",
    23940 => x"00000000", 23941 => x"00000000", 23942 => x"00000000",
    23943 => x"00000000", 23944 => x"00000000", 23945 => x"00000000",
    23946 => x"00000000", 23947 => x"00000000", 23948 => x"00000000",
    23949 => x"00000000", 23950 => x"00000000", 23951 => x"00000000",
    23952 => x"00000000", 23953 => x"00000000", 23954 => x"00000000",
    23955 => x"00000000", 23956 => x"00000000", 23957 => x"00000000",
    23958 => x"00000000", 23959 => x"00000000", 23960 => x"00000000",
    23961 => x"00000000", 23962 => x"00000000", 23963 => x"00000000",
    23964 => x"00000000", 23965 => x"00000000", 23966 => x"00000000",
    23967 => x"00000000", 23968 => x"00000000", 23969 => x"00000000",
    23970 => x"00000000", 23971 => x"00000000", 23972 => x"00000000",
    23973 => x"00000000", 23974 => x"00000000", 23975 => x"00000000",
    23976 => x"00000000", 23977 => x"00000000", 23978 => x"00000000",
    23979 => x"00000000", 23980 => x"00000000", 23981 => x"00000000",
    23982 => x"00000000", 23983 => x"00000000", 23984 => x"00000000",
    23985 => x"00000000", 23986 => x"00000000", 23987 => x"00000000",
    23988 => x"00000000", 23989 => x"00000000", 23990 => x"00000000",
    23991 => x"00000000", 23992 => x"00000000", 23993 => x"00000000",
    23994 => x"00000000", 23995 => x"00000000", 23996 => x"00000000",
    23997 => x"00000000", 23998 => x"00000000", 23999 => x"00000000",
    24000 => x"00000000", 24001 => x"00000000", 24002 => x"00000000",
    24003 => x"00000000", 24004 => x"00000000", 24005 => x"00000000",
    24006 => x"00000000", 24007 => x"00000000", 24008 => x"00000000",
    24009 => x"00000000", 24010 => x"00000000", 24011 => x"00000000",
    24012 => x"00000000", 24013 => x"00000000", 24014 => x"00000000",
    24015 => x"00000000", 24016 => x"00000000", 24017 => x"00000000",
    24018 => x"00000000", 24019 => x"00000000", 24020 => x"00000000",
    24021 => x"00000000", 24022 => x"00000000", 24023 => x"00000000",
    24024 => x"00000000", 24025 => x"00000000", 24026 => x"00000000",
    24027 => x"00000000", 24028 => x"00000000", 24029 => x"00000000",
    24030 => x"00000000", 24031 => x"00000000", 24032 => x"00000000",
    24033 => x"00000000", 24034 => x"00000000", 24035 => x"00000000",
    24036 => x"00000000", 24037 => x"00000000", 24038 => x"00000000",
    24039 => x"00000000", 24040 => x"00000000", 24041 => x"00000000",
    24042 => x"00000000", 24043 => x"00000000", 24044 => x"00000000",
    24045 => x"00000000", 24046 => x"00000000", 24047 => x"00000000",
    24048 => x"00000000", 24049 => x"00000000", 24050 => x"00000000",
    24051 => x"00000000", 24052 => x"00000000", 24053 => x"00000000",
    24054 => x"00000000", 24055 => x"00000000", 24056 => x"00000000",
    24057 => x"00000000", 24058 => x"00000000", 24059 => x"00000000",
    24060 => x"00000000", 24061 => x"00000000", 24062 => x"00000000",
    24063 => x"00000000", 24064 => x"00000000", 24065 => x"00000000",
    24066 => x"00000000", 24067 => x"00000000", 24068 => x"00000000",
    24069 => x"00000000", 24070 => x"00000000", 24071 => x"00000000",
    24072 => x"00000000", 24073 => x"00000000", 24074 => x"00000000",
    24075 => x"00000000", 24076 => x"00000000", 24077 => x"00000000",
    24078 => x"00000000", 24079 => x"00000000", 24080 => x"00000000",
    24081 => x"00000000", 24082 => x"00000000", 24083 => x"00000000",
    24084 => x"00000000", 24085 => x"00000000", 24086 => x"00000000",
    24087 => x"00000000", 24088 => x"00000000", 24089 => x"00000000",
    24090 => x"00000000", 24091 => x"00000000", 24092 => x"00000000",
    24093 => x"00000000", 24094 => x"00000000", 24095 => x"00000000",
    24096 => x"00000000", 24097 => x"00000000", 24098 => x"00000000",
    24099 => x"00000000", 24100 => x"00000000", 24101 => x"00000000",
    24102 => x"00000000", 24103 => x"00000000", 24104 => x"00000000",
    24105 => x"00000000", 24106 => x"00000000", 24107 => x"00000000",
    24108 => x"00000000", 24109 => x"00000000", 24110 => x"00000000",
    24111 => x"00000000", 24112 => x"00000000", 24113 => x"00000000",
    24114 => x"00000000", 24115 => x"00000000", 24116 => x"00000000",
    24117 => x"00000000", 24118 => x"00000000", 24119 => x"00000000",
    24120 => x"00000000", 24121 => x"00000000", 24122 => x"00000000",
    24123 => x"00000000", 24124 => x"00000000", 24125 => x"00000000",
    24126 => x"00000000", 24127 => x"00000000", 24128 => x"00000000",
    24129 => x"00000000", 24130 => x"00000000", 24131 => x"00000000",
    24132 => x"00000000", 24133 => x"00000000", 24134 => x"00000000",
    24135 => x"00000000", 24136 => x"00000000", 24137 => x"00000000",
    24138 => x"00000000", 24139 => x"00000000", 24140 => x"00000000",
    24141 => x"00000000", 24142 => x"00000000", 24143 => x"00000000",
    24144 => x"00000000", 24145 => x"00000000", 24146 => x"00000000",
    24147 => x"00000000", 24148 => x"00000000", 24149 => x"00000000",
    24150 => x"00000000", 24151 => x"00000000", 24152 => x"00000000",
    24153 => x"00000000", 24154 => x"00000000", 24155 => x"00000000",
    24156 => x"00000000", 24157 => x"00000000", 24158 => x"00000000",
    24159 => x"00000000", 24160 => x"00000000", 24161 => x"00000000",
    24162 => x"00000000", 24163 => x"00000000", 24164 => x"00000000",
    24165 => x"00000000", 24166 => x"00000000", 24167 => x"00000000",
    24168 => x"00000000", 24169 => x"00000000", 24170 => x"00000000",
    24171 => x"00000000", 24172 => x"00000000", 24173 => x"00000000",
    24174 => x"00000000", 24175 => x"00000000", 24176 => x"00000000",
    24177 => x"00000000", 24178 => x"00000000", 24179 => x"00000000",
    24180 => x"00000000", 24181 => x"00000000", 24182 => x"00000000",
    24183 => x"00000000", 24184 => x"00000000", 24185 => x"00000000",
    24186 => x"00000000", 24187 => x"00000000", 24188 => x"00000000",
    24189 => x"00000000", 24190 => x"00000000", 24191 => x"00000000",
    24192 => x"00000000", 24193 => x"00000000", 24194 => x"00000000",
    24195 => x"00000000", 24196 => x"00000000", 24197 => x"00000000",
    24198 => x"00000000", 24199 => x"00000000", 24200 => x"00000000",
    24201 => x"00000000", 24202 => x"00000000", 24203 => x"00000000",
    24204 => x"00000000", 24205 => x"00000000", 24206 => x"00000000",
    24207 => x"00000000", 24208 => x"00000000", 24209 => x"00000000",
    24210 => x"00000000", 24211 => x"00000000", 24212 => x"00000000",
    24213 => x"00000000", 24214 => x"00000000", 24215 => x"00000000",
    24216 => x"00000000", 24217 => x"00000000", 24218 => x"00000000",
    24219 => x"00000000", 24220 => x"00000000", 24221 => x"00000000",
    24222 => x"00000000", 24223 => x"00000000", 24224 => x"00000000",
    24225 => x"00000000", 24226 => x"00000000", 24227 => x"00000000",
    24228 => x"00000000", 24229 => x"00000000", 24230 => x"00000000",
    24231 => x"00000000", 24232 => x"00000000", 24233 => x"00000000",
    24234 => x"00000000", 24235 => x"00000000", 24236 => x"00000000",
    24237 => x"00000000", 24238 => x"00000000", 24239 => x"00000000",
    24240 => x"00000000", 24241 => x"00000000", 24242 => x"00000000",
    24243 => x"00000000", 24244 => x"00000000", 24245 => x"00000000",
    24246 => x"00000000", 24247 => x"00000000", 24248 => x"00000000",
    24249 => x"00000000", 24250 => x"00000000", 24251 => x"00000000",
    24252 => x"00000000", 24253 => x"00000000", 24254 => x"00000000",
    24255 => x"00000000", 24256 => x"00000000", 24257 => x"00000000",
    24258 => x"00000000", 24259 => x"00000000", 24260 => x"00000000",
    24261 => x"00000000", 24262 => x"00000000", 24263 => x"00000000",
    24264 => x"00000000", 24265 => x"00000000", 24266 => x"00000000",
    24267 => x"00000000", 24268 => x"00000000", 24269 => x"00000000",
    24270 => x"00000000", 24271 => x"00000000", 24272 => x"00000000",
    24273 => x"00000000", 24274 => x"00000000", 24275 => x"00000000",
    24276 => x"00000000", 24277 => x"00000000", 24278 => x"00000000",
    24279 => x"00000000", 24280 => x"00000000", 24281 => x"00000000",
    24282 => x"00000000", 24283 => x"00000000", 24284 => x"00000000",
    24285 => x"00000000", 24286 => x"00000000", 24287 => x"00000000",
    24288 => x"00000000", 24289 => x"00000000", 24290 => x"00000000",
    24291 => x"00000000", 24292 => x"00000000", 24293 => x"00000000",
    24294 => x"00000000", 24295 => x"00000000", 24296 => x"00000000",
    24297 => x"00000000", 24298 => x"00000000", 24299 => x"00000000",
    24300 => x"00000000", 24301 => x"00000000", 24302 => x"00000000",
    24303 => x"00000000", 24304 => x"00000000", 24305 => x"00000000",
    24306 => x"00000000", 24307 => x"00000000", 24308 => x"00000000",
    24309 => x"00000000", 24310 => x"00000000", 24311 => x"00000000",
    24312 => x"00000000", 24313 => x"00000000", 24314 => x"00000000",
    24315 => x"00000000", 24316 => x"00000000", 24317 => x"00000000",
    24318 => x"00000000", 24319 => x"00000000", 24320 => x"00000000",
    24321 => x"00000000", 24322 => x"00000000", 24323 => x"00000000",
    24324 => x"00000000", 24325 => x"00000000", 24326 => x"00000000",
    24327 => x"00000000", 24328 => x"00000000", 24329 => x"00000000",
    24330 => x"00000000", 24331 => x"00000000", 24332 => x"00000000",
    24333 => x"00000000", 24334 => x"00000000", 24335 => x"00000000",
    24336 => x"00000000", 24337 => x"00000000", 24338 => x"00000000",
    24339 => x"00000000", 24340 => x"00000000", 24341 => x"00000000",
    24342 => x"00000000", 24343 => x"00000000", 24344 => x"00000000",
    24345 => x"00000000", 24346 => x"00000000", 24347 => x"00000000",
    24348 => x"00000000", 24349 => x"00000000", 24350 => x"00000000",
    24351 => x"00000000", 24352 => x"00000000", 24353 => x"00000000",
    24354 => x"00000000", 24355 => x"00000000", 24356 => x"00000000",
    24357 => x"00000000", 24358 => x"00000000", 24359 => x"00000000",
    24360 => x"00000000", 24361 => x"00000000", 24362 => x"00000000",
    24363 => x"00000000", 24364 => x"00000000", 24365 => x"00000000",
    24366 => x"00000000", 24367 => x"00000000", 24368 => x"00000000",
    24369 => x"00000000", 24370 => x"00000000", 24371 => x"00000000",
    24372 => x"00000000", 24373 => x"00000000", 24374 => x"00000000",
    24375 => x"00000000", 24376 => x"00000000", 24377 => x"00000000",
    24378 => x"00000000", 24379 => x"00000000", 24380 => x"00000000",
    24381 => x"00000000", 24382 => x"00000000", 24383 => x"00000000",
    24384 => x"00000000", 24385 => x"00000000", 24386 => x"00000000",
    24387 => x"00000000", 24388 => x"00000000", 24389 => x"00000000",
    24390 => x"00000000", 24391 => x"00000000", 24392 => x"00000000",
    24393 => x"00000000", 24394 => x"00000000", 24395 => x"00000000",
    24396 => x"00000000", 24397 => x"00000000", 24398 => x"00000000",
    24399 => x"00000000", 24400 => x"00000000", 24401 => x"00000000",
    24402 => x"00000000", 24403 => x"00000000", 24404 => x"00000000",
    24405 => x"00000000", 24406 => x"00000000", 24407 => x"00000000",
    24408 => x"00000000", 24409 => x"00000000", 24410 => x"00000000",
    24411 => x"00000000", 24412 => x"00000000", 24413 => x"00000000",
    24414 => x"00000000", 24415 => x"00000000", 24416 => x"00000000",
    24417 => x"00000000", 24418 => x"00000000", 24419 => x"00000000",
    24420 => x"00000000", 24421 => x"00000000", 24422 => x"00000000",
    24423 => x"00000000", 24424 => x"00000000", 24425 => x"00000000",
    24426 => x"00000000", 24427 => x"00000000", 24428 => x"00000000",
    24429 => x"00000000", 24430 => x"00000000", 24431 => x"00000000",
    24432 => x"00000000", 24433 => x"00000000", 24434 => x"00000000",
    24435 => x"00000000", 24436 => x"00000000", 24437 => x"00000000",
    24438 => x"00000000", 24439 => x"00000000", 24440 => x"00000000",
    24441 => x"00000000", 24442 => x"00000000", 24443 => x"00000000",
    24444 => x"00000000", 24445 => x"00000000", 24446 => x"00000000",
    24447 => x"00000000", 24448 => x"00000000", 24449 => x"00000000",
    24450 => x"00000000", 24451 => x"00000000", 24452 => x"00000000",
    24453 => x"00000000", 24454 => x"00000000", 24455 => x"00000000",
    24456 => x"00000000", 24457 => x"00000000", 24458 => x"00000000",
    24459 => x"00000000", 24460 => x"00000000", 24461 => x"00000000",
    24462 => x"00000000", 24463 => x"00000000", 24464 => x"00000000",
    24465 => x"00000000", 24466 => x"00000000", 24467 => x"00000000",
    24468 => x"00000000", 24469 => x"00000000", 24470 => x"00000000",
    24471 => x"00000000", 24472 => x"00000000", 24473 => x"00000000",
    24474 => x"00000000", 24475 => x"00000000", 24476 => x"00000000",
    24477 => x"00000000", 24478 => x"00000000", 24479 => x"00000000",
    24480 => x"00000000", 24481 => x"00000000", 24482 => x"00000000",
    24483 => x"00000000", 24484 => x"00000000", 24485 => x"00000000",
    24486 => x"00000000", 24487 => x"00000000", 24488 => x"00000000",
    24489 => x"00000000", 24490 => x"00000000", 24491 => x"00000000",
    24492 => x"00000000", 24493 => x"00000000", 24494 => x"00000000",
    24495 => x"00000000", 24496 => x"00000000", 24497 => x"00000000",
    24498 => x"00000000", 24499 => x"00000000", 24500 => x"00000000",
    24501 => x"00000000", 24502 => x"00000000", 24503 => x"00000000",
    24504 => x"00000000", 24505 => x"00000000", 24506 => x"00000000",
    24507 => x"00000000", 24508 => x"00000000", 24509 => x"00000000",
    24510 => x"00000000", 24511 => x"00000000", 24512 => x"00000000",
    24513 => x"00000000", 24514 => x"00000000", 24515 => x"00000000",
    24516 => x"00000000", 24517 => x"00000000", 24518 => x"00000000",
    24519 => x"00000000", 24520 => x"00000000", 24521 => x"00000000",
    24522 => x"00000000", 24523 => x"00000000", 24524 => x"00000000",
    24525 => x"00000000", 24526 => x"00000000", 24527 => x"00000000",
    24528 => x"00000000", 24529 => x"00000000", 24530 => x"00000000",
    24531 => x"00000000", 24532 => x"00000000", 24533 => x"00000000",
    24534 => x"00000000", 24535 => x"00000000", 24536 => x"00000000",
    24537 => x"00000000", 24538 => x"00000000", 24539 => x"00000000",
    24540 => x"00000000", 24541 => x"00000000", 24542 => x"00000000",
    24543 => x"00000000", 24544 => x"00000000", 24545 => x"00000000",
    24546 => x"00000000", 24547 => x"00000000", 24548 => x"00000000",
    24549 => x"00000000", 24550 => x"00000000", 24551 => x"00000000",
    24552 => x"00000000", 24553 => x"00000000", 24554 => x"00000000",
    24555 => x"00000000", 24556 => x"00000000", 24557 => x"00000000",
    24558 => x"00000000", 24559 => x"00000000", 24560 => x"00000000",
    24561 => x"00000000", 24562 => x"00000000", 24563 => x"00000000",
    24564 => x"00000000", 24565 => x"00000000", 24566 => x"00000000",
    24567 => x"00000000", 24568 => x"00000000", 24569 => x"00000000",
    24570 => x"00000000", 24571 => x"00000000", 24572 => x"00000000",
    24573 => x"00000000", 24574 => x"00000000", 24575 => x"00000000",
    24576 => x"00000000", 24577 => x"00000000", 24578 => x"00000000",
    24579 => x"00000000", 24580 => x"00000000", 24581 => x"00000000",
    24582 => x"00000000", 24583 => x"00000000", 24584 => x"00000000",
    24585 => x"00000000", 24586 => x"00000000", 24587 => x"00000000",
    24588 => x"00000000", 24589 => x"00000000", 24590 => x"00000000",
    24591 => x"00000000", 24592 => x"00000000", 24593 => x"00000000",
    24594 => x"00000000", 24595 => x"00000000", 24596 => x"00000000",
    24597 => x"00000000", 24598 => x"00000000", 24599 => x"00000000",
    24600 => x"00000000", 24601 => x"00000000", 24602 => x"00000000",
    24603 => x"00000000", 24604 => x"00000000", 24605 => x"00000000",
    24606 => x"00000000", 24607 => x"00000000", 24608 => x"00000000",
    24609 => x"00000000", 24610 => x"00000000", 24611 => x"00000000",
    24612 => x"00000000", 24613 => x"00000000", 24614 => x"00000000",
    24615 => x"00000000", 24616 => x"00000000", 24617 => x"00000000",
    24618 => x"00000000", 24619 => x"00000000", 24620 => x"00000000",
    24621 => x"00000000", 24622 => x"00000000", 24623 => x"00000000",
    24624 => x"00000000", 24625 => x"00000000", 24626 => x"00000000",
    24627 => x"00000000", 24628 => x"00000000", 24629 => x"00000000",
    24630 => x"00000000", 24631 => x"00000000", 24632 => x"00000000",
    24633 => x"00000000", 24634 => x"00000000", 24635 => x"00000000",
    24636 => x"00000000", 24637 => x"00000000", 24638 => x"00000000",
    24639 => x"00000000", 24640 => x"00000000", 24641 => x"00000000",
    24642 => x"00000000", 24643 => x"00000000", 24644 => x"00000000",
    24645 => x"00000000", 24646 => x"00000000", 24647 => x"00000000",
    24648 => x"00000000", 24649 => x"00000000", 24650 => x"00000000",
    24651 => x"00000000", 24652 => x"00000000", 24653 => x"00000000",
    24654 => x"00000000", 24655 => x"00000000", 24656 => x"00000000",
    24657 => x"00000000", 24658 => x"00000000", 24659 => x"00000000",
    24660 => x"00000000", 24661 => x"00000000", 24662 => x"00000000",
    24663 => x"00000000", 24664 => x"00000000", 24665 => x"00000000",
    24666 => x"00000000", 24667 => x"00000000", 24668 => x"00000000",
    24669 => x"00000000", 24670 => x"00000000", 24671 => x"00000000",
    24672 => x"00000000", 24673 => x"00000000", 24674 => x"00000000",
    24675 => x"00000000", 24676 => x"00000000", 24677 => x"00000000",
    24678 => x"00000000", 24679 => x"00000000", 24680 => x"00000000",
    24681 => x"00000000", 24682 => x"00000000", 24683 => x"00000000",
    24684 => x"00000000", 24685 => x"00000000", 24686 => x"00000000",
    24687 => x"00000000", 24688 => x"00000000", 24689 => x"00000000",
    24690 => x"00000000", 24691 => x"00000000", 24692 => x"00000000",
    24693 => x"00000000", 24694 => x"00000000", 24695 => x"00000000",
    24696 => x"00000000", 24697 => x"00000000", 24698 => x"00000000",
    24699 => x"00000000", 24700 => x"00000000", 24701 => x"00000000",
    24702 => x"00000000", 24703 => x"00000000", 24704 => x"00000000",
    24705 => x"00000000", 24706 => x"00000000", 24707 => x"00000000",
    24708 => x"00000000", 24709 => x"00000000", 24710 => x"00000000",
    24711 => x"00000000", 24712 => x"00000000", 24713 => x"00000000",
    24714 => x"00000000", 24715 => x"00000000", 24716 => x"00000000",
    24717 => x"00000000", 24718 => x"00000000", 24719 => x"00000000",
    24720 => x"00000000", 24721 => x"00000000", 24722 => x"00000000",
    24723 => x"00000000", 24724 => x"00000000", 24725 => x"00000000",
    24726 => x"00000000", 24727 => x"00000000", 24728 => x"00000000",
    24729 => x"00000000", 24730 => x"00000000", 24731 => x"00000000",
    24732 => x"00000000", 24733 => x"00000000", 24734 => x"00000000",
    24735 => x"00000000", 24736 => x"00000000", 24737 => x"00000000",
    24738 => x"00000000", 24739 => x"00000000", 24740 => x"00000000",
    24741 => x"00000000", 24742 => x"00000000", 24743 => x"00000000",
    24744 => x"00000000", 24745 => x"00000000", 24746 => x"00000000",
    24747 => x"00000000", 24748 => x"00000000", 24749 => x"00000000",
    24750 => x"00000000", 24751 => x"00000000", 24752 => x"00000000",
    24753 => x"00000000", 24754 => x"00000000", 24755 => x"00000000",
    24756 => x"00000000", 24757 => x"00000000", 24758 => x"00000000",
    24759 => x"00000000", 24760 => x"00000000", 24761 => x"00000000",
    24762 => x"00000000", 24763 => x"00000000", 24764 => x"00000000",
    24765 => x"00000000", 24766 => x"00000000", 24767 => x"00000000",
    24768 => x"00000000", 24769 => x"00000000", 24770 => x"00000000",
    24771 => x"00000000", 24772 => x"00000000", 24773 => x"00000000",
    24774 => x"00000000", 24775 => x"00000000", 24776 => x"00000000",
    24777 => x"00000000", 24778 => x"00000000", 24779 => x"00000000",
    24780 => x"00000000", 24781 => x"00000000", 24782 => x"00000000",
    24783 => x"00000000", 24784 => x"00000000", 24785 => x"00000000",
    24786 => x"00000000", 24787 => x"00000000", 24788 => x"00000000",
    24789 => x"00000000", 24790 => x"00000000", 24791 => x"00000000",
    24792 => x"00000000", 24793 => x"00000000", 24794 => x"00000000",
    24795 => x"00000000", 24796 => x"00000000", 24797 => x"00000000",
    24798 => x"00000000", 24799 => x"00000000", 24800 => x"00000000",
    24801 => x"00000000", 24802 => x"00000000", 24803 => x"00000000",
    24804 => x"00000000", 24805 => x"00000000", 24806 => x"00000000",
    24807 => x"00000000", 24808 => x"00000000", 24809 => x"00000000",
    24810 => x"00000000", 24811 => x"00000000", 24812 => x"00000000",
    24813 => x"00000000", 24814 => x"00000000", 24815 => x"00000000",
    24816 => x"00000000", 24817 => x"00000000", 24818 => x"00000000",
    24819 => x"00000000", 24820 => x"00000000", 24821 => x"00000000",
    24822 => x"00000000", 24823 => x"00000000", 24824 => x"00000000",
    24825 => x"00000000", 24826 => x"00000000", 24827 => x"00000000",
    24828 => x"00000000", 24829 => x"00000000", 24830 => x"00000000",
    24831 => x"00000000", 24832 => x"00000000", 24833 => x"00000000",
    24834 => x"00000000", 24835 => x"00000000", 24836 => x"00000000",
    24837 => x"00000000", 24838 => x"00000000", 24839 => x"00000000",
    24840 => x"00000000", 24841 => x"00000000", 24842 => x"00000000",
    24843 => x"00000000", 24844 => x"00000000", 24845 => x"00000000",
    24846 => x"00000000", 24847 => x"00000000", 24848 => x"00000000",
    24849 => x"00000000", 24850 => x"00000000", 24851 => x"00000000",
    24852 => x"00000000", 24853 => x"00000000", 24854 => x"00000000",
    24855 => x"00000000", 24856 => x"00000000", 24857 => x"00000000",
    24858 => x"00000000", 24859 => x"00000000", 24860 => x"00000000",
    24861 => x"00000000", 24862 => x"00000000", 24863 => x"00000000",
    24864 => x"00000000", 24865 => x"00000000", 24866 => x"00000000",
    24867 => x"00000000", 24868 => x"00000000", 24869 => x"00000000",
    24870 => x"00000000", 24871 => x"00000000", 24872 => x"00000000",
    24873 => x"00000000", 24874 => x"00000000", 24875 => x"00000000",
    24876 => x"00000000", 24877 => x"00000000", 24878 => x"00000000",
    24879 => x"00000000", 24880 => x"00000000", 24881 => x"00000000",
    24882 => x"00000000", 24883 => x"00000000", 24884 => x"00000000",
    24885 => x"00000000", 24886 => x"00000000", 24887 => x"00000000",
    24888 => x"00000000", 24889 => x"00000000", 24890 => x"00000000",
    24891 => x"00000000", 24892 => x"00000000", 24893 => x"00000000",
    24894 => x"00000000", 24895 => x"00000000", 24896 => x"00000000",
    24897 => x"00000000", 24898 => x"00000000", 24899 => x"00000000",
    24900 => x"00000000", 24901 => x"00000000", 24902 => x"00000000",
    24903 => x"00000000", 24904 => x"00000000", 24905 => x"00000000",
    24906 => x"00000000", 24907 => x"00000000", 24908 => x"00000000",
    24909 => x"00000000", 24910 => x"00000000", 24911 => x"00000000",
    24912 => x"00000000", 24913 => x"00000000", 24914 => x"00000000",
    24915 => x"00000000", 24916 => x"00000000", 24917 => x"00000000",
    24918 => x"00000000", 24919 => x"00000000", 24920 => x"00000000",
    24921 => x"00000000", 24922 => x"00000000", 24923 => x"00000000",
    24924 => x"00000000", 24925 => x"00000000", 24926 => x"00000000",
    24927 => x"00000000", 24928 => x"00000000", 24929 => x"00000000",
    24930 => x"00000000", 24931 => x"00000000", 24932 => x"00000000",
    24933 => x"00000000", 24934 => x"00000000", 24935 => x"00000000",
    24936 => x"00000000", 24937 => x"00000000", 24938 => x"00000000",
    24939 => x"00000000", 24940 => x"00000000", 24941 => x"00000000",
    24942 => x"00000000", 24943 => x"00000000", 24944 => x"00000000",
    24945 => x"00000000", 24946 => x"00000000", 24947 => x"00000000",
    24948 => x"00000000", 24949 => x"00000000", 24950 => x"00000000",
    24951 => x"00000000", 24952 => x"00000000", 24953 => x"00000000",
    24954 => x"00000000", 24955 => x"00000000", 24956 => x"00000000",
    24957 => x"00000000", 24958 => x"00000000", 24959 => x"00000000",
    24960 => x"00000000", 24961 => x"00000000", 24962 => x"00000000",
    24963 => x"00000000", 24964 => x"00000000", 24965 => x"00000000",
    24966 => x"00000000", 24967 => x"00000000", 24968 => x"00000000",
    24969 => x"00000000", 24970 => x"00000000", 24971 => x"00000000",
    24972 => x"00000000", 24973 => x"00000000", 24974 => x"00000000",
    24975 => x"00000000", 24976 => x"00000000", 24977 => x"00000000",
    24978 => x"00000000", 24979 => x"00000000", 24980 => x"00000000",
    24981 => x"00000000", 24982 => x"00000000", 24983 => x"00000000",
    24984 => x"00000000", 24985 => x"00000000", 24986 => x"00000000",
    24987 => x"00000000", 24988 => x"00000000", 24989 => x"00000000",
    24990 => x"00000000", 24991 => x"00000000", 24992 => x"00000000",
    24993 => x"00000000", 24994 => x"00000000", 24995 => x"00000000",
    24996 => x"00000000", 24997 => x"00000000", 24998 => x"00000000",
    24999 => x"00000000", 25000 => x"00000000", 25001 => x"00000000",
    25002 => x"00000000", 25003 => x"00000000", 25004 => x"00000000",
    25005 => x"00000000", 25006 => x"00000000", 25007 => x"00000000",
    25008 => x"00000000", 25009 => x"00000000", 25010 => x"00000000",
    25011 => x"00000000", 25012 => x"00000000", 25013 => x"00000000",
    25014 => x"00000000", 25015 => x"00000000", 25016 => x"00000000",
    25017 => x"00000000", 25018 => x"00000000", 25019 => x"00000000",
    25020 => x"00000000", 25021 => x"00000000", 25022 => x"00000000",
    25023 => x"00000000", 25024 => x"00000000", 25025 => x"00000000",
    25026 => x"00000000", 25027 => x"00000000", 25028 => x"00000000",
    25029 => x"00000000", 25030 => x"00000000", 25031 => x"00000000",
    25032 => x"00000000", 25033 => x"00000000", 25034 => x"00000000",
    25035 => x"00000000", 25036 => x"00000000", 25037 => x"00000000",
    25038 => x"00000000", 25039 => x"00000000", 25040 => x"00000000",
    25041 => x"00000000", 25042 => x"00000000", 25043 => x"00000000",
    25044 => x"00000000", 25045 => x"00000000", 25046 => x"00000000",
    25047 => x"00000000", 25048 => x"00000000", 25049 => x"00000000",
    25050 => x"00000000", 25051 => x"00000000", 25052 => x"00000000",
    25053 => x"00000000", 25054 => x"00000000", 25055 => x"00000000",
    25056 => x"00000000", 25057 => x"00000000", 25058 => x"00000000",
    25059 => x"00000000", 25060 => x"00000000", 25061 => x"00000000",
    25062 => x"00000000", 25063 => x"00000000", 25064 => x"00000000",
    25065 => x"00000000", 25066 => x"00000000", 25067 => x"00000000",
    25068 => x"00000000", 25069 => x"00000000", 25070 => x"00000000",
    25071 => x"00000000", 25072 => x"00000000", 25073 => x"00000000",
    25074 => x"00000000", 25075 => x"00000000", 25076 => x"00000000",
    25077 => x"00000000", 25078 => x"00000000", 25079 => x"00000000",
    25080 => x"00000000", 25081 => x"00000000", 25082 => x"00000000",
    25083 => x"00000000", 25084 => x"00000000", 25085 => x"00000000",
    25086 => x"00000000", 25087 => x"00000000", 25088 => x"00000000",
    25089 => x"00000000", 25090 => x"00000000", 25091 => x"00000000",
    25092 => x"00000000", 25093 => x"00000000", 25094 => x"00000000",
    25095 => x"00000000", 25096 => x"00000000", 25097 => x"00000000",
    25098 => x"00000000", 25099 => x"00000000", 25100 => x"00000000",
    25101 => x"00000000", 25102 => x"00000000", 25103 => x"00000000",
    25104 => x"00000000", 25105 => x"00000000", 25106 => x"00000000",
    25107 => x"00000000", 25108 => x"00000000", 25109 => x"00000000",
    25110 => x"00000000", 25111 => x"00000000", 25112 => x"00000000",
    25113 => x"00000000", 25114 => x"00000000", 25115 => x"00000000",
    25116 => x"00000000", 25117 => x"00000000", 25118 => x"00000000",
    25119 => x"00000000", 25120 => x"00000000", 25121 => x"00000000",
    25122 => x"00000000", 25123 => x"00000000", 25124 => x"00000000",
    25125 => x"00000000", 25126 => x"00000000", 25127 => x"00000000",
    25128 => x"00000000", 25129 => x"00000000", 25130 => x"00000000",
    25131 => x"00000000", 25132 => x"00000000", 25133 => x"00000000",
    25134 => x"00000000", 25135 => x"00000000", 25136 => x"00000000",
    25137 => x"00000000", 25138 => x"00000000", 25139 => x"00000000",
    25140 => x"00000000", 25141 => x"00000000", 25142 => x"00000000",
    25143 => x"00000000", 25144 => x"00000000", 25145 => x"00000000",
    25146 => x"00000000", 25147 => x"00000000", 25148 => x"00000000",
    25149 => x"00000000", 25150 => x"00000000", 25151 => x"00000000",
    25152 => x"00000000", 25153 => x"00000000", 25154 => x"00000000",
    25155 => x"00000000", 25156 => x"00000000", 25157 => x"00000000",
    25158 => x"00000000", 25159 => x"00000000", 25160 => x"00000000",
    25161 => x"00000000", 25162 => x"00000000", 25163 => x"00000000",
    25164 => x"00000000", 25165 => x"00000000", 25166 => x"00000000",
    25167 => x"00000000", 25168 => x"00000000", 25169 => x"00000000",
    25170 => x"00000000", 25171 => x"00000000", 25172 => x"00000000",
    25173 => x"00000000", 25174 => x"00000000", 25175 => x"00000000",
    25176 => x"00000000", 25177 => x"00000000", 25178 => x"00000000",
    25179 => x"00000000", 25180 => x"00000000", 25181 => x"00000000",
    25182 => x"00000000", 25183 => x"00000000", 25184 => x"00000000",
    25185 => x"00000000", 25186 => x"00000000", 25187 => x"00000000",
    25188 => x"00000000", 25189 => x"00000000", 25190 => x"00000000",
    25191 => x"00000000", 25192 => x"00000000", 25193 => x"00000000",
    25194 => x"00000000", 25195 => x"00000000", 25196 => x"00000000",
    25197 => x"00000000", 25198 => x"00000000", 25199 => x"00000000",
    25200 => x"00000000", 25201 => x"00000000", 25202 => x"00000000",
    25203 => x"00000000", 25204 => x"00000000", 25205 => x"00000000",
    25206 => x"00000000", 25207 => x"00000000", 25208 => x"00000000",
    25209 => x"00000000", 25210 => x"00000000", 25211 => x"00000000",
    25212 => x"00000000", 25213 => x"00000000", 25214 => x"00000000",
    25215 => x"00000000", 25216 => x"00000000", 25217 => x"00000000",
    25218 => x"00000000", 25219 => x"00000000", 25220 => x"00000000",
    25221 => x"00000000", 25222 => x"00000000", 25223 => x"00000000",
    25224 => x"00000000", 25225 => x"00000000", 25226 => x"00000000",
    25227 => x"00000000", 25228 => x"00000000", 25229 => x"00000000",
    25230 => x"00000000", 25231 => x"00000000", 25232 => x"00000000",
    25233 => x"00000000", 25234 => x"00000000", 25235 => x"00000000",
    25236 => x"00000000", 25237 => x"00000000", 25238 => x"00000000",
    25239 => x"00000000", 25240 => x"00000000", 25241 => x"00000000",
    25242 => x"00000000", 25243 => x"00000000", 25244 => x"00000000",
    25245 => x"00000000", 25246 => x"00000000", 25247 => x"00000000",
    25248 => x"00000000", 25249 => x"00000000", 25250 => x"00000000",
    25251 => x"00000000", 25252 => x"00000000", 25253 => x"00000000",
    25254 => x"00000000", 25255 => x"00000000", 25256 => x"00000000",
    25257 => x"00000000", 25258 => x"00000000", 25259 => x"00000000",
    25260 => x"00000000", 25261 => x"00000000", 25262 => x"00000000",
    25263 => x"00000000", 25264 => x"00000000", 25265 => x"00000000",
    25266 => x"00000000", 25267 => x"00000000", 25268 => x"00000000",
    25269 => x"00000000", 25270 => x"00000000", 25271 => x"00000000",
    25272 => x"00000000", 25273 => x"00000000", 25274 => x"00000000",
    25275 => x"00000000", 25276 => x"00000000", 25277 => x"00000000",
    25278 => x"00000000", 25279 => x"00000000", 25280 => x"00000000",
    25281 => x"00000000", 25282 => x"00000000", 25283 => x"00000000",
    25284 => x"00000000", 25285 => x"00000000", 25286 => x"00000000",
    25287 => x"00000000", 25288 => x"00000000", 25289 => x"00000000",
    25290 => x"00000000", 25291 => x"00000000", 25292 => x"00000000",
    25293 => x"00000000", 25294 => x"00000000", 25295 => x"00000000",
    25296 => x"00000000", 25297 => x"00000000", 25298 => x"00000000",
    25299 => x"00000000", 25300 => x"00000000", 25301 => x"00000000",
    25302 => x"00000000", 25303 => x"00000000", 25304 => x"00000000",
    25305 => x"00000000", 25306 => x"00000000", 25307 => x"00000000",
    25308 => x"00000000", 25309 => x"00000000", 25310 => x"00000000",
    25311 => x"00000000", 25312 => x"00000000", 25313 => x"00000000",
    25314 => x"00000000", 25315 => x"00000000", 25316 => x"00000000",
    25317 => x"00000000", 25318 => x"00000000", 25319 => x"00000000",
    25320 => x"00000000", 25321 => x"00000000", 25322 => x"00000000",
    25323 => x"00000000", 25324 => x"00000000", 25325 => x"00000000",
    25326 => x"00000000", 25327 => x"00000000", 25328 => x"00000000",
    25329 => x"00000000", 25330 => x"00000000", 25331 => x"00000000",
    25332 => x"00000000", 25333 => x"00000000", 25334 => x"00000000",
    25335 => x"00000000", 25336 => x"00000000", 25337 => x"00000000",
    25338 => x"00000000", 25339 => x"00000000", 25340 => x"00000000",
    25341 => x"00000000", 25342 => x"00000000", 25343 => x"00000000",
    25344 => x"00000000", 25345 => x"00000000", 25346 => x"00000000",
    25347 => x"00000000", 25348 => x"00000000", 25349 => x"00000000",
    25350 => x"00000000", 25351 => x"00000000", 25352 => x"00000000",
    25353 => x"00000000", 25354 => x"00000000", 25355 => x"00000000",
    25356 => x"00000000", 25357 => x"00000000", 25358 => x"00000000",
    25359 => x"00000000", 25360 => x"00000000", 25361 => x"00000000",
    25362 => x"00000000", 25363 => x"00000000", 25364 => x"00000000",
    25365 => x"00000000", 25366 => x"00000000", 25367 => x"00000000",
    25368 => x"00000000", 25369 => x"00000000", 25370 => x"00000000",
    25371 => x"00000000", 25372 => x"00000000", 25373 => x"00000000",
    25374 => x"00000000", 25375 => x"00000000", 25376 => x"00000000",
    25377 => x"00000000", 25378 => x"00000000", 25379 => x"00000000",
    25380 => x"00000000", 25381 => x"00000000", 25382 => x"00000000",
    25383 => x"00000000", 25384 => x"00000000", 25385 => x"00000000",
    25386 => x"00000000", 25387 => x"00000000", 25388 => x"00000000",
    25389 => x"00000000", 25390 => x"00000000", 25391 => x"00000000",
    25392 => x"00000000", 25393 => x"00000000", 25394 => x"00000000",
    25395 => x"00000000", 25396 => x"00000000", 25397 => x"00000000",
    25398 => x"00000000", 25399 => x"00000000", 25400 => x"00000000",
    25401 => x"00000000", 25402 => x"00000000", 25403 => x"00000000",
    25404 => x"00000000", 25405 => x"00000000", 25406 => x"00000000",
    25407 => x"00000000", 25408 => x"00000000", 25409 => x"00000000",
    25410 => x"00000000", 25411 => x"00000000", 25412 => x"00000000",
    25413 => x"00000000", 25414 => x"00000000", 25415 => x"00000000",
    25416 => x"00000000", 25417 => x"00000000", 25418 => x"00000000",
    25419 => x"00000000", 25420 => x"00000000", 25421 => x"00000000",
    25422 => x"00000000", 25423 => x"00000000", 25424 => x"00000000",
    25425 => x"00000000", 25426 => x"00000000", 25427 => x"00000000",
    25428 => x"00000000", 25429 => x"00000000", 25430 => x"00000000",
    25431 => x"00000000", 25432 => x"00000000", 25433 => x"00000000",
    25434 => x"00000000", 25435 => x"00000000", 25436 => x"00000000",
    25437 => x"00000000", 25438 => x"00000000", 25439 => x"00000000",
    25440 => x"00000000", 25441 => x"00000000", 25442 => x"00000000",
    25443 => x"00000000", 25444 => x"00000000", 25445 => x"00000000",
    25446 => x"00000000", 25447 => x"00000000", 25448 => x"00000000",
    25449 => x"00000000", 25450 => x"00000000", 25451 => x"00000000",
    25452 => x"00000000", 25453 => x"00000000", 25454 => x"00000000",
    25455 => x"00000000", 25456 => x"00000000", 25457 => x"00000000",
    25458 => x"00000000", 25459 => x"00000000", 25460 => x"00000000",
    25461 => x"00000000", 25462 => x"00000000", 25463 => x"00000000",
    25464 => x"00000000", 25465 => x"00000000", 25466 => x"00000000",
    25467 => x"00000000", 25468 => x"00000000", 25469 => x"00000000",
    25470 => x"00000000", 25471 => x"00000000", 25472 => x"00000000",
    25473 => x"00000000", 25474 => x"00000000", 25475 => x"00000000",
    25476 => x"00000000", 25477 => x"00000000", 25478 => x"00000000",
    25479 => x"00000000", 25480 => x"00000000", 25481 => x"00000000",
    25482 => x"00000000", 25483 => x"00000000", 25484 => x"00000000",
    25485 => x"00000000", 25486 => x"00000000", 25487 => x"00000000",
    25488 => x"00000000", 25489 => x"00000000", 25490 => x"00000000",
    25491 => x"00000000", 25492 => x"00000000", 25493 => x"00000000",
    25494 => x"00000000", 25495 => x"00000000", 25496 => x"00000000",
    25497 => x"00000000", 25498 => x"00000000", 25499 => x"00000000",
    25500 => x"00000000", 25501 => x"00000000", 25502 => x"00000000",
    25503 => x"00000000", 25504 => x"00000000", 25505 => x"00000000",
    25506 => x"00000000", 25507 => x"00000000", 25508 => x"00000000",
    25509 => x"00000000", 25510 => x"00000000", 25511 => x"00000000",
    25512 => x"00000000", 25513 => x"00000000", 25514 => x"00000000",
    25515 => x"00000000", 25516 => x"00000000", 25517 => x"00000000",
    25518 => x"00000000", 25519 => x"00000000", 25520 => x"00000000",
    25521 => x"00000000", 25522 => x"00000000", 25523 => x"00000000",
    25524 => x"00000000", 25525 => x"00000000", 25526 => x"00000000",
    25527 => x"00000000", 25528 => x"00000000", 25529 => x"00000000",
    25530 => x"00000000", 25531 => x"00000000", 25532 => x"00000000",
    25533 => x"00000000", 25534 => x"00000000", 25535 => x"00000000",
    25536 => x"00000000", 25537 => x"00000000", 25538 => x"00000000",
    25539 => x"00000000", 25540 => x"00000000", 25541 => x"00000000",
    25542 => x"00000000", 25543 => x"00000000", 25544 => x"00000000",
    25545 => x"00000000", 25546 => x"00000000", 25547 => x"00000000",
    25548 => x"00000000", 25549 => x"00000000", 25550 => x"00000000",
    25551 => x"00000000", 25552 => x"00000000", 25553 => x"00000000",
    25554 => x"00000000", 25555 => x"00000000", 25556 => x"00000000",
    25557 => x"00000000", 25558 => x"00000000", 25559 => x"00000000",
    25560 => x"00000000", 25561 => x"00000000", 25562 => x"00000000",
    25563 => x"00000000", 25564 => x"00000000", 25565 => x"00000000",
    25566 => x"00000000", 25567 => x"00000000", 25568 => x"00000000",
    25569 => x"00000000", 25570 => x"00000000", 25571 => x"00000000",
    25572 => x"00000000", 25573 => x"00000000", 25574 => x"00000000",
    25575 => x"00000000", 25576 => x"00000000", 25577 => x"00000000",
    25578 => x"00000000", 25579 => x"00000000", 25580 => x"00000000",
    25581 => x"00000000", 25582 => x"00000000", 25583 => x"00000000",
    25584 => x"00000000", 25585 => x"00000000", 25586 => x"00000000",
    25587 => x"00000000", 25588 => x"00000000", 25589 => x"00000000",
    25590 => x"00000000", 25591 => x"00000000", 25592 => x"00000000",
    25593 => x"00000000", 25594 => x"00000000", 25595 => x"00000000",
    25596 => x"00000000", 25597 => x"00000000", 25598 => x"00000000",
    25599 => x"00000000", 25600 => x"00000000", 25601 => x"00000000",
    25602 => x"00000000", 25603 => x"00000000", 25604 => x"00000000",
    25605 => x"00000000", 25606 => x"00000000", 25607 => x"00000000",
    25608 => x"00000000", 25609 => x"00000000", 25610 => x"00000000",
    25611 => x"00000000", 25612 => x"00000000", 25613 => x"00000000",
    25614 => x"00000000", 25615 => x"00000000", 25616 => x"00000000",
    25617 => x"00000000", 25618 => x"00000000", 25619 => x"00000000",
    25620 => x"00000000", 25621 => x"00000000", 25622 => x"00000000",
    25623 => x"00000000", 25624 => x"00000000", 25625 => x"00000000",
    25626 => x"00000000", 25627 => x"00000000", 25628 => x"00000000",
    25629 => x"00000000", 25630 => x"00000000", 25631 => x"00000000",
    25632 => x"00000000", 25633 => x"00000000", 25634 => x"00000000",
    25635 => x"00000000", 25636 => x"00000000", 25637 => x"00000000",
    25638 => x"00000000", 25639 => x"00000000", 25640 => x"00000000",
    25641 => x"00000000", 25642 => x"00000000", 25643 => x"00000000",
    25644 => x"00000000", 25645 => x"00000000", 25646 => x"00000000",
    25647 => x"00000000", 25648 => x"00000000", 25649 => x"00000000",
    25650 => x"00000000", 25651 => x"00000000", 25652 => x"00000000",
    25653 => x"00000000", 25654 => x"00000000", 25655 => x"00000000",
    25656 => x"00000000", 25657 => x"00000000", 25658 => x"00000000",
    25659 => x"00000000", 25660 => x"00000000", 25661 => x"00000000",
    25662 => x"00000000", 25663 => x"00000000", 25664 => x"00000000",
    25665 => x"00000000", 25666 => x"00000000", 25667 => x"00000000",
    25668 => x"00000000", 25669 => x"00000000", 25670 => x"00000000",
    25671 => x"00000000", 25672 => x"00000000", 25673 => x"00000000",
    25674 => x"00000000", 25675 => x"00000000", 25676 => x"00000000",
    25677 => x"00000000", 25678 => x"00000000", 25679 => x"00000000",
    25680 => x"00000000", 25681 => x"00000000", 25682 => x"00000000",
    25683 => x"00000000", 25684 => x"00000000", 25685 => x"00000000",
    25686 => x"00000000", 25687 => x"00000000", 25688 => x"00000000",
    25689 => x"00000000", 25690 => x"00000000", 25691 => x"00000000",
    25692 => x"00000000", 25693 => x"00000000", 25694 => x"00000000",
    25695 => x"00000000", 25696 => x"00000000", 25697 => x"00000000",
    25698 => x"00000000", 25699 => x"00000000", 25700 => x"00000000",
    25701 => x"00000000", 25702 => x"00000000", 25703 => x"00000000",
    25704 => x"00000000", 25705 => x"00000000", 25706 => x"00000000",
    25707 => x"00000000", 25708 => x"00000000", 25709 => x"00000000",
    25710 => x"00000000", 25711 => x"00000000", 25712 => x"00000000",
    25713 => x"00000000", 25714 => x"00000000", 25715 => x"00000000",
    25716 => x"00000000", 25717 => x"00000000", 25718 => x"00000000",
    25719 => x"00000000", 25720 => x"00000000", 25721 => x"00000000",
    25722 => x"00000000", 25723 => x"00000000", 25724 => x"00000000",
    25725 => x"00000000", 25726 => x"00000000", 25727 => x"00000000",
    25728 => x"00000000", 25729 => x"00000000", 25730 => x"00000000",
    25731 => x"00000000", 25732 => x"00000000", 25733 => x"00000000",
    25734 => x"00000000", 25735 => x"00000000", 25736 => x"00000000",
    25737 => x"00000000", 25738 => x"00000000", 25739 => x"00000000",
    25740 => x"00000000", 25741 => x"00000000", 25742 => x"00000000",
    25743 => x"00000000", 25744 => x"00000000", 25745 => x"00000000",
    25746 => x"00000000", 25747 => x"00000000", 25748 => x"00000000",
    25749 => x"00000000", 25750 => x"00000000", 25751 => x"00000000",
    25752 => x"00000000", 25753 => x"00000000", 25754 => x"00000000",
    25755 => x"00000000", 25756 => x"00000000", 25757 => x"00000000",
    25758 => x"00000000", 25759 => x"00000000", 25760 => x"00000000",
    25761 => x"00000000", 25762 => x"00000000", 25763 => x"00000000",
    25764 => x"00000000", 25765 => x"00000000", 25766 => x"00000000",
    25767 => x"00000000", 25768 => x"00000000", 25769 => x"00000000",
    25770 => x"00000000", 25771 => x"00000000", 25772 => x"00000000",
    25773 => x"00000000", 25774 => x"00000000", 25775 => x"00000000",
    25776 => x"00000000", 25777 => x"00000000", 25778 => x"00000000",
    25779 => x"00000000", 25780 => x"00000000", 25781 => x"00000000",
    25782 => x"00000000", 25783 => x"00000000", 25784 => x"00000000",
    25785 => x"00000000", 25786 => x"00000000", 25787 => x"00000000",
    25788 => x"00000000", 25789 => x"00000000", 25790 => x"00000000",
    25791 => x"00000000", 25792 => x"00000000", 25793 => x"00000000",
    25794 => x"00000000", 25795 => x"00000000", 25796 => x"00000000",
    25797 => x"00000000", 25798 => x"00000000", 25799 => x"00000000",
    25800 => x"00000000", 25801 => x"00000000", 25802 => x"00000000",
    25803 => x"00000000", 25804 => x"00000000", 25805 => x"00000000",
    25806 => x"00000000", 25807 => x"00000000", 25808 => x"00000000",
    25809 => x"00000000", 25810 => x"00000000", 25811 => x"00000000",
    25812 => x"00000000", 25813 => x"00000000", 25814 => x"00000000",
    25815 => x"00000000", 25816 => x"00000000", 25817 => x"00000000",
    25818 => x"00000000", 25819 => x"00000000", 25820 => x"00000000",
    25821 => x"00000000", 25822 => x"00000000", 25823 => x"00000000",
    25824 => x"00000000", 25825 => x"00000000", 25826 => x"00000000",
    25827 => x"00000000", 25828 => x"00000000", 25829 => x"00000000",
    25830 => x"00000000", 25831 => x"00000000", 25832 => x"00000000",
    25833 => x"00000000", 25834 => x"00000000", 25835 => x"00000000",
    25836 => x"00000000", 25837 => x"00000000", 25838 => x"00000000",
    25839 => x"00000000", 25840 => x"00000000", 25841 => x"00000000",
    25842 => x"00000000", 25843 => x"00000000", 25844 => x"00000000",
    25845 => x"00000000", 25846 => x"00000000", 25847 => x"00000000",
    25848 => x"00000000", 25849 => x"00000000", 25850 => x"00000000",
    25851 => x"00000000", 25852 => x"00000000", 25853 => x"00000000",
    25854 => x"00000000", 25855 => x"00000000", 25856 => x"00000000",
    25857 => x"00000000", 25858 => x"00000000", 25859 => x"00000000",
    25860 => x"00000000", 25861 => x"00000000", 25862 => x"00000000",
    25863 => x"00000000", 25864 => x"00000000", 25865 => x"00000000",
    25866 => x"00000000", 25867 => x"00000000", 25868 => x"00000000",
    25869 => x"00000000", 25870 => x"00000000", 25871 => x"00000000",
    25872 => x"00000000", 25873 => x"00000000", 25874 => x"00000000",
    25875 => x"00000000", 25876 => x"00000000", 25877 => x"00000000",
    25878 => x"00000000", 25879 => x"00000000", 25880 => x"00000000",
    25881 => x"00000000", 25882 => x"00000000", 25883 => x"00000000",
    25884 => x"00000000", 25885 => x"00000000", 25886 => x"00000000",
    25887 => x"00000000", 25888 => x"00000000", 25889 => x"00000000",
    25890 => x"00000000", 25891 => x"00000000", 25892 => x"00000000",
    25893 => x"00000000", 25894 => x"00000000", 25895 => x"00000000",
    25896 => x"00000000", 25897 => x"00000000", 25898 => x"00000000",
    25899 => x"00000000", 25900 => x"00000000", 25901 => x"00000000",
    25902 => x"00000000", 25903 => x"00000000", 25904 => x"00000000",
    25905 => x"00000000", 25906 => x"00000000", 25907 => x"00000000",
    25908 => x"00000000", 25909 => x"00000000", 25910 => x"00000000",
    25911 => x"00000000", 25912 => x"00000000", 25913 => x"00000000",
    25914 => x"00000000", 25915 => x"00000000", 25916 => x"00000000",
    25917 => x"00000000", 25918 => x"00000000", 25919 => x"00000000",
    25920 => x"00000000", 25921 => x"00000000", 25922 => x"00000000",
    25923 => x"00000000", 25924 => x"00000000", 25925 => x"00000000",
    25926 => x"00000000", 25927 => x"00000000", 25928 => x"00000000",
    25929 => x"00000000", 25930 => x"00000000", 25931 => x"00000000",
    25932 => x"00000000", 25933 => x"00000000", 25934 => x"00000000",
    25935 => x"00000000", 25936 => x"00000000", 25937 => x"00000000",
    25938 => x"00000000", 25939 => x"00000000", 25940 => x"00000000",
    25941 => x"00000000", 25942 => x"00000000", 25943 => x"00000000",
    25944 => x"00000000", 25945 => x"00000000", 25946 => x"00000000",
    25947 => x"00000000", 25948 => x"00000000", 25949 => x"00000000",
    25950 => x"00000000", 25951 => x"00000000", 25952 => x"00000000",
    25953 => x"00000000", 25954 => x"00000000", 25955 => x"00000000",
    25956 => x"00000000", 25957 => x"00000000", 25958 => x"00000000",
    25959 => x"00000000", 25960 => x"00000000", 25961 => x"00000000",
    25962 => x"00000000", 25963 => x"00000000", 25964 => x"00000000",
    25965 => x"00000000", 25966 => x"00000000", 25967 => x"00000000",
    25968 => x"00000000", 25969 => x"00000000", 25970 => x"00000000",
    25971 => x"00000000", 25972 => x"00000000", 25973 => x"00000000",
    25974 => x"00000000", 25975 => x"00000000", 25976 => x"00000000",
    25977 => x"00000000", 25978 => x"00000000", 25979 => x"00000000",
    25980 => x"00000000", 25981 => x"00000000", 25982 => x"00000000",
    25983 => x"00000000", 25984 => x"00000000", 25985 => x"00000000",
    25986 => x"00000000", 25987 => x"00000000", 25988 => x"00000000",
    25989 => x"00000000", 25990 => x"00000000", 25991 => x"00000000",
    25992 => x"00000000", 25993 => x"00000000", 25994 => x"00000000",
    25995 => x"00000000", 25996 => x"00000000", 25997 => x"00000000",
    25998 => x"00000000", 25999 => x"00000000", 26000 => x"00000000",
    26001 => x"00000000", 26002 => x"00000000", 26003 => x"00000000",
    26004 => x"00000000", 26005 => x"00000000", 26006 => x"00000000",
    26007 => x"00000000", 26008 => x"00000000", 26009 => x"00000000",
    26010 => x"00000000", 26011 => x"00000000", 26012 => x"00000000",
    26013 => x"00000000", 26014 => x"00000000", 26015 => x"00000000",
    26016 => x"00000000", 26017 => x"00000000", 26018 => x"00000000",
    26019 => x"00000000", 26020 => x"00000000", 26021 => x"00000000",
    26022 => x"00000000", 26023 => x"00000000", 26024 => x"00000000",
    26025 => x"00000000", 26026 => x"00000000", 26027 => x"00000000",
    26028 => x"00000000", 26029 => x"00000000", 26030 => x"00000000",
    26031 => x"00000000", 26032 => x"00000000", 26033 => x"00000000",
    26034 => x"00000000", 26035 => x"00000000", 26036 => x"00000000",
    26037 => x"00000000", 26038 => x"00000000", 26039 => x"00000000",
    26040 => x"00000000", 26041 => x"00000000", 26042 => x"00000000",
    26043 => x"00000000", 26044 => x"00000000", 26045 => x"00000000",
    26046 => x"00000000", 26047 => x"00000000", 26048 => x"00000000",
    26049 => x"00000000", 26050 => x"00000000", 26051 => x"00000000",
    26052 => x"00000000", 26053 => x"00000000", 26054 => x"00000000",
    26055 => x"00000000", 26056 => x"00000000", 26057 => x"00000000",
    26058 => x"00000000", 26059 => x"00000000", 26060 => x"00000000",
    26061 => x"00000000", 26062 => x"00000000", 26063 => x"00000000",
    26064 => x"00000000", 26065 => x"00000000", 26066 => x"00000000",
    26067 => x"00000000", 26068 => x"00000000", 26069 => x"00000000",
    26070 => x"00000000", 26071 => x"00000000", 26072 => x"00000000",
    26073 => x"00000000", 26074 => x"00000000", 26075 => x"00000000",
    26076 => x"00000000", 26077 => x"00000000", 26078 => x"00000000",
    26079 => x"00000000", 26080 => x"00000000", 26081 => x"00000000",
    26082 => x"00000000", 26083 => x"00000000", 26084 => x"00000000",
    26085 => x"00000000", 26086 => x"00000000", 26087 => x"00000000",
    26088 => x"00000000", 26089 => x"00000000", 26090 => x"00000000",
    26091 => x"00000000", 26092 => x"00000000", 26093 => x"00000000",
    26094 => x"00000000", 26095 => x"00000000", 26096 => x"00000000",
    26097 => x"00000000", 26098 => x"00000000", 26099 => x"00000000",
    26100 => x"00000000", 26101 => x"00000000", 26102 => x"00000000",
    26103 => x"00000000", 26104 => x"00000000", 26105 => x"00000000",
    26106 => x"00000000", 26107 => x"00000000", 26108 => x"00000000",
    26109 => x"00000000", 26110 => x"00000000", 26111 => x"00000000",
    26112 => x"00000000", 26113 => x"00000000", 26114 => x"00000000",
    26115 => x"00000000", 26116 => x"00000000", 26117 => x"00000000",
    26118 => x"00000000", 26119 => x"00000000", 26120 => x"00000000",
    26121 => x"00000000", 26122 => x"00000000", 26123 => x"00000000",
    26124 => x"00000000", 26125 => x"00000000", 26126 => x"00000000",
    26127 => x"00000000", 26128 => x"00000000", 26129 => x"00000000",
    26130 => x"00000000", 26131 => x"00000000", 26132 => x"00000000",
    26133 => x"00000000", 26134 => x"00000000", 26135 => x"00000000",
    26136 => x"00000000", 26137 => x"00000000", 26138 => x"00000000",
    26139 => x"00000000", 26140 => x"00000000", 26141 => x"00000000",
    26142 => x"00000000", 26143 => x"00000000", 26144 => x"00000000",
    26145 => x"00000000", 26146 => x"00000000", 26147 => x"00000000",
    26148 => x"00000000", 26149 => x"00000000", 26150 => x"00000000",
    26151 => x"00000000", 26152 => x"00000000", 26153 => x"00000000",
    26154 => x"00000000", 26155 => x"00000000", 26156 => x"00000000",
    26157 => x"00000000", 26158 => x"00000000", 26159 => x"00000000",
    26160 => x"00000000", 26161 => x"00000000", 26162 => x"00000000",
    26163 => x"00000000", 26164 => x"00000000", 26165 => x"00000000",
    26166 => x"00000000", 26167 => x"00000000", 26168 => x"00000000",
    26169 => x"00000000", 26170 => x"00000000", 26171 => x"00000000",
    26172 => x"00000000", 26173 => x"00000000", 26174 => x"00000000",
    26175 => x"00000000", 26176 => x"00000000", 26177 => x"00000000",
    26178 => x"00000000", 26179 => x"00000000", 26180 => x"00000000",
    26181 => x"00000000", 26182 => x"00000000", 26183 => x"00000000",
    26184 => x"00000000", 26185 => x"00000000", 26186 => x"00000000",
    26187 => x"00000000", 26188 => x"00000000", 26189 => x"00000000",
    26190 => x"00000000", 26191 => x"00000000", 26192 => x"00000000",
    26193 => x"00000000", 26194 => x"00000000", 26195 => x"00000000",
    26196 => x"00000000", 26197 => x"00000000", 26198 => x"00000000",
    26199 => x"00000000", 26200 => x"00000000", 26201 => x"00000000",
    26202 => x"00000000", 26203 => x"00000000", 26204 => x"00000000",
    26205 => x"00000000", 26206 => x"00000000", 26207 => x"00000000",
    26208 => x"00000000", 26209 => x"00000000", 26210 => x"00000000",
    26211 => x"00000000", 26212 => x"00000000", 26213 => x"00000000",
    26214 => x"00000000", 26215 => x"00000000", 26216 => x"00000000",
    26217 => x"00000000", 26218 => x"00000000", 26219 => x"00000000",
    26220 => x"00000000", 26221 => x"00000000", 26222 => x"00000000",
    26223 => x"00000000", 26224 => x"00000000", 26225 => x"00000000",
    26226 => x"00000000", 26227 => x"00000000", 26228 => x"00000000",
    26229 => x"00000000", 26230 => x"00000000", 26231 => x"00000000",
    26232 => x"00000000", 26233 => x"00000000", 26234 => x"00000000",
    26235 => x"00000000", 26236 => x"00000000", 26237 => x"00000000",
    26238 => x"00000000", 26239 => x"00000000", 26240 => x"00000000",
    26241 => x"00000000", 26242 => x"00000000", 26243 => x"00000000",
    26244 => x"00000000", 26245 => x"00000000", 26246 => x"00000000",
    26247 => x"00000000", 26248 => x"00000000", 26249 => x"00000000",
    26250 => x"00000000", 26251 => x"00000000", 26252 => x"00000000",
    26253 => x"00000000", 26254 => x"00000000", 26255 => x"00000000",
    26256 => x"00000000", 26257 => x"00000000", 26258 => x"00000000",
    26259 => x"00000000", 26260 => x"00000000", 26261 => x"00000000",
    26262 => x"00000000", 26263 => x"00000000", 26264 => x"00000000",
    26265 => x"00000000", 26266 => x"00000000", 26267 => x"00000000",
    26268 => x"00000000", 26269 => x"00000000", 26270 => x"00000000",
    26271 => x"00000000", 26272 => x"00000000", 26273 => x"00000000",
    26274 => x"00000000", 26275 => x"00000000", 26276 => x"00000000",
    26277 => x"00000000", 26278 => x"00000000", 26279 => x"00000000",
    26280 => x"00000000", 26281 => x"00000000", 26282 => x"00000000",
    26283 => x"00000000", 26284 => x"00000000", 26285 => x"00000000",
    26286 => x"00000000", 26287 => x"00000000", 26288 => x"00000000",
    26289 => x"00000000", 26290 => x"00000000", 26291 => x"00000000",
    26292 => x"00000000", 26293 => x"00000000", 26294 => x"00000000",
    26295 => x"00000000", 26296 => x"00000000", 26297 => x"00000000",
    26298 => x"00000000", 26299 => x"00000000", 26300 => x"00000000",
    26301 => x"00000000", 26302 => x"00000000", 26303 => x"00000000",
    26304 => x"00000000", 26305 => x"00000000", 26306 => x"00000000",
    26307 => x"00000000", 26308 => x"00000000", 26309 => x"00000000",
    26310 => x"00000000", 26311 => x"00000000", 26312 => x"00000000",
    26313 => x"00000000", 26314 => x"00000000", 26315 => x"00000000",
    26316 => x"00000000", 26317 => x"00000000", 26318 => x"00000000",
    26319 => x"00000000", 26320 => x"00000000", 26321 => x"00000000",
    26322 => x"00000000", 26323 => x"00000000", 26324 => x"00000000",
    26325 => x"00000000", 26326 => x"00000000", 26327 => x"00000000",
    26328 => x"00000000", 26329 => x"00000000", 26330 => x"00000000",
    26331 => x"00000000", 26332 => x"00000000", 26333 => x"00000000",
    26334 => x"00000000", 26335 => x"00000000", 26336 => x"00000000",
    26337 => x"00000000", 26338 => x"00000000", 26339 => x"00000000",
    26340 => x"00000000", 26341 => x"00000000", 26342 => x"00000000",
    26343 => x"00000000", 26344 => x"00000000", 26345 => x"00000000",
    26346 => x"00000000", 26347 => x"00000000", 26348 => x"00000000",
    26349 => x"00000000", 26350 => x"00000000", 26351 => x"00000000",
    26352 => x"00000000", 26353 => x"00000000", 26354 => x"00000000",
    26355 => x"00000000", 26356 => x"00000000", 26357 => x"00000000",
    26358 => x"00000000", 26359 => x"00000000", 26360 => x"00000000",
    26361 => x"00000000", 26362 => x"00000000", 26363 => x"00000000",
    26364 => x"00000000", 26365 => x"00000000", 26366 => x"00000000",
    26367 => x"00000000", 26368 => x"00000000", 26369 => x"00000000",
    26370 => x"00000000", 26371 => x"00000000", 26372 => x"00000000",
    26373 => x"00000000", 26374 => x"00000000", 26375 => x"00000000",
    26376 => x"00000000", 26377 => x"00000000", 26378 => x"00000000",
    26379 => x"00000000", 26380 => x"00000000", 26381 => x"00000000",
    26382 => x"00000000", 26383 => x"00000000", 26384 => x"00000000",
    26385 => x"00000000", 26386 => x"00000000", 26387 => x"00000000",
    26388 => x"00000000", 26389 => x"00000000", 26390 => x"00000000",
    26391 => x"00000000", 26392 => x"00000000", 26393 => x"00000000",
    26394 => x"00000000", 26395 => x"00000000", 26396 => x"00000000",
    26397 => x"00000000", 26398 => x"00000000", 26399 => x"00000000",
    26400 => x"00000000", 26401 => x"00000000", 26402 => x"00000000",
    26403 => x"00000000", 26404 => x"00000000", 26405 => x"00000000",
    26406 => x"00000000", 26407 => x"00000000", 26408 => x"00000000",
    26409 => x"00000000", 26410 => x"00000000", 26411 => x"00000000",
    26412 => x"00000000", 26413 => x"00000000", 26414 => x"00000000",
    26415 => x"00000000", 26416 => x"00000000", 26417 => x"00000000",
    26418 => x"00000000", 26419 => x"00000000", 26420 => x"00000000",
    26421 => x"00000000", 26422 => x"00000000", 26423 => x"00000000",
    26424 => x"00000000", 26425 => x"00000000", 26426 => x"00000000",
    26427 => x"00000000", 26428 => x"00000000", 26429 => x"00000000",
    26430 => x"00000000", 26431 => x"00000000", 26432 => x"00000000",
    26433 => x"00000000", 26434 => x"00000000", 26435 => x"00000000",
    26436 => x"00000000", 26437 => x"00000000", 26438 => x"00000000",
    26439 => x"00000000", 26440 => x"00000000", 26441 => x"00000000",
    26442 => x"00000000", 26443 => x"00000000", 26444 => x"00000000",
    26445 => x"00000000", 26446 => x"00000000", 26447 => x"00000000",
    26448 => x"00000000", 26449 => x"00000000", 26450 => x"00000000",
    26451 => x"00000000", 26452 => x"00000000", 26453 => x"00000000",
    26454 => x"00000000", 26455 => x"00000000", 26456 => x"00000000",
    26457 => x"00000000", 26458 => x"00000000", 26459 => x"00000000",
    26460 => x"00000000", 26461 => x"00000000", 26462 => x"00000000",
    26463 => x"00000000", 26464 => x"00000000", 26465 => x"00000000",
    26466 => x"00000000", 26467 => x"00000000", 26468 => x"00000000",
    26469 => x"00000000", 26470 => x"00000000", 26471 => x"00000000",
    26472 => x"00000000", 26473 => x"00000000", 26474 => x"00000000",
    26475 => x"00000000", 26476 => x"00000000", 26477 => x"00000000",
    26478 => x"00000000", 26479 => x"00000000", 26480 => x"00000000",
    26481 => x"00000000", 26482 => x"00000000", 26483 => x"00000000",
    26484 => x"00000000", 26485 => x"00000000", 26486 => x"00000000",
    26487 => x"00000000", 26488 => x"00000000", 26489 => x"00000000",
    26490 => x"00000000", 26491 => x"00000000", 26492 => x"00000000",
    26493 => x"00000000", 26494 => x"00000000", 26495 => x"00000000",
    26496 => x"00000000", 26497 => x"00000000", 26498 => x"00000000",
    26499 => x"00000000", 26500 => x"00000000", 26501 => x"00000000",
    26502 => x"00000000", 26503 => x"00000000", 26504 => x"00000000",
    26505 => x"00000000", 26506 => x"00000000", 26507 => x"00000000",
    26508 => x"00000000", 26509 => x"00000000", 26510 => x"00000000",
    26511 => x"00000000", 26512 => x"00000000", 26513 => x"00000000",
    26514 => x"00000000", 26515 => x"00000000", 26516 => x"00000000",
    26517 => x"00000000", 26518 => x"00000000", 26519 => x"00000000",
    26520 => x"00000000", 26521 => x"00000000", 26522 => x"00000000",
    26523 => x"00000000", 26524 => x"00000000", 26525 => x"00000000",
    26526 => x"00000000", 26527 => x"00000000", 26528 => x"00000000",
    26529 => x"00000000", 26530 => x"00000000", 26531 => x"00000000",
    26532 => x"00000000", 26533 => x"00000000", 26534 => x"00000000",
    26535 => x"00000000", 26536 => x"00000000", 26537 => x"00000000",
    26538 => x"00000000", 26539 => x"00000000", 26540 => x"00000000",
    26541 => x"00000000", 26542 => x"00000000", 26543 => x"00000000",
    26544 => x"00000000", 26545 => x"00000000", 26546 => x"00000000",
    26547 => x"00000000", 26548 => x"00000000", 26549 => x"00000000",
    26550 => x"00000000", 26551 => x"00000000", 26552 => x"00000000",
    26553 => x"00000000", 26554 => x"00000000", 26555 => x"00000000",
    26556 => x"00000000", 26557 => x"00000000", 26558 => x"00000000",
    26559 => x"00000000", 26560 => x"00000000", 26561 => x"00000000",
    26562 => x"00000000", 26563 => x"00000000", 26564 => x"00000000",
    26565 => x"00000000", 26566 => x"00000000", 26567 => x"00000000",
    26568 => x"00000000", 26569 => x"00000000", 26570 => x"00000000",
    26571 => x"00000000", 26572 => x"00000000", 26573 => x"00000000",
    26574 => x"00000000", 26575 => x"00000000", 26576 => x"00000000",
    26577 => x"00000000", 26578 => x"00000000", 26579 => x"00000000",
    26580 => x"00000000", 26581 => x"00000000", 26582 => x"00000000",
    26583 => x"00000000", 26584 => x"00000000", 26585 => x"00000000",
    26586 => x"00000000", 26587 => x"00000000", 26588 => x"00000000",
    26589 => x"00000000", 26590 => x"00000000", 26591 => x"00000000",
    26592 => x"00000000", 26593 => x"00000000", 26594 => x"00000000",
    26595 => x"00000000", 26596 => x"00000000", 26597 => x"00000000",
    26598 => x"00000000", 26599 => x"00000000", 26600 => x"00000000",
    26601 => x"00000000", 26602 => x"00000000", 26603 => x"00000000",
    26604 => x"00000000", 26605 => x"00000000", 26606 => x"00000000",
    26607 => x"00000000", 26608 => x"00000000", 26609 => x"00000000",
    26610 => x"00000000", 26611 => x"00000000", 26612 => x"00000000",
    26613 => x"00000000", 26614 => x"00000000", 26615 => x"00000000",
    26616 => x"00000000", 26617 => x"00000000", 26618 => x"00000000",
    26619 => x"00000000", 26620 => x"00000000", 26621 => x"00000000",
    26622 => x"00000000", 26623 => x"00000000", 26624 => x"00000000",
    26625 => x"00000000", 26626 => x"00000000", 26627 => x"00000000",
    26628 => x"00000000", 26629 => x"00000000", 26630 => x"00000000",
    26631 => x"00000000", 26632 => x"00000000", 26633 => x"00000000",
    26634 => x"00000000", 26635 => x"00000000", 26636 => x"00000000",
    26637 => x"00000000", 26638 => x"00000000", 26639 => x"00000000",
    26640 => x"00000000", 26641 => x"00000000", 26642 => x"00000000",
    26643 => x"00000000", 26644 => x"00000000", 26645 => x"00000000",
    26646 => x"00000000", 26647 => x"00000000", 26648 => x"00000000",
    26649 => x"00000000", 26650 => x"00000000", 26651 => x"00000000",
    26652 => x"00000000", 26653 => x"00000000", 26654 => x"00000000",
    26655 => x"00000000", 26656 => x"00000000", 26657 => x"00000000",
    26658 => x"00000000", 26659 => x"00000000", 26660 => x"00000000",
    26661 => x"00000000", 26662 => x"00000000", 26663 => x"00000000",
    26664 => x"00000000", 26665 => x"00000000", 26666 => x"00000000",
    26667 => x"00000000", 26668 => x"00000000", 26669 => x"00000000",
    26670 => x"00000000", 26671 => x"00000000", 26672 => x"00000000",
    26673 => x"00000000", 26674 => x"00000000", 26675 => x"00000000",
    26676 => x"00000000", 26677 => x"00000000", 26678 => x"00000000",
    26679 => x"00000000", 26680 => x"00000000", 26681 => x"00000000",
    26682 => x"00000000", 26683 => x"00000000", 26684 => x"00000000",
    26685 => x"00000000", 26686 => x"00000000", 26687 => x"00000000",
    26688 => x"00000000", 26689 => x"00000000", 26690 => x"00000000",
    26691 => x"00000000", 26692 => x"00000000", 26693 => x"00000000",
    26694 => x"00000000", 26695 => x"00000000", 26696 => x"00000000",
    26697 => x"00000000", 26698 => x"00000000", 26699 => x"00000000",
    26700 => x"00000000", 26701 => x"00000000", 26702 => x"00000000",
    26703 => x"00000000", 26704 => x"00000000", 26705 => x"00000000",
    26706 => x"00000000", 26707 => x"00000000", 26708 => x"00000000",
    26709 => x"00000000", 26710 => x"00000000", 26711 => x"00000000",
    26712 => x"00000000", 26713 => x"00000000", 26714 => x"00000000",
    26715 => x"00000000", 26716 => x"00000000", 26717 => x"00000000",
    26718 => x"00000000", 26719 => x"00000000", 26720 => x"00000000",
    26721 => x"00000000", 26722 => x"00000000", 26723 => x"00000000",
    26724 => x"00000000", 26725 => x"00000000", 26726 => x"00000000",
    26727 => x"00000000", 26728 => x"00000000", 26729 => x"00000000",
    26730 => x"00000000", 26731 => x"00000000", 26732 => x"00000000",
    26733 => x"00000000", 26734 => x"00000000", 26735 => x"00000000",
    26736 => x"00000000", 26737 => x"00000000", 26738 => x"00000000",
    26739 => x"00000000", 26740 => x"00000000", 26741 => x"00000000",
    26742 => x"00000000", 26743 => x"00000000", 26744 => x"00000000",
    26745 => x"00000000", 26746 => x"00000000", 26747 => x"00000000",
    26748 => x"00000000", 26749 => x"00000000", 26750 => x"00000000",
    26751 => x"00000000", 26752 => x"00000000", 26753 => x"00000000",
    26754 => x"00000000", 26755 => x"00000000", 26756 => x"00000000",
    26757 => x"00000000", 26758 => x"00000000", 26759 => x"00000000",
    26760 => x"00000000", 26761 => x"00000000", 26762 => x"00000000",
    26763 => x"00000000", 26764 => x"00000000", 26765 => x"00000000",
    26766 => x"00000000", 26767 => x"00000000", 26768 => x"00000000",
    26769 => x"00000000", 26770 => x"00000000", 26771 => x"00000000",
    26772 => x"00000000", 26773 => x"00000000", 26774 => x"00000000",
    26775 => x"00000000", 26776 => x"00000000", 26777 => x"00000000",
    26778 => x"00000000", 26779 => x"00000000", 26780 => x"00000000",
    26781 => x"00000000", 26782 => x"00000000", 26783 => x"00000000",
    26784 => x"00000000", 26785 => x"00000000", 26786 => x"00000000",
    26787 => x"00000000", 26788 => x"00000000", 26789 => x"00000000",
    26790 => x"00000000", 26791 => x"00000000", 26792 => x"00000000",
    26793 => x"00000000", 26794 => x"00000000", 26795 => x"00000000",
    26796 => x"00000000", 26797 => x"00000000", 26798 => x"00000000",
    26799 => x"00000000", 26800 => x"00000000", 26801 => x"00000000",
    26802 => x"00000000", 26803 => x"00000000", 26804 => x"00000000",
    26805 => x"00000000", 26806 => x"00000000", 26807 => x"00000000",
    26808 => x"00000000", 26809 => x"00000000", 26810 => x"00000000",
    26811 => x"00000000", 26812 => x"00000000", 26813 => x"00000000",
    26814 => x"00000000", 26815 => x"00000000", 26816 => x"00000000",
    26817 => x"00000000", 26818 => x"00000000", 26819 => x"00000000",
    26820 => x"00000000", 26821 => x"00000000", 26822 => x"00000000",
    26823 => x"00000000", 26824 => x"00000000", 26825 => x"00000000",
    26826 => x"00000000", 26827 => x"00000000", 26828 => x"00000000",
    26829 => x"00000000", 26830 => x"00000000", 26831 => x"00000000",
    26832 => x"00000000", 26833 => x"00000000", 26834 => x"00000000",
    26835 => x"00000000", 26836 => x"00000000", 26837 => x"00000000",
    26838 => x"00000000", 26839 => x"00000000", 26840 => x"00000000",
    26841 => x"00000000", 26842 => x"00000000", 26843 => x"00000000",
    26844 => x"00000000", 26845 => x"00000000", 26846 => x"00000000",
    26847 => x"00000000", 26848 => x"00000000", 26849 => x"00000000",
    26850 => x"00000000", 26851 => x"00000000", 26852 => x"00000000",
    26853 => x"00000000", 26854 => x"00000000", 26855 => x"00000000",
    26856 => x"00000000", 26857 => x"00000000", 26858 => x"00000000",
    26859 => x"00000000", 26860 => x"00000000", 26861 => x"00000000",
    26862 => x"00000000", 26863 => x"00000000", 26864 => x"00000000",
    26865 => x"00000000", 26866 => x"00000000", 26867 => x"00000000",
    26868 => x"00000000", 26869 => x"00000000", 26870 => x"00000000",
    26871 => x"00000000", 26872 => x"00000000", 26873 => x"00000000",
    26874 => x"00000000", 26875 => x"00000000", 26876 => x"00000000",
    26877 => x"00000000", 26878 => x"00000000", 26879 => x"00000000",
    26880 => x"00000000", 26881 => x"00000000", 26882 => x"00000000",
    26883 => x"00000000", 26884 => x"00000000", 26885 => x"00000000",
    26886 => x"00000000", 26887 => x"00000000", 26888 => x"00000000",
    26889 => x"00000000", 26890 => x"00000000", 26891 => x"00000000",
    26892 => x"00000000", 26893 => x"00000000", 26894 => x"00000000",
    26895 => x"00000000", 26896 => x"00000000", 26897 => x"00000000",
    26898 => x"00000000", 26899 => x"00000000", 26900 => x"00000000",
    26901 => x"00000000", 26902 => x"00000000", 26903 => x"00000000",
    26904 => x"00000000", 26905 => x"00000000", 26906 => x"00000000",
    26907 => x"00000000", 26908 => x"00000000", 26909 => x"00000000",
    26910 => x"00000000", 26911 => x"00000000", 26912 => x"00000000",
    26913 => x"00000000", 26914 => x"00000000", 26915 => x"00000000",
    26916 => x"00000000", 26917 => x"00000000", 26918 => x"00000000",
    26919 => x"00000000", 26920 => x"00000000", 26921 => x"00000000",
    26922 => x"00000000", 26923 => x"00000000", 26924 => x"00000000",
    26925 => x"00000000", 26926 => x"00000000", 26927 => x"00000000",
    26928 => x"00000000", 26929 => x"00000000", 26930 => x"00000000",
    26931 => x"00000000", 26932 => x"00000000", 26933 => x"00000000",
    26934 => x"00000000", 26935 => x"00000000", 26936 => x"00000000",
    26937 => x"00000000", 26938 => x"00000000", 26939 => x"00000000",
    26940 => x"00000000", 26941 => x"00000000", 26942 => x"00000000",
    26943 => x"00000000", 26944 => x"00000000", 26945 => x"00000000",
    26946 => x"00000000", 26947 => x"00000000", 26948 => x"00000000",
    26949 => x"00000000", 26950 => x"00000000", 26951 => x"00000000",
    26952 => x"00000000", 26953 => x"00000000", 26954 => x"00000000",
    26955 => x"00000000", 26956 => x"00000000", 26957 => x"00000000",
    26958 => x"00000000", 26959 => x"00000000", 26960 => x"00000000",
    26961 => x"00000000", 26962 => x"00000000", 26963 => x"00000000",
    26964 => x"00000000", 26965 => x"00000000", 26966 => x"00000000",
    26967 => x"00000000", 26968 => x"00000000", 26969 => x"00000000",
    26970 => x"00000000", 26971 => x"00000000", 26972 => x"00000000",
    26973 => x"00000000", 26974 => x"00000000", 26975 => x"00000000",
    26976 => x"00000000", 26977 => x"00000000", 26978 => x"00000000",
    26979 => x"00000000", 26980 => x"00000000", 26981 => x"00000000",
    26982 => x"00000000", 26983 => x"00000000", 26984 => x"00000000",
    26985 => x"00000000", 26986 => x"00000000", 26987 => x"00000000",
    26988 => x"00000000", 26989 => x"00000000", 26990 => x"00000000",
    26991 => x"00000000", 26992 => x"00000000", 26993 => x"00000000",
    26994 => x"00000000", 26995 => x"00000000", 26996 => x"00000000",
    26997 => x"00000000", 26998 => x"00000000", 26999 => x"00000000",
    27000 => x"00000000", 27001 => x"00000000", 27002 => x"00000000",
    27003 => x"00000000", 27004 => x"00000000", 27005 => x"00000000",
    27006 => x"00000000", 27007 => x"00000000", 27008 => x"00000000",
    27009 => x"00000000", 27010 => x"00000000", 27011 => x"00000000",
    27012 => x"00000000", 27013 => x"00000000", 27014 => x"00000000",
    27015 => x"00000000", 27016 => x"00000000", 27017 => x"00000000",
    27018 => x"00000000", 27019 => x"00000000", 27020 => x"00000000",
    27021 => x"00000000", 27022 => x"00000000", 27023 => x"00000000",
    27024 => x"00000000", 27025 => x"00000000", 27026 => x"00000000",
    27027 => x"00000000", 27028 => x"00000000", 27029 => x"00000000",
    27030 => x"00000000", 27031 => x"00000000", 27032 => x"00000000",
    27033 => x"00000000", 27034 => x"00000000", 27035 => x"00000000",
    27036 => x"00000000", 27037 => x"00000000", 27038 => x"00000000",
    27039 => x"00000000", 27040 => x"00000000", 27041 => x"00000000",
    27042 => x"00000000", 27043 => x"00000000", 27044 => x"00000000",
    27045 => x"00000000", 27046 => x"00000000", 27047 => x"00000000",
    27048 => x"00000000", 27049 => x"00000000", 27050 => x"00000000",
    27051 => x"00000000", 27052 => x"00000000", 27053 => x"00000000",
    27054 => x"00000000", 27055 => x"00000000", 27056 => x"00000000",
    27057 => x"00000000", 27058 => x"00000000", 27059 => x"00000000",
    27060 => x"00000000", 27061 => x"00000000", 27062 => x"00000000",
    27063 => x"00000000", 27064 => x"00000000", 27065 => x"00000000",
    27066 => x"00000000", 27067 => x"00000000", 27068 => x"00000000",
    27069 => x"00000000", 27070 => x"00000000", 27071 => x"00000000",
    27072 => x"00000000", 27073 => x"00000000", 27074 => x"00000000",
    27075 => x"00000000", 27076 => x"00000000", 27077 => x"00000000",
    27078 => x"00000000", 27079 => x"00000000", 27080 => x"00000000",
    27081 => x"00000000", 27082 => x"00000000", 27083 => x"00000000",
    27084 => x"00000000", 27085 => x"00000000", 27086 => x"00000000",
    27087 => x"00000000", 27088 => x"00000000", 27089 => x"00000000",
    27090 => x"00000000", 27091 => x"00000000", 27092 => x"00000000",
    27093 => x"00000000", 27094 => x"00000000", 27095 => x"00000000",
    27096 => x"00000000", 27097 => x"00000000", 27098 => x"00000000",
    27099 => x"00000000", 27100 => x"00000000", 27101 => x"00000000",
    27102 => x"00000000", 27103 => x"00000000", 27104 => x"00000000",
    27105 => x"00000000", 27106 => x"00000000", 27107 => x"00000000",
    27108 => x"00000000", 27109 => x"00000000", 27110 => x"00000000",
    27111 => x"00000000", 27112 => x"00000000", 27113 => x"00000000",
    27114 => x"00000000", 27115 => x"00000000", 27116 => x"00000000",
    27117 => x"00000000", 27118 => x"00000000", 27119 => x"00000000",
    27120 => x"00000000", 27121 => x"00000000", 27122 => x"00000000",
    27123 => x"00000000", 27124 => x"00000000", 27125 => x"00000000",
    27126 => x"00000000", 27127 => x"00000000", 27128 => x"00000000",
    27129 => x"00000000", 27130 => x"00000000", 27131 => x"00000000",
    27132 => x"00000000", 27133 => x"00000000", 27134 => x"00000000",
    27135 => x"00000000", 27136 => x"00000000", 27137 => x"00000000",
    27138 => x"00000000", 27139 => x"00000000", 27140 => x"00000000",
    27141 => x"00000000", 27142 => x"00000000", 27143 => x"00000000",
    27144 => x"00000000", 27145 => x"00000000", 27146 => x"00000000",
    27147 => x"00000000", 27148 => x"00000000", 27149 => x"00000000",
    27150 => x"00000000", 27151 => x"00000000", 27152 => x"00000000",
    27153 => x"00000000", 27154 => x"00000000", 27155 => x"00000000",
    27156 => x"00000000", 27157 => x"00000000", 27158 => x"00000000",
    27159 => x"00000000", 27160 => x"00000000", 27161 => x"00000000",
    27162 => x"00000000", 27163 => x"00000000", 27164 => x"00000000",
    27165 => x"00000000", 27166 => x"00000000", 27167 => x"00000000",
    27168 => x"00000000", 27169 => x"00000000", 27170 => x"00000000",
    27171 => x"00000000", 27172 => x"00000000", 27173 => x"00000000",
    27174 => x"00000000", 27175 => x"00000000", 27176 => x"00000000",
    27177 => x"00000000", 27178 => x"00000000", 27179 => x"00000000",
    27180 => x"00000000", 27181 => x"00000000", 27182 => x"00000000",
    27183 => x"00000000", 27184 => x"00000000", 27185 => x"00000000",
    27186 => x"00000000", 27187 => x"00000000", 27188 => x"00000000",
    27189 => x"00000000", 27190 => x"00000000", 27191 => x"00000000",
    27192 => x"00000000", 27193 => x"00000000", 27194 => x"00000000",
    27195 => x"00000000", 27196 => x"00000000", 27197 => x"00000000",
    27198 => x"00000000", 27199 => x"00000000", 27200 => x"00000000",
    27201 => x"00000000", 27202 => x"00000000", 27203 => x"00000000",
    27204 => x"00000000", 27205 => x"00000000", 27206 => x"00000000",
    27207 => x"00000000", 27208 => x"00000000", 27209 => x"00000000",
    27210 => x"00000000", 27211 => x"00000000", 27212 => x"00000000",
    27213 => x"00000000", 27214 => x"00000000", 27215 => x"00000000",
    27216 => x"00000000", 27217 => x"00000000", 27218 => x"00000000",
    27219 => x"00000000", 27220 => x"00000000", 27221 => x"00000000",
    27222 => x"00000000", 27223 => x"00000000", 27224 => x"00000000",
    27225 => x"00000000", 27226 => x"00000000", 27227 => x"00000000",
    27228 => x"00000000", 27229 => x"00000000", 27230 => x"00000000",
    27231 => x"00000000", 27232 => x"00000000", 27233 => x"00000000",
    27234 => x"00000000", 27235 => x"00000000", 27236 => x"00000000",
    27237 => x"00000000", 27238 => x"00000000", 27239 => x"00000000",
    27240 => x"00000000", 27241 => x"00000000", 27242 => x"00000000",
    27243 => x"00000000", 27244 => x"00000000", 27245 => x"00000000",
    27246 => x"00000000", 27247 => x"00000000", 27248 => x"00000000",
    27249 => x"00000000", 27250 => x"00000000", 27251 => x"00000000",
    27252 => x"00000000", 27253 => x"00000000", 27254 => x"00000000",
    27255 => x"00000000", 27256 => x"00000000", 27257 => x"00000000",
    27258 => x"00000000", 27259 => x"00000000", 27260 => x"00000000",
    27261 => x"00000000", 27262 => x"00000000", 27263 => x"00000000",
    27264 => x"00000000", 27265 => x"00000000", 27266 => x"00000000",
    27267 => x"00000000", 27268 => x"00000000", 27269 => x"00000000",
    27270 => x"00000000", 27271 => x"00000000", 27272 => x"00000000",
    27273 => x"00000000", 27274 => x"00000000", 27275 => x"00000000",
    27276 => x"00000000", 27277 => x"00000000", 27278 => x"00000000",
    27279 => x"00000000", 27280 => x"00000000", 27281 => x"00000000",
    27282 => x"00000000", 27283 => x"00000000", 27284 => x"00000000",
    27285 => x"00000000", 27286 => x"00000000", 27287 => x"00000000",
    27288 => x"00000000", 27289 => x"00000000", 27290 => x"00000000",
    27291 => x"00000000", 27292 => x"00000000", 27293 => x"00000000",
    27294 => x"00000000", 27295 => x"00000000", 27296 => x"00000000",
    27297 => x"00000000", 27298 => x"00000000", 27299 => x"00000000",
    27300 => x"00000000", 27301 => x"00000000", 27302 => x"00000000",
    27303 => x"00000000", 27304 => x"00000000", 27305 => x"00000000",
    27306 => x"00000000", 27307 => x"00000000", 27308 => x"00000000",
    27309 => x"00000000", 27310 => x"00000000", 27311 => x"00000000",
    27312 => x"00000000", 27313 => x"00000000", 27314 => x"00000000",
    27315 => x"00000000", 27316 => x"00000000", 27317 => x"00000000",
    27318 => x"00000000", 27319 => x"00000000", 27320 => x"00000000",
    27321 => x"00000000", 27322 => x"00000000", 27323 => x"00000000",
    27324 => x"00000000", 27325 => x"00000000", 27326 => x"00000000",
    27327 => x"00000000", 27328 => x"00000000", 27329 => x"00000000",
    27330 => x"00000000", 27331 => x"00000000", 27332 => x"00000000",
    27333 => x"00000000", 27334 => x"00000000", 27335 => x"00000000",
    27336 => x"00000000", 27337 => x"00000000", 27338 => x"00000000",
    27339 => x"00000000", 27340 => x"00000000", 27341 => x"00000000",
    27342 => x"00000000", 27343 => x"00000000", 27344 => x"00000000",
    27345 => x"00000000", 27346 => x"00000000", 27347 => x"00000000",
    27348 => x"00000000", 27349 => x"00000000", 27350 => x"00000000",
    27351 => x"00000000", 27352 => x"00000000", 27353 => x"00000000",
    27354 => x"00000000", 27355 => x"00000000", 27356 => x"00000000",
    27357 => x"00000000", 27358 => x"00000000", 27359 => x"00000000",
    27360 => x"00000000", 27361 => x"00000000", 27362 => x"00000000",
    27363 => x"00000000", 27364 => x"00000000", 27365 => x"00000000",
    27366 => x"00000000", 27367 => x"00000000", 27368 => x"00000000",
    27369 => x"00000000", 27370 => x"00000000", 27371 => x"00000000",
    27372 => x"00000000", 27373 => x"00000000", 27374 => x"00000000",
    27375 => x"00000000", 27376 => x"00000000", 27377 => x"00000000",
    27378 => x"00000000", 27379 => x"00000000", 27380 => x"00000000",
    27381 => x"00000000", 27382 => x"00000000", 27383 => x"00000000",
    27384 => x"00000000", 27385 => x"00000000", 27386 => x"00000000",
    27387 => x"00000000", 27388 => x"00000000", 27389 => x"00000000",
    27390 => x"00000000", 27391 => x"00000000", 27392 => x"00000000",
    27393 => x"00000000", 27394 => x"00000000", 27395 => x"00000000",
    27396 => x"00000000", 27397 => x"00000000", 27398 => x"00000000",
    27399 => x"00000000", 27400 => x"00000000", 27401 => x"00000000",
    27402 => x"00000000", 27403 => x"00000000", 27404 => x"00000000",
    27405 => x"00000000", 27406 => x"00000000", 27407 => x"00000000",
    27408 => x"00000000", 27409 => x"00000000", 27410 => x"00000000",
    27411 => x"00000000", 27412 => x"00000000", 27413 => x"00000000",
    27414 => x"00000000", 27415 => x"00000000", 27416 => x"00000000",
    27417 => x"00000000", 27418 => x"00000000", 27419 => x"00000000",
    27420 => x"00000000", 27421 => x"00000000", 27422 => x"00000000",
    27423 => x"00000000", 27424 => x"00000000", 27425 => x"00000000",
    27426 => x"00000000", 27427 => x"00000000", 27428 => x"00000000",
    27429 => x"00000000", 27430 => x"00000000", 27431 => x"00000000",
    27432 => x"00000000", 27433 => x"00000000", 27434 => x"00000000",
    27435 => x"00000000", 27436 => x"00000000", 27437 => x"00000000",
    27438 => x"00000000", 27439 => x"00000000", 27440 => x"00000000",
    27441 => x"00000000", 27442 => x"00000000", 27443 => x"00000000",
    27444 => x"00000000", 27445 => x"00000000", 27446 => x"00000000",
    27447 => x"00000000", 27448 => x"00000000", 27449 => x"00000000",
    27450 => x"00000000", 27451 => x"00000000", 27452 => x"00000000",
    27453 => x"00000000", 27454 => x"00000000", 27455 => x"00000000",
    27456 => x"00000000", 27457 => x"00000000", 27458 => x"00000000",
    27459 => x"00000000", 27460 => x"00000000", 27461 => x"00000000",
    27462 => x"00000000", 27463 => x"00000000", 27464 => x"00000000",
    27465 => x"00000000", 27466 => x"00000000", 27467 => x"00000000",
    27468 => x"00000000", 27469 => x"00000000", 27470 => x"00000000",
    27471 => x"00000000", 27472 => x"00000000", 27473 => x"00000000",
    27474 => x"00000000", 27475 => x"00000000", 27476 => x"00000000",
    27477 => x"00000000", 27478 => x"00000000", 27479 => x"00000000",
    27480 => x"00000000", 27481 => x"00000000", 27482 => x"00000000",
    27483 => x"00000000", 27484 => x"00000000", 27485 => x"00000000",
    27486 => x"00000000", 27487 => x"00000000", 27488 => x"00000000",
    27489 => x"00000000", 27490 => x"00000000", 27491 => x"00000000",
    27492 => x"00000000", 27493 => x"00000000", 27494 => x"00000000",
    27495 => x"00000000", 27496 => x"00000000", 27497 => x"00000000",
    27498 => x"00000000", 27499 => x"00000000", 27500 => x"00000000",
    27501 => x"00000000", 27502 => x"00000000", 27503 => x"00000000",
    27504 => x"00000000", 27505 => x"00000000", 27506 => x"00000000",
    27507 => x"00000000", 27508 => x"00000000", 27509 => x"00000000",
    27510 => x"00000000", 27511 => x"00000000", 27512 => x"00000000",
    27513 => x"00000000", 27514 => x"00000000", 27515 => x"00000000",
    27516 => x"00000000", 27517 => x"00000000", 27518 => x"00000000",
    27519 => x"00000000", 27520 => x"00000000", 27521 => x"00000000",
    27522 => x"00000000", 27523 => x"00000000", 27524 => x"00000000",
    27525 => x"00000000", 27526 => x"00000000", 27527 => x"00000000",
    27528 => x"00000000", 27529 => x"00000000", 27530 => x"00000000",
    27531 => x"00000000", 27532 => x"00000000", 27533 => x"00000000",
    27534 => x"00000000", 27535 => x"00000000", 27536 => x"00000000",
    27537 => x"00000000", 27538 => x"00000000", 27539 => x"00000000",
    27540 => x"00000000", 27541 => x"00000000", 27542 => x"00000000",
    27543 => x"00000000", 27544 => x"00000000", 27545 => x"00000000",
    27546 => x"00000000", 27547 => x"00000000", 27548 => x"00000000",
    27549 => x"00000000", 27550 => x"00000000", 27551 => x"00000000",
    27552 => x"00000000", 27553 => x"00000000", 27554 => x"00000000",
    27555 => x"00000000", 27556 => x"00000000", 27557 => x"00000000",
    27558 => x"00000000", 27559 => x"00000000", 27560 => x"00000000",
    27561 => x"00000000", 27562 => x"00000000", 27563 => x"00000000",
    27564 => x"00000000", 27565 => x"00000000", 27566 => x"00000000",
    27567 => x"00000000", 27568 => x"00000000", 27569 => x"00000000",
    27570 => x"00000000", 27571 => x"00000000", 27572 => x"00000000",
    27573 => x"00000000", 27574 => x"00000000", 27575 => x"00000000",
    27576 => x"00000000", 27577 => x"00000000", 27578 => x"00000000",
    27579 => x"00000000", 27580 => x"00000000", 27581 => x"00000000",
    27582 => x"00000000", 27583 => x"00000000", 27584 => x"00000000",
    27585 => x"00000000", 27586 => x"00000000", 27587 => x"00000000",
    27588 => x"00000000", 27589 => x"00000000", 27590 => x"00000000",
    27591 => x"00000000", 27592 => x"00000000", 27593 => x"00000000",
    27594 => x"00000000", 27595 => x"00000000", 27596 => x"00000000",
    27597 => x"00000000", 27598 => x"00000000", 27599 => x"00000000",
    27600 => x"00000000", 27601 => x"00000000", 27602 => x"00000000",
    27603 => x"00000000", 27604 => x"00000000", 27605 => x"00000000",
    27606 => x"00000000", 27607 => x"00000000", 27608 => x"00000000",
    27609 => x"00000000", 27610 => x"00000000", 27611 => x"00000000",
    27612 => x"00000000", 27613 => x"00000000", 27614 => x"00000000",
    27615 => x"00000000", 27616 => x"00000000", 27617 => x"00000000",
    27618 => x"00000000", 27619 => x"00000000", 27620 => x"00000000",
    27621 => x"00000000", 27622 => x"00000000", 27623 => x"00000000",
    27624 => x"00000000", 27625 => x"00000000", 27626 => x"00000000",
    27627 => x"00000000", 27628 => x"00000000", 27629 => x"00000000",
    27630 => x"00000000", 27631 => x"00000000", 27632 => x"00000000",
    27633 => x"00000000", 27634 => x"00000000", 27635 => x"00000000",
    27636 => x"00000000", 27637 => x"00000000", 27638 => x"00000000",
    27639 => x"00000000", 27640 => x"00000000", 27641 => x"00000000",
    27642 => x"00000000", 27643 => x"00000000", 27644 => x"00000000",
    27645 => x"00000000", 27646 => x"00000000", 27647 => x"00000000",
    27648 => x"00000000", 27649 => x"00000000", 27650 => x"00000000",
    27651 => x"00000000", 27652 => x"00000000", 27653 => x"00000000",
    27654 => x"00000000", 27655 => x"00000000", 27656 => x"00000000",
    27657 => x"00000000", 27658 => x"00000000", 27659 => x"00000000",
    27660 => x"00000000", 27661 => x"00000000", 27662 => x"00000000",
    27663 => x"00000000", 27664 => x"00000000", 27665 => x"00000000",
    27666 => x"00000000", 27667 => x"00000000", 27668 => x"00000000",
    27669 => x"00000000", 27670 => x"00000000", 27671 => x"00000000",
    27672 => x"00000000", 27673 => x"00000000", 27674 => x"00000000",
    27675 => x"00000000", 27676 => x"00000000", 27677 => x"00000000",
    27678 => x"00000000", 27679 => x"00000000", 27680 => x"00000000",
    27681 => x"00000000", 27682 => x"00000000", 27683 => x"00000000",
    27684 => x"00000000", 27685 => x"00000000", 27686 => x"00000000",
    27687 => x"00000000", 27688 => x"00000000", 27689 => x"00000000",
    27690 => x"00000000", 27691 => x"00000000", 27692 => x"00000000",
    27693 => x"00000000", 27694 => x"00000000", 27695 => x"00000000",
    27696 => x"00000000", 27697 => x"00000000", 27698 => x"00000000",
    27699 => x"00000000", 27700 => x"00000000", 27701 => x"00000000",
    27702 => x"00000000", 27703 => x"00000000", 27704 => x"00000000",
    27705 => x"00000000", 27706 => x"00000000", 27707 => x"00000000",
    27708 => x"00000000", 27709 => x"00000000", 27710 => x"00000000",
    27711 => x"00000000", 27712 => x"00000000", 27713 => x"00000000",
    27714 => x"00000000", 27715 => x"00000000", 27716 => x"00000000",
    27717 => x"00000000", 27718 => x"00000000", 27719 => x"00000000",
    27720 => x"00000000", 27721 => x"00000000", 27722 => x"00000000",
    27723 => x"00000000", 27724 => x"00000000", 27725 => x"00000000",
    27726 => x"00000000", 27727 => x"00000000", 27728 => x"00000000",
    27729 => x"00000000", 27730 => x"00000000", 27731 => x"00000000",
    27732 => x"00000000", 27733 => x"00000000", 27734 => x"00000000",
    27735 => x"00000000", 27736 => x"00000000", 27737 => x"00000000",
    27738 => x"00000000", 27739 => x"00000000", 27740 => x"00000000",
    27741 => x"00000000", 27742 => x"00000000", 27743 => x"00000000",
    27744 => x"00000000", 27745 => x"00000000", 27746 => x"00000000",
    27747 => x"00000000", 27748 => x"00000000", 27749 => x"00000000",
    27750 => x"00000000", 27751 => x"00000000", 27752 => x"00000000",
    27753 => x"00000000", 27754 => x"00000000", 27755 => x"00000000",
    27756 => x"00000000", 27757 => x"00000000", 27758 => x"00000000",
    27759 => x"00000000", 27760 => x"00000000", 27761 => x"00000000",
    27762 => x"00000000", 27763 => x"00000000", 27764 => x"00000000",
    27765 => x"00000000", 27766 => x"00000000", 27767 => x"00000000",
    27768 => x"00000000", 27769 => x"00000000", 27770 => x"00000000",
    27771 => x"00000000", 27772 => x"00000000", 27773 => x"00000000",
    27774 => x"00000000", 27775 => x"00000000", 27776 => x"00000000",
    27777 => x"00000000", 27778 => x"00000000", 27779 => x"00000000",
    27780 => x"00000000", 27781 => x"00000000", 27782 => x"00000000",
    27783 => x"00000000", 27784 => x"00000000", 27785 => x"00000000",
    27786 => x"00000000", 27787 => x"00000000", 27788 => x"00000000",
    27789 => x"00000000", 27790 => x"00000000", 27791 => x"00000000",
    27792 => x"00000000", 27793 => x"00000000", 27794 => x"00000000",
    27795 => x"00000000", 27796 => x"00000000", 27797 => x"00000000",
    27798 => x"00000000", 27799 => x"00000000", 27800 => x"00000000",
    27801 => x"00000000", 27802 => x"00000000", 27803 => x"00000000",
    27804 => x"00000000", 27805 => x"00000000", 27806 => x"00000000",
    27807 => x"00000000", 27808 => x"00000000", 27809 => x"00000000",
    27810 => x"00000000", 27811 => x"00000000", 27812 => x"00000000",
    27813 => x"00000000", 27814 => x"00000000", 27815 => x"00000000",
    27816 => x"00000000", 27817 => x"00000000", 27818 => x"00000000",
    27819 => x"00000000", 27820 => x"00000000", 27821 => x"00000000",
    27822 => x"00000000", 27823 => x"00000000", 27824 => x"00000000",
    27825 => x"00000000", 27826 => x"00000000", 27827 => x"00000000",
    27828 => x"00000000", 27829 => x"00000000", 27830 => x"00000000",
    27831 => x"00000000", 27832 => x"00000000", 27833 => x"00000000",
    27834 => x"00000000", 27835 => x"00000000", 27836 => x"00000000",
    27837 => x"00000000", 27838 => x"00000000", 27839 => x"00000000",
    27840 => x"00000000", 27841 => x"00000000", 27842 => x"00000000",
    27843 => x"00000000", 27844 => x"00000000", 27845 => x"00000000",
    27846 => x"00000000", 27847 => x"00000000", 27848 => x"00000000",
    27849 => x"00000000", 27850 => x"00000000", 27851 => x"00000000",
    27852 => x"00000000", 27853 => x"00000000", 27854 => x"00000000",
    27855 => x"00000000", 27856 => x"00000000", 27857 => x"00000000",
    27858 => x"00000000", 27859 => x"00000000", 27860 => x"00000000",
    27861 => x"00000000", 27862 => x"00000000", 27863 => x"00000000",
    27864 => x"00000000", 27865 => x"00000000", 27866 => x"00000000",
    27867 => x"00000000", 27868 => x"00000000", 27869 => x"00000000",
    27870 => x"00000000", 27871 => x"00000000", 27872 => x"00000000",
    27873 => x"00000000", 27874 => x"00000000", 27875 => x"00000000",
    27876 => x"00000000", 27877 => x"00000000", 27878 => x"00000000",
    27879 => x"00000000", 27880 => x"00000000", 27881 => x"00000000",
    27882 => x"00000000", 27883 => x"00000000", 27884 => x"00000000",
    27885 => x"00000000", 27886 => x"00000000", 27887 => x"00000000",
    27888 => x"00000000", 27889 => x"00000000", 27890 => x"00000000",
    27891 => x"00000000", 27892 => x"00000000", 27893 => x"00000000",
    27894 => x"00000000", 27895 => x"00000000", 27896 => x"00000000",
    27897 => x"00000000", 27898 => x"00000000", 27899 => x"00000000",
    27900 => x"00000000", 27901 => x"00000000", 27902 => x"00000000",
    27903 => x"00000000", 27904 => x"00000000", 27905 => x"00000000",
    27906 => x"00000000", 27907 => x"00000000", 27908 => x"00000000",
    27909 => x"00000000", 27910 => x"00000000", 27911 => x"00000000",
    27912 => x"00000000", 27913 => x"00000000", 27914 => x"00000000",
    27915 => x"00000000", 27916 => x"00000000", 27917 => x"00000000",
    27918 => x"00000000", 27919 => x"00000000", 27920 => x"00000000",
    27921 => x"00000000", 27922 => x"00000000", 27923 => x"00000000",
    27924 => x"00000000", 27925 => x"00000000", 27926 => x"00000000",
    27927 => x"00000000", 27928 => x"00000000", 27929 => x"00000000",
    27930 => x"00000000", 27931 => x"00000000", 27932 => x"00000000",
    27933 => x"00000000", 27934 => x"00000000", 27935 => x"00000000",
    27936 => x"00000000", 27937 => x"00000000", 27938 => x"00000000",
    27939 => x"00000000", 27940 => x"00000000", 27941 => x"00000000",
    27942 => x"00000000", 27943 => x"00000000", 27944 => x"00000000",
    27945 => x"00000000", 27946 => x"00000000", 27947 => x"00000000",
    27948 => x"00000000", 27949 => x"00000000", 27950 => x"00000000",
    27951 => x"00000000", 27952 => x"00000000", 27953 => x"00000000",
    27954 => x"00000000", 27955 => x"00000000", 27956 => x"00000000",
    27957 => x"00000000", 27958 => x"00000000", 27959 => x"00000000",
    27960 => x"00000000", 27961 => x"00000000", 27962 => x"00000000",
    27963 => x"00000000", 27964 => x"00000000", 27965 => x"00000000",
    27966 => x"00000000", 27967 => x"00000000", 27968 => x"00000000",
    27969 => x"00000000", 27970 => x"00000000", 27971 => x"00000000",
    27972 => x"00000000", 27973 => x"00000000", 27974 => x"00000000",
    27975 => x"00000000", 27976 => x"00000000", 27977 => x"00000000",
    27978 => x"00000000", 27979 => x"00000000", 27980 => x"00000000",
    27981 => x"00000000", 27982 => x"00000000", 27983 => x"00000000",
    27984 => x"00000000", 27985 => x"00000000", 27986 => x"00000000",
    27987 => x"00000000", 27988 => x"00000000", 27989 => x"00000000",
    27990 => x"00000000", 27991 => x"00000000", 27992 => x"00000000",
    27993 => x"00000000", 27994 => x"00000000", 27995 => x"00000000",
    27996 => x"00000000", 27997 => x"00000000", 27998 => x"00000000",
    27999 => x"00000000", 28000 => x"00000000", 28001 => x"00000000",
    28002 => x"00000000", 28003 => x"00000000", 28004 => x"00000000",
    28005 => x"00000000", 28006 => x"00000000", 28007 => x"00000000",
    28008 => x"00000000", 28009 => x"00000000", 28010 => x"00000000",
    28011 => x"00000000", 28012 => x"00000000", 28013 => x"00000000",
    28014 => x"00000000", 28015 => x"00000000", 28016 => x"00000000",
    28017 => x"00000000", 28018 => x"00000000", 28019 => x"00000000",
    28020 => x"00000000", 28021 => x"00000000", 28022 => x"00000000",
    28023 => x"00000000", 28024 => x"00000000", 28025 => x"00000000",
    28026 => x"00000000", 28027 => x"00000000", 28028 => x"00000000",
    28029 => x"00000000", 28030 => x"00000000", 28031 => x"00000000",
    28032 => x"00000000", 28033 => x"00000000", 28034 => x"00000000",
    28035 => x"00000000", 28036 => x"00000000", 28037 => x"00000000",
    28038 => x"00000000", 28039 => x"00000000", 28040 => x"00000000",
    28041 => x"00000000", 28042 => x"00000000", 28043 => x"00000000",
    28044 => x"00000000", 28045 => x"00000000", 28046 => x"00000000",
    28047 => x"00000000", 28048 => x"00000000", 28049 => x"00000000",
    28050 => x"00000000", 28051 => x"00000000", 28052 => x"00000000",
    28053 => x"00000000", 28054 => x"00000000", 28055 => x"00000000",
    28056 => x"00000000", 28057 => x"00000000", 28058 => x"00000000",
    28059 => x"00000000", 28060 => x"00000000", 28061 => x"00000000",
    28062 => x"00000000", 28063 => x"00000000", 28064 => x"00000000",
    28065 => x"00000000", 28066 => x"00000000", 28067 => x"00000000",
    28068 => x"00000000", 28069 => x"00000000", 28070 => x"00000000",
    28071 => x"00000000", 28072 => x"00000000", 28073 => x"00000000",
    28074 => x"00000000", 28075 => x"00000000", 28076 => x"00000000",
    28077 => x"00000000", 28078 => x"00000000", 28079 => x"00000000",
    28080 => x"00000000", 28081 => x"00000000", 28082 => x"00000000",
    28083 => x"00000000", 28084 => x"00000000", 28085 => x"00000000",
    28086 => x"00000000", 28087 => x"00000000", 28088 => x"00000000",
    28089 => x"00000000", 28090 => x"00000000", 28091 => x"00000000",
    28092 => x"00000000", 28093 => x"00000000", 28094 => x"00000000",
    28095 => x"00000000", 28096 => x"00000000", 28097 => x"00000000",
    28098 => x"00000000", 28099 => x"00000000", 28100 => x"00000000",
    28101 => x"00000000", 28102 => x"00000000", 28103 => x"00000000",
    28104 => x"00000000", 28105 => x"00000000", 28106 => x"00000000",
    28107 => x"00000000", 28108 => x"00000000", 28109 => x"00000000",
    28110 => x"00000000", 28111 => x"00000000", 28112 => x"00000000",
    28113 => x"00000000", 28114 => x"00000000", 28115 => x"00000000",
    28116 => x"00000000", 28117 => x"00000000", 28118 => x"00000000",
    28119 => x"00000000", 28120 => x"00000000", 28121 => x"00000000",
    28122 => x"00000000", 28123 => x"00000000", 28124 => x"00000000",
    28125 => x"00000000", 28126 => x"00000000", 28127 => x"00000000",
    28128 => x"00000000", 28129 => x"00000000", 28130 => x"00000000",
    28131 => x"00000000", 28132 => x"00000000", 28133 => x"00000000",
    28134 => x"00000000", 28135 => x"00000000", 28136 => x"00000000",
    28137 => x"00000000", 28138 => x"00000000", 28139 => x"00000000",
    28140 => x"00000000", 28141 => x"00000000", 28142 => x"00000000",
    28143 => x"00000000", 28144 => x"00000000", 28145 => x"00000000",
    28146 => x"00000000", 28147 => x"00000000", 28148 => x"00000000",
    28149 => x"00000000", 28150 => x"00000000", 28151 => x"00000000",
    28152 => x"00000000", 28153 => x"00000000", 28154 => x"00000000",
    28155 => x"00000000", 28156 => x"00000000", 28157 => x"00000000",
    28158 => x"00000000", 28159 => x"00000000", 28160 => x"00000000",
    28161 => x"00000000", 28162 => x"00000000", 28163 => x"00000000",
    28164 => x"00000000", 28165 => x"00000000", 28166 => x"00000000",
    28167 => x"00000000", 28168 => x"00000000", 28169 => x"00000000",
    28170 => x"00000000", 28171 => x"00000000", 28172 => x"00000000",
    28173 => x"00000000", 28174 => x"00000000", 28175 => x"00000000",
    28176 => x"00000000", 28177 => x"00000000", 28178 => x"00000000",
    28179 => x"00000000", 28180 => x"00000000", 28181 => x"00000000",
    28182 => x"00000000", 28183 => x"00000000", 28184 => x"00000000",
    28185 => x"00000000", 28186 => x"00000000", 28187 => x"00000000",
    28188 => x"00000000", 28189 => x"00000000", 28190 => x"00000000",
    28191 => x"00000000", 28192 => x"00000000", 28193 => x"00000000",
    28194 => x"00000000", 28195 => x"00000000", 28196 => x"00000000",
    28197 => x"00000000", 28198 => x"00000000", 28199 => x"00000000",
    28200 => x"00000000", 28201 => x"00000000", 28202 => x"00000000",
    28203 => x"00000000", 28204 => x"00000000", 28205 => x"00000000",
    28206 => x"00000000", 28207 => x"00000000", 28208 => x"00000000",
    28209 => x"00000000", 28210 => x"00000000", 28211 => x"00000000",
    28212 => x"00000000", 28213 => x"00000000", 28214 => x"00000000",
    28215 => x"00000000", 28216 => x"00000000", 28217 => x"00000000",
    28218 => x"00000000", 28219 => x"00000000", 28220 => x"00000000",
    28221 => x"00000000", 28222 => x"00000000", 28223 => x"00000000",
    28224 => x"00000000", 28225 => x"00000000", 28226 => x"00000000",
    28227 => x"00000000", 28228 => x"00000000", 28229 => x"00000000",
    28230 => x"00000000", 28231 => x"00000000", 28232 => x"00000000",
    28233 => x"00000000", 28234 => x"00000000", 28235 => x"00000000",
    28236 => x"00000000", 28237 => x"00000000", 28238 => x"00000000",
    28239 => x"00000000", 28240 => x"00000000", 28241 => x"00000000",
    28242 => x"00000000", 28243 => x"00000000", 28244 => x"00000000",
    28245 => x"00000000", 28246 => x"00000000", 28247 => x"00000000",
    28248 => x"00000000", 28249 => x"00000000", 28250 => x"00000000",
    28251 => x"00000000", 28252 => x"00000000", 28253 => x"00000000",
    28254 => x"00000000", 28255 => x"00000000", 28256 => x"00000000",
    28257 => x"00000000", 28258 => x"00000000", 28259 => x"00000000",
    28260 => x"00000000", 28261 => x"00000000", 28262 => x"00000000",
    28263 => x"00000000", 28264 => x"00000000", 28265 => x"00000000",
    28266 => x"00000000", 28267 => x"00000000", 28268 => x"00000000",
    28269 => x"00000000", 28270 => x"00000000", 28271 => x"00000000",
    28272 => x"00000000", 28273 => x"00000000", 28274 => x"00000000",
    28275 => x"00000000", 28276 => x"00000000", 28277 => x"00000000",
    28278 => x"00000000", 28279 => x"00000000", 28280 => x"00000000",
    28281 => x"00000000", 28282 => x"00000000", 28283 => x"00000000",
    28284 => x"00000000", 28285 => x"00000000", 28286 => x"00000000",
    28287 => x"00000000", 28288 => x"00000000", 28289 => x"00000000",
    28290 => x"00000000", 28291 => x"00000000", 28292 => x"00000000",
    28293 => x"00000000", 28294 => x"00000000", 28295 => x"00000000",
    28296 => x"00000000", 28297 => x"00000000", 28298 => x"00000000",
    28299 => x"00000000", 28300 => x"00000000", 28301 => x"00000000",
    28302 => x"00000000", 28303 => x"00000000", 28304 => x"00000000",
    28305 => x"00000000", 28306 => x"00000000", 28307 => x"00000000",
    28308 => x"00000000", 28309 => x"00000000", 28310 => x"00000000",
    28311 => x"00000000", 28312 => x"00000000", 28313 => x"00000000",
    28314 => x"00000000", 28315 => x"00000000", 28316 => x"00000000",
    28317 => x"00000000", 28318 => x"00000000", 28319 => x"00000000",
    28320 => x"00000000", 28321 => x"00000000", 28322 => x"00000000",
    28323 => x"00000000", 28324 => x"00000000", 28325 => x"00000000",
    28326 => x"00000000", 28327 => x"00000000", 28328 => x"00000000",
    28329 => x"00000000", 28330 => x"00000000", 28331 => x"00000000",
    28332 => x"00000000", 28333 => x"00000000", 28334 => x"00000000",
    28335 => x"00000000", 28336 => x"00000000", 28337 => x"00000000",
    28338 => x"00000000", 28339 => x"00000000", 28340 => x"00000000",
    28341 => x"00000000", 28342 => x"00000000", 28343 => x"00000000",
    28344 => x"00000000", 28345 => x"00000000", 28346 => x"00000000",
    28347 => x"00000000", 28348 => x"00000000", 28349 => x"00000000",
    28350 => x"00000000", 28351 => x"00000000", 28352 => x"00000000",
    28353 => x"00000000", 28354 => x"00000000", 28355 => x"00000000",
    28356 => x"00000000", 28357 => x"00000000", 28358 => x"00000000",
    28359 => x"00000000", 28360 => x"00000000", 28361 => x"00000000",
    28362 => x"00000000", 28363 => x"00000000", 28364 => x"00000000",
    28365 => x"00000000", 28366 => x"00000000", 28367 => x"00000000",
    28368 => x"00000000", 28369 => x"00000000", 28370 => x"00000000",
    28371 => x"00000000", 28372 => x"00000000", 28373 => x"00000000",
    28374 => x"00000000", 28375 => x"00000000", 28376 => x"00000000",
    28377 => x"00000000", 28378 => x"00000000", 28379 => x"00000000",
    28380 => x"00000000", 28381 => x"00000000", 28382 => x"00000000",
    28383 => x"00000000", 28384 => x"00000000", 28385 => x"00000000",
    28386 => x"00000000", 28387 => x"00000000", 28388 => x"00000000",
    28389 => x"00000000", 28390 => x"00000000", 28391 => x"00000000",
    28392 => x"00000000", 28393 => x"00000000", 28394 => x"00000000",
    28395 => x"00000000", 28396 => x"00000000", 28397 => x"00000000",
    28398 => x"00000000", 28399 => x"00000000", 28400 => x"00000000",
    28401 => x"00000000", 28402 => x"00000000", 28403 => x"00000000",
    28404 => x"00000000", 28405 => x"00000000", 28406 => x"00000000",
    28407 => x"00000000", 28408 => x"00000000", 28409 => x"00000000",
    28410 => x"00000000", 28411 => x"00000000", 28412 => x"00000000",
    28413 => x"00000000", 28414 => x"00000000", 28415 => x"00000000",
    28416 => x"00000000", 28417 => x"00000000", 28418 => x"00000000",
    28419 => x"00000000", 28420 => x"00000000", 28421 => x"00000000",
    28422 => x"00000000", 28423 => x"00000000", 28424 => x"00000000",
    28425 => x"00000000", 28426 => x"00000000", 28427 => x"00000000",
    28428 => x"00000000", 28429 => x"00000000", 28430 => x"00000000",
    28431 => x"00000000", 28432 => x"00000000", 28433 => x"00000000",
    28434 => x"00000000", 28435 => x"00000000", 28436 => x"00000000",
    28437 => x"00000000", 28438 => x"00000000", 28439 => x"00000000",
    28440 => x"00000000", 28441 => x"00000000", 28442 => x"00000000",
    28443 => x"00000000", 28444 => x"00000000", 28445 => x"00000000",
    28446 => x"00000000", 28447 => x"00000000", 28448 => x"00000000",
    28449 => x"00000000", 28450 => x"00000000", 28451 => x"00000000",
    28452 => x"00000000", 28453 => x"00000000", 28454 => x"00000000",
    28455 => x"00000000", 28456 => x"00000000", 28457 => x"00000000",
    28458 => x"00000000", 28459 => x"00000000", 28460 => x"00000000",
    28461 => x"00000000", 28462 => x"00000000", 28463 => x"00000000",
    28464 => x"00000000", 28465 => x"00000000", 28466 => x"00000000",
    28467 => x"00000000", 28468 => x"00000000", 28469 => x"00000000",
    28470 => x"00000000", 28471 => x"00000000", 28472 => x"00000000",
    28473 => x"00000000", 28474 => x"00000000", 28475 => x"00000000",
    28476 => x"00000000", 28477 => x"00000000", 28478 => x"00000000",
    28479 => x"00000000", 28480 => x"00000000", 28481 => x"00000000",
    28482 => x"00000000", 28483 => x"00000000", 28484 => x"00000000",
    28485 => x"00000000", 28486 => x"00000000", 28487 => x"00000000",
    28488 => x"00000000", 28489 => x"00000000", 28490 => x"00000000",
    28491 => x"00000000", 28492 => x"00000000", 28493 => x"00000000",
    28494 => x"00000000", 28495 => x"00000000", 28496 => x"00000000",
    28497 => x"00000000", 28498 => x"00000000", 28499 => x"00000000",
    28500 => x"00000000", 28501 => x"00000000", 28502 => x"00000000",
    28503 => x"00000000", 28504 => x"00000000", 28505 => x"00000000",
    28506 => x"00000000", 28507 => x"00000000", 28508 => x"00000000",
    28509 => x"00000000", 28510 => x"00000000", 28511 => x"00000000",
    28512 => x"00000000", 28513 => x"00000000", 28514 => x"00000000",
    28515 => x"00000000", 28516 => x"00000000", 28517 => x"00000000",
    28518 => x"00000000", 28519 => x"00000000", 28520 => x"00000000",
    28521 => x"00000000", 28522 => x"00000000", 28523 => x"00000000",
    28524 => x"00000000", 28525 => x"00000000", 28526 => x"00000000",
    28527 => x"00000000", 28528 => x"00000000", 28529 => x"00000000",
    28530 => x"00000000", 28531 => x"00000000", 28532 => x"00000000",
    28533 => x"00000000", 28534 => x"00000000", 28535 => x"00000000",
    28536 => x"00000000", 28537 => x"00000000", 28538 => x"00000000",
    28539 => x"00000000", 28540 => x"00000000", 28541 => x"00000000",
    28542 => x"00000000", 28543 => x"00000000", 28544 => x"00000000",
    28545 => x"00000000", 28546 => x"00000000", 28547 => x"00000000",
    28548 => x"00000000", 28549 => x"00000000", 28550 => x"00000000",
    28551 => x"00000000", 28552 => x"00000000", 28553 => x"00000000",
    28554 => x"00000000", 28555 => x"00000000", 28556 => x"00000000",
    28557 => x"00000000", 28558 => x"00000000", 28559 => x"00000000",
    28560 => x"00000000", 28561 => x"00000000", 28562 => x"00000000",
    28563 => x"00000000", 28564 => x"00000000", 28565 => x"00000000",
    28566 => x"00000000", 28567 => x"00000000", 28568 => x"00000000",
    28569 => x"00000000", 28570 => x"00000000", 28571 => x"00000000",
    28572 => x"00000000", 28573 => x"00000000", 28574 => x"00000000",
    28575 => x"00000000", 28576 => x"00000000", 28577 => x"00000000",
    28578 => x"00000000", 28579 => x"00000000", 28580 => x"00000000",
    28581 => x"00000000", 28582 => x"00000000", 28583 => x"00000000",
    28584 => x"00000000", 28585 => x"00000000", 28586 => x"00000000",
    28587 => x"00000000", 28588 => x"00000000", 28589 => x"00000000",
    28590 => x"00000000", 28591 => x"00000000", 28592 => x"00000000",
    28593 => x"00000000", 28594 => x"00000000", 28595 => x"00000000",
    28596 => x"00000000", 28597 => x"00000000", 28598 => x"00000000",
    28599 => x"00000000", 28600 => x"00000000", 28601 => x"00000000",
    28602 => x"00000000", 28603 => x"00000000", 28604 => x"00000000",
    28605 => x"00000000", 28606 => x"00000000", 28607 => x"00000000",
    28608 => x"00000000", 28609 => x"00000000", 28610 => x"00000000",
    28611 => x"00000000", 28612 => x"00000000", 28613 => x"00000000",
    28614 => x"00000000", 28615 => x"00000000", 28616 => x"00000000",
    28617 => x"00000000", 28618 => x"00000000", 28619 => x"00000000",
    28620 => x"00000000", 28621 => x"00000000", 28622 => x"00000000",
    28623 => x"00000000", 28624 => x"00000000", 28625 => x"00000000",
    28626 => x"00000000", 28627 => x"00000000", 28628 => x"00000000",
    28629 => x"00000000", 28630 => x"00000000", 28631 => x"00000000",
    28632 => x"00000000", 28633 => x"00000000", 28634 => x"00000000",
    28635 => x"00000000", 28636 => x"00000000", 28637 => x"00000000",
    28638 => x"00000000", 28639 => x"00000000", 28640 => x"00000000",
    28641 => x"00000000", 28642 => x"00000000", 28643 => x"00000000",
    28644 => x"00000000", 28645 => x"00000000", 28646 => x"00000000",
    28647 => x"00000000", 28648 => x"00000000", 28649 => x"00000000",
    28650 => x"00000000", 28651 => x"00000000", 28652 => x"00000000",
    28653 => x"00000000", 28654 => x"00000000", 28655 => x"00000000",
    28656 => x"00000000", 28657 => x"00000000", 28658 => x"00000000",
    28659 => x"00000000", 28660 => x"00000000", 28661 => x"00000000",
    28662 => x"00000000", 28663 => x"00000000", 28664 => x"00000000",
    28665 => x"00000000", 28666 => x"00000000", 28667 => x"00000000",
    28668 => x"00000000", 28669 => x"00000000", 28670 => x"00000000",
    28671 => x"00000000", 28672 => x"00000000", 28673 => x"00000000",
    28674 => x"00000000", 28675 => x"00000000", 28676 => x"00000000",
    28677 => x"00000000", 28678 => x"00000000", 28679 => x"00000000",
    28680 => x"00000000", 28681 => x"00000000", 28682 => x"00000000",
    28683 => x"00000000", 28684 => x"00000000", 28685 => x"00000000",
    28686 => x"00000000", 28687 => x"00000000", 28688 => x"00000000",
    28689 => x"00000000", 28690 => x"00000000", 28691 => x"00000000",
    28692 => x"00000000", 28693 => x"00000000", 28694 => x"00000000",
    28695 => x"00000000", 28696 => x"00000000", 28697 => x"00000000",
    28698 => x"00000000", 28699 => x"00000000", 28700 => x"00000000",
    28701 => x"00000000", 28702 => x"00000000", 28703 => x"00000000",
    28704 => x"00000000", 28705 => x"00000000", 28706 => x"00000000",
    28707 => x"00000000", 28708 => x"00000000", 28709 => x"00000000",
    28710 => x"00000000", 28711 => x"00000000", 28712 => x"00000000",
    28713 => x"00000000", 28714 => x"00000000", 28715 => x"00000000",
    28716 => x"00000000", 28717 => x"00000000", 28718 => x"00000000",
    28719 => x"00000000", 28720 => x"00000000", 28721 => x"00000000",
    28722 => x"00000000", 28723 => x"00000000", 28724 => x"00000000",
    28725 => x"00000000", 28726 => x"00000000", 28727 => x"00000000",
    28728 => x"00000000", 28729 => x"00000000", 28730 => x"00000000",
    28731 => x"00000000", 28732 => x"00000000", 28733 => x"00000000",
    28734 => x"00000000", 28735 => x"00000000", 28736 => x"00000000",
    28737 => x"00000000", 28738 => x"00000000", 28739 => x"00000000",
    28740 => x"00000000", 28741 => x"00000000", 28742 => x"00000000",
    28743 => x"00000000", 28744 => x"00000000", 28745 => x"00000000",
    28746 => x"00000000", 28747 => x"00000000", 28748 => x"00000000",
    28749 => x"00000000", 28750 => x"00000000", 28751 => x"00000000",
    28752 => x"00000000", 28753 => x"00000000", 28754 => x"00000000",
    28755 => x"00000000", 28756 => x"00000000", 28757 => x"00000000",
    28758 => x"00000000", 28759 => x"00000000", 28760 => x"00000000",
    28761 => x"00000000", 28762 => x"00000000", 28763 => x"00000000",
    28764 => x"00000000", 28765 => x"00000000", 28766 => x"00000000",
    28767 => x"00000000", 28768 => x"00000000", 28769 => x"00000000",
    28770 => x"00000000", 28771 => x"00000000", 28772 => x"00000000",
    28773 => x"00000000", 28774 => x"00000000", 28775 => x"00000000",
    28776 => x"00000000", 28777 => x"00000000", 28778 => x"00000000",
    28779 => x"00000000", 28780 => x"00000000", 28781 => x"00000000",
    28782 => x"00000000", 28783 => x"00000000", 28784 => x"00000000",
    28785 => x"00000000", 28786 => x"00000000", 28787 => x"00000000",
    28788 => x"00000000", 28789 => x"00000000", 28790 => x"00000000",
    28791 => x"00000000", 28792 => x"00000000", 28793 => x"00000000",
    28794 => x"00000000", 28795 => x"00000000", 28796 => x"00000000",
    28797 => x"00000000", 28798 => x"00000000", 28799 => x"00000000",
    28800 => x"00000000", 28801 => x"00000000", 28802 => x"00000000",
    28803 => x"00000000", 28804 => x"00000000", 28805 => x"00000000",
    28806 => x"00000000", 28807 => x"00000000", 28808 => x"00000000",
    28809 => x"00000000", 28810 => x"00000000", 28811 => x"00000000",
    28812 => x"00000000", 28813 => x"00000000", 28814 => x"00000000",
    28815 => x"00000000", 28816 => x"00000000", 28817 => x"00000000",
    28818 => x"00000000", 28819 => x"00000000", 28820 => x"00000000",
    28821 => x"00000000", 28822 => x"00000000", 28823 => x"00000000",
    28824 => x"00000000", 28825 => x"00000000", 28826 => x"00000000",
    28827 => x"00000000", 28828 => x"00000000", 28829 => x"00000000",
    28830 => x"00000000", 28831 => x"00000000", 28832 => x"00000000",
    28833 => x"00000000", 28834 => x"00000000", 28835 => x"00000000",
    28836 => x"00000000", 28837 => x"00000000", 28838 => x"00000000",
    28839 => x"00000000", 28840 => x"00000000", 28841 => x"00000000",
    28842 => x"00000000", 28843 => x"00000000", 28844 => x"00000000",
    28845 => x"00000000", 28846 => x"00000000", 28847 => x"00000000",
    28848 => x"00000000", 28849 => x"00000000", 28850 => x"00000000",
    28851 => x"00000000", 28852 => x"00000000", 28853 => x"00000000",
    28854 => x"00000000", 28855 => x"00000000", 28856 => x"00000000",
    28857 => x"00000000", 28858 => x"00000000", 28859 => x"00000000",
    28860 => x"00000000", 28861 => x"00000000", 28862 => x"00000000",
    28863 => x"00000000", 28864 => x"00000000", 28865 => x"00000000",
    28866 => x"00000000", 28867 => x"00000000", 28868 => x"00000000",
    28869 => x"00000000", 28870 => x"00000000", 28871 => x"00000000",
    28872 => x"00000000", 28873 => x"00000000", 28874 => x"00000000",
    28875 => x"00000000", 28876 => x"00000000", 28877 => x"00000000",
    28878 => x"00000000", 28879 => x"00000000", 28880 => x"00000000",
    28881 => x"00000000", 28882 => x"00000000", 28883 => x"00000000",
    28884 => x"00000000", 28885 => x"00000000", 28886 => x"00000000",
    28887 => x"00000000", 28888 => x"00000000", 28889 => x"00000000",
    28890 => x"00000000", 28891 => x"00000000", 28892 => x"00000000",
    28893 => x"00000000", 28894 => x"00000000", 28895 => x"00000000",
    28896 => x"00000000", 28897 => x"00000000", 28898 => x"00000000",
    28899 => x"00000000", 28900 => x"00000000", 28901 => x"00000000",
    28902 => x"00000000", 28903 => x"00000000", 28904 => x"00000000",
    28905 => x"00000000", 28906 => x"00000000", 28907 => x"00000000",
    28908 => x"00000000", 28909 => x"00000000", 28910 => x"00000000",
    28911 => x"00000000", 28912 => x"00000000", 28913 => x"00000000",
    28914 => x"00000000", 28915 => x"00000000", 28916 => x"00000000",
    28917 => x"00000000", 28918 => x"00000000", 28919 => x"00000000",
    28920 => x"00000000", 28921 => x"00000000", 28922 => x"00000000",
    28923 => x"00000000", 28924 => x"00000000", 28925 => x"00000000",
    28926 => x"00000000", 28927 => x"00000000", 28928 => x"00000000",
    28929 => x"00000000", 28930 => x"00000000", 28931 => x"00000000",
    28932 => x"00000000", 28933 => x"00000000", 28934 => x"00000000",
    28935 => x"00000000", 28936 => x"00000000", 28937 => x"00000000",
    28938 => x"00000000", 28939 => x"00000000", 28940 => x"00000000",
    28941 => x"00000000", 28942 => x"00000000", 28943 => x"00000000",
    28944 => x"00000000", 28945 => x"00000000", 28946 => x"00000000",
    28947 => x"00000000", 28948 => x"00000000", 28949 => x"00000000",
    28950 => x"00000000", 28951 => x"00000000", 28952 => x"00000000",
    28953 => x"00000000", 28954 => x"00000000", 28955 => x"00000000",
    28956 => x"00000000", 28957 => x"00000000", 28958 => x"00000000",
    28959 => x"00000000", 28960 => x"00000000", 28961 => x"00000000",
    28962 => x"00000000", 28963 => x"00000000", 28964 => x"00000000",
    28965 => x"00000000", 28966 => x"00000000", 28967 => x"00000000",
    28968 => x"00000000", 28969 => x"00000000", 28970 => x"00000000",
    28971 => x"00000000", 28972 => x"00000000", 28973 => x"00000000",
    28974 => x"00000000", 28975 => x"00000000", 28976 => x"00000000",
    28977 => x"00000000", 28978 => x"00000000", 28979 => x"00000000",
    28980 => x"00000000", 28981 => x"00000000", 28982 => x"00000000",
    28983 => x"00000000", 28984 => x"00000000", 28985 => x"00000000",
    28986 => x"00000000", 28987 => x"00000000", 28988 => x"00000000",
    28989 => x"00000000", 28990 => x"00000000", 28991 => x"00000000",
    28992 => x"00000000", 28993 => x"00000000", 28994 => x"00000000",
    28995 => x"00000000", 28996 => x"00000000", 28997 => x"00000000",
    28998 => x"00000000", 28999 => x"00000000", 29000 => x"00000000",
    29001 => x"00000000", 29002 => x"00000000", 29003 => x"00000000",
    29004 => x"00000000", 29005 => x"00000000", 29006 => x"00000000",
    29007 => x"00000000", 29008 => x"00000000", 29009 => x"00000000",
    29010 => x"00000000", 29011 => x"00000000", 29012 => x"00000000",
    29013 => x"00000000", 29014 => x"00000000", 29015 => x"00000000",
    29016 => x"00000000", 29017 => x"00000000", 29018 => x"00000000",
    29019 => x"00000000", 29020 => x"00000000", 29021 => x"00000000",
    29022 => x"00000000", 29023 => x"00000000", 29024 => x"00000000",
    29025 => x"00000000", 29026 => x"00000000", 29027 => x"00000000",
    29028 => x"00000000", 29029 => x"00000000", 29030 => x"00000000",
    29031 => x"00000000", 29032 => x"00000000", 29033 => x"00000000",
    29034 => x"00000000", 29035 => x"00000000", 29036 => x"00000000",
    29037 => x"00000000", 29038 => x"00000000", 29039 => x"00000000",
    29040 => x"00000000", 29041 => x"00000000", 29042 => x"00000000",
    29043 => x"00000000", 29044 => x"00000000", 29045 => x"00000000",
    29046 => x"00000000", 29047 => x"00000000", 29048 => x"00000000",
    29049 => x"00000000", 29050 => x"00000000", 29051 => x"00000000",
    29052 => x"00000000", 29053 => x"00000000", 29054 => x"00000000",
    29055 => x"00000000", 29056 => x"00000000", 29057 => x"00000000",
    29058 => x"00000000", 29059 => x"00000000", 29060 => x"00000000",
    29061 => x"00000000", 29062 => x"00000000", 29063 => x"00000000",
    29064 => x"00000000", 29065 => x"00000000", 29066 => x"00000000",
    29067 => x"00000000", 29068 => x"00000000", 29069 => x"00000000",
    29070 => x"00000000", 29071 => x"00000000", 29072 => x"00000000",
    29073 => x"00000000", 29074 => x"00000000", 29075 => x"00000000",
    29076 => x"00000000", 29077 => x"00000000", 29078 => x"00000000",
    29079 => x"00000000", 29080 => x"00000000", 29081 => x"00000000",
    29082 => x"00000000", 29083 => x"00000000", 29084 => x"00000000",
    29085 => x"00000000", 29086 => x"00000000", 29087 => x"00000000",
    29088 => x"00000000", 29089 => x"00000000", 29090 => x"00000000",
    29091 => x"00000000", 29092 => x"00000000", 29093 => x"00000000",
    29094 => x"00000000", 29095 => x"00000000", 29096 => x"00000000",
    29097 => x"00000000", 29098 => x"00000000", 29099 => x"00000000",
    29100 => x"00000000", 29101 => x"00000000", 29102 => x"00000000",
    29103 => x"00000000", 29104 => x"00000000", 29105 => x"00000000",
    29106 => x"00000000", 29107 => x"00000000", 29108 => x"00000000",
    29109 => x"00000000", 29110 => x"00000000", 29111 => x"00000000",
    29112 => x"00000000", 29113 => x"00000000", 29114 => x"00000000",
    29115 => x"00000000", 29116 => x"00000000", 29117 => x"00000000",
    29118 => x"00000000", 29119 => x"00000000", 29120 => x"00000000",
    29121 => x"00000000", 29122 => x"00000000", 29123 => x"00000000",
    29124 => x"00000000", 29125 => x"00000000", 29126 => x"00000000",
    29127 => x"00000000", 29128 => x"00000000", 29129 => x"00000000",
    29130 => x"00000000", 29131 => x"00000000", 29132 => x"00000000",
    29133 => x"00000000", 29134 => x"00000000", 29135 => x"00000000",
    29136 => x"00000000", 29137 => x"00000000", 29138 => x"00000000",
    29139 => x"00000000", 29140 => x"00000000", 29141 => x"00000000",
    29142 => x"00000000", 29143 => x"00000000", 29144 => x"00000000",
    29145 => x"00000000", 29146 => x"00000000", 29147 => x"00000000",
    29148 => x"00000000", 29149 => x"00000000", 29150 => x"00000000",
    29151 => x"00000000", 29152 => x"00000000", 29153 => x"00000000",
    29154 => x"00000000", 29155 => x"00000000", 29156 => x"00000000",
    29157 => x"00000000", 29158 => x"00000000", 29159 => x"00000000",
    29160 => x"00000000", 29161 => x"00000000", 29162 => x"00000000",
    29163 => x"00000000", 29164 => x"00000000", 29165 => x"00000000",
    29166 => x"00000000", 29167 => x"00000000", 29168 => x"00000000",
    29169 => x"00000000", 29170 => x"00000000", 29171 => x"00000000",
    29172 => x"00000000", 29173 => x"00000000", 29174 => x"00000000",
    29175 => x"00000000", 29176 => x"00000000", 29177 => x"00000000",
    29178 => x"00000000", 29179 => x"00000000", 29180 => x"00000000",
    29181 => x"00000000", 29182 => x"00000000", 29183 => x"00000000",
    29184 => x"00000000", 29185 => x"00000000", 29186 => x"00000000",
    29187 => x"00000000", 29188 => x"00000000", 29189 => x"00000000",
    29190 => x"00000000", 29191 => x"00000000", 29192 => x"00000000",
    29193 => x"00000000", 29194 => x"00000000", 29195 => x"00000000",
    29196 => x"00000000", 29197 => x"00000000", 29198 => x"00000000",
    29199 => x"00000000", 29200 => x"00000000", 29201 => x"00000000",
    29202 => x"00000000", 29203 => x"00000000", 29204 => x"00000000",
    29205 => x"00000000", 29206 => x"00000000", 29207 => x"00000000",
    29208 => x"00000000", 29209 => x"00000000", 29210 => x"00000000",
    29211 => x"00000000", 29212 => x"00000000", 29213 => x"00000000",
    29214 => x"00000000", 29215 => x"00000000", 29216 => x"00000000",
    29217 => x"00000000", 29218 => x"00000000", 29219 => x"00000000",
    29220 => x"00000000", 29221 => x"00000000", 29222 => x"00000000",
    29223 => x"00000000", 29224 => x"00000000", 29225 => x"00000000",
    29226 => x"00000000", 29227 => x"00000000", 29228 => x"00000000",
    29229 => x"00000000", 29230 => x"00000000", 29231 => x"00000000",
    29232 => x"00000000", 29233 => x"00000000", 29234 => x"00000000",
    29235 => x"00000000", 29236 => x"00000000", 29237 => x"00000000",
    29238 => x"00000000", 29239 => x"00000000", 29240 => x"00000000",
    29241 => x"00000000", 29242 => x"00000000", 29243 => x"00000000",
    29244 => x"00000000", 29245 => x"00000000", 29246 => x"00000000",
    29247 => x"00000000", 29248 => x"00000000", 29249 => x"00000000",
    29250 => x"00000000", 29251 => x"00000000", 29252 => x"00000000",
    29253 => x"00000000", 29254 => x"00000000", 29255 => x"00000000",
    29256 => x"00000000", 29257 => x"00000000", 29258 => x"00000000",
    29259 => x"00000000", 29260 => x"00000000", 29261 => x"00000000",
    29262 => x"00000000", 29263 => x"00000000", 29264 => x"00000000",
    29265 => x"00000000", 29266 => x"00000000", 29267 => x"00000000",
    29268 => x"00000000", 29269 => x"00000000", 29270 => x"00000000",
    29271 => x"00000000", 29272 => x"00000000", 29273 => x"00000000",
    29274 => x"00000000", 29275 => x"00000000", 29276 => x"00000000",
    29277 => x"00000000", 29278 => x"00000000", 29279 => x"00000000",
    29280 => x"00000000", 29281 => x"00000000", 29282 => x"00000000",
    29283 => x"00000000", 29284 => x"00000000", 29285 => x"00000000",
    29286 => x"00000000", 29287 => x"00000000", 29288 => x"00000000",
    29289 => x"00000000", 29290 => x"00000000", 29291 => x"00000000",
    29292 => x"00000000", 29293 => x"00000000", 29294 => x"00000000",
    29295 => x"00000000", 29296 => x"00000000", 29297 => x"00000000",
    29298 => x"00000000", 29299 => x"00000000", 29300 => x"00000000",
    29301 => x"00000000", 29302 => x"00000000", 29303 => x"00000000",
    29304 => x"00000000", 29305 => x"00000000", 29306 => x"00000000",
    29307 => x"00000000", 29308 => x"00000000", 29309 => x"00000000",
    29310 => x"00000000", 29311 => x"00000000", 29312 => x"00000000",
    29313 => x"00000000", 29314 => x"00000000", 29315 => x"00000000",
    29316 => x"00000000", 29317 => x"00000000", 29318 => x"00000000",
    29319 => x"00000000", 29320 => x"00000000", 29321 => x"00000000",
    29322 => x"00000000", 29323 => x"00000000", 29324 => x"00000000",
    29325 => x"00000000", 29326 => x"00000000", 29327 => x"00000000",
    29328 => x"00000000", 29329 => x"00000000", 29330 => x"00000000",
    29331 => x"00000000", 29332 => x"00000000", 29333 => x"00000000",
    29334 => x"00000000", 29335 => x"00000000", 29336 => x"00000000",
    29337 => x"00000000", 29338 => x"00000000", 29339 => x"00000000",
    29340 => x"00000000", 29341 => x"00000000", 29342 => x"00000000",
    29343 => x"00000000", 29344 => x"00000000", 29345 => x"00000000",
    29346 => x"00000000", 29347 => x"00000000", 29348 => x"00000000",
    29349 => x"00000000", 29350 => x"00000000", 29351 => x"00000000",
    29352 => x"00000000", 29353 => x"00000000", 29354 => x"00000000",
    29355 => x"00000000", 29356 => x"00000000", 29357 => x"00000000",
    29358 => x"00000000", 29359 => x"00000000", 29360 => x"00000000",
    29361 => x"00000000", 29362 => x"00000000", 29363 => x"00000000",
    29364 => x"00000000", 29365 => x"00000000", 29366 => x"00000000",
    29367 => x"00000000", 29368 => x"00000000", 29369 => x"00000000",
    29370 => x"00000000", 29371 => x"00000000", 29372 => x"00000000",
    29373 => x"00000000", 29374 => x"00000000", 29375 => x"00000000",
    29376 => x"00000000", 29377 => x"00000000", 29378 => x"00000000",
    29379 => x"00000000", 29380 => x"00000000", 29381 => x"00000000",
    29382 => x"00000000", 29383 => x"00000000", 29384 => x"00000000",
    29385 => x"00000000", 29386 => x"00000000", 29387 => x"00000000",
    29388 => x"00000000", 29389 => x"00000000", 29390 => x"00000000",
    29391 => x"00000000", 29392 => x"00000000", 29393 => x"00000000",
    29394 => x"00000000", 29395 => x"00000000", 29396 => x"00000000",
    29397 => x"00000000", 29398 => x"00000000", 29399 => x"00000000",
    29400 => x"00000000", 29401 => x"00000000", 29402 => x"00000000",
    29403 => x"00000000", 29404 => x"00000000", 29405 => x"00000000",
    29406 => x"00000000", 29407 => x"00000000", 29408 => x"00000000",
    29409 => x"00000000", 29410 => x"00000000", 29411 => x"00000000",
    29412 => x"00000000", 29413 => x"00000000", 29414 => x"00000000",
    29415 => x"00000000", 29416 => x"00000000", 29417 => x"00000000",
    29418 => x"00000000", 29419 => x"00000000", 29420 => x"00000000",
    29421 => x"00000000", 29422 => x"00000000", 29423 => x"00000000",
    29424 => x"00000000", 29425 => x"00000000", 29426 => x"00000000",
    29427 => x"00000000", 29428 => x"00000000", 29429 => x"00000000",
    29430 => x"00000000", 29431 => x"00000000", 29432 => x"00000000",
    29433 => x"00000000", 29434 => x"00000000", 29435 => x"00000000",
    29436 => x"00000000", 29437 => x"00000000", 29438 => x"00000000",
    29439 => x"00000000", 29440 => x"00000000", 29441 => x"00000000",
    29442 => x"00000000", 29443 => x"00000000", 29444 => x"00000000",
    29445 => x"00000000", 29446 => x"00000000", 29447 => x"00000000",
    29448 => x"00000000", 29449 => x"00000000", 29450 => x"00000000",
    29451 => x"00000000", 29452 => x"00000000", 29453 => x"00000000",
    29454 => x"00000000", 29455 => x"00000000", 29456 => x"00000000",
    29457 => x"00000000", 29458 => x"00000000", 29459 => x"00000000",
    29460 => x"00000000", 29461 => x"00000000", 29462 => x"00000000",
    29463 => x"00000000", 29464 => x"00000000", 29465 => x"00000000",
    29466 => x"00000000", 29467 => x"00000000", 29468 => x"00000000",
    29469 => x"00000000", 29470 => x"00000000", 29471 => x"00000000",
    29472 => x"00000000", 29473 => x"00000000", 29474 => x"00000000",
    29475 => x"00000000", 29476 => x"00000000", 29477 => x"00000000",
    29478 => x"00000000", 29479 => x"00000000", 29480 => x"00000000",
    29481 => x"00000000", 29482 => x"00000000", 29483 => x"00000000",
    29484 => x"00000000", 29485 => x"00000000", 29486 => x"00000000",
    29487 => x"00000000", 29488 => x"00000000", 29489 => x"00000000",
    29490 => x"00000000", 29491 => x"00000000", 29492 => x"00000000",
    29493 => x"00000000", 29494 => x"00000000", 29495 => x"00000000",
    29496 => x"00000000", 29497 => x"00000000", 29498 => x"00000000",
    29499 => x"00000000", 29500 => x"00000000", 29501 => x"00000000",
    29502 => x"00000000", 29503 => x"00000000", 29504 => x"00000000",
    29505 => x"00000000", 29506 => x"00000000", 29507 => x"00000000",
    29508 => x"00000000", 29509 => x"00000000", 29510 => x"00000000",
    29511 => x"00000000", 29512 => x"00000000", 29513 => x"00000000",
    29514 => x"00000000", 29515 => x"00000000", 29516 => x"00000000",
    29517 => x"00000000", 29518 => x"00000000", 29519 => x"00000000",
    29520 => x"00000000", 29521 => x"00000000", 29522 => x"00000000",
    29523 => x"00000000", 29524 => x"00000000", 29525 => x"00000000",
    29526 => x"00000000", 29527 => x"00000000", 29528 => x"00000000",
    29529 => x"00000000", 29530 => x"00000000", 29531 => x"00000000",
    29532 => x"00000000", 29533 => x"00000000", 29534 => x"00000000",
    29535 => x"00000000", 29536 => x"00000000", 29537 => x"00000000",
    29538 => x"00000000", 29539 => x"00000000", 29540 => x"00000000",
    29541 => x"00000000", 29542 => x"00000000", 29543 => x"00000000",
    29544 => x"00000000", 29545 => x"00000000", 29546 => x"00000000",
    29547 => x"00000000", 29548 => x"00000000", 29549 => x"00000000",
    29550 => x"00000000", 29551 => x"00000000", 29552 => x"00000000",
    29553 => x"00000000", 29554 => x"00000000", 29555 => x"00000000",
    29556 => x"00000000", 29557 => x"00000000", 29558 => x"00000000",
    29559 => x"00000000", 29560 => x"00000000", 29561 => x"00000000",
    29562 => x"00000000", 29563 => x"00000000", 29564 => x"00000000",
    29565 => x"00000000", 29566 => x"00000000", 29567 => x"00000000",
    29568 => x"00000000", 29569 => x"00000000", 29570 => x"00000000",
    29571 => x"00000000", 29572 => x"00000000", 29573 => x"00000000",
    29574 => x"00000000", 29575 => x"00000000", 29576 => x"00000000",
    29577 => x"00000000", 29578 => x"00000000", 29579 => x"00000000",
    29580 => x"00000000", 29581 => x"00000000", 29582 => x"00000000",
    29583 => x"00000000", 29584 => x"00000000", 29585 => x"00000000",
    29586 => x"00000000", 29587 => x"00000000", 29588 => x"00000000",
    29589 => x"00000000", 29590 => x"00000000", 29591 => x"00000000",
    29592 => x"00000000", 29593 => x"00000000", 29594 => x"00000000",
    29595 => x"00000000", 29596 => x"00000000", 29597 => x"00000000",
    29598 => x"00000000", 29599 => x"00000000", 29600 => x"00000000",
    29601 => x"00000000", 29602 => x"00000000", 29603 => x"00000000",
    29604 => x"00000000", 29605 => x"00000000", 29606 => x"00000000",
    29607 => x"00000000", 29608 => x"00000000", 29609 => x"00000000",
    29610 => x"00000000", 29611 => x"00000000", 29612 => x"00000000",
    29613 => x"00000000", 29614 => x"00000000", 29615 => x"00000000",
    29616 => x"00000000", 29617 => x"00000000", 29618 => x"00000000",
    29619 => x"00000000", 29620 => x"00000000", 29621 => x"00000000",
    29622 => x"00000000", 29623 => x"00000000", 29624 => x"00000000",
    29625 => x"00000000", 29626 => x"00000000", 29627 => x"00000000",
    29628 => x"00000000", 29629 => x"00000000", 29630 => x"00000000",
    29631 => x"00000000", 29632 => x"00000000", 29633 => x"00000000",
    29634 => x"00000000", 29635 => x"00000000", 29636 => x"00000000",
    29637 => x"00000000", 29638 => x"00000000", 29639 => x"00000000",
    29640 => x"00000000", 29641 => x"00000000", 29642 => x"00000000",
    29643 => x"00000000", 29644 => x"00000000", 29645 => x"00000000",
    29646 => x"00000000", 29647 => x"00000000", 29648 => x"00000000",
    29649 => x"00000000", 29650 => x"00000000", 29651 => x"00000000",
    29652 => x"00000000", 29653 => x"00000000", 29654 => x"00000000",
    29655 => x"00000000", 29656 => x"00000000", 29657 => x"00000000",
    29658 => x"00000000", 29659 => x"00000000", 29660 => x"00000000",
    29661 => x"00000000", 29662 => x"00000000", 29663 => x"00000000",
    29664 => x"00000000", 29665 => x"00000000", 29666 => x"00000000",
    29667 => x"00000000", 29668 => x"00000000", 29669 => x"00000000",
    29670 => x"00000000", 29671 => x"00000000", 29672 => x"00000000",
    29673 => x"00000000", 29674 => x"00000000", 29675 => x"00000000",
    29676 => x"00000000", 29677 => x"00000000", 29678 => x"00000000",
    29679 => x"00000000", 29680 => x"00000000", 29681 => x"00000000",
    29682 => x"00000000", 29683 => x"00000000", 29684 => x"00000000",
    29685 => x"00000000", 29686 => x"00000000", 29687 => x"00000000",
    29688 => x"00000000", 29689 => x"00000000", 29690 => x"00000000",
    29691 => x"00000000", 29692 => x"00000000", 29693 => x"00000000",
    29694 => x"00000000", 29695 => x"00000000", 29696 => x"00000000",
    29697 => x"00000000", 29698 => x"00000000", 29699 => x"00000000",
    29700 => x"00000000", 29701 => x"00000000", 29702 => x"00000000",
    29703 => x"00000000", 29704 => x"00000000", 29705 => x"00000000",
    29706 => x"00000000", 29707 => x"00000000", 29708 => x"00000000",
    29709 => x"00000000", 29710 => x"00000000", 29711 => x"00000000",
    29712 => x"00000000", 29713 => x"00000000", 29714 => x"00000000",
    29715 => x"00000000", 29716 => x"00000000", 29717 => x"00000000",
    29718 => x"00000000", 29719 => x"00000000", 29720 => x"00000000",
    29721 => x"00000000", 29722 => x"00000000", 29723 => x"00000000",
    29724 => x"00000000", 29725 => x"00000000", 29726 => x"00000000",
    29727 => x"00000000", 29728 => x"00000000", 29729 => x"00000000",
    29730 => x"00000000", 29731 => x"00000000", 29732 => x"00000000",
    29733 => x"00000000", 29734 => x"00000000", 29735 => x"00000000",
    29736 => x"00000000", 29737 => x"00000000", 29738 => x"00000000",
    29739 => x"00000000", 29740 => x"00000000", 29741 => x"00000000",
    29742 => x"00000000", 29743 => x"00000000", 29744 => x"00000000",
    29745 => x"00000000", 29746 => x"00000000", 29747 => x"00000000",
    29748 => x"00000000", 29749 => x"00000000", 29750 => x"00000000",
    29751 => x"00000000", 29752 => x"00000000", 29753 => x"00000000",
    29754 => x"00000000", 29755 => x"00000000", 29756 => x"00000000",
    29757 => x"00000000", 29758 => x"00000000", 29759 => x"00000000",
    29760 => x"00000000", 29761 => x"00000000", 29762 => x"00000000",
    29763 => x"00000000", 29764 => x"00000000", 29765 => x"00000000",
    29766 => x"00000000", 29767 => x"00000000", 29768 => x"00000000",
    29769 => x"00000000", 29770 => x"00000000", 29771 => x"00000000",
    29772 => x"00000000", 29773 => x"00000000", 29774 => x"00000000",
    29775 => x"00000000", 29776 => x"00000000", 29777 => x"00000000",
    29778 => x"00000000", 29779 => x"00000000", 29780 => x"00000000",
    29781 => x"00000000", 29782 => x"00000000", 29783 => x"00000000",
    29784 => x"00000000", 29785 => x"00000000", 29786 => x"00000000",
    29787 => x"00000000", 29788 => x"00000000", 29789 => x"00000000",
    29790 => x"00000000", 29791 => x"00000000", 29792 => x"00000000",
    29793 => x"00000000", 29794 => x"00000000", 29795 => x"00000000",
    29796 => x"00000000", 29797 => x"00000000", 29798 => x"00000000",
    29799 => x"00000000", 29800 => x"00000000", 29801 => x"00000000",
    29802 => x"00000000", 29803 => x"00000000", 29804 => x"00000000",
    29805 => x"00000000", 29806 => x"00000000", 29807 => x"00000000",
    29808 => x"00000000", 29809 => x"00000000", 29810 => x"00000000",
    29811 => x"00000000", 29812 => x"00000000", 29813 => x"00000000",
    29814 => x"00000000", 29815 => x"00000000", 29816 => x"00000000",
    29817 => x"00000000", 29818 => x"00000000", 29819 => x"00000000",
    29820 => x"00000000", 29821 => x"00000000", 29822 => x"00000000",
    29823 => x"00000000", 29824 => x"00000000", 29825 => x"00000000",
    29826 => x"00000000", 29827 => x"00000000", 29828 => x"00000000",
    29829 => x"00000000", 29830 => x"00000000", 29831 => x"00000000",
    29832 => x"00000000", 29833 => x"00000000", 29834 => x"00000000",
    29835 => x"00000000", 29836 => x"00000000", 29837 => x"00000000",
    29838 => x"00000000", 29839 => x"00000000", 29840 => x"00000000",
    29841 => x"00000000", 29842 => x"00000000", 29843 => x"00000000",
    29844 => x"00000000", 29845 => x"00000000", 29846 => x"00000000",
    29847 => x"00000000", 29848 => x"00000000", 29849 => x"00000000",
    29850 => x"00000000", 29851 => x"00000000", 29852 => x"00000000",
    29853 => x"00000000", 29854 => x"00000000", 29855 => x"00000000",
    29856 => x"00000000", 29857 => x"00000000", 29858 => x"00000000",
    29859 => x"00000000", 29860 => x"00000000", 29861 => x"00000000",
    29862 => x"00000000", 29863 => x"00000000", 29864 => x"00000000",
    29865 => x"00000000", 29866 => x"00000000", 29867 => x"00000000",
    29868 => x"00000000", 29869 => x"00000000", 29870 => x"00000000",
    29871 => x"00000000", 29872 => x"00000000", 29873 => x"00000000",
    29874 => x"00000000", 29875 => x"00000000", 29876 => x"00000000",
    29877 => x"00000000", 29878 => x"00000000", 29879 => x"00000000",
    29880 => x"00000000", 29881 => x"00000000", 29882 => x"00000000",
    29883 => x"00000000", 29884 => x"00000000", 29885 => x"00000000",
    29886 => x"00000000", 29887 => x"00000000", 29888 => x"00000000",
    29889 => x"00000000", 29890 => x"00000000", 29891 => x"00000000",
    29892 => x"00000000", 29893 => x"00000000", 29894 => x"00000000",
    29895 => x"00000000", 29896 => x"00000000", 29897 => x"00000000",
    29898 => x"00000000", 29899 => x"00000000", 29900 => x"00000000",
    29901 => x"00000000", 29902 => x"00000000", 29903 => x"00000000",
    29904 => x"00000000", 29905 => x"00000000", 29906 => x"00000000",
    29907 => x"00000000", 29908 => x"00000000", 29909 => x"00000000",
    29910 => x"00000000", 29911 => x"00000000", 29912 => x"00000000",
    29913 => x"00000000", 29914 => x"00000000", 29915 => x"00000000",
    29916 => x"00000000", 29917 => x"00000000", 29918 => x"00000000",
    29919 => x"00000000", 29920 => x"00000000", 29921 => x"00000000",
    29922 => x"00000000", 29923 => x"00000000", 29924 => x"00000000",
    29925 => x"00000000", 29926 => x"00000000", 29927 => x"00000000",
    29928 => x"00000000", 29929 => x"00000000", 29930 => x"00000000",
    29931 => x"00000000", 29932 => x"00000000", 29933 => x"00000000",
    29934 => x"00000000", 29935 => x"00000000", 29936 => x"00000000",
    29937 => x"00000000", 29938 => x"00000000", 29939 => x"00000000",
    29940 => x"00000000", 29941 => x"00000000", 29942 => x"00000000",
    29943 => x"00000000", 29944 => x"00000000", 29945 => x"00000000",
    29946 => x"00000000", 29947 => x"00000000", 29948 => x"00000000",
    29949 => x"00000000", 29950 => x"00000000", 29951 => x"00000000",
    29952 => x"00000000", 29953 => x"00000000", 29954 => x"00000000",
    29955 => x"00000000", 29956 => x"00000000", 29957 => x"00000000",
    29958 => x"00000000", 29959 => x"00000000", 29960 => x"00000000",
    29961 => x"00000000", 29962 => x"00000000", 29963 => x"00000000",
    29964 => x"00000000", 29965 => x"00000000", 29966 => x"00000000",
    29967 => x"00000000", 29968 => x"00000000", 29969 => x"00000000",
    29970 => x"00000000", 29971 => x"00000000", 29972 => x"00000000",
    29973 => x"00000000", 29974 => x"00000000", 29975 => x"00000000",
    29976 => x"00000000", 29977 => x"00000000", 29978 => x"00000000",
    29979 => x"00000000", 29980 => x"00000000", 29981 => x"00000000",
    29982 => x"00000000", 29983 => x"00000000", 29984 => x"00000000",
    29985 => x"00000000", 29986 => x"00000000", 29987 => x"00000000",
    29988 => x"00000000", 29989 => x"00000000", 29990 => x"00000000",
    29991 => x"00000000", 29992 => x"00000000", 29993 => x"00000000",
    29994 => x"00000000", 29995 => x"00000000", 29996 => x"00000000",
    29997 => x"00000000", 29998 => x"00000000", 29999 => x"00000000",
    30000 => x"00000000", 30001 => x"00000000", 30002 => x"00000000",
    30003 => x"00000000", 30004 => x"00000000", 30005 => x"00000000",
    30006 => x"00000000", 30007 => x"00000000", 30008 => x"00000000",
    30009 => x"00000000", 30010 => x"00000000", 30011 => x"00000000",
    30012 => x"00000000", 30013 => x"00000000", 30014 => x"00000000",
    30015 => x"00000000", 30016 => x"00000000", 30017 => x"00000000",
    30018 => x"00000000", 30019 => x"00000000", 30020 => x"00000000",
    30021 => x"00000000", 30022 => x"00000000", 30023 => x"00000000",
    30024 => x"00000000", 30025 => x"00000000", 30026 => x"00000000",
    30027 => x"00000000", 30028 => x"00000000", 30029 => x"00000000",
    30030 => x"00000000", 30031 => x"00000000", 30032 => x"00000000",
    30033 => x"00000000", 30034 => x"00000000", 30035 => x"00000000",
    30036 => x"00000000", 30037 => x"00000000", 30038 => x"00000000",
    30039 => x"00000000", 30040 => x"00000000", 30041 => x"00000000",
    30042 => x"00000000", 30043 => x"00000000", 30044 => x"00000000",
    30045 => x"00000000", 30046 => x"00000000", 30047 => x"00000000",
    30048 => x"00000000", 30049 => x"00000000", 30050 => x"00000000",
    30051 => x"00000000", 30052 => x"00000000", 30053 => x"00000000",
    30054 => x"00000000", 30055 => x"00000000", 30056 => x"00000000",
    30057 => x"00000000", 30058 => x"00000000", 30059 => x"00000000",
    30060 => x"00000000", 30061 => x"00000000", 30062 => x"00000000",
    30063 => x"00000000", 30064 => x"00000000", 30065 => x"00000000",
    30066 => x"00000000", 30067 => x"00000000", 30068 => x"00000000",
    30069 => x"00000000", 30070 => x"00000000", 30071 => x"00000000",
    30072 => x"00000000", 30073 => x"00000000", 30074 => x"00000000",
    30075 => x"00000000", 30076 => x"00000000", 30077 => x"00000000",
    30078 => x"00000000", 30079 => x"00000000", 30080 => x"00000000",
    30081 => x"00000000", 30082 => x"00000000", 30083 => x"00000000",
    30084 => x"00000000", 30085 => x"00000000", 30086 => x"00000000",
    30087 => x"00000000", 30088 => x"00000000", 30089 => x"00000000",
    30090 => x"00000000", 30091 => x"00000000", 30092 => x"00000000",
    30093 => x"00000000", 30094 => x"00000000", 30095 => x"00000000",
    30096 => x"00000000", 30097 => x"00000000", 30098 => x"00000000",
    30099 => x"00000000", 30100 => x"00000000", 30101 => x"00000000",
    30102 => x"00000000", 30103 => x"00000000", 30104 => x"00000000",
    30105 => x"00000000", 30106 => x"00000000", 30107 => x"00000000",
    30108 => x"00000000", 30109 => x"00000000", 30110 => x"00000000",
    30111 => x"00000000", 30112 => x"00000000", 30113 => x"00000000",
    30114 => x"00000000", 30115 => x"00000000", 30116 => x"00000000",
    30117 => x"00000000", 30118 => x"00000000", 30119 => x"00000000",
    30120 => x"00000000", 30121 => x"00000000", 30122 => x"00000000",
    30123 => x"00000000", 30124 => x"00000000", 30125 => x"00000000",
    30126 => x"00000000", 30127 => x"00000000", 30128 => x"00000000",
    30129 => x"00000000", 30130 => x"00000000", 30131 => x"00000000",
    30132 => x"00000000", 30133 => x"00000000", 30134 => x"00000000",
    30135 => x"00000000", 30136 => x"00000000", 30137 => x"00000000",
    30138 => x"00000000", 30139 => x"00000000", 30140 => x"00000000",
    30141 => x"00000000", 30142 => x"00000000", 30143 => x"00000000",
    30144 => x"00000000", 30145 => x"00000000", 30146 => x"00000000",
    30147 => x"00000000", 30148 => x"00000000", 30149 => x"00000000",
    30150 => x"00000000", 30151 => x"00000000", 30152 => x"00000000",
    30153 => x"00000000", 30154 => x"00000000", 30155 => x"00000000",
    30156 => x"00000000", 30157 => x"00000000", 30158 => x"00000000",
    30159 => x"00000000", 30160 => x"00000000", 30161 => x"00000000",
    30162 => x"00000000", 30163 => x"00000000", 30164 => x"00000000",
    30165 => x"00000000", 30166 => x"00000000", 30167 => x"00000000",
    30168 => x"00000000", 30169 => x"00000000", 30170 => x"00000000",
    30171 => x"00000000", 30172 => x"00000000", 30173 => x"00000000",
    30174 => x"00000000", 30175 => x"00000000", 30176 => x"00000000",
    30177 => x"00000000", 30178 => x"00000000", 30179 => x"00000000",
    30180 => x"00000000", 30181 => x"00000000", 30182 => x"00000000",
    30183 => x"00000000", 30184 => x"00000000", 30185 => x"00000000",
    30186 => x"00000000", 30187 => x"00000000", 30188 => x"00000000",
    30189 => x"00000000", 30190 => x"00000000", 30191 => x"00000000",
    30192 => x"00000000", 30193 => x"00000000", 30194 => x"00000000",
    30195 => x"00000000", 30196 => x"00000000", 30197 => x"00000000",
    30198 => x"00000000", 30199 => x"00000000", 30200 => x"00000000",
    30201 => x"00000000", 30202 => x"00000000", 30203 => x"00000000",
    30204 => x"00000000", 30205 => x"00000000", 30206 => x"00000000",
    30207 => x"00000000", 30208 => x"00000000", 30209 => x"00000000",
    30210 => x"00000000", 30211 => x"00000000", 30212 => x"00000000",
    30213 => x"00000000", 30214 => x"00000000", 30215 => x"00000000",
    30216 => x"00000000", 30217 => x"00000000", 30218 => x"00000000",
    30219 => x"00000000", 30220 => x"00000000", 30221 => x"00000000",
    30222 => x"00000000", 30223 => x"00000000", 30224 => x"00000000",
    30225 => x"00000000", 30226 => x"00000000", 30227 => x"00000000",
    30228 => x"00000000", 30229 => x"00000000", 30230 => x"00000000",
    30231 => x"00000000", 30232 => x"00000000", 30233 => x"00000000",
    30234 => x"00000000", 30235 => x"00000000", 30236 => x"00000000",
    30237 => x"00000000", 30238 => x"00000000", 30239 => x"00000000",
    30240 => x"00000000", 30241 => x"00000000", 30242 => x"00000000",
    30243 => x"00000000", 30244 => x"00000000", 30245 => x"00000000",
    30246 => x"00000000", 30247 => x"00000000", 30248 => x"00000000",
    30249 => x"00000000", 30250 => x"00000000", 30251 => x"00000000",
    30252 => x"00000000", 30253 => x"00000000", 30254 => x"00000000",
    30255 => x"00000000", 30256 => x"00000000", 30257 => x"00000000",
    30258 => x"00000000", 30259 => x"00000000", 30260 => x"00000000",
    30261 => x"00000000", 30262 => x"00000000", 30263 => x"00000000",
    30264 => x"00000000", 30265 => x"00000000", 30266 => x"00000000",
    30267 => x"00000000", 30268 => x"00000000", 30269 => x"00000000",
    30270 => x"00000000", 30271 => x"00000000", 30272 => x"00000000",
    30273 => x"00000000", 30274 => x"00000000", 30275 => x"00000000",
    30276 => x"00000000", 30277 => x"00000000", 30278 => x"00000000",
    30279 => x"00000000", 30280 => x"00000000", 30281 => x"00000000",
    30282 => x"00000000", 30283 => x"00000000", 30284 => x"00000000",
    30285 => x"00000000", 30286 => x"00000000", 30287 => x"00000000",
    30288 => x"00000000", 30289 => x"00000000", 30290 => x"00000000",
    30291 => x"00000000", 30292 => x"00000000", 30293 => x"00000000",
    30294 => x"00000000", 30295 => x"00000000", 30296 => x"00000000",
    30297 => x"00000000", 30298 => x"00000000", 30299 => x"00000000",
    30300 => x"00000000", 30301 => x"00000000", 30302 => x"00000000",
    30303 => x"00000000", 30304 => x"00000000", 30305 => x"00000000",
    30306 => x"00000000", 30307 => x"00000000", 30308 => x"00000000",
    30309 => x"00000000", 30310 => x"00000000", 30311 => x"00000000",
    30312 => x"00000000", 30313 => x"00000000", 30314 => x"00000000",
    30315 => x"00000000", 30316 => x"00000000", 30317 => x"00000000",
    30318 => x"00000000", 30319 => x"00000000", 30320 => x"00000000",
    30321 => x"00000000", 30322 => x"00000000", 30323 => x"00000000",
    30324 => x"00000000", 30325 => x"00000000", 30326 => x"00000000",
    30327 => x"00000000", 30328 => x"00000000", 30329 => x"00000000",
    30330 => x"00000000", 30331 => x"00000000", 30332 => x"00000000",
    30333 => x"00000000", 30334 => x"00000000", 30335 => x"00000000",
    30336 => x"00000000", 30337 => x"00000000", 30338 => x"00000000",
    30339 => x"00000000", 30340 => x"00000000", 30341 => x"00000000",
    30342 => x"00000000", 30343 => x"00000000", 30344 => x"00000000",
    30345 => x"00000000", 30346 => x"00000000", 30347 => x"00000000",
    30348 => x"00000000", 30349 => x"00000000", 30350 => x"00000000",
    30351 => x"00000000", 30352 => x"00000000", 30353 => x"00000000",
    30354 => x"00000000", 30355 => x"00000000", 30356 => x"00000000",
    30357 => x"00000000", 30358 => x"00000000", 30359 => x"00000000",
    30360 => x"00000000", 30361 => x"00000000", 30362 => x"00000000",
    30363 => x"00000000", 30364 => x"00000000", 30365 => x"00000000",
    30366 => x"00000000", 30367 => x"00000000", 30368 => x"00000000",
    30369 => x"00000000", 30370 => x"00000000", 30371 => x"00000000",
    30372 => x"00000000", 30373 => x"00000000", 30374 => x"00000000",
    30375 => x"00000000", 30376 => x"00000000", 30377 => x"00000000",
    30378 => x"00000000", 30379 => x"00000000", 30380 => x"00000000",
    30381 => x"00000000", 30382 => x"00000000", 30383 => x"00000000",
    30384 => x"00000000", 30385 => x"00000000", 30386 => x"00000000",
    30387 => x"00000000", 30388 => x"00000000", 30389 => x"00000000",
    30390 => x"00000000", 30391 => x"00000000", 30392 => x"00000000",
    30393 => x"00000000", 30394 => x"00000000", 30395 => x"00000000",
    30396 => x"00000000", 30397 => x"00000000", 30398 => x"00000000",
    30399 => x"00000000", 30400 => x"00000000", 30401 => x"00000000",
    30402 => x"00000000", 30403 => x"00000000", 30404 => x"00000000",
    30405 => x"00000000", 30406 => x"00000000", 30407 => x"00000000",
    30408 => x"00000000", 30409 => x"00000000", 30410 => x"00000000",
    30411 => x"00000000", 30412 => x"00000000", 30413 => x"00000000",
    30414 => x"00000000", 30415 => x"00000000", 30416 => x"00000000",
    30417 => x"00000000", 30418 => x"00000000", 30419 => x"00000000",
    30420 => x"00000000", 30421 => x"00000000", 30422 => x"00000000",
    30423 => x"00000000", 30424 => x"00000000", 30425 => x"00000000",
    30426 => x"00000000", 30427 => x"00000000", 30428 => x"00000000",
    30429 => x"00000000", 30430 => x"00000000", 30431 => x"00000000",
    30432 => x"00000000", 30433 => x"00000000", 30434 => x"00000000",
    30435 => x"00000000", 30436 => x"00000000", 30437 => x"00000000",
    30438 => x"00000000", 30439 => x"00000000", 30440 => x"00000000",
    30441 => x"00000000", 30442 => x"00000000", 30443 => x"00000000",
    30444 => x"00000000", 30445 => x"00000000", 30446 => x"00000000",
    30447 => x"00000000", 30448 => x"00000000", 30449 => x"00000000",
    30450 => x"00000000", 30451 => x"00000000", 30452 => x"00000000",
    30453 => x"00000000", 30454 => x"00000000", 30455 => x"00000000",
    30456 => x"00000000", 30457 => x"00000000", 30458 => x"00000000",
    30459 => x"00000000", 30460 => x"00000000", 30461 => x"00000000",
    30462 => x"00000000", 30463 => x"00000000", 30464 => x"00000000",
    30465 => x"00000000", 30466 => x"00000000", 30467 => x"00000000",
    30468 => x"00000000", 30469 => x"00000000", 30470 => x"00000000",
    30471 => x"00000000", 30472 => x"00000000", 30473 => x"00000000",
    30474 => x"00000000", 30475 => x"00000000", 30476 => x"00000000",
    30477 => x"00000000", 30478 => x"00000000", 30479 => x"00000000",
    30480 => x"00000000", 30481 => x"00000000", 30482 => x"00000000",
    30483 => x"00000000", 30484 => x"00000000", 30485 => x"00000000",
    30486 => x"00000000", 30487 => x"00000000", 30488 => x"00000000",
    30489 => x"00000000", 30490 => x"00000000", 30491 => x"00000000",
    30492 => x"00000000", 30493 => x"00000000", 30494 => x"00000000",
    30495 => x"00000000", 30496 => x"00000000", 30497 => x"00000000",
    30498 => x"00000000", 30499 => x"00000000", 30500 => x"00000000",
    30501 => x"00000000", 30502 => x"00000000", 30503 => x"00000000",
    30504 => x"00000000", 30505 => x"00000000", 30506 => x"00000000",
    30507 => x"00000000", 30508 => x"00000000", 30509 => x"00000000",
    30510 => x"00000000", 30511 => x"00000000", 30512 => x"00000000",
    30513 => x"00000000", 30514 => x"00000000", 30515 => x"00000000",
    30516 => x"00000000", 30517 => x"00000000", 30518 => x"00000000",
    30519 => x"00000000", 30520 => x"00000000", 30521 => x"00000000",
    30522 => x"00000000", 30523 => x"00000000", 30524 => x"00000000",
    30525 => x"00000000", 30526 => x"00000000", 30527 => x"00000000",
    30528 => x"00000000", 30529 => x"00000000", 30530 => x"00000000",
    30531 => x"00000000", 30532 => x"00000000", 30533 => x"00000000",
    30534 => x"00000000", 30535 => x"00000000", 30536 => x"00000000",
    30537 => x"00000000", 30538 => x"00000000", 30539 => x"00000000",
    30540 => x"00000000", 30541 => x"00000000", 30542 => x"00000000",
    30543 => x"00000000", 30544 => x"00000000", 30545 => x"00000000",
    30546 => x"00000000", 30547 => x"00000000", 30548 => x"00000000",
    30549 => x"00000000", 30550 => x"00000000", 30551 => x"00000000",
    30552 => x"00000000", 30553 => x"00000000", 30554 => x"00000000",
    30555 => x"00000000", 30556 => x"00000000", 30557 => x"00000000",
    30558 => x"00000000", 30559 => x"00000000", 30560 => x"00000000",
    30561 => x"00000000", 30562 => x"00000000", 30563 => x"00000000",
    30564 => x"00000000", 30565 => x"00000000", 30566 => x"00000000",
    30567 => x"00000000", 30568 => x"00000000", 30569 => x"00000000",
    30570 => x"00000000", 30571 => x"00000000", 30572 => x"00000000",
    30573 => x"00000000", 30574 => x"00000000", 30575 => x"00000000",
    30576 => x"00000000", 30577 => x"00000000", 30578 => x"00000000",
    30579 => x"00000000", 30580 => x"00000000", 30581 => x"00000000",
    30582 => x"00000000", 30583 => x"00000000", 30584 => x"00000000",
    30585 => x"00000000", 30586 => x"00000000", 30587 => x"00000000",
    30588 => x"00000000", 30589 => x"00000000", 30590 => x"00000000",
    30591 => x"00000000", 30592 => x"00000000", 30593 => x"00000000",
    30594 => x"00000000", 30595 => x"00000000", 30596 => x"00000000",
    30597 => x"00000000", 30598 => x"00000000", 30599 => x"00000000",
    30600 => x"00000000", 30601 => x"00000000", 30602 => x"00000000",
    30603 => x"00000000", 30604 => x"00000000", 30605 => x"00000000",
    30606 => x"00000000", 30607 => x"00000000", 30608 => x"00000000",
    30609 => x"00000000", 30610 => x"00000000", 30611 => x"00000000",
    30612 => x"00000000", 30613 => x"00000000", 30614 => x"00000000",
    30615 => x"00000000", 30616 => x"00000000", 30617 => x"00000000",
    30618 => x"00000000", 30619 => x"00000000", 30620 => x"00000000",
    30621 => x"00000000", 30622 => x"00000000", 30623 => x"00000000",
    30624 => x"00000000", 30625 => x"00000000", 30626 => x"00000000",
    30627 => x"00000000", 30628 => x"00000000", 30629 => x"00000000",
    30630 => x"00000000", 30631 => x"00000000", 30632 => x"00000000",
    30633 => x"00000000", 30634 => x"00000000", 30635 => x"00000000",
    30636 => x"00000000", 30637 => x"00000000", 30638 => x"00000000",
    30639 => x"00000000", 30640 => x"00000000", 30641 => x"00000000",
    30642 => x"00000000", 30643 => x"00000000", 30644 => x"00000000",
    30645 => x"00000000", 30646 => x"00000000", 30647 => x"00000000",
    30648 => x"00000000", 30649 => x"00000000", 30650 => x"00000000",
    30651 => x"00000000", 30652 => x"00000000", 30653 => x"00000000",
    30654 => x"00000000", 30655 => x"00000000", 30656 => x"00000000",
    30657 => x"00000000", 30658 => x"00000000", 30659 => x"00000000",
    30660 => x"00000000", 30661 => x"00000000", 30662 => x"00000000",
    30663 => x"00000000", 30664 => x"00000000", 30665 => x"00000000",
    30666 => x"00000000", 30667 => x"00000000", 30668 => x"00000000",
    30669 => x"00000000", 30670 => x"00000000", 30671 => x"00000000",
    30672 => x"00000000", 30673 => x"00000000", 30674 => x"00000000",
    30675 => x"00000000", 30676 => x"00000000", 30677 => x"00000000",
    30678 => x"00000000", 30679 => x"00000000", 30680 => x"00000000",
    30681 => x"00000000", 30682 => x"00000000", 30683 => x"00000000",
    30684 => x"00000000", 30685 => x"00000000", 30686 => x"00000000",
    30687 => x"00000000", 30688 => x"00000000", 30689 => x"00000000",
    30690 => x"00000000", 30691 => x"00000000", 30692 => x"00000000",
    30693 => x"00000000", 30694 => x"00000000", 30695 => x"00000000",
    30696 => x"00000000", 30697 => x"00000000", 30698 => x"00000000",
    30699 => x"00000000", 30700 => x"00000000", 30701 => x"00000000",
    30702 => x"00000000", 30703 => x"00000000", 30704 => x"00000000",
    30705 => x"00000000", 30706 => x"00000000", 30707 => x"00000000",
    30708 => x"00000000", 30709 => x"00000000", 30710 => x"00000000",
    30711 => x"00000000", 30712 => x"00000000", 30713 => x"00000000",
    30714 => x"00000000", 30715 => x"00000000", 30716 => x"00000000",
    30717 => x"00000000", 30718 => x"00000000", 30719 => x"00000000",
    30720 => x"00000000", 30721 => x"00000000", 30722 => x"00000000",
    30723 => x"00000000", 30724 => x"00000000", 30725 => x"00000000",
    30726 => x"00000000", 30727 => x"00000000", 30728 => x"00000000",
    30729 => x"00000000", 30730 => x"00000000", 30731 => x"00000000",
    30732 => x"00000000", 30733 => x"00000000", 30734 => x"00000000",
    30735 => x"00000000", 30736 => x"00000000", 30737 => x"00000000",
    30738 => x"00000000", 30739 => x"00000000", 30740 => x"00000000",
    30741 => x"00000000", 30742 => x"00000000", 30743 => x"00000000",
    30744 => x"00000000", 30745 => x"00000000", 30746 => x"00000000",
    30747 => x"00000000", 30748 => x"00000000", 30749 => x"00000000",
    30750 => x"00000000", 30751 => x"00000000", 30752 => x"00000000",
    30753 => x"00000000", 30754 => x"00000000", 30755 => x"00000000",
    30756 => x"00000000", 30757 => x"00000000", 30758 => x"00000000",
    30759 => x"00000000", 30760 => x"00000000", 30761 => x"00000000",
    30762 => x"00000000", 30763 => x"00000000", 30764 => x"00000000",
    30765 => x"00000000", 30766 => x"00000000", 30767 => x"00000000",
    30768 => x"00000000", 30769 => x"00000000", 30770 => x"00000000",
    30771 => x"00000000", 30772 => x"00000000", 30773 => x"00000000",
    30774 => x"00000000", 30775 => x"00000000", 30776 => x"00000000",
    30777 => x"00000000", 30778 => x"00000000", 30779 => x"00000000",
    30780 => x"00000000", 30781 => x"00000000", 30782 => x"00000000",
    30783 => x"00000000", 30784 => x"00000000", 30785 => x"00000000",
    30786 => x"00000000", 30787 => x"00000000", 30788 => x"00000000",
    30789 => x"00000000", 30790 => x"00000000", 30791 => x"00000000",
    30792 => x"00000000", 30793 => x"00000000", 30794 => x"00000000",
    30795 => x"00000000", 30796 => x"00000000", 30797 => x"00000000",
    30798 => x"00000000", 30799 => x"00000000", 30800 => x"00000000",
    30801 => x"00000000", 30802 => x"00000000", 30803 => x"00000000",
    30804 => x"00000000", 30805 => x"00000000", 30806 => x"00000000",
    30807 => x"00000000", 30808 => x"00000000", 30809 => x"00000000",
    30810 => x"00000000", 30811 => x"00000000", 30812 => x"00000000",
    30813 => x"00000000", 30814 => x"00000000", 30815 => x"00000000",
    30816 => x"00000000", 30817 => x"00000000", 30818 => x"00000000",
    30819 => x"00000000", 30820 => x"00000000", 30821 => x"00000000",
    30822 => x"00000000", 30823 => x"00000000", 30824 => x"00000000",
    30825 => x"00000000", 30826 => x"00000000", 30827 => x"00000000",
    30828 => x"00000000", 30829 => x"00000000", 30830 => x"00000000",
    30831 => x"00000000", 30832 => x"00000000", 30833 => x"00000000",
    30834 => x"00000000", 30835 => x"00000000", 30836 => x"00000000",
    30837 => x"00000000", 30838 => x"00000000", 30839 => x"00000000",
    30840 => x"00000000", 30841 => x"00000000", 30842 => x"00000000",
    30843 => x"00000000", 30844 => x"00000000", 30845 => x"00000000",
    30846 => x"00000000", 30847 => x"00000000", 30848 => x"00000000",
    30849 => x"00000000", 30850 => x"00000000", 30851 => x"00000000",
    30852 => x"00000000", 30853 => x"00000000", 30854 => x"00000000",
    30855 => x"00000000", 30856 => x"00000000", 30857 => x"00000000",
    30858 => x"00000000", 30859 => x"00000000", 30860 => x"00000000",
    30861 => x"00000000", 30862 => x"00000000", 30863 => x"00000000",
    30864 => x"00000000", 30865 => x"00000000", 30866 => x"00000000",
    30867 => x"00000000", 30868 => x"00000000", 30869 => x"00000000",
    30870 => x"00000000", 30871 => x"00000000", 30872 => x"00000000",
    30873 => x"00000000", 30874 => x"00000000", 30875 => x"00000000",
    30876 => x"00000000", 30877 => x"00000000", 30878 => x"00000000",
    30879 => x"00000000", 30880 => x"00000000", 30881 => x"00000000",
    30882 => x"00000000", 30883 => x"00000000", 30884 => x"00000000",
    30885 => x"00000000", 30886 => x"00000000", 30887 => x"00000000",
    30888 => x"00000000", 30889 => x"00000000", 30890 => x"00000000",
    30891 => x"00000000", 30892 => x"00000000", 30893 => x"00000000",
    30894 => x"00000000", 30895 => x"00000000", 30896 => x"00000000",
    30897 => x"00000000", 30898 => x"00000000", 30899 => x"00000000",
    30900 => x"00000000", 30901 => x"00000000", 30902 => x"00000000",
    30903 => x"00000000", 30904 => x"00000000", 30905 => x"00000000",
    30906 => x"00000000", 30907 => x"00000000", 30908 => x"00000000",
    30909 => x"00000000", 30910 => x"00000000", 30911 => x"00000000",
    30912 => x"00000000", 30913 => x"00000000", 30914 => x"00000000",
    30915 => x"00000000", 30916 => x"00000000", 30917 => x"00000000",
    30918 => x"00000000", 30919 => x"00000000", 30920 => x"00000000",
    30921 => x"00000000", 30922 => x"00000000", 30923 => x"00000000",
    30924 => x"00000000", 30925 => x"00000000", 30926 => x"00000000",
    30927 => x"00000000", 30928 => x"00000000", 30929 => x"00000000",
    30930 => x"00000000", 30931 => x"00000000", 30932 => x"00000000",
    30933 => x"00000000", 30934 => x"00000000", 30935 => x"00000000",
    30936 => x"00000000", 30937 => x"00000000", 30938 => x"00000000",
    30939 => x"00000000", 30940 => x"00000000", 30941 => x"00000000",
    30942 => x"00000000", 30943 => x"00000000", 30944 => x"00000000",
    30945 => x"00000000", 30946 => x"00000000", 30947 => x"00000000",
    30948 => x"00000000", 30949 => x"00000000", 30950 => x"00000000",
    30951 => x"00000000", 30952 => x"00000000", 30953 => x"00000000",
    30954 => x"00000000", 30955 => x"00000000", 30956 => x"00000000",
    30957 => x"00000000", 30958 => x"00000000", 30959 => x"00000000",
    30960 => x"00000000", 30961 => x"00000000", 30962 => x"00000000",
    30963 => x"00000000", 30964 => x"00000000", 30965 => x"00000000",
    30966 => x"00000000", 30967 => x"00000000", 30968 => x"00000000",
    30969 => x"00000000", 30970 => x"00000000", 30971 => x"00000000",
    30972 => x"00000000", 30973 => x"00000000", 30974 => x"00000000",
    30975 => x"00000000", 30976 => x"00000000", 30977 => x"00000000",
    30978 => x"00000000", 30979 => x"00000000", 30980 => x"00000000",
    30981 => x"00000000", 30982 => x"00000000", 30983 => x"00000000",
    30984 => x"00000000", 30985 => x"00000000", 30986 => x"00000000",
    30987 => x"00000000", 30988 => x"00000000", 30989 => x"00000000",
    30990 => x"00000000", 30991 => x"00000000", 30992 => x"00000000",
    30993 => x"00000000", 30994 => x"00000000", 30995 => x"00000000",
    30996 => x"00000000", 30997 => x"00000000", 30998 => x"00000000",
    30999 => x"00000000", 31000 => x"00000000", 31001 => x"00000000",
    31002 => x"00000000", 31003 => x"00000000", 31004 => x"00000000",
    31005 => x"00000000", 31006 => x"00000000", 31007 => x"00000000",
    31008 => x"00000000", 31009 => x"00000000", 31010 => x"00000000",
    31011 => x"00000000", 31012 => x"00000000", 31013 => x"00000000",
    31014 => x"00000000", 31015 => x"00000000", 31016 => x"00000000",
    31017 => x"00000000", 31018 => x"00000000", 31019 => x"00000000",
    31020 => x"00000000", 31021 => x"00000000", 31022 => x"00000000",
    31023 => x"00000000", 31024 => x"00000000", 31025 => x"00000000",
    31026 => x"00000000", 31027 => x"00000000", 31028 => x"00000000",
    31029 => x"00000000", 31030 => x"00000000", 31031 => x"00000000",
    31032 => x"00000000", 31033 => x"00000000", 31034 => x"00000000",
    31035 => x"00000000", 31036 => x"00000000", 31037 => x"00000000",
    31038 => x"00000000", 31039 => x"00000000", 31040 => x"00000000",
    31041 => x"00000000", 31042 => x"00000000", 31043 => x"00000000",
    31044 => x"00000000", 31045 => x"00000000", 31046 => x"00000000",
    31047 => x"00000000", 31048 => x"00000000", 31049 => x"00000000",
    31050 => x"00000000", 31051 => x"00000000", 31052 => x"00000000",
    31053 => x"00000000", 31054 => x"00000000", 31055 => x"00000000",
    31056 => x"00000000", 31057 => x"00000000", 31058 => x"00000000",
    31059 => x"00000000", 31060 => x"00000000", 31061 => x"00000000",
    31062 => x"00000000", 31063 => x"00000000", 31064 => x"00000000",
    31065 => x"00000000", 31066 => x"00000000", 31067 => x"00000000",
    31068 => x"00000000", 31069 => x"00000000", 31070 => x"00000000",
    31071 => x"00000000", 31072 => x"00000000", 31073 => x"00000000",
    31074 => x"00000000", 31075 => x"00000000", 31076 => x"00000000",
    31077 => x"00000000", 31078 => x"00000000", 31079 => x"00000000",
    31080 => x"00000000", 31081 => x"00000000", 31082 => x"00000000",
    31083 => x"00000000", 31084 => x"00000000", 31085 => x"00000000",
    31086 => x"00000000", 31087 => x"00000000", 31088 => x"00000000",
    31089 => x"00000000", 31090 => x"00000000", 31091 => x"00000000",
    31092 => x"00000000", 31093 => x"00000000", 31094 => x"00000000",
    31095 => x"00000000", 31096 => x"00000000", 31097 => x"00000000",
    31098 => x"00000000", 31099 => x"00000000", 31100 => x"00000000",
    31101 => x"00000000", 31102 => x"00000000", 31103 => x"00000000",
    31104 => x"00000000", 31105 => x"00000000", 31106 => x"00000000",
    31107 => x"00000000", 31108 => x"00000000", 31109 => x"00000000",
    31110 => x"00000000", 31111 => x"00000000", 31112 => x"00000000",
    31113 => x"00000000", 31114 => x"00000000", 31115 => x"00000000",
    31116 => x"00000000", 31117 => x"00000000", 31118 => x"00000000",
    31119 => x"00000000", 31120 => x"00000000", 31121 => x"00000000",
    31122 => x"00000000", 31123 => x"00000000", 31124 => x"00000000",
    31125 => x"00000000", 31126 => x"00000000", 31127 => x"00000000",
    31128 => x"00000000", 31129 => x"00000000", 31130 => x"00000000",
    31131 => x"00000000", 31132 => x"00000000", 31133 => x"00000000",
    31134 => x"00000000", 31135 => x"00000000", 31136 => x"00000000",
    31137 => x"00000000", 31138 => x"00000000", 31139 => x"00000000",
    31140 => x"00000000", 31141 => x"00000000", 31142 => x"00000000",
    31143 => x"00000000", 31144 => x"00000000", 31145 => x"00000000",
    31146 => x"00000000", 31147 => x"00000000", 31148 => x"00000000",
    31149 => x"00000000", 31150 => x"00000000", 31151 => x"00000000",
    31152 => x"00000000", 31153 => x"00000000", 31154 => x"00000000",
    31155 => x"00000000", 31156 => x"00000000", 31157 => x"00000000",
    31158 => x"00000000", 31159 => x"00000000", 31160 => x"00000000",
    31161 => x"00000000", 31162 => x"00000000", 31163 => x"00000000",
    31164 => x"00000000", 31165 => x"00000000", 31166 => x"00000000",
    31167 => x"00000000", 31168 => x"00000000", 31169 => x"00000000",
    31170 => x"00000000", 31171 => x"00000000", 31172 => x"00000000",
    31173 => x"00000000", 31174 => x"00000000", 31175 => x"00000000",
    31176 => x"00000000", 31177 => x"00000000", 31178 => x"00000000",
    31179 => x"00000000", 31180 => x"00000000", 31181 => x"00000000",
    31182 => x"00000000", 31183 => x"00000000", 31184 => x"00000000",
    31185 => x"00000000", 31186 => x"00000000", 31187 => x"00000000",
    31188 => x"00000000", 31189 => x"00000000", 31190 => x"00000000",
    31191 => x"00000000", 31192 => x"00000000", 31193 => x"00000000",
    31194 => x"00000000", 31195 => x"00000000", 31196 => x"00000000",
    31197 => x"00000000", 31198 => x"00000000", 31199 => x"00000000",
    31200 => x"00000000", 31201 => x"00000000", 31202 => x"00000000",
    31203 => x"00000000", 31204 => x"00000000", 31205 => x"00000000",
    31206 => x"00000000", 31207 => x"00000000", 31208 => x"00000000",
    31209 => x"00000000", 31210 => x"00000000", 31211 => x"00000000",
    31212 => x"00000000", 31213 => x"00000000", 31214 => x"00000000",
    31215 => x"00000000", 31216 => x"00000000", 31217 => x"00000000",
    31218 => x"00000000", 31219 => x"00000000", 31220 => x"00000000",
    31221 => x"00000000", 31222 => x"00000000", 31223 => x"00000000",
    31224 => x"00000000", 31225 => x"00000000", 31226 => x"00000000",
    31227 => x"00000000", 31228 => x"00000000", 31229 => x"00000000",
    31230 => x"00000000", 31231 => x"00000000", 31232 => x"00000000",
    31233 => x"00000000", 31234 => x"00000000", 31235 => x"00000000",
    31236 => x"00000000", 31237 => x"00000000", 31238 => x"00000000",
    31239 => x"00000000", 31240 => x"00000000", 31241 => x"00000000",
    31242 => x"00000000", 31243 => x"00000000", 31244 => x"00000000",
    31245 => x"00000000", 31246 => x"00000000", 31247 => x"00000000",
    31248 => x"00000000", 31249 => x"00000000", 31250 => x"00000000",
    31251 => x"00000000", 31252 => x"00000000", 31253 => x"00000000",
    31254 => x"00000000", 31255 => x"00000000", 31256 => x"00000000",
    31257 => x"00000000", 31258 => x"00000000", 31259 => x"00000000",
    31260 => x"00000000", 31261 => x"00000000", 31262 => x"00000000",
    31263 => x"00000000", 31264 => x"00000000", 31265 => x"00000000",
    31266 => x"00000000", 31267 => x"00000000", 31268 => x"00000000",
    31269 => x"00000000", 31270 => x"00000000", 31271 => x"00000000",
    31272 => x"00000000", 31273 => x"00000000", 31274 => x"00000000",
    31275 => x"00000000", 31276 => x"00000000", 31277 => x"00000000",
    31278 => x"00000000", 31279 => x"00000000", 31280 => x"00000000",
    31281 => x"00000000", 31282 => x"00000000", 31283 => x"00000000",
    31284 => x"00000000", 31285 => x"00000000", 31286 => x"00000000",
    31287 => x"00000000", 31288 => x"00000000", 31289 => x"00000000",
    31290 => x"00000000", 31291 => x"00000000", 31292 => x"00000000",
    31293 => x"00000000", 31294 => x"00000000", 31295 => x"00000000",
    31296 => x"00000000", 31297 => x"00000000", 31298 => x"00000000",
    31299 => x"00000000", 31300 => x"00000000", 31301 => x"00000000",
    31302 => x"00000000", 31303 => x"00000000", 31304 => x"00000000",
    31305 => x"00000000", 31306 => x"00000000", 31307 => x"00000000",
    31308 => x"00000000", 31309 => x"00000000", 31310 => x"00000000",
    31311 => x"00000000", 31312 => x"00000000", 31313 => x"00000000",
    31314 => x"00000000", 31315 => x"00000000", 31316 => x"00000000",
    31317 => x"00000000", 31318 => x"00000000", 31319 => x"00000000",
    31320 => x"00000000", 31321 => x"00000000", 31322 => x"00000000",
    31323 => x"00000000", 31324 => x"00000000", 31325 => x"00000000",
    31326 => x"00000000", 31327 => x"00000000", 31328 => x"00000000",
    31329 => x"00000000", 31330 => x"00000000", 31331 => x"00000000",
    31332 => x"00000000", 31333 => x"00000000", 31334 => x"00000000",
    31335 => x"00000000", 31336 => x"00000000", 31337 => x"00000000",
    31338 => x"00000000", 31339 => x"00000000", 31340 => x"00000000",
    31341 => x"00000000", 31342 => x"00000000", 31343 => x"00000000",
    31344 => x"00000000", 31345 => x"00000000", 31346 => x"00000000",
    31347 => x"00000000", 31348 => x"00000000", 31349 => x"00000000",
    31350 => x"00000000", 31351 => x"00000000", 31352 => x"00000000",
    31353 => x"00000000", 31354 => x"00000000", 31355 => x"00000000",
    31356 => x"00000000", 31357 => x"00000000", 31358 => x"00000000",
    31359 => x"00000000", 31360 => x"00000000", 31361 => x"00000000",
    31362 => x"00000000", 31363 => x"00000000", 31364 => x"00000000",
    31365 => x"00000000", 31366 => x"00000000", 31367 => x"00000000",
    31368 => x"00000000", 31369 => x"00000000", 31370 => x"00000000",
    31371 => x"00000000", 31372 => x"00000000", 31373 => x"00000000",
    31374 => x"00000000", 31375 => x"00000000", 31376 => x"00000000",
    31377 => x"00000000", 31378 => x"00000000", 31379 => x"00000000",
    31380 => x"00000000", 31381 => x"00000000", 31382 => x"00000000",
    31383 => x"00000000", 31384 => x"00000000", 31385 => x"00000000",
    31386 => x"00000000", 31387 => x"00000000", 31388 => x"00000000",
    31389 => x"00000000", 31390 => x"00000000", 31391 => x"00000000",
    31392 => x"00000000", 31393 => x"00000000", 31394 => x"00000000",
    31395 => x"00000000", 31396 => x"00000000", 31397 => x"00000000",
    31398 => x"00000000", 31399 => x"00000000", 31400 => x"00000000",
    31401 => x"00000000", 31402 => x"00000000", 31403 => x"00000000",
    31404 => x"00000000", 31405 => x"00000000", 31406 => x"00000000",
    31407 => x"00000000", 31408 => x"00000000", 31409 => x"00000000",
    31410 => x"00000000", 31411 => x"00000000", 31412 => x"00000000",
    31413 => x"00000000", 31414 => x"00000000", 31415 => x"00000000",
    31416 => x"00000000", 31417 => x"00000000", 31418 => x"00000000",
    31419 => x"00000000", 31420 => x"00000000", 31421 => x"00000000",
    31422 => x"00000000", 31423 => x"00000000", 31424 => x"00000000",
    31425 => x"00000000", 31426 => x"00000000", 31427 => x"00000000",
    31428 => x"00000000", 31429 => x"00000000", 31430 => x"00000000",
    31431 => x"00000000", 31432 => x"00000000", 31433 => x"00000000",
    31434 => x"00000000", 31435 => x"00000000", 31436 => x"00000000",
    31437 => x"00000000", 31438 => x"00000000", 31439 => x"00000000",
    31440 => x"00000000", 31441 => x"00000000", 31442 => x"00000000",
    31443 => x"00000000", 31444 => x"00000000", 31445 => x"00000000",
    31446 => x"00000000", 31447 => x"00000000", 31448 => x"00000000",
    31449 => x"00000000", 31450 => x"00000000", 31451 => x"00000000",
    31452 => x"00000000", 31453 => x"00000000", 31454 => x"00000000",
    31455 => x"00000000", 31456 => x"00000000", 31457 => x"00000000",
    31458 => x"00000000", 31459 => x"00000000", 31460 => x"00000000",
    31461 => x"00000000", 31462 => x"00000000", 31463 => x"00000000",
    31464 => x"00000000", 31465 => x"00000000", 31466 => x"00000000",
    31467 => x"00000000", 31468 => x"00000000", 31469 => x"00000000",
    31470 => x"00000000", 31471 => x"00000000", 31472 => x"00000000",
    31473 => x"00000000", 31474 => x"00000000", 31475 => x"00000000",
    31476 => x"00000000", 31477 => x"00000000", 31478 => x"00000000",
    31479 => x"00000000", 31480 => x"00000000", 31481 => x"00000000",
    31482 => x"00000000", 31483 => x"00000000", 31484 => x"00000000",
    31485 => x"00000000", 31486 => x"00000000", 31487 => x"00000000",
    31488 => x"00000000", 31489 => x"00000000", 31490 => x"00000000",
    31491 => x"00000000", 31492 => x"00000000", 31493 => x"00000000",
    31494 => x"00000000", 31495 => x"00000000", 31496 => x"00000000",
    31497 => x"00000000", 31498 => x"00000000", 31499 => x"00000000",
    31500 => x"00000000", 31501 => x"00000000", 31502 => x"00000000",
    31503 => x"00000000", 31504 => x"00000000", 31505 => x"00000000",
    31506 => x"00000000", 31507 => x"00000000", 31508 => x"00000000",
    31509 => x"00000000", 31510 => x"00000000", 31511 => x"00000000",
    31512 => x"00000000", 31513 => x"00000000", 31514 => x"00000000",
    31515 => x"00000000", 31516 => x"00000000", 31517 => x"00000000",
    31518 => x"00000000", 31519 => x"00000000", 31520 => x"00000000",
    31521 => x"00000000", 31522 => x"00000000", 31523 => x"00000000",
    31524 => x"00000000", 31525 => x"00000000", 31526 => x"00000000",
    31527 => x"00000000", 31528 => x"00000000", 31529 => x"00000000",
    31530 => x"00000000", 31531 => x"00000000", 31532 => x"00000000",
    31533 => x"00000000", 31534 => x"00000000", 31535 => x"00000000",
    31536 => x"00000000", 31537 => x"00000000", 31538 => x"00000000",
    31539 => x"00000000", 31540 => x"00000000", 31541 => x"00000000",
    31542 => x"00000000", 31543 => x"00000000", 31544 => x"00000000",
    31545 => x"00000000", 31546 => x"00000000", 31547 => x"00000000",
    31548 => x"00000000", 31549 => x"00000000", 31550 => x"00000000",
    31551 => x"00000000", 31552 => x"00000000", 31553 => x"00000000",
    31554 => x"00000000", 31555 => x"00000000", 31556 => x"00000000",
    31557 => x"00000000", 31558 => x"00000000", 31559 => x"00000000",
    31560 => x"00000000", 31561 => x"00000000", 31562 => x"00000000",
    31563 => x"00000000", 31564 => x"00000000", 31565 => x"00000000",
    31566 => x"00000000", 31567 => x"00000000", 31568 => x"00000000",
    31569 => x"00000000", 31570 => x"00000000", 31571 => x"00000000",
    31572 => x"00000000", 31573 => x"00000000", 31574 => x"00000000",
    31575 => x"00000000", 31576 => x"00000000", 31577 => x"00000000",
    31578 => x"00000000", 31579 => x"00000000", 31580 => x"00000000",
    31581 => x"00000000", 31582 => x"00000000", 31583 => x"00000000",
    31584 => x"00000000", 31585 => x"00000000", 31586 => x"00000000",
    31587 => x"00000000", 31588 => x"00000000", 31589 => x"00000000",
    31590 => x"00000000", 31591 => x"00000000", 31592 => x"00000000",
    31593 => x"00000000", 31594 => x"00000000", 31595 => x"00000000",
    31596 => x"00000000", 31597 => x"00000000", 31598 => x"00000000",
    31599 => x"00000000", 31600 => x"00000000", 31601 => x"00000000",
    31602 => x"00000000", 31603 => x"00000000", 31604 => x"00000000",
    31605 => x"00000000", 31606 => x"00000000", 31607 => x"00000000",
    31608 => x"00000000", 31609 => x"00000000", 31610 => x"00000000",
    31611 => x"00000000", 31612 => x"00000000", 31613 => x"00000000",
    31614 => x"00000000", 31615 => x"00000000", 31616 => x"00000000",
    31617 => x"00000000", 31618 => x"00000000", 31619 => x"00000000",
    31620 => x"00000000", 31621 => x"00000000", 31622 => x"00000000",
    31623 => x"00000000", 31624 => x"00000000", 31625 => x"00000000",
    31626 => x"00000000", 31627 => x"00000000", 31628 => x"00000000",
    31629 => x"00000000", 31630 => x"00000000", 31631 => x"00000000",
    31632 => x"00000000", 31633 => x"00000000", 31634 => x"00000000",
    31635 => x"00000000", 31636 => x"00000000", 31637 => x"00000000",
    31638 => x"00000000", 31639 => x"00000000", 31640 => x"00000000",
    31641 => x"00000000", 31642 => x"00000000", 31643 => x"00000000",
    31644 => x"00000000", 31645 => x"00000000", 31646 => x"00000000",
    31647 => x"00000000", 31648 => x"00000000", 31649 => x"00000000",
    31650 => x"00000000", 31651 => x"00000000", 31652 => x"00000000",
    31653 => x"00000000", 31654 => x"00000000", 31655 => x"00000000",
    31656 => x"00000000", 31657 => x"00000000", 31658 => x"00000000",
    31659 => x"00000000", 31660 => x"00000000", 31661 => x"00000000",
    31662 => x"00000000", 31663 => x"00000000", 31664 => x"00000000",
    31665 => x"00000000", 31666 => x"00000000", 31667 => x"00000000",
    31668 => x"00000000", 31669 => x"00000000", 31670 => x"00000000",
    31671 => x"00000000", 31672 => x"00000000", 31673 => x"00000000",
    31674 => x"00000000", 31675 => x"00000000", 31676 => x"00000000",
    31677 => x"00000000", 31678 => x"00000000", 31679 => x"00000000",
    31680 => x"00000000", 31681 => x"00000000", 31682 => x"00000000",
    31683 => x"00000000", 31684 => x"00000000", 31685 => x"00000000",
    31686 => x"00000000", 31687 => x"00000000", 31688 => x"00000000",
    31689 => x"00000000", 31690 => x"00000000", 31691 => x"00000000",
    31692 => x"00000000", 31693 => x"00000000", 31694 => x"00000000",
    31695 => x"00000000", 31696 => x"00000000", 31697 => x"00000000",
    31698 => x"00000000", 31699 => x"00000000", 31700 => x"00000000",
    31701 => x"00000000", 31702 => x"00000000", 31703 => x"00000000",
    31704 => x"00000000", 31705 => x"00000000", 31706 => x"00000000",
    31707 => x"00000000", 31708 => x"00000000", 31709 => x"00000000",
    31710 => x"00000000", 31711 => x"00000000", 31712 => x"00000000",
    31713 => x"00000000", 31714 => x"00000000", 31715 => x"00000000",
    31716 => x"00000000", 31717 => x"00000000", 31718 => x"00000000",
    31719 => x"00000000", 31720 => x"00000000", 31721 => x"00000000",
    31722 => x"00000000", 31723 => x"00000000", 31724 => x"00000000",
    31725 => x"00000000", 31726 => x"00000000", 31727 => x"00000000",
    31728 => x"00000000", 31729 => x"00000000", 31730 => x"00000000",
    31731 => x"00000000", 31732 => x"00000000", 31733 => x"00000000",
    31734 => x"00000000", 31735 => x"00000000", 31736 => x"00000000",
    31737 => x"00000000", 31738 => x"00000000", 31739 => x"00000000",
    31740 => x"00000000", 31741 => x"00000000", 31742 => x"00000000",
    31743 => x"00000000", 31744 => x"00000000", 31745 => x"00000000",
    31746 => x"00000000", 31747 => x"00000000", 31748 => x"00000000",
    31749 => x"00000000", 31750 => x"00000000", 31751 => x"00000000",
    31752 => x"00000000", 31753 => x"00000000", 31754 => x"00000000",
    31755 => x"00000000", 31756 => x"00000000", 31757 => x"00000000",
    31758 => x"00000000", 31759 => x"00000000", 31760 => x"00000000",
    31761 => x"00000000", 31762 => x"00000000", 31763 => x"00000000",
    31764 => x"00000000", 31765 => x"00000000", 31766 => x"00000000",
    31767 => x"00000000", 31768 => x"00000000", 31769 => x"00000000",
    31770 => x"00000000", 31771 => x"00000000", 31772 => x"00000000",
    31773 => x"00000000", 31774 => x"00000000", 31775 => x"00000000",
    31776 => x"00000000", 31777 => x"00000000", 31778 => x"00000000",
    31779 => x"00000000", 31780 => x"00000000", 31781 => x"00000000",
    31782 => x"00000000", 31783 => x"00000000", 31784 => x"00000000",
    31785 => x"00000000", 31786 => x"00000000", 31787 => x"00000000",
    31788 => x"00000000", 31789 => x"00000000", 31790 => x"00000000",
    31791 => x"00000000", 31792 => x"00000000", 31793 => x"00000000",
    31794 => x"00000000", 31795 => x"00000000", 31796 => x"00000000",
    31797 => x"00000000", 31798 => x"00000000", 31799 => x"00000000",
    31800 => x"00000000", 31801 => x"00000000", 31802 => x"00000000",
    31803 => x"00000000", 31804 => x"00000000", 31805 => x"00000000",
    31806 => x"00000000", 31807 => x"00000000", 31808 => x"00000000",
    31809 => x"00000000", 31810 => x"00000000", 31811 => x"00000000",
    31812 => x"00000000", 31813 => x"00000000", 31814 => x"00000000",
    31815 => x"00000000", 31816 => x"00000000", 31817 => x"00000000",
    31818 => x"00000000", 31819 => x"00000000", 31820 => x"00000000",
    31821 => x"00000000", 31822 => x"00000000", 31823 => x"00000000",
    31824 => x"00000000", 31825 => x"00000000", 31826 => x"00000000",
    31827 => x"00000000", 31828 => x"00000000", 31829 => x"00000000",
    31830 => x"00000000", 31831 => x"00000000", 31832 => x"00000000",
    31833 => x"00000000", 31834 => x"00000000", 31835 => x"00000000",
    31836 => x"00000000", 31837 => x"00000000", 31838 => x"00000000",
    31839 => x"00000000", 31840 => x"00000000", 31841 => x"00000000",
    31842 => x"00000000", 31843 => x"00000000", 31844 => x"00000000",
    31845 => x"00000000", 31846 => x"00000000", 31847 => x"00000000",
    31848 => x"00000000", 31849 => x"00000000", 31850 => x"00000000",
    31851 => x"00000000", 31852 => x"00000000", 31853 => x"00000000",
    31854 => x"00000000", 31855 => x"00000000", 31856 => x"00000000",
    31857 => x"00000000", 31858 => x"00000000", 31859 => x"00000000",
    31860 => x"00000000", 31861 => x"00000000", 31862 => x"00000000",
    31863 => x"00000000", 31864 => x"00000000", 31865 => x"00000000",
    31866 => x"00000000", 31867 => x"00000000", 31868 => x"00000000",
    31869 => x"00000000", 31870 => x"00000000", 31871 => x"00000000",
    31872 => x"00000000", 31873 => x"00000000", 31874 => x"00000000",
    31875 => x"00000000", 31876 => x"00000000", 31877 => x"00000000",
    31878 => x"00000000", 31879 => x"00000000", 31880 => x"00000000",
    31881 => x"00000000", 31882 => x"00000000", 31883 => x"00000000",
    31884 => x"00000000", 31885 => x"00000000", 31886 => x"00000000",
    31887 => x"00000000", 31888 => x"00000000", 31889 => x"00000000",
    31890 => x"00000000", 31891 => x"00000000", 31892 => x"00000000",
    31893 => x"00000000", 31894 => x"00000000", 31895 => x"00000000",
    31896 => x"00000000", 31897 => x"00000000", 31898 => x"00000000",
    31899 => x"00000000", 31900 => x"00000000", 31901 => x"00000000",
    31902 => x"00000000", 31903 => x"00000000", 31904 => x"00000000",
    31905 => x"00000000", 31906 => x"00000000", 31907 => x"00000000",
    31908 => x"00000000", 31909 => x"00000000", 31910 => x"00000000",
    31911 => x"00000000", 31912 => x"00000000", 31913 => x"00000000",
    31914 => x"00000000", 31915 => x"00000000", 31916 => x"00000000",
    31917 => x"00000000", 31918 => x"00000000", 31919 => x"00000000",
    31920 => x"00000000", 31921 => x"00000000", 31922 => x"00000000",
    31923 => x"00000000", 31924 => x"00000000", 31925 => x"00000000",
    31926 => x"00000000", 31927 => x"00000000", 31928 => x"00000000",
    31929 => x"00000000", 31930 => x"00000000", 31931 => x"00000000",
    31932 => x"00000000", 31933 => x"00000000", 31934 => x"00000000",
    31935 => x"00000000", 31936 => x"00000000", 31937 => x"00000000",
    31938 => x"00000000", 31939 => x"00000000", 31940 => x"00000000",
    31941 => x"00000000", 31942 => x"00000000", 31943 => x"00000000",
    31944 => x"00000000", 31945 => x"00000000", 31946 => x"00000000",
    31947 => x"00000000", 31948 => x"00000000", 31949 => x"00000000",
    31950 => x"00000000", 31951 => x"00000000", 31952 => x"00000000",
    31953 => x"00000000", 31954 => x"00000000", 31955 => x"00000000",
    31956 => x"00000000", 31957 => x"00000000", 31958 => x"00000000",
    31959 => x"00000000", 31960 => x"00000000", 31961 => x"00000000",
    31962 => x"00000000", 31963 => x"00000000", 31964 => x"00000000",
    31965 => x"00000000", 31966 => x"00000000", 31967 => x"00000000",
    31968 => x"00000000", 31969 => x"00000000", 31970 => x"00000000",
    31971 => x"00000000", 31972 => x"00000000", 31973 => x"00000000",
    31974 => x"00000000", 31975 => x"00000000", 31976 => x"00000000",
    31977 => x"00000000", 31978 => x"00000000", 31979 => x"00000000",
    31980 => x"00000000", 31981 => x"00000000", 31982 => x"00000000",
    31983 => x"00000000", 31984 => x"00000000", 31985 => x"00000000",
    31986 => x"00000000", 31987 => x"00000000", 31988 => x"00000000",
    31989 => x"00000000", 31990 => x"00000000", 31991 => x"00000000",
    31992 => x"00000000", 31993 => x"00000000", 31994 => x"00000000",
    31995 => x"00000000", 31996 => x"00000000", 31997 => x"00000000",
    31998 => x"00000000", 31999 => x"00000000", 32000 => x"00000000",
    32001 => x"00000000", 32002 => x"00000000", 32003 => x"00000000",
    32004 => x"00000000", 32005 => x"00000000", 32006 => x"00000000",
    32007 => x"00000000", 32008 => x"00000000", 32009 => x"00000000",
    32010 => x"00000000", 32011 => x"00000000", 32012 => x"00000000",
    32013 => x"00000000", 32014 => x"00000000", 32015 => x"00000000",
    32016 => x"00000000", 32017 => x"00000000", 32018 => x"00000000",
    32019 => x"00000000", 32020 => x"00000000", 32021 => x"00000000",
    32022 => x"00000000", 32023 => x"00000000", 32024 => x"00000000",
    32025 => x"00000000", 32026 => x"00000000", 32027 => x"00000000",
    32028 => x"00000000", 32029 => x"00000000", 32030 => x"00000000",
    32031 => x"00000000", 32032 => x"00000000", 32033 => x"00000000",
    32034 => x"00000000", 32035 => x"00000000", 32036 => x"00000000",
    32037 => x"00000000", 32038 => x"00000000", 32039 => x"00000000",
    32040 => x"00000000", 32041 => x"00000000", 32042 => x"00000000",
    32043 => x"00000000", 32044 => x"00000000", 32045 => x"00000000",
    32046 => x"00000000", 32047 => x"00000000", 32048 => x"00000000",
    32049 => x"00000000", 32050 => x"00000000", 32051 => x"00000000",
    32052 => x"00000000", 32053 => x"00000000", 32054 => x"00000000",
    32055 => x"00000000", 32056 => x"00000000", 32057 => x"00000000",
    32058 => x"00000000", 32059 => x"00000000", 32060 => x"00000000",
    32061 => x"00000000", 32062 => x"00000000", 32063 => x"00000000",
    32064 => x"00000000", 32065 => x"00000000", 32066 => x"00000000",
    32067 => x"00000000", 32068 => x"00000000", 32069 => x"00000000",
    32070 => x"00000000", 32071 => x"00000000", 32072 => x"00000000",
    32073 => x"00000000", 32074 => x"00000000", 32075 => x"00000000",
    32076 => x"00000000", 32077 => x"00000000", 32078 => x"00000000",
    32079 => x"00000000", 32080 => x"00000000", 32081 => x"00000000",
    32082 => x"00000000", 32083 => x"00000000", 32084 => x"00000000",
    32085 => x"00000000", 32086 => x"00000000", 32087 => x"00000000",
    32088 => x"00000000", 32089 => x"00000000", 32090 => x"00000000",
    32091 => x"00000000", 32092 => x"00000000", 32093 => x"00000000",
    32094 => x"00000000", 32095 => x"00000000", 32096 => x"00000000",
    32097 => x"00000000", 32098 => x"00000000", 32099 => x"00000000",
    32100 => x"00000000", 32101 => x"00000000", 32102 => x"00000000",
    32103 => x"00000000", 32104 => x"00000000", 32105 => x"00000000",
    32106 => x"00000000", 32107 => x"00000000", 32108 => x"00000000",
    32109 => x"00000000", 32110 => x"00000000", 32111 => x"00000000",
    32112 => x"00000000", 32113 => x"00000000", 32114 => x"00000000",
    32115 => x"00000000", 32116 => x"00000000", 32117 => x"00000000",
    32118 => x"00000000", 32119 => x"00000000", 32120 => x"00000000",
    32121 => x"00000000", 32122 => x"00000000", 32123 => x"00000000",
    32124 => x"00000000", 32125 => x"00000000", 32126 => x"00000000",
    32127 => x"00000000", 32128 => x"00000000", 32129 => x"00000000",
    32130 => x"00000000", 32131 => x"00000000", 32132 => x"00000000",
    32133 => x"00000000", 32134 => x"00000000", 32135 => x"00000000",
    32136 => x"00000000", 32137 => x"00000000", 32138 => x"00000000",
    32139 => x"00000000", 32140 => x"00000000", 32141 => x"00000000",
    32142 => x"00000000", 32143 => x"00000000", 32144 => x"00000000",
    32145 => x"00000000", 32146 => x"00000000", 32147 => x"00000000",
    32148 => x"00000000", 32149 => x"00000000", 32150 => x"00000000",
    32151 => x"00000000", 32152 => x"00000000", 32153 => x"00000000",
    32154 => x"00000000", 32155 => x"00000000", 32156 => x"00000000",
    32157 => x"00000000", 32158 => x"00000000", 32159 => x"00000000",
    32160 => x"00000000", 32161 => x"00000000", 32162 => x"00000000",
    32163 => x"00000000", 32164 => x"00000000", 32165 => x"00000000",
    32166 => x"00000000", 32167 => x"00000000", 32168 => x"00000000",
    32169 => x"00000000", 32170 => x"00000000", 32171 => x"00000000",
    32172 => x"00000000", 32173 => x"00000000", 32174 => x"00000000",
    32175 => x"00000000", 32176 => x"00000000", 32177 => x"00000000",
    32178 => x"00000000", 32179 => x"00000000", 32180 => x"00000000",
    32181 => x"00000000", 32182 => x"00000000", 32183 => x"00000000",
    32184 => x"00000000", 32185 => x"00000000", 32186 => x"00000000",
    32187 => x"00000000", 32188 => x"00000000", 32189 => x"00000000",
    32190 => x"00000000", 32191 => x"00000000", 32192 => x"00000000",
    32193 => x"00000000", 32194 => x"00000000", 32195 => x"00000000",
    32196 => x"00000000", 32197 => x"00000000", 32198 => x"00000000",
    32199 => x"00000000", 32200 => x"00000000", 32201 => x"00000000",
    32202 => x"00000000", 32203 => x"00000000", 32204 => x"00000000",
    32205 => x"00000000", 32206 => x"00000000", 32207 => x"00000000",
    32208 => x"00000000", 32209 => x"00000000", 32210 => x"00000000",
    32211 => x"00000000", 32212 => x"00000000", 32213 => x"00000000",
    32214 => x"00000000", 32215 => x"00000000", 32216 => x"00000000",
    32217 => x"00000000", 32218 => x"00000000", 32219 => x"00000000",
    32220 => x"00000000", 32221 => x"00000000", 32222 => x"00000000",
    32223 => x"00000000", 32224 => x"00000000", 32225 => x"00000000",
    32226 => x"00000000", 32227 => x"00000000", 32228 => x"00000000",
    32229 => x"00000000", 32230 => x"00000000", 32231 => x"00000000",
    32232 => x"00000000", 32233 => x"00000000", 32234 => x"00000000",
    32235 => x"00000000", 32236 => x"00000000", 32237 => x"00000000",
    32238 => x"00000000", 32239 => x"00000000", 32240 => x"00000000",
    32241 => x"00000000", 32242 => x"00000000", 32243 => x"00000000",
    32244 => x"00000000", 32245 => x"00000000", 32246 => x"00000000",
    32247 => x"00000000", 32248 => x"00000000", 32249 => x"00000000",
    32250 => x"00000000", 32251 => x"00000000", 32252 => x"00000000",
    32253 => x"00000000", 32254 => x"00000000", 32255 => x"00000000",
    32256 => x"00000000", 32257 => x"00000000", 32258 => x"00000000",
    32259 => x"00000000", 32260 => x"00000000", 32261 => x"00000000",
    32262 => x"00000000", 32263 => x"00000000", 32264 => x"00000000",
    32265 => x"00000000", 32266 => x"00000000", 32267 => x"00000000",
    32268 => x"00000000", 32269 => x"00000000", 32270 => x"00000000",
    32271 => x"00000000", 32272 => x"00000000", 32273 => x"00000000",
    32274 => x"00000000", 32275 => x"00000000", 32276 => x"00000000",
    32277 => x"00000000", 32278 => x"00000000", 32279 => x"00000000",
    32280 => x"00000000", 32281 => x"00000000", 32282 => x"00000000",
    32283 => x"00000000", 32284 => x"00000000", 32285 => x"00000000",
    32286 => x"00000000", 32287 => x"00000000", 32288 => x"00000000",
    32289 => x"00000000", 32290 => x"00000000", 32291 => x"00000000",
    32292 => x"00000000", 32293 => x"00000000", 32294 => x"00000000",
    32295 => x"00000000", 32296 => x"00000000", 32297 => x"00000000",
    32298 => x"00000000", 32299 => x"00000000", 32300 => x"00000000",
    32301 => x"00000000", 32302 => x"00000000", 32303 => x"00000000",
    32304 => x"00000000", 32305 => x"00000000", 32306 => x"00000000",
    32307 => x"00000000", 32308 => x"00000000", 32309 => x"00000000",
    32310 => x"00000000", 32311 => x"00000000", 32312 => x"00000000",
    32313 => x"00000000", 32314 => x"00000000", 32315 => x"00000000",
    32316 => x"00000000", 32317 => x"00000000", 32318 => x"00000000",
    32319 => x"00000000", 32320 => x"00000000", 32321 => x"00000000",
    32322 => x"00000000", 32323 => x"00000000", 32324 => x"00000000",
    32325 => x"00000000", 32326 => x"00000000", 32327 => x"00000000",
    32328 => x"00000000", 32329 => x"00000000", 32330 => x"00000000",
    32331 => x"00000000", 32332 => x"00000000", 32333 => x"00000000",
    32334 => x"00000000", 32335 => x"00000000", 32336 => x"00000000",
    32337 => x"00000000", 32338 => x"00000000", 32339 => x"00000000",
    32340 => x"00000000", 32341 => x"00000000", 32342 => x"00000000",
    32343 => x"00000000", 32344 => x"00000000", 32345 => x"00000000",
    32346 => x"00000000", 32347 => x"00000000", 32348 => x"00000000",
    32349 => x"00000000", 32350 => x"00000000", 32351 => x"00000000",
    32352 => x"00000000", 32353 => x"00000000", 32354 => x"00000000",
    32355 => x"00000000", 32356 => x"00000000", 32357 => x"00000000",
    32358 => x"00000000", 32359 => x"00000000", 32360 => x"00000000",
    32361 => x"00000000", 32362 => x"00000000", 32363 => x"00000000",
    32364 => x"00000000", 32365 => x"00000000", 32366 => x"00000000",
    32367 => x"00000000", 32368 => x"00000000", 32369 => x"00000000",
    32370 => x"00000000", 32371 => x"00000000", 32372 => x"00000000",
    32373 => x"00000000", 32374 => x"00000000", 32375 => x"00000000",
    32376 => x"00000000", 32377 => x"00000000", 32378 => x"00000000",
    32379 => x"00000000", 32380 => x"00000000", 32381 => x"00000000",
    32382 => x"00000000", 32383 => x"00000000", 32384 => x"00000000",
    32385 => x"00000000", 32386 => x"00000000", 32387 => x"00000000",
    32388 => x"00000000", 32389 => x"00000000", 32390 => x"00000000",
    32391 => x"00000000", 32392 => x"00000000", 32393 => x"00000000",
    32394 => x"00000000", 32395 => x"00000000", 32396 => x"00000000",
    32397 => x"00000000", 32398 => x"00000000", 32399 => x"00000000",
    32400 => x"00000000", 32401 => x"00000000", 32402 => x"00000000",
    32403 => x"00000000", 32404 => x"00000000", 32405 => x"00000000",
    32406 => x"00000000", 32407 => x"00000000", 32408 => x"00000000",
    32409 => x"00000000", 32410 => x"00000000", 32411 => x"00000000",
    32412 => x"00000000", 32413 => x"00000000", 32414 => x"00000000",
    32415 => x"00000000", 32416 => x"00000000", 32417 => x"00000000",
    32418 => x"00000000", 32419 => x"00000000", 32420 => x"00000000",
    32421 => x"00000000", 32422 => x"00000000", 32423 => x"00000000",
    32424 => x"00000000", 32425 => x"00000000", 32426 => x"00000000",
    32427 => x"00000000", 32428 => x"00000000", 32429 => x"00000000",
    32430 => x"00000000", 32431 => x"00000000", 32432 => x"00000000",
    32433 => x"00000000", 32434 => x"00000000", 32435 => x"00000000",
    32436 => x"00000000", 32437 => x"00000000", 32438 => x"00000000",
    32439 => x"00000000", 32440 => x"00000000", 32441 => x"00000000",
    32442 => x"00000000", 32443 => x"00000000", 32444 => x"00000000",
    32445 => x"00000000", 32446 => x"00000000", 32447 => x"00000000",
    32448 => x"00000000", 32449 => x"00000000", 32450 => x"00000000",
    32451 => x"00000000", 32452 => x"00000000", 32453 => x"00000000",
    32454 => x"00000000", 32455 => x"00000000", 32456 => x"00000000",
    32457 => x"00000000", 32458 => x"00000000", 32459 => x"00000000",
    32460 => x"00000000", 32461 => x"00000000", 32462 => x"00000000",
    32463 => x"00000000", 32464 => x"00000000", 32465 => x"00000000",
    32466 => x"00000000", 32467 => x"00000000", 32468 => x"00000000",
    32469 => x"00000000", 32470 => x"00000000", 32471 => x"00000000",
    32472 => x"00000000", 32473 => x"00000000", 32474 => x"00000000",
    32475 => x"00000000", 32476 => x"00000000", 32477 => x"00000000",
    32478 => x"00000000", 32479 => x"00000000", 32480 => x"00000000",
    32481 => x"00000000", 32482 => x"00000000", 32483 => x"00000000",
    32484 => x"00000000", 32485 => x"00000000", 32486 => x"00000000",
    32487 => x"00000000", 32488 => x"00000000", 32489 => x"00000000",
    32490 => x"00000000", 32491 => x"00000000", 32492 => x"00000000",
    32493 => x"00000000", 32494 => x"00000000", 32495 => x"00000000",
    32496 => x"00000000", 32497 => x"00000000", 32498 => x"00000000",
    32499 => x"00000000", 32500 => x"00000000", 32501 => x"00000000",
    32502 => x"00000000", 32503 => x"00000000", 32504 => x"00000000",
    32505 => x"00000000", 32506 => x"00000000", 32507 => x"00000000",
    32508 => x"00000000", 32509 => x"00000000", 32510 => x"00000000",
    32511 => x"00000000", 32512 => x"00000000", 32513 => x"00000000",
    32514 => x"00000000", 32515 => x"00000000", 32516 => x"00000000",
    32517 => x"00000000", 32518 => x"00000000", 32519 => x"00000000",
    32520 => x"00000000", 32521 => x"00000000", 32522 => x"00000000",
    32523 => x"00000000", 32524 => x"00000000", 32525 => x"00000000",
    32526 => x"00000000", 32527 => x"00000000", 32528 => x"00000000",
    32529 => x"00000000", 32530 => x"00000000", 32531 => x"00000000",
    32532 => x"00000000", 32533 => x"00000000", 32534 => x"00000000",
    32535 => x"00000000", 32536 => x"00000000", 32537 => x"00000000",
    32538 => x"00000000", 32539 => x"00000000", 32540 => x"00000000",
    32541 => x"00000000", 32542 => x"00000000", 32543 => x"00000000",
    32544 => x"00000000", 32545 => x"00000000", 32546 => x"00000000",
    32547 => x"00000000", 32548 => x"00000000", 32549 => x"00000000",
    32550 => x"00000000", 32551 => x"00000000", 32552 => x"00000000",
    32553 => x"00000000", 32554 => x"00000000", 32555 => x"00000000",
    32556 => x"00000000", 32557 => x"00000000", 32558 => x"00000000",
    32559 => x"00000000", 32560 => x"00000000", 32561 => x"00000000",
    32562 => x"00000000", 32563 => x"00000000", 32564 => x"00000000",
    32565 => x"00000000", 32566 => x"00000000", 32567 => x"00000000",
    32568 => x"00000000", 32569 => x"00000000", 32570 => x"00000000",
    32571 => x"00000000", 32572 => x"00000000", 32573 => x"00000000",
    32574 => x"00000000", 32575 => x"00000000", 32576 => x"00000000",
    32577 => x"00000000", 32578 => x"00000000", 32579 => x"00000000",
    32580 => x"00000000", 32581 => x"00000000", 32582 => x"00000000",
    32583 => x"00000000", 32584 => x"00000000", 32585 => x"00000000",
    32586 => x"00000000", 32587 => x"00000000", 32588 => x"00000000",
    32589 => x"00000000", 32590 => x"00000000", 32591 => x"00000000",
    32592 => x"00000000", 32593 => x"00000000", 32594 => x"00000000",
    32595 => x"00000000", 32596 => x"00000000", 32597 => x"00000000",
    32598 => x"00000000", 32599 => x"00000000", 32600 => x"00000000",
    32601 => x"00000000", 32602 => x"00000000", 32603 => x"00000000",
    32604 => x"00000000", 32605 => x"00000000", 32606 => x"00000000",
    32607 => x"00000000", 32608 => x"00000000", 32609 => x"00000000",
    32610 => x"00000000", 32611 => x"00000000", 32612 => x"00000000",
    32613 => x"00000000", 32614 => x"00000000", 32615 => x"00000000",
    32616 => x"00000000", 32617 => x"00000000", 32618 => x"00000000",
    32619 => x"00000000", 32620 => x"00000000", 32621 => x"00000000",
    32622 => x"00000000", 32623 => x"00000000", 32624 => x"00000000",
    32625 => x"00000000", 32626 => x"00000000", 32627 => x"00000000",
    32628 => x"00000000", 32629 => x"00000000", 32630 => x"00000000",
    32631 => x"00000000", 32632 => x"00000000", 32633 => x"00000000",
    32634 => x"00000000", 32635 => x"00000000", 32636 => x"00000000",
    32637 => x"00000000", 32638 => x"00000000", 32639 => x"00000000",
    32640 => x"00000000", 32641 => x"00000000", 32642 => x"00000000",
    32643 => x"00000000", 32644 => x"00000000", 32645 => x"00000000",
    32646 => x"00000000", 32647 => x"00000000", 32648 => x"00000000",
    32649 => x"00000000", 32650 => x"00000000", 32651 => x"00000000",
    32652 => x"00000000", 32653 => x"00000000", 32654 => x"00000000",
    32655 => x"00000000", 32656 => x"00000000", 32657 => x"00000000",
    32658 => x"00000000", 32659 => x"00000000", 32660 => x"00000000",
    32661 => x"00000000", 32662 => x"00000000", 32663 => x"00000000",
    32664 => x"00000000", 32665 => x"00000000", 32666 => x"00000000",
    32667 => x"00000000", 32668 => x"00000000", 32669 => x"00000000",
    32670 => x"00000000", 32671 => x"00000000", 32672 => x"00000000",
    32673 => x"00000000", 32674 => x"00000000", 32675 => x"00000000",
    32676 => x"00000000", 32677 => x"00000000", 32678 => x"00000000",
    32679 => x"00000000", 32680 => x"00000000", 32681 => x"00000000",
    32682 => x"00000000", 32683 => x"00000000", 32684 => x"00000000",
    32685 => x"00000000", 32686 => x"00000000", 32687 => x"00000000",
    32688 => x"00000000", 32689 => x"00000000", 32690 => x"00000000",
    32691 => x"00000000", 32692 => x"00000000", 32693 => x"00000000",
    32694 => x"00000000", 32695 => x"00000000", 32696 => x"00000000",
    32697 => x"00000000", 32698 => x"00000000", 32699 => x"00000000",
    32700 => x"00000000", 32701 => x"00000000", 32702 => x"00000000",
    32703 => x"00000000", 32704 => x"00000000", 32705 => x"00000000",
    32706 => x"00000000", 32707 => x"00000000", 32708 => x"00000000",
    32709 => x"00000000", 32710 => x"00000000", 32711 => x"00000000",
    32712 => x"00000000", 32713 => x"00000000", 32714 => x"00000000",
    32715 => x"00000000", 32716 => x"00000000", 32717 => x"00000000",
    32718 => x"00000000", 32719 => x"00000000", 32720 => x"00000000",
    32721 => x"00000000", 32722 => x"00000000", 32723 => x"00000000",
    32724 => x"00000000", 32725 => x"00000000", 32726 => x"00000000",
    32727 => x"00000000", 32728 => x"00000000", 32729 => x"00000000",
    32730 => x"00000000", 32731 => x"00000000", 32732 => x"00000000",
    32733 => x"00000000", 32734 => x"00000000", 32735 => x"00000000",
    32736 => x"00000000", 32737 => x"00000000", 32738 => x"00000000",
    32739 => x"00000000", 32740 => x"00000000", 32741 => x"00000000",
    32742 => x"00000000", 32743 => x"00000000", 32744 => x"00000000",
    32745 => x"00000000", 32746 => x"00000000", 32747 => x"00000000",
    32748 => x"00000000", 32749 => x"00000000", 32750 => x"00000000",
    32751 => x"00000000", 32752 => x"00000000", 32753 => x"00000000",
    32754 => x"00000000", 32755 => x"00000000", 32756 => x"00000000",
    32757 => x"00000000", 32758 => x"00000000", 32759 => x"00000000",
    32760 => x"00000000", 32761 => x"00000000", 32762 => x"00000000",
    32763 => x"00000000", 32764 => x"00000000", 32765 => x"00000000",
    32766 => x"00000000", 32767 => x"00000000");
end wrc_bin_pkg;

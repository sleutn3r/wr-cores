// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
POPle66HqaoOXQZ3DKTqT4p8NcOE204ogvyCSnK1YUt9YpOhwdRcU3bntmQJb2nJ
0tiC/hCRkazZhsbIEiI/6IX085SA2dPk5G2RMNiQ4UthgEHWfAg8aNXDD57MBD8B
dE+t6o5deScd8ho7QkhT76UfnYNAcBZPEDa6Jlbmkpc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3712)
Sw5HM0AJ1aXg8aDQSLCceeqjaA3lUBCFrX/KHWMEsOgSsx0BHPz7x0KMJthjTUEq
JEaSElgVXbJ6XVWih9v2SpxtuoZedTvlRxgkOvTW4GnDvq3onNOrstHaaTmNW2zp
dpNFkyZPo0XTJ6BXhAOdffn+4Lrw3/Ouc+xvYSGdcPtj5Q4Ye0yPuSsh0YOL+By3
7whoHVlGrQdbLYPlaQvrNUzDl/OcyMmXsm+8wtaB18+/EB83CLJJ3p5x9SY1BHiF
ymeVSfGbQw4LEBkzIHP4EBD30XViRhjivxIkUNJVzgIGqf3hOlHE6xi1VVjq5ibS
VZf7ujhPyPYgp1iC/RavdTaLtdPJ/agQJTa1BjapvfnR+1J03E/Y2zswV4pml5M6
N+yPPaB+xtQ1iHYo9GZD3ikqQ/U62GYdK36/IaJDXgM0z63CtOW3vw4vUceglud9
OUE+HaLbhvBabYGp901x2nSyISQ+0zYehmkzs2m3OC/w/BysDqMbu5q6RDo8GGlz
Dj0yfRBeUWXq09FZXC/PQkMZAYkGp02/jURxCv6+pA+D9UKVJHlAYKIllnj+V/BD
5vaIQnj4jdi0iPpdCMiqBkKNt8ENLllQyO6+Ll5XBy+9XS3WA6u/uzjU9nf7UVv5
C+p99tlGpVhq1uowG7uIusF+lztMSbXwphYmN4zVx8npdFNzn1HAcqmOVhOQ2T4d
1Hy6xaD5sg/DcakPxPnSIKzJTbM87jXxHFCVz5QfCu7S8w6cfVR6kUEoWZCpi6Wj
FkpQksRWjzk58c+ft04+ZGjiTUmS5bxXe0cZg5NbshGu/lmfnl98CGMZs414mQ33
fuIHhC/AESvR7PDTJRJ5WiDuVfdqFpcK5L1aiWzNQIUa0TxMIvMaPB4GKcCWMrkU
gN0UjAcanwQwTCmi65zNlyofxiJkq6tJVlaHpcS5fj24/58wgilBnQ1h5p0V/5v/
W7/mP94fxyPin+VBlXh6NZMIWtaHKU+Oa8gFB6B+5kerPc5Hrmani+F+tMbnDoS7
RWW+n51eWVwWAS+fsNqrsyzBcWfaijiD+O/Lk9qhbTH3w9n+eEiNvFez268ZbwUp
YRDIDd3h2/lpkfP+gbOdnk7Jsoi5szQLCaSX0wS/a1QnqRaPF4KIjoGawaPMC4da
kWljWZpDMB6X3RSxWhl+WHqM39/v+3lOhdvGqmh3FUi0YcQXP4rFVg5hpr3YlY9C
eJyMSkCVjYjh9zb4T9MpAZ9zu0oKX8ySLJkg9TVXIdtpLOt7fRPZpXOTiBrf7PTF
8LTe0nwmuyAqNp0I03cIByjuD8qIhjPXQKQvmDNjS71jW5jttwFMv4unpRf8YZVX
To8mJafurYx0rTgoz4kOLxAGHCWJtrgCnBiFIEegXKhDjs9YUjoasGIpw4DwOGo/
LiCfmgm+LRqdLyu6mqC1Qqr0+IWKfjDQ9TghPCculZML/VUdmRPgM9fl8hKO5qFE
FHrQqONDcHbwIU8vIeV25OFTpBcvAhxq6PeDCMIEybQedOvYkMGUN8ILGFgJPljB
QYx/MWu6MpOk2YeCmfHkihhilgdCVi3SzVXtqASsNOWmoou8etijOURG/PSjxoBn
AWgTO0rAqM4tU1HqfoBcPYe55u395BiAsuZeiB4wmd0TcNC8nuaMFEU11tWRG3VJ
o7VqS899ri1VmjhAJGlK7St57cotLqmuh07f/9bUitvzOSz+Mu1Iktur0V6O+mqK
X168anXQaL85IrHx92seNoU4lUxd8qWFGoIDW3qKeBRDSHh3YiicOQw/uPDBSRPx
5WItVCzONAtZoC/MY9cZvXWRjARXMGbu6GdqjEXGjcnlD9m21oM+03cwTWtZxdZ3
ZNRd6srulSE8ALE4d86Q2CSqv1UOTjhe+bh5Fl1VZysrxOlGvEaq7WqHdQ0Dy/q2
Q27hygxYdDfo/p0XXm5IXngT9f5qDxnt5YjF1VK48TqfuKTUfOqAgWej4c1/xJW+
5jxpMS9Hche8tYujeFQl/bykIHM3LLXAkXE5nJBVPmYAqE3Y0LD/TDPsXjbzZrvj
pFt3mgbWqEG+fpUTPuZW6B2zXkMWnRtlNQG0bVJXCdsitrzoO6g6bRBbvpBemh9X
lSmXPOFgSY/21ctXBNk4miaxbS/Yrs8z5G70rb3wI2VFM8+xT4xZ5YTK7GTqFB3a
h0BlmLbcM0Ib27ohE3rbP0SVywZ4jc8rQdwCB1dpWyZKGLCHq5PZvHeaFZytcZdQ
JvI2JYbtDhatIhqrnxpL0Yd86AMd57TXXDQ0D/bnIDRWUel4Y/Zm80HFSJBZALoo
N5VlfUFK25pu7NIzttLHrjVEFvEGpDWAUbJTsuf7LI4orsdRVKtTnIze70bvCBzq
7rL8XJEg6A1kPCrH83fxZYWAoZdAL1aXIGsk/udPRbdRyVPUDiquz65RU3/WDfR4
ZJVuoAuJI0go1WemaMMBjG4tu+6ff5rnJfc3CTZGM0vzUzOAN/y9YhJM3ZtVuKo+
CDmlYfvZZD8FmpYIEykfHqg73j/vlnHfRqoye5IAAtTKKssR52pm79PXZRGCB1yJ
qC/Vwk9x4h7xasqMsrvdfDfC6LIqUVqBOL326rb1agdIEp7Er3Yozp55urvZqroC
uvm4yBBtBoUf+tstkUBial0FoOIJFNnU/A7ncZL8pafoKLQnx6puxEd6hvOchOa2
coah+ntx8mPAtzRXr/Cctytqi6kZg9+S/j1+TiBXguBQ3Cl2Zm/fqIcGeNxvMzEv
nhKNpQj1qUlBaMg4aZixvAAbaAPv433GMohgtwKIiapyHWiRIPjw7gp+tCi+sPJ6
fhUnkZN1J+iMFbT/MI+duz0iHbv3I0lRNNpYOnbilZtSkLIoGBGYqY9tSRi1BZ3x
1bCQTiQlvW8P9BcuRLBjydj+z9SwDiiLzIaCThZkNEkUfhMFSujsBela6xFHjora
/C1sjqOGEq2J9IS+N9Kn5zwwRoJo2HeksN+ppRfXRe1uEGboUmobMoSLrxVEzjtC
LSSAqYMIAeAaYSw1wShNUgaxPt8lDAYZrviHHUtpKpCPNpRjlI4NycoNbZ3v81dp
UpsfALKk72zChvPtsNYYpq7kUg6gBFXkxPC0Sa3qB9q3HrhSsUVwr7awK/LkuK6R
lza/LqEAUI5VYle4sjmudGAzfl/0nO0ImT3Yjz+mv8JrZ872VTSw+uXwhxhiSlUP
6a7rfiaPw/NDdR/fDwiPZcDCXIHgHbIbpdH4iTSIrSB6138gFIZVvs+yYG0Wyd23
tGjRAF6xoIQEoA3UmzK+1StLfZbdWLVKXtwcK/NmBVZv+yhDySKf3KCo3X5dlktN
JwJCrwTma6x0NDxApBqFgYMlGhzagnaF318KH/aFK71XVV1g45SZUsc2+jggWKnJ
BrB31BHDaJBFHa81W6efkDlrjUaezpvfKs6dQwAcz9YxnxG2movKn3uBprw39owV
Ov8mXtoxLUIioHIUE3BVQ1j+WcNg5GGl/7bYOK5gd/H8mUS5Wg03IUPmgGbZ82Hx
2pWrTgvJGdnFtvHcoyio4iSlnT9eXvJUXw/9iITO4HunUHZgsxy6YuvZ8W6j9td9
aku502I6G3C1fspreV2bacV7/aa21QsNrVpFNA+8r2bcRLNNGn6Dg1j9vq17HwPO
Z/G5GDx6LM4AQteAsQpGkU3q792iJ4WdPOM5jPVhl+c8GDKyXRPYM6i8oe3Z5DyU
CdSjS8fnJkT0v037pSIUH4w+1LMg6JwoRy2JlEJdOKd6urS02O2EvcvMEPHzh+MX
zTQP13MIZlVBMXrpJalfCtCZuUiPjUeO1csl5TJFSlStdmOBxbSoLXrIjEBPtOaT
CcaM0OvzW0OYhVwh+ZXX78daFW3OHFDmF1cMX+7nedSCq3f9pxSihBiMGENCBw3P
Msm3LPBQur1RXvOanNdvg4S17SaVXhWN8NbMAxIFwnMXMemtvnWTAArJ24iyJF8O
QpZZFSClhoa7wTIFQUOrU/ezR6RVxtPkO44mGH2bgRDjDdPpAZF8FYRJY6V79fpE
Yh6ADf1Mwxr3kxw5lhgaeDylplHmLvP747s0yew6zCV/L3lzhME/my0Z67Q+J1qy
etarSOoCBjsenn58u7yfMv7t5jclvX3SFRpIqmUB4O/ATdvHgz/1tlgQwvWripLG
xJax3qQG9gkY/lYhp2n4qspbZLzcPVxfSHP+IH3HUM9rnQWrDWUnFNbWqKw4e2we
ENWg9yoW5ggpaS4qQogw+aTz1fOspfnstl5dCs3y+md/3h9fBNDiD5LgJhO2ZGWj
ET4KCA8IRqVZEGXzvI5TXjybd0qjyslIq4sghqBaYBthtVf6n966CblUgU9jVfzh
Mn6chYn34taz61+kgc4TN8XUuSzZ2i9xcML1SzA+AeZYDB0OtS1PSQK+FCyHqq7R
cZQqiPej40TVhTfntGhlCE4aTaO/wSkWjisiSwjpik9ivwse/K1anqvrg30Gn0h1
jYtKelQbUw48knF29O79gc5EgtwW9fFAg3ZM1Rze/BbErOdpICvvwzUTk7sNoldp
AEcqXVlZXXbftKz7fUJqk4gctaAU2ZajWyf7i0HEw5izLHzQSggWlrOsM9jlcvXU
FWZXubxWXOHbLbPDdQAi2Y5Dc2GxX6sbWnwcs+/fz6/ID4RrcBsOjUehD03+2owo
0KlaVIkYjjSP+X8UpGcfYmXlEoakXu/qprIez6dM8rzd+X10HgDeIInvI5kOwqYi
O3tzmUD/3C3Ovp1kZW0a1HOdpaHXCgdP3D1owk5YgWbdudmLmrA2pbRluf6pHsh6
e6Uo62n69/EvVEFFT0bE/0ipbNxsHa19S0Bx406u0n6Q8XpKVL6+bHqzzgsEBgcu
B/PCnfc9GDXN1SQ89ZVkOzaH9ALFiOLNU77D4L11GJ07LSuWKmLxSPPmn3rRGqAY
rf/3Av76JHrI+c29DC8zHA==
`pragma protect end_protected

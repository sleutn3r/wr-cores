// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DhhtcJfOOAqZuznirymxac5nBEJ0EpSMWEqFkVFQZcMdnDu+KF8/AXMh5hNSMCXI
VkTCnFYw5xBq98xIDzk42mHzW1W3PAMzzfMzB/eTmeeFik4OvSYWgz+QAgwH1ZIG
i8V39mRhu8Hwq7i6+xbtKS8Zc7svfDzO9uyU7PM121g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 70016)
gHWZ7/qzou5/szi72yzv4//1f6kiesTtnP2TmEsWxki/3n4MDXeAdbsVqmEsqh01
+t+4t0TxP6y+uQLHrADHOOrJ861qSwxVWEj2zBnTo9ww9ZY3wzw4QGkBxuoaDmDX
eqeJaFyZ1NEZ2JN07GuXa0SEEF7KkXkoU/fI2ddOrGWl6wN1m6nR3F8jsqd9BsPM
HXNJbAinTBsmzhZ8688VUfHWy0J0wZX6F0BRASmUf+MW1FYF2QpgJXy1KAZ0uVzC
A+JIedtlsdGJ6w4p+GX2od35Elnwprw1vFMi8X1T4BdDYbF47wj+3FzqYP2LCWj/
dUkxsW9ftttR8NLmz+3Z80cjun7Azpis74vge2xBJB90Hk2pQs2Ag6TRKubsjG0f
lv2vCfeL9EBMxXF3BmnViEC+LcrBrsSBvg9WchEnPSh0fJiYYpkYKsMb9kbKjmcj
7luV610KPGdXsb3K+s1UTgJLz2nw4pTvfpqsmDJ2GQkrubr9WfwF3vvb8mRbuIQ/
jh24oZbz41CD2V4slnnFPTaB1MgfRbrv+D1gt1rbRNNX8okwnyXQfi8MOs6qR8QS
Dor+Cqts+sT/Cqv31lqk5ajIOnANaJkTgQFOStCvWOTIxZwnANnYHzyNAhF5fvEl
DQobD3rEAFlt4kd+6VQNECcgQw5Z3/8qDLPDcI5FdlKnIJoNlqVFbZeydrTTx3TZ
A+m+SVgUr7yhU7hV5+ISo1Sx1csHFdHepmF3EAIyrMcZZEUYWWw4BtEt6ZkqufwE
iFRRaEt/5g8274kPnXGx+KIWYv3Z6pKft9c1V4JZ4mD6TQOF6Ypazsq4OAJzqRHi
AFjWjdJGrNwJxfhGCDasyvRTnzoEH/Sdy10xaB8/PgmTfk3q+YndPebyqMyLfw0v
MVGQ95htpiEv45C3u9QSSmeXufDupvyMLicFGgphdGKNM2ZeVTGxAd1Mk049D/To
H87Q7jKBogQJAjSkfbIlPiztBbZLKvIwhIPrRt0MorqwUaEBGzUjBfPyOy8Mnobq
CelCheyA052zw7PvHts4Xib1ddn+Ag0yBHjzL+PGbrO+2VsFS2jwIxjaCEvKP+IS
ywugK6MbXPQuQVnQeDpbl+aarpU8uTsbji/SPr/UceWoh3mTXGrUlTQwGuos2WzD
97yQ0WkwL0FV748k1TqldFluuwwaB6YlgOEAnJQlYeS03uwBDrBSuZJWkQjZ82q/
R+1HNfBd4b8KD9UueGpsG0JZPaTcL91Awz1Wrm/QKuQeqHM1p81c6uhHo3veonbr
rpm+2auL4TWCHu5Rr3LO60zuDOeW9nd61dtKLDNmWAxALNIYlxTyM/h9DbGtttsi
G0tOjTbZ2XMenE066sWVZUOaQgJ241XyQvxkz02cO7/zUSVYXw7O03WtbwuU8J9Q
+qze+0fgIbdQ4yoR3EwkVU8fNxv3nnZuxi7dJ6IpT2qwXYiARFJ1VuXx/ttu8qez
cyE2N0cE4RQQ5Fr8xfHW+VemwKLFEwTFB3Lt0AMjmqfFHLzIXfsFW7lG/vKqcsi1
GKsGDMhouvwZSExRsbpamMQ3SIkQT5X2qqNYG9krI2BRHPjjGaMERo3eQpvVADup
fSRVwwwMbY/ZPkwmM9OIndcDodQBK/21HU74BJxz00XPwSgw/UbGivqd0juIGK94
xDWI/Y8iIzimbgAXkT3MSCsm6JjouzzUPdaMq/5riuCFP4tWzEuTEC7blcWCzqGq
Hugt8Mn0ZU9YOKKbY2+dR2bYJi1VnRmSo0hF37kpgDRYIJSUWoxAusLthzwO1nEE
++6e5tQq0Jdxg4iFmfZNTS03kVsH3n/F/9NUM7uxBC3wMpb5odI6dkTPs3TMTYVz
aGyby2CCFnzdJ0ykp6uedg3qStEWTrjueTXle/W7yepwn81kCWPtYKazJX0rUpRD
wmKTVF0V+VwtCjx1oN9F2rXuINv1uGqrFWkYF5urmvGp24iBhdSuqTDsu1CiQX/l
4nZUU5fNCwKrma3khvkp/R24uU91jo3YiB5habIHPnuWdQsNSILKg2zNbtYTJAjc
9hMwrus96fn60VUabuEd5f0WpStn0jCFqnN+U/ZD45sIcCSolFkIUOLvy9l/WpZd
7QjU9EB2GUqcRIFziNvr9R2xMCApQNeo7p83IbeEyuB1Dfs3WKFNGhp7vATsl21x
Idc7RChmFgBHyZibmaY9NozjiJIQ5TcEgFpa5xsbwYsj4HQOg8sk8t66YYQV2938
jqIKibZGbe5rTro9DPT2rCnLFzz3UM4m+VJOOqkf8kaPq6I2Gl8aGIighuVXOKHi
gD6Cnm6xtcX7eftHSmvftZBlQpyYjAQBqni9fGpB3EWVH1/Somd3BS87xlYSej5i
uDR70ISRBcFYzvzdPDs6HLRIHiyH3hiofzEV+TWD4L9/sDkAzORvnBbDNtMR3wCE
L2OUzlUoFfbWpjyJIWqFczyKRpwJPkWn4N4MfBm0bLKGDLdvihTDW587IYGIraM4
xKBdqK98DLXrnZKvPFQjZXClMdpguIcG5v6KsiqXp4R7Pquuv7ZiUX2VxlIHz2Dd
BwNalSBw+ZyddowJXCt68WIg2+yGQWOas1CjafOT5B1dZt+QqdMnOUR35hVw3UEt
g1wpdrtCogMSEXQhirea4RcZ1Jyua0LDrTb9PZkGMmFjnwJugwltU0Fme3HYaeKa
rJUlC1twK9rII2zQ4HXyiOGuYGV6V9k37UgHgDtSM3WcxxTkbF7gIMDj//MKu7dk
2L/1bflgio34ZlI0cMkh9vJgPUPIqkEH+JgShAmsiK464+3SwBZm4oYnowaC7xLu
geRXzYHUNZ6d6AugyZymeC8hORVdLlgdUXNvYDyupwIraVeErM/WbXSThqMDfUab
1MvnpoOjatrA3aEBHrr64orq0ZBhwd9wMR6UC/sKPAqmi6OEovR1dBHrUQoN1TmN
xhcLT3LpF6RAKxCYdiQDQjhkVWFfH2ozyGbKq09NKyNvKUC86AwBW2AqV/ektkRP
1fd3QqwS0YhQ4RMaOgoGhSoMlfr1ZBMjHMv5Y6DWECQ/+ADhRoIvPz6BjGNx70iW
yw3boOraFbPeBTH8GzPorQ61FHpKnOiDUVC2u33ruuaPmbIvu4C6/slFpRR+bgIM
LP9Rjf2OL6HfJHubaVAiqVTbKVAqL0/qIL2v//NRh+SpqPipD2EsQ08UY2iI6/80
48/WXaRcvaoLqPb1C9Q+MEOXQagxtCFjzi6sh6n+vswnGcI0SxmAqWbgXABxRYhp
S/9PuvKSwqCNzP7tnddg+NqScoLhCkwsKFJ81tEpCJ69OdCz4coMyoIl1O6fMWsg
XK+sgWOUjeT3HpydYGRuLITWQSHxHkqJdipaVNSLQQmqmwuNv6oZm2PCjXuRKmoy
hls2zWPhNBXEj8ll7JrnoV4b2JjHfYeN2Vua2/mZ0gYrMu5TxulRpji+dyr7aFs5
fuXGLJhA62ryk1fBHo9u0oCRR9+RRPPf7Tu1kTWL/5aq885zHaad/EDa9ahlJVKE
2jzHtGV9oBx71MlFYkWIbV8qwOdkDWZZCXik8ScEbuCzbsVXmTtkRkeQijtHU7df
L9+9AiGAJ3xIMqMFl2Mal9Uy6FnUlhru5+3XEI+xyyIF0rV998iXOIyPaDvpZ+d8
RRCJwZMIL19/fcaO7w2MhG+h6nVT/uQ/w9ckJygTRso2ZIrtv//oWT8hvISyruQU
9rh+SWHcxNs/ZEEFaiQFbwW/UjU4Am3lF1QP7h+Qbwgue3XhOvDmsRNe3J84cBBN
OwzpLEhazRcXt/Jc45sdu2Mp6pyS4dgAxSi/3x7CtG3n8AUm0V/FlQ5leE6ZVIIK
7AWA+IOYod2bKZNwtg98BM7bx/CeqMmFBwDNT3hJuZ2syIEnOSgO7qjMLWgerILF
2FMsYv4jWm58YFi91+iOrBU6BV3PHwb9SkgHLpIp92XXWbrDt4OJ/H3RK5316LXW
AZJ4HysnSEfwvPTo8I7W1WzU88xlIRNSwqSjqara9Yyq1R5Zn+BiB6hDKVlncHhd
8JgetJNPcRdp39lRe5zjFFE72FJgruE/mpJgYbM6q1q4lph2BCge/aw1UB9kT8Ic
Gq4uJ4LrbGQx/hwG+Ov6w6asw7kGfNVLJ84M4odPd2PWomvt4flkMIup2Fww7lyx
5eNnNdzhlOzU+uufuOLsjG1SlN/Eav+YNViB+B6KBZKJEwljC+9kV0eGU65sUz5Z
YkaHVgyRADVMZqdqkGTnHfOmE4Oh7r16pY7zuGwBIGkJgKSYEz/BMfjzFxPCJZyT
w9ILsucgVK4kt6WhTVRDQE9LhsODRfOrGo8ezbwS9NBH9On+MMOo6Ku5j+VZoUtp
3eGOq80n76x9qjZGG1qcjnDkTe3xYALuHFcxWEahjbC0JbDxr7Cgg884Hf8DTiUt
HE24Y4v/9vM39jj4JuZkZW5//6BYSs+SLdxvObdfbO8k/YuIDsctys/9IfPI05/v
FEsFl9VX3xFybZfIAGcU4aXzRrd8X8EDufj5zlp1yNT4Y8HT5y1dNe/OeXCl3mPt
wxIRKKOwigvMG5nWwrr2RxWy9xuaVnwNzhf4DVrutxYCL5fnBr9PhHdZoYcd3QHv
okh24Xl742g+GpDzwvfqFhPYyMVOMYwQnKy2YnxKnOzY/rd6f17nzaFykc7+TI/F
h75ep8pqWdI3CC1AO6WrZfd5MIm7nvtwFrTKRUn/XqkThoWGbxG0I2B9zkSycSnb
HpZO/RhMk9PnSjgX7hIkhQseOJpphCNriS1nuX+z7teNHmbVqraznN8U/5Ktm4kq
vaj6RBdM2vMgi6NrcZ0AVgeTE0n9lDhSb8nlfVSPPoZxHZhIJbX1JhURh8psSX1v
+zl1bxXcDyzOzl2AKbHfw+tUHTjXIX8B6XrOLb3OTzqbP1P7S/9zBMBDy6lxd42W
zX8Zj50/fkmqaYeDpB3ARt2ghUvOea6B76qBpIeJ0hUM+ISRZp3NWIZPtFgPxtis
6Oq5krEelsmrU6oDhmY8RVcRSXyciT75tLAYkdTYbL0A045G32t5dP6rwdWIgdei
sRwepcyLdTpWz+jGZRU3lK72VS522H2W3k3LvvQLWZDfFmxtCx2oIcFPnjTi8sXo
d/GYQAdF1fe8nqCaDGiIyO+ds/zGBNWB0ciwY0tiDgf0hZ7ud7OBn/XPD5/ns5vf
Jzs5Yk6cHcVQAyhUTAfvIzyfadsM8IjInmQbRDr688wpyiN9LhCgZP1g+uOtX5L2
MJJ5zaWGdTZOEvrqKrbmZxSEx25JIFEUvN7NfhBJVIyUbPBiS415+f2D9PGoQcV6
GRiLKAITHJLjbeEBDjnqqv5cGu+dpnFIf2iv9OfOLc7qey8+ozdtSzA/mqnQOmik
MubPetSthNYYfkm7/NV3y9UD0+4D/jup85YT+edgl8Nw3VjivZQEoC4wimpJIPvd
noDZs10y8nAfonUqxcqV6FG4HC+h7kQwnmKRSP+lL5dhO+QoErIgvomv8UZNcOfy
1NthnE4UF1755Fi1U2Vw4VIo9TbUYI5cUXHTkGYLEz05+CvnWIoSx8qFpiGfwaKA
6nU1t7g/WRXZZT4wU+/OV+W67sCD1LXL4nWr9TjUhD0QoJTgoQggA32Y6+pB1LEh
Jjc0mbk1dKmiwn8EGnnY49PNAahDsdcW9C4zvj4LbD3Sd5Em/4RtLDIY6MiGB0os
J0RooHamFtzCAfhCX1PuGT5pvHZ8PWEoq7apUEkO2o+YJSKFn8n1gWVvCrb92X8A
wsXSCIhqZ0vLkDaIeQ/ZvKlxMyv+0b7VjeRdx9raJuWB98nl2xRe2a8PMxouUEm5
nWDCZluD7BIij7QTpb5KLgrCI57g47GslXG+HtykDfdmR871M9BcxCGTzEQQY+lA
6IIVvPY30XJQtlb/G4g249r+Dw6jd9S5Fbow60KwtfhlKYQ8flfLSlLFKS9g4PNl
Q6xyB8Kw+Y4XY9cQTseC/5OyMMtDCwhyPMgoNVKFOA3REG3t60JFh6FzxF/Ji0Mm
txbnlgiauIByToB7FX+ZMtTG74JSC4hZwSby8FkAzc4VvzdZ4SDurmJCys6hN8iq
cyjchugy9pS2LhKDu35HjSyiZim9Bvsn/RezKvhbNVXw5Qc6R2dyRaTJazCSddq9
PN1Ym8l01mVyAyK4EFHGQMVtP02e75JsNSAvBIdt0hTfsS9kguA8nvdmGUIsPpQC
qyi0cdcl3V0jeUGPlG1TyufrR7uizRjNlIbjjECZrGcv6bIBFT8OfUBs9xxO4HUB
6zfmZKevcYJ3e71o8dxNi5G6yLt1QtqrnK9xe/xyspViZ2QU8jVbiok5H3UTwP6D
Q3Wm/Fluv1fytprDw1QiXti+Pp1hetB7quJCNQhzqrXaPon+nJxF3LLr6x5POtVt
P6OJV1rqgGKqTpmPj3r5GGPIu256ZA/JKVsumikgYi8pZyD0kyvn+kyddThlenrv
Ed0TA4p+AETlnhRTrnyrDSYYGBv1VgzW32WPkLsFq2luxK10DQOIudD+FeZMN4jr
Z37/dEla0mNYO8153tbb09Cf7SReQVspIWDE4fGLhsDetPajCQ6AVMRr8S/+fsZF
rQF2ugjIw4RRh6VqRf3h9qwMLWjXQ5y/ZzhnkLSQI3WmJ76bpHRV+BSVnrPUsiX3
ryATfWnmIRfgW0ZDxQodGLWPQcL0xi51fZq7aZdhGG0iFaw522Mebn0BT6NbTRGk
NRKYZNuSqWyAbWYT4gJLphnAaZa+DbEcKqsmnY0QB9SYvDcpURxwady+O59Ypnzx
f0WHC3dadX2UibH+ubAQx6TubDELOkoTjUlBEXEnPDPYvLfCpdhVh7iZI5q2BEgp
4t+3y0H4tnwJy/edBnf0BsavTr2qWCb+rZyrJCtj64h+WUGuFbEc2DmoMmiVLPAj
WQU+ASBjTfYenWPlNyJf/FW3X50sXOGvnbWhyTnBQxFv6gHn2v+36ssUIl8stxBd
A3fRniw+w2VeKbVi9sUxJpyadIivpck+Nqag5rLsNt1r79Cifgw9GS4IstbXVqvv
DuBLX2AWkFbLVHN01T6g6HzdECPap0IoflXV+xIJLTeDLRl0ARz7diKfKzh3ESEq
Ug4isru0tMAfR3kttscF/xdJdzymkEULUWuts14zzaisTCK0fzt3P2ANgdnUotns
Tshoxc/ne1tkHeRlselM6bSJ+Kqq80OJ+m5Oxipm+OguwsfNBgkRYeWzsw+Nu3+v
cHmxn8wtVDBnZvHlY5Sippr3Q08HhVc4APRSRGl2PjljGCg1V9BPi8JZPukVDcjT
R8BYKafUnRpbkRzIj686EmqOS5NM5AKREfL12Qkv1BSnacv0n6ydrE1Pgz+hXAwy
iKlAdA1VDA9TiKALrGSD+CxT3AOM/fz6UHSeWNgw4Q6nL46eP/BqiMeL/o0vzp3D
UNQ4lhhivvdu+btg6jfwzpwtxKTrQw2d0Tl5tGljOFzLAscBHEgFGkI3yk0zWqOx
TK8oylJE9xHBOX5nqcvtrF4vgxTvN7m03iAuXbKs3WD52Me2fsk6zrMcmoVL4uIW
m9G2WMxScLVTZG+XYWmJZaXG8At1Qo2xCWc/0leXQIrS26pcJ8XDCy3654t7wxaP
TJAIUYMgotQLHqrJr/8Vrsp4sE9kTi4CyUbvX2XIEdZhoDlQGJVJCO1hH2G/KnSs
VP16uaIGS8QoB5jBQgA6hZABNj/XI/ouuQmuBgop3+PUaMxV5MtCD09iZ1GsXUEL
JGcomI6uW/MwZs5AdKSk3uqBicmnfEZQm2PRpxGL6qhOilKMQNCnv+omMy1LnqXu
7AED3i/jWI9aPqSuOlf+O9HRB18Q2LiHfKYihVjU7eKh08UpnmXSH34w4g3DYWlO
xVms9lrgfS+IGqfrMvlzZksYAlxYYaRZgflsiFxHFTKW8kvSnpcLXB4iz5+0h4gv
c/rfpq8oIPMFw8oivayJeHvXgOpo8cWHIqEd/vrYUEG5etYf5Nua2rO0KKSQHIny
Dir1hdCI/08pE5DH+InJZIIMAqmK139c+9BuPTbOmzA2HjuL3F/5xLLLhFtWG4w9
oCtWBUnCFEE9P6OxQqkpsHMSSkfFJRf24FEpsa/CyoLSnxbl6QUqgDuwbQHnXlB2
DUw/fWLA5I9QcWMSLjTOZ4IgM3LLHsQQR8PPqjEyT0oC7nchCMMW/eVrL+sVASe3
lu3vsla+5+qVmEv/zLDFCJurnx0oRijHiQpz+aCeXN40G5fejyD9DK3xjX38oLi9
BKEvvnqrHdmzGrEXd+SxTTITFD007vD3zI3dLQXKq6URzRneQKWBHQiCbw27Sp71
Xm/BZbqQQjsquZVvnv/ERmWBofIU1pa1u3qYd3H85KgC2wdbzi6jFIItXTT3dcqb
k18aDK4/JzISURnXDMAgA3hcX5FzqJL6AY3JJxuGKSyK3k/1oYaPKgQP5wax6WY9
Q5O1j4Jzqche9Uj+/Oi3XPfTtdjlaY25/6Ai9OZ/GB5PXauPRvGSe/PtGinknQXR
4wNSQXrozcRNZ9bBw9P57wBn1ILxAmby/zzevkTeGAf1kT0TlWaohYyTFalswAuO
yOBrhe0bl7dTKTdbtkkWR+qJ3ub60W3pJvmeAMpgUa0be+xfFq6JT6LVqn7ocq2l
4LMOZZNqJ0C47I7eNjQFkUdu/8lRNhFNL5DwbFtrFM3xjJzbBH3DJVdSwRTx1aFI
ZVV6B4n3Mz8ZZhf8TZqx2h3p56fKkgYKnBsd31lGgKnwWjMJT2hKkzYpCgpBR4mt
TKVABBybrfsMI/z8yh8t0gdLs+hRiqfQw2KgaIOSCbeIJ7vtDZ5jQFzF6IVOqQFU
98QlIz7KEs5BKidtjHTDNH2oW+bjVxt0ycqXKMn9N9nbucsdT6RB1NvexnbX3wfd
XAjBKeZiSyBk0sVYx+lQlzLPbVAxbz7nGb1vsUmJPQqgS7cYgk7q2XmE9pC1+E0t
xYRSQECFkT3YQergULPm2M0K23i07QH+wdAb3qszuojsmb2OKcDfLK+otb1oWJXs
HdfaifgyBQjO4M80EmoDoactfuF5Hl7oJvgrXpC2B43pem3rPanztMfhTx1m6JhN
GQ4avlprqKys6b1en8RHv3tWUk7QqsWhP3H3MjTH3rKlQwTP0rzgboLnUAUHHgzt
IdYwxo6Nt9g9GgJ5this4w2qtGlDddT7Hp+GDzCzNp4Txfu7FJzKcGehFqkPwhcp
MnPPSVpS8J6TfZHCo2cmbbQGtBvevSlFqIXcx1iUa4WnmXqUXapf69phKuW0kudO
Al0/oL8/JSynEWQFUF/lIRMc94hDnOTSYHqcRMi3qB0NNMs9lCe48O9PfK0zAUVd
AgwYVxPAEs7BOyg4Exrl6bgKOHmCmvDyEa+THB15fau3J1ajP8PsjIUxREnLV2nw
K8+gTWxDOadgX5eZTDcwAhNvK9UsKo3iYTz9jHTKOUd68VqhElszbWexQizafwtU
CYGLapcGJbkENTA/ORQBiT9vau56M56BJHGMe06zktUQsMKoku5H+HtowrALT1Wn
8umK45Ferw9R38PDaX7kYcR2BMHqyJI8NLaorORW5GmwMF3q5W2VIH88q1nGmbWE
u1RxQXAL5rmzWRGz3WXbppnAconSatq6IFKZLePuideyC+Qi2JIo5zfGSeT9fLDU
fAVX/u/rFJww9RmBrQBc+4tbgGiHFTvefGxjhabstHO3TxamgseSg3FtuSrNrg3M
WbMh7G0FKvrCUU6zKSPUq0ElbvFy+r9GjB413mtxrH3sjrbe0Y/UH1k9KKr1a97b
w1MqpyOXYFKL50YOz2LRdnNOjBDVbBiQU0C7CfzTcp2IfvQD9kNXgj2SSm4mzZOd
RqQ5eG69tKimKZ5C4rhVnz8yCcp9NfM52iOafaMzCB5makZMK0U2zRKqHC878Hsq
UBWlXQ2jS6ziPHf8kPHt0OWeafOkqBjgIvMHPFYr2ENjgda0TKuJ5ljPYJnjbj7f
YgM4I1zW04SN9ABYf6/Lecl5JRDf7isSTvn60Jnr2/ybIYHSu3dcnlce68V2LOde
d3mS0vF3ScdgM2RMlO8FS+Iw/UdxBmErwny+6UlTlWm6CCMDWxFXdOSh1mMawp8y
lkQxnoFIGOm5yKtemAgZlLHh5qk1j96p7slsB49Cugi2adMQiuCdC4DzZY92N3kd
8Y2xaRlqql7EHmk93oI/JBXn1FuZyb+rmNNCRig+CBo4u0WREcsbWxkHitOLHlwp
FQ9UZFGPCxZ/oX/vhvFnF2xz+7TIRlSAaIjl5MWSjgX7HaiLWmW0++ZNvcDyiTft
JIhAZANB89ppK4aFyjrG47i1aL7VNk6McAkhtoWrkoZD7dBPUm5tsEvUUHhGUxpv
RAOzHOJRrn986viYQBaH5RZRgIAeLIQJJCjP0ntA11aIhS3eTWWsxa9x1JEUoggq
lPP5DikuA37zBnPp05jHZZCu+Hel5JEgB9Q6gL2e79v4GaGONn2hbqAt8MVuGZgm
afZNpuok4tZuAf+0dmYTBX9zdavjX73rH9hXnHCyyskuk6bCosdUoG+zsZz+xkpp
EfHUhiE3FFuI3DKFJ41sYPNHBwBFTi6mpdO9o0/M2WbHUEpqA2oUbcVQjMAclGat
rhRRUIQjSP6gWatTpa/IwznRKWTYFVwwSJFPbEWMgtxbjqDHW/a/KRpoF1coVdLF
beeW/Xr5BlduplZt1OBzr9Uq7dXsFic8PxsLgJb9TE1U0aqw/6Tfm5oR58HqlZZ1
R80zKSd73m9YXu2ubbeX87xZHv+WrbBu+k8wTR2+dhKip5G4MAHRBOf8KCypL/6B
Sy1WpJHnqCuB2n+/ar5dCwzH9PGw6F3oa+x4h97Oq2UMnTOcf07Sjmnim1raaq4M
XFYqyvnT9Zx3AvSWtW/QN3kdt/Jl1t0dFZf+2Jf4Q4KmZm3g8jepa9MEbVTyouE7
ayWXxxIsufvNjumy8Epb8YCDWIDRnFmlRzsTkjLSo/q3QMowpK1kYQxkTW6RTsmW
6Gj5WDskkmj7j1uG5DtMbrs+G6EEi6kF5ijr952PMKaEdLkDVPbiyr7fpeVWaNBS
0tbFTmZJ9g0swMkoNlduCywwBJJ0eWfEnRZp08tCa+9gxitlzaUR9Tbq4XwpB4Jr
J7poUHXyC8B49K+wt4KE/GJQyNANcpBZUZuAF21/EFIZeaT5Oko+UmO7jcopyII8
5JEtXWch/GyYbMBlrt4J/jTHczNayGeLfsjSJMw0ONG0Gco2CLFx/8bHFdgRF9+P
6Xlq+xgrDXCr3cYTThbi/erMIQKB/w8xsZxVr2d0gSBDAJsXBdflNRqoOUQrYsJD
G9vYUDWfRCy5+Vy+oJY8Q3Fl2TXhE8zlXC5G09Y+3RjM5SP1LfjsVpzF6jrQXnnu
y/Ip21EBSjgRhQYJt6LZnbOaQMo/uWLTcc5F2/PiRahFtCl2K6iu/JvPkXGe3GYk
sPC6WbNl17k+nsUiA3KY5S6YDcbTyNPfWWVP6AQ/zL4QU9VkqTXqJ2FQNT+6emuy
ADa/KmG0CMpmx1T68+sl8T6cFmwBSoGKieU3yF0AV+7nczzHoAbFtK4jY3AoYgfj
ORUs7NaIe2akaXQoIRC7xbyWhAOA+qKvQWuiluA7PfXrGuZIcJiuHkbn8B/AO2/P
SgC/NVJlumHlG6wzMSxid1oOLU1LMZ7h7zBsjYcmOe2afq4cHFpvtMqUEIL8eSCJ
sXaQL5vqM+Ammcm7e0CvfdyGa5ws5ZWjspOCLtKBHisQDhF2hEejKtmkjdmEdpt4
MENBzn/IUnmTRZBSXBtCO8uwn1fyJ5h+pb8LZ/EP/WNfCrV3kBCGAN11VhbJKLjr
ijydZyYFt9mB/ZixzXwa8Bl6EamNp5Mo2napGsXM9oWsdhZufbCfeLbTHftJHyEf
q5E3cPadGqq3Vvfbaa+vriGxzBVVRm1yMQsYqFmo2bPbthH1Oz3L5aMbk9aV/Z50
ZB6SuyHjJkgjS/VgJT+PNko/ZM11HiJ+Ypeior8x0hARvenTx3Wnw8mLpweK8qYo
VN42oTZxVZSZTdYLOH81zyjQ3EvWcipJz5H7j6O6wqshmoknyFPazcXHyLKVca1r
wzp1SbOQ3Yd6bQg8fmQXSLDsTnEUuGTOERhLI8iBsMkNwvHIyTXMO7sHaXPnOzWl
9Xkpf4509Dq5gywqdEgVr/0D+Yh+EPKWzwOW7FBbpeBWSz9/+lrQfNK0IPy40PYK
bYAMw4OmFxsUZWVWgWs21pHzD8dofvWfq5VHhA2SYo1DasLSBkZe9+WJav5vm/p7
MhMLB12IDCQR++wngTX81ChyneB3DS9Z0Gc082rjBU92pBKedtaAkR6ygLcalIsY
8SrymeB83tGOUs1EnF1fLelj0aGVYGVs8iirkLmhccp2N3R3p4flaxKD/rvxPhFa
eTt+ogY2rTzwD9UbsWNflw79INvyHE3uA/26G87DHfHJI/Su1KRZSP48gZ2+pwJ7
VNduc3mPKLd6+Gcm9RHWXycRYmsXt+ImR+aIcBu5ABJy1CsBdf3SWMqCrPrRAAXs
6adiGQDnROiOrC2GHyMi59/IaYiV5MHJryoqDGoa2I3HrPCTBRTciTxffapGlpfV
pZt69A1/lOFxkf0vSAz9LZPOsJJohmKCwLAkSzmzsFKjfL30MtiGi+biQkEITIS8
1mpiSNWXIqlUVzvvHtotEkvNLThmSh+6Q49fQDJoNiKlA8ZRW2rqelP+fD5mEztD
fSYgOmpJPf59C6fhn0DEwoHlzPIuIFKhBj7+IfAB+kgu/Xqzl+xDU5znLSTxq4Ix
KRZUG/KR0Hw6SPx+6idtRGBY3PTl1rFJIkTCdgWFoUtiuwCj9zIlIm6dwGKlRejN
9rRP+Z4/bW4xAlb2Y4ryVFZEkKY6c4V815LYRkCm16Agxz/7osjXY0JvYfggYKz1
gGTHPsHpGnJEsNmEX0uPQLQ20InDXWDJR9GNIvCZoNFcHoTEFsmEbQ7O9uWxKzIb
0tAWuarnAEi7/s7iS2xLuMg6r28pM1hN0ouJUt2okSs9KPxjtpK9hWTLxMvJUZLB
1Rg8gK7s5fVLT0ygf/oPj8NgSWyiu3Q/bEbq8t+l3LaCjdDcYZPQgD02dyKWISjn
L7smxux4QGNYu2DoeqU9kIpg/5F4EeEWIOqDN2UFxd47Kt173VRjI/3CuhbXfDEa
2zRuEJTFkEvrW4G65rW61ilWc8Atzt6uzfkExkV0riLokpcNRisJrbut8+nIWGvo
2P+zYDNSDcNxWKe+kkuMcfwz3Emn9eDOlOGhSdVVpuFZG2iQJq5em+gZZEkr9vSq
pVxTJiolq5p+189q7XPlCy1du69sEPnX8GywnGpwfefWkMwZp7JHRMRdl7PA79r+
efuy0hz5WzZS8SUDC9LhCtacjYPnQkTXv3JCq5HqU7oa4mQDtYnaKgRfOttXY7Fc
AdfRppcEjKCu5lLoFGTlY+NKp+7hXVZB/Qv+5avZcptQVL+ebaOOaPWu36vCJ/ot
TlsautdEJuUH0ATxnHiplVLF8C6wPbht5a4G/UdlHyoUHf1WY7anjrAIeJiwQEFn
2y9m4L/VWGvSe53RkdlQv8VUe5iuii8X5NduInykrlrKoIwsq9ZJyIJsK4Nsv1e3
byXvWHnOEyKm6EXEe1mnMU9el2Q6ESm9hnhKWO8zTfdQG/O8XJqqNdF+6GvO1kVD
Or9z3+i9GyCuRw4QCoC+i1ZMopUGUi6JRZzUSXVx1RYEPvly+/SZ11IbNR1eHR4d
86SRpCwG9Ko+EK0+qEBxlpZLBTXugxsqadr21oHDa0aFhguMduMUv63XHXuOTpLb
Uuh//liCZfbn8JasDH7/sOWSb1eADrPhOb67yp8wFQzW6r0nZsOuecp3g9jhljzl
4EW4g5oM1aXZmhuwfsnTN8DWS2Oxssoys/d/wxwIytZ3yk1hLhaGeHi8Fg22D8JL
eo17Ioq5vXaoAS/sUhMeE2oOTgLJOuz4FnaqNzp2YkxecgBLvNr50Dm84AYiTpwE
7XZktMMXSHHwQstX01dZ30THXof2v5JwfOCPwlzqgJnND7h9vJHogbPtPXIAhtUv
WWX1mkG623I7gp14TOndSDBSc6g2+Xa4pj7tSnbG2bDkUEnDkAS1ePszzpWVVCwi
ve5b71gU4FQx0/ZMZdel+vjCJKRRFF20VuMJQUjdztJmLIvcCExo6ojON1ryboeQ
o3u93nmDxLzArqaKZRaX5aF+KRO0k3s5ZaXeR35U7o05XzUESeiK+9+qF4LNZngG
Vmsz5D3n9tsXv9SvCH0fcqc+zu/DLy8DBm31+jIP5pxzNaCFmnklPrb4DQGSGONg
bcXLF31lWjKMJAhpbkv54h/CXQi8NvESAwXtfzR8YOGLLW4cgrakV6L3dVCXgSnJ
3TVY8DmkaGdDo5Q4ANskjeClYZDFDlqXRDVTqdJSTVpyOH4aWVXrMEyzHOppqJ0L
UdftI9hM/1Q7eCU2OQvPrgb5O1hX0HpP/OgRXPiDXhUMIvY273wmFrZVj3MEpPW0
HKbpx4Es3LyrMVkCQ/YuyBJ5KyfoX+oyXpAgPRfvlONTkhuKBwHlZrZoqFryKJVC
PH0HTXAbIHN3NuAn5WlsoH9b2cTyoETYANjKCq5KqcFedna+SgTvWgnB6l4FOYBj
g/0w5WSoZDPYMp2YUNksF6fHQAZRjGEggCCz4kZvuu/TGhmksNOeKMlGuu+MUYf+
74j9R1jsdOFA9AOQXBGmV1wzOxSVLPzaW0q17JZdKdd9mT6iOemcw6KYmie4gTiD
YMQBdqMshcyLnPMamTL91mBDDjvx4+XNFg8JSljzVfhIxS3DEgdIBamQDu9ZZiWe
/vjASGPMKg8u9lNDpo2JRyeHwpzYf0JZdaZtDWZK6JiTa8efUJloHbk1SS/v/R+f
C7hZbdvu62WNTV8qP9WjMIqYvQS64M4KuMkQ6mXwsbYzvef5gWWso9HqPs0JUTsO
pk9ix/dwcPw+XbPY6yN0nleY1HYbKxQFdVjuGhTXf0J6nqyLruL4NlQwPnIOpsIA
uoei+pXodf5bVrUslDILsZVddxY507RB4HHAuSYpzzWlsDnsLRl9Usc3gDv/ZxNn
J91SvKM7GZHzBu7YylE2eYkbHrIAEPXR1ndHL29MRl1eGeRSX37Aa1DSb0XsiWH4
LrQrSK2aUd21GIiVn2xttrKROsAST7/cwMDxO82OGQjNkOx+tySnKPss4JfKcwYh
Gq8eioiU6OBn+DcDrnFQhBdC/flHaYOXICwoyA6/+1Cr+cMF+tRULW7ulKRDqE/W
cStfC763mA8zwxCm1wV4RAuSP7lVfWJArfAoscalweLP3KidpGqYg7mpmxoxiji7
8TJLDAwu+OQs1xs1Qz9vWQ5RwoNdSSBhd85JsCmtt9rJ6R/5PWYuURFwvTaImERm
9zZ1ZPgYQ8b05j4nPW+yTqe7pwlu5FaTvke+zDRYp5hoW1n1Pn0rMjMmtNdc5x5q
KUMY70LiXUs2ooX2zLsxnLg6/TTRbUFbIi3vw25rG4LHQaOGQczUwmzj2W9pGVFr
Sf28K5OZtPWDK1dnV7MEgyPWJwX/mx/v+HUhxF5jfry510f+N6OOWf7ZLHJNx1P1
+aSAPVWGodScdAF1Qe/u/F33DfygwqESBxdBad+w6LYsS1NPh8S3xZ0p1+fhPXLE
77hUtVl5HQIiIzGiP5YAPxzLy9DA95p7ivDVws5zEFxQ1LL6siwqJbhuR75m/Bs/
f7qMcPeB6IvbFIp2orK5NPXR9MAiwGdqYw5x+F/1Bcq6TubkPNaGmdAbTID9wkLu
vZbqcwcXtnY+p9Rqc6SGTg2WA/Bm+sukxY+32gpa58E9tV6ze6SWyM4Vys1clKAa
22d/94ijNHp/71NqX8x+0/QPosEU6GErGhdE7rQ47h9DHpwarOAsY4dEqC54+zih
k2HirDFWm7sa13ty3w0LWMgmCUn80UU/HRoNxJwa0waTAZIT792VphgDu79OjwXX
agg9DXMbWCL6voaSTHyLfzmmfEUuVcFS/6AEE3WJf7HY1Do3veoU4DgobwrCjKgb
Nq0vrPECZxeI8njs07haBS7set3RRvCXZt5xeP/RC2bx9886Ve+82QtQBLNCzg4S
b+e2Slq7rTdRHzmFpWkWc4xHhFmnodqBHUachBUOucQkNsge0AD1DexC/RxFZcBK
K6vPjWDLVjmc5gVVe8LC/988tneLByQ1kfrXpSqjI9T+IRzC8zlDEdObAx4/214W
l6O5QG8M9k0RzZnyBYJPZ/h8hdelIeOKbpyRefucQv3BvXUNigs2kMYOQq/FfwuK
VszK9+zSGZ3Ej177TI//Q2HgGNwTSniQX3MC+ThFOng+tD34MH+ckAjMnG6o6+m8
h/PJGQ1UqPi60gUV6WRvDZ3t1S4DQ2cBG7LlH/MvgCX+OynrT/Ef7vJj0Es7JlN0
ZOJHO+6IKTzlIkFU6rjBAqbtVT+1UjSkR3s7km5QDsGjKi/z52sB9ebL6Z2Namhn
SWtWNBMxKdv/zRz9h7MTBrRnKx8Wb5wQURu0pdFQ5PBVCxZ3w8psFgh0XVwQ9sIw
uWZwf4nXWNokkzjSOZ7nfUfS2S3aEDGfntu/1k39WZaJePQsodBkB9mgSMKHQw0u
08JqskBqBekIW1jMcGFNeCZK/MVuj0u8pPjjFY5+FKE7k4DMKB7IV47xocsKndbJ
deqI69/5+YFp5CD+AYbiE4bAgNZznIwYZv799fWnQBx3pWIZWyNVi07wdYCZtzBm
I8K8C6qmi/DbJQq/DMVLUgqW/InQ2jpJkOjK8aa+y1UjO0mmJJNJOZCke359OkaR
0tCkY+OyTFJU4FY8/UzIkeTRZpEMVo61J7eoPi190FKmfXi881yEqc82sISdztc8
5pVF0rqo8XF5WX4Z/EW5xPM152biRIjzgLNyG+iB2hPSL0L/1B93Nerj0FWAZx62
gIqFTOqCZHYU8wtNbDDkWwcxqCN+Fyr24zcDDBY5AmYUuCMz4lMCa9qfCiP4x7Fp
OY36MlG9AFBqewDBpP1aT7fWpS+z+IEs3EB9ymqnzAi/ZXl7yRe0ijWIHQ1fZSNE
+lLGXzT3j5l3vd1Oh0Cwj8Z1IkWoAgzLbMGBpue2EssMm5Twpqc2fXesiM97gvo6
ZzCDIrY2gCQijq7iQ1yMAf/zduK0a5Uj2vnITyvvpsQChiDtsu7VpkiJka3IHkvR
xUECmUSHJbHN8xjnw6RAntFwcojmzGO0AzsdQI7uVa8YGGRRHQatB2454PXQDr9+
PFyNvf3aQxpZDGIOz96+nCgbTWhSpZ48oNbdGE8DtbnEmOSMLr4UTLeeFmFVA6QG
45NxIhJCfMGbxi7kvSyuZaGZov4Fw0SwJ3nlGMZwqVAqRFC/TunkH/Yh/E7FXIQh
WWd5YAPSnyhYdw+rvLhG6/NZKzjo+fzu+MAHnY5IArrgmBw5pCMl1VIIC/r0iISy
bZg1f/z+Ti/5DvqDeN8DRUweHKZMsXnDJaEVFTeFysdtaF63n5Ishrtd/l6Nr36t
69sRbtPQ+BTWW7ul0tI9VshfmT2OSM6wr1CVfQjnoNuWh8CylCJmDRcYhFHDAfbF
T6eQaDGKnYuj6Ge05sEfQLeX2qyMOVPi5vzQPV4kcp8zp4uNENvA2kH5PR5ICNpu
oWIpob6Q49iJDuaXGM1V7ergflpX79uqSDbjKpCwhyGc2wPwhJ74jK4a8Up72tST
DdneRFXKiwlF8osx6cvzVnM0lJw2xVHfisCxnEyoeC+j9PGd2QY9nrjuHtsAOQcf
csk+uq/F+Blp9OhcsMadd4RuekkLG0jm9+XqcvgI6H2zXN5/+KFLG2joS/ivhiuv
K40kZog9wCxma4x7I1xsGp9q2ZG+yijIZIEuWS6FubkSBlmBkl9lCydJaoPCuvzM
QwD3kHux3GvqCHMPo7nliDWyjv3pUvg9VO0kD0t44C087lGJ6A3CbFRPkvfAgXZi
S1RXdglViV/KTG3Bs4HJe9cd7zzUBOAtWmFT8alg1PL1OKVJ7/wiwjDe9BcHA1Xj
W/QPrWxSNAYQtHHSZqG7x6gWg0cYQI08+sb4WgliN9LB4nvDzykElhfVfxqBJv1p
LQok4U8nNP/wZpf4bUpxLlZKTQgMjl9JR7F9erQWS7a1Cu8kTNsJuBtCO/4DVjOg
0JJCqnXcNiiJ+KDyo5zs5JHad20SOPOCEBDqJTmDff2lyMSQt9ZO7xIRgcb0O+wx
GHbzJuX1stR8GRPIpnT/F/OSZ6j2DAC37lxWYOkD/VpuFnUz4PxPBQxR+XHkxNAY
U+fXDjDtuAOiHyvU9M8EjCvjhsSjXWy3Koy1tIlhVtEnGh/je4JPoKy2jq2RpnHz
6H3vIeX+lhQ4ECYfJ1HU1eDqftaFnuvXtop+p3F/QZhP1T1SJpVDnnGDHjQVyjj9
NtnoiSYsmL6hmIaE18ZNHpsJj5nuVOEUfOoNoG23R4i5OXHtb56iK3ZfBQ/2NYNe
+uvYnxSlRbBl+31ORa/0YP7vPohdRCjQ7/kxmTH6WiV+35nlLAT1gS+tUJ21slsH
Lb89v/aF1lIXlTUCEUSrdpdok3wQz7mpo1+U+3AjjhsyPwZ1doyjOHdzVdDHWlsy
AG595ViWgfWIz7gygb7b1ThcPBaoGGj1iUaAYtR8b6r9SSerEC0QDw5Vj4r9+sym
vtGBqRnik+iA6FVhkTYq6aXPWHb8J9OfKenT93WD5vDDNlduqSRY0U0ZXAHCAsbC
BlSyQ6G8Rp+08Id0SHQI0ObvOJg2rb8KOKbJvhS0CG09hhi9akJrEmQoxBK5/ar/
Vqc67lMTZMQlVZcLE7q4uJCf9NKcjYRNK061eHU6mz8q9WyL+pCSDIEjpyqxrcKo
S+hnkfNW9w2DbG+7uhWguBo1whvsGzcOp5ZI2S37GO94enrC7eeRwSegHp6wS2vm
MCd36E2SVltxia6PHH/HwoGJCXY4aVVuZ06qifqbhyeNCagfs9bdnPA1tftseg5G
0HfFxXTlNHvAjbnS7/Kg1ygzIBzP1IPG3l1AcTdC5W/0JEvwnRuj9Uib6DcfBJjS
QxALWV6GcQ91rF8Vazz6qnepzXzi46bvzrTa9aJ6gY6JDLJhT3TK9tR+f70dDECE
vE6YEUYKu6kUG92KU+ZpgePAAbn0fPRkCuFGx+uCwVD7pieq6XLitX7hRUd4u+1p
+K2xM/IyyBYH8Nw8g17W0cn1dAiTxmm9D9Ptot4TKVOWwSBXPq63xFHJkQNWmlf9
InzELT9AAxWtm2ru5JVV5o51GHSLFKZh74Yo8bnvbvQOSscXrcbraD6NZMNYBLNt
w0vizxU5YCMUi/htnVBuAODAZ8xeSJ3ezEhAevkp70JkFQy+xUNli/tCCT6KS9n3
l5/10to9mcOgJPm3pfaV+PU1bnuRzvVs6KjWnWR1dNdj4uX5KQIJL6KmNPfUd7Y7
mbFlerBFTBMpcxYKszKZuffRQATOE3/vAV64/M8grolWuRZso0PaYz+d0R4E/pJM
pWbRtEXPc8GOqL/vrQXjEXRelgsQ9DFL0BkNoML+BH4Uft67awXTmeZfNwOON3LS
ryceXkcsqLn7pkb99VpRJDErMTt3OEEyC3CqLF3tYUXZKbR6nH++ZEzb3adkQtJS
8vB20uMzJmvYKWIguZZ8h9lV9L3RV8v+IASY01I5Ff1cewidGyVCzoKi0g23MEUz
uwrNcoBczLi0Ks/bReIUh3+wdA8+z+wMPe+LXsi4puEFF04Ok6O9TIbC+9HPzx8x
Ku9A7zbw+JHuXYMycW0b4XL6+2Y9bKgJuqntPph9FRWaYZ5QbPUS4ud7JGTG5yip
TD3d4KFfAs9l8P9avpEcPTSLhgWigrCSNX2yM6zu0StJZcPJg6Q6kSPp+cOtay1t
YGYvWtGvCaU9j3yNohpdJxG8OVmhL21aGlMJkQLjUrgg+SKLj0fdXSgGcPiSaSPf
cYdBNMgf19QsBanOUGvVXcMC535k9IlVrPASQdhaeCPWIhxEfXfp4s/p7d2eN9Gc
EY0N+ebZ05UHsVUy5uJNun6aQmIx48DG/T2rTily+4QnJcIIfJomOw2Es/NlhBE+
cHNxTRGcBefMB4ko6cTim+Zf7Gg5dsK1giEFLXxMZ2TV8pgZlZSPHOYgbYSazHFt
c48U8ZKv2bRtaN5OBgy9AOfFUEraNy9pCQpKxCsYmTPggqSlkeu+VJDFRyBy5hjZ
VxsIQ7FjTs2IWyhQWs69ic/rx+eP/jJBmx0mYfRQ17aaMCr/uhH2Y78H9ZaNu48p
IKpOC7nbzEryMfbEE9sQCR+Lz5LaSdddS/ncE/zMNSEgsrkKMfQD2kzQ9ZAYErkj
M+dZOI+oXkQ2JVEeHDtImkVuUGdHjIIK1PDA8XJa3gxOs9ZyE+l3FF4shcYBzzG5
WsuxASLRWtdpqwtpjd0Ckoeid/D4W+5vU/DTJ0VXl19v3tTZ3T/2V0jeZBPeTA4X
y0p98MknSCnUxgl55hU3sfTVDzy/IAqkSu421k/Qmb+bSshl/2VLrzls08nF3xVn
kgzN4lE+VQgkVQlFdySwxlUuvGGho6X93mgKxzdarnai/M0snotprARjSj5vmUrM
Bh9GJYfwPZ7OHNCB0rP2OYAxTzWu4bpnGSbKb9vKi51gNdU8+p7lfWQvAAnq87qK
a1HqfdD02MN4DSVYf+9g1wYGk39cVtcFUNNFB2TNZ6jSna2v3Vq39xgf2FpuZAkz
jddTeoe+24O2W+w/x0CVzAhQBitQZ+wR11au++1HiwEPLq0YteJo3zWI/IEmRbjr
WToYlCbKDk0ZwroDpiCFDF8GKoLqdHXsiXwhf8ltDQ5Q0iU4s6j5kgJMEpTRipQW
tD4kl9i5QW9wWM8lwBuN6ibfXlgWxGHM+a4iyPTvwr5xKVDIRgtIAD/ohc/DshI0
qvn8uwbE8eKvjDYaZE0wx3MuwccWY6EfBFWGOokIcxWXVazAxrdQUT7HBxjw08e6
Wc2ZUzNG+22iOzn942bqkudFerBUJmAQ5dPFIN/5Xk//S57GX0EJUiigl8UHZj5C
Puw7R96HDqNtZs4xm36NSwrePEIVZ+wioMjUdEs2dhd3svIeNqE9+l3+A9K/8XsN
GyVtGLPhfAACr+OKorv3LbP8QsbBHwiJiENvZL4C3m0FQARg76TK3D/mCBgwZKae
4jcEMnhydT35Lf9AvuEp/y+Lu46CFyMQwc565wjg4/ah4MRBVbSzropbctbgZ9/H
RuQG5p7cKeSwWA/TEAgvzmAS/K/w1GwFxui30TL+bRBpT+ar6uFheY01Bd9hc3Cr
xD+8qlQ2ZMRFynhHQGVD4MsTE9/FFiRAQgXxXgcSIT6tybcA+8sXTMalz1Wb6G2s
ozOoM2+YXJxySWSi1K5CUIq/cGx3Vl97lVylBGJ1m7gN9TFVCp/bNpfdTREL/hvX
Hmlj8msTv3s/ngwFwI/UyUIHil1Tczv3E7t4Y8zqXnUH1m1Pe+tnF3Zn9muaYk9t
IgPivT8jh+v6rZHA85CtowAbIjt4Teu6Pj8lMN5kr9FxjySlmulsizAGMt6R/b8T
YbVY274WdrCOJX28YpDD5WuTG0o/sMBg7OYegPLTGK0DcZnDiuCXYybf7R0ulxY4
OmAQCyN4p3Ql18kQhvnfALoMTeuuhfsi+bssJXAH/EddxCLjExo9HJ8gR+CIT8Bj
CVu6j1kQLXuZw8UET8j9FRa9bKQV8ADN3HC4hFNajLP8JtSxpmWMl0EvHM/FxpKR
l6yoL5VU+5QRlJglpF9PWGm2+OAlECk8CoSRUlrAYTBcegD7++lZRf6c7LbrguU8
suFCTTi0RhgjoTv5jQ2HpQnGVJYnGdXyKZPW4bL9eaaihbiSBW7uCs9Lm0s9uoQd
UVLvWcn2VRtp02PiICSdT5PKGSgSBkPjPOTU+EbrkxAT4mL7Cl0A/UqYwTPKcdoX
p2EDnan3qNMeg1NoBWUJvj0X5eSLBgPwRO/Co0DYm3DGaG0nzsKJ5dLtbeXNFNrd
d8fRXjMwzpkhU6K8AeP0GtrsuyhfvYSFa6OArugySQLeXMC3AjdKJZmMvWAsitNI
PQNbgpKx7LEnmTCWkUNw4SSk/ou5IIsSpRntm5T3MqP92wGjOPjH6suwvx19BhZr
tvxF0sNGfxg2YXHbEvxKX5czNfDKZHB12j25IeMsWjAfOmrdSCrfnFaZEr81Y2Ap
ceUGuebznblWS+716OW3/Pvx938y3a6z33Xwv6AluEDnrYYX44Ry5mDIYoXZUg2n
wi1WXQwBi8CeTaihDbHRXJvDGfwVjm4RJxDYXGmGAqRwYWea+DGvCQDiqA0USIWg
Qr7E9ZdHmpj4UtXLfdGsIuNskvNKgv5+Rtni8B5cOMRLVNt+zdHuq4CVzx9Bfsws
hcQuWqRALI9ERYLfFhUw8jTtY3OdnbQofBKj52rxBU8Aukhg56aw0LVKoGgwUGUQ
p0zaNagz4J5oj+WRh4GCSoVlNTz2JDBJbSQbf35eLtotnzMwQStYURgDtpIansN3
S3/7GVS1XhaHULDvs1l2zYcFgwqr7Bwng/akw5bCjR0WthkQpjHaysqKZT1JAY7L
ToIte4/ZBu2y7LNw3p1IYqF7K9dtdY9htb0IdiiGDlRsXKGaq1k406K6jWmlj8Zr
rdbYec+4UDiQypCgNosRBVavXPNMk6zNWodZ7aPAHgcEtdRLpJPIjLwm+ZQhScnt
FjtLcbi5XWDzXtbiYByVDwjVsjh+h7op7CqDYMHYNNjDhI1QjzrzVdQZ6rl+EDsV
Sv6kiQN5+9aUDab5K9y+V5QWFfVp9kKoCAePIcP5WlJEwHwB6ERGHjRg5czH2ed2
0vdGzTt+SJm+jvSK2D7kUmRJrBiLnRcH9TcSr5xeLfEtkP5DZxvcEZ1OiN6F22b+
MyD+A2hoODPqhhp7wzjqrHIiBO+cMeWXku9lO4BRUcuQE0nsUAs4fQGumr+WIJ02
ILC4Psr8qOdrCiB85ZuxbC2OORPbQzDTmtDb9flKGZIG8sjKYgHJQV+N2kUNTfTg
qzg4uRRrVgPoVcpQOf5jTSQAWWPHQSk70AxQtfHo7uC6IGoxWa8RIFwzfp5uKPaa
m+w+dsGJ1s4O1JalGfLiSuuSsFS0B/dso7WXK8BCQxw+tdBILqvUZZYSuQk5gOJd
r+3qXfe0Fyf5OnbFdMN1F3PO0LQjBp/K9HwxUYDiBc6LRTN22rAS1bq1EoEhpsrQ
2t2yebzIa0tvLjifhhDZljNgh2IvkxUwO6/IbXGC7BEnMDHzvm379fxoBLEiPojd
yWQgCzRWG8OTpBrJJ+QS0ixwzLEfpyvb03FK/4yk7DDWya/hLDDPs5/ev5Lq8KsC
j1YJwfPXznvnwthH0dQ6qIlwgxyHAvlGG7MOsK7y2ogrUlzMhcC6JK3UGOeW2t3j
zOd8yCNc8wCOGkeTwPXldSgYGgoiq3JFSCpCHMpi7OKFQfdOagov2oa+u/PaP0oL
XXkloGko+CgRhMfwNExByYIFyQloCkQoSXoBe/MUAy5jJNV7mdHxOCtzKlMYg5bX
BCx1tnkpy/sZh83MTIkXsYlsOQ7wa8+1MyYAErUuBbeBrsXQZNsfpHra0d2q0RAN
RzvFu5OURpkW+rS+j4ZR4jJfB/T++J2jtIy+d3dj9OMPA1snP89JTxsHbaPgifjF
H3bRdBLmDsXXg8qi9BAcY5thSnHije23nglpV1nTCJ5aaC1mZBqLTsTAEN/uOPJ/
JLHcH4U71xEKihAY7mwmxjwkK1b7Mu8nuUB1y17OOiv40ymnN0pks6F21yB4iY56
CeVakltHxjYP3D8Kk3LWrQwBAl1+GP34MgM0L5z9qQCKfc8RzoZ5QQc5B9qLOov+
rtYWVFUXju8StH2Mede+uFjAi9UwSN4X++cEPnvCD7klZrb6LZ4EvaoUJmlm2hH1
VLX8Ufl47lBasbIW27RS33cMF70/K3D9W4P8XsLX8GAmBc6RGHZ2uPq6HZVkG3Io
I6ZWY7Brx/Gewx83kLTF72kGBp4q1fWnk9aNw6Eayv1c+jrhsngv465veRkTzyvI
H78PTX/3jD8K9zZTtlQ2dYZhBoWraGtSgJrsKHjtJzxkiKVX81B+2fM0F25FZV3z
hnnY5fioWZC4u77uyhO9H/kLTSn25oQQGwCSa7q66YaTDnI/Gx+llOv+T7fS+BFn
rEjHJxzv1iRLe1bVPee3PiSEPa53jdJIVkl9FnB2U1oeMHPfr3+29Hicb/rkkhHI
og8a7V8ktSJrqJEQGWcobaTIsthYNBBC+xxSFTI1U9xg5JmG+KS0BIjQFtwExjP2
GcBRIOihlW4fmWRSpJihyCcUdFkW7Qff+OBUZb+D6wq/wmcFQN8fffNOS7HHZegK
AUjTGKL4LpXpN2maAximSLdd0aqtPDcw9HNVT+jatUyEMKu6iVau6dokanD6BO6l
taGntKeMu/4kluWkVCJycBJknGvPJtla1P7dYxHFRsPrc1zizfvB1te8AEnuOh4I
l2yw2lvtWEQzujD52Ntj3NuCA0A60SwkF5n2W3+5R5g1MEfRaH7caa6WxVcdE1zf
T7VwDPUUNLQp9DOqIXCgAuqLSzmjPvyEUI/rjexP5NL4huxcXDpNafZEAAWBxcWV
2e2qJgFPPZvF8j6uDP3nIh86mu1wxRiL1NqrZFaNeFX9bJEdr6XHGVVDVcm/ujv+
VoFYA+Vgnu/8+W1fByMRIYxKpleup9aAwT7X+ORTU/zqEcUTF32jqhiL/4aqhu4W
1hMhJCOwVeOTu2sCBZYYcbhulwXeN/XZaS4jq6sTFpm8PGvpj4bZYHEHpJV6FCpc
8DaTx+Zq6Ye91CTZLlIbeJkk8TRtXf3vaa4JGEgPSl4D+J7dHQAm3DoxqLGpeJSD
sEG5zc/3kk1ovGf6liHk0yJdJguQgEumifejZsClz693GToUF2I1v5fZPVo6y/aW
KYiV10oM+Qtn6QxiZrwOrQaVjrgHIzDglMT0vj1g0f70HHrRKTanYMrmlDZUFH6c
u1CT0glHCaVc7L7F549y2w1H5oWELQVS5fPzZt9xJvAeku4fJ71C9lqdjxHqPugG
VxXq2ZPzJ5OZuaf8VtWl/a0rxnatn/7ntG/6RZR0Y1TlPOQ6S21Fyp+PukziS1Ly
TkmgYL3C6ODV1boFHWLv80gxSsx8tIs6530jO1YBHEl/tQ25TBt8l/TbAzMCtKup
vDwfI4cOCDfuLa4KECZv6rdjpdgkzg84Dwmqv2pF9/dvMYJ4dgzamr/CEi4SvXMH
DbMG5Jy8CHXQsemF5KsguytoVkKhINoL++1oO+XsYpja1tpLnIpTILQSy66p3u9C
yBPW3yLi3h7N9m9MZwwaQftn1Kh2yvgG0wbhAKcaeXyuqr0e2JRZ3BVPv9V7StOi
i6Ee09hUzsK9zaLoYlbfO96/FZVw+FZFfHfm6oh8c5lKPIPcxCIDzA/5poKJPO0u
QD6FjdcDsG7TQcRwvI/nSK/KDLWabnZV/BZyvC52AvLAj5I4b4x/pmkB4qzgWqB1
GDAeXFVlll28UDwPQW2y1GxnXU2YUNfX6/fZp9/sqLGWVexSxOjB7ks17mG9fWRb
zz1f97Vv400eTsGWdMSmcAYz87f7OVeVG8TZ7YJEX7uEjDyqxUhvYAWVyNFfQ+GP
r4xyAcJjj02MZ8rDb2MvlS1pb9b4a1ci3I8i10SadkcHDeu//opiiJCYpf6lJLdx
uD0B0l3KcAULtzlGsI+rMezNGHyDqJTlWpbQdFoK09AgofMvJO7liVNoYizscHCH
xxUVP/OAJT7q48CM/83WPXAGCfwfEQ5KgkfAfQieKtr2UCqggE3SJ9fRJsE/q38H
q1kAOheh8dT3e5QoniiwGtAu8xA8sjkN9ADJzSWhCTehYxpQel8EK0mHwDGkyvxq
sZHAI2BDMHixr0PUXOkAEPxLgeIrYuFb5ar0+SotA4RTrKgdwvXo6vFrm4Ga4mW+
l5wTXcDJV6d0RRc+RTlsVkSmUzxCMDWPCdxp5K4Wo+R0dn00VSoSKqxVYDPo00S0
x6y9ItYEVOQAYjI8PTBJ+bEiLAEFgp+2OqJ/pLcuOS+k9oYPiOmBqVWL9hCqmQus
JMhXu13cUUH15olL6SYRUwb1aPp1r1/23rjCeF7no9shOsdlKBc0WJGdw57HqpVq
oGRO+77qmy92+Kqh6gAAS1fwP7ND7nEtSh0fA9+Z23QH/TnDSeIzCctiNfYSCLmb
bZadAYQkgelq4atU4OiYTLd7J2B3DpDIWtTpgFWTGsrc5400a8YBni46J6hfeMZo
F2fDKkkz/G67SQ34V1+guJeG2Bou/cwBEppm7hr/d3zix8JFXGYI1sstWwB7BU2c
O5t1qRa1/8bfrBqf9FY5VbPogntabAKkDnFHdGUcDIvxA34TQ4HVr/Hl5f+CvXOL
8bpeX6gDKnFCZETJ2KCkSeau3MoUaOeMZSUVHvgM4CpjeSm7CUjcDg6mwUDC6I5w
IgJ8Lu5w17qRJhlxijv9WZsP12q4AU0gc8eAVgqmVRnWHPnnw6KbeHCCcQJSIhRZ
JW4WPRqGeH7kgx+p5b6bII/7ysXegPwBnZxWD6YkEe3OXwtKGEM3ehH43L5IF6/x
67Wpvp8m5uPaaajZb3+x+hF8TiBSU5gam0KaTHqv+/rvGIPwgzM8H7S9TZzyjpaZ
ZiUf/mF9GP0Lmlir5F8q6ENOOrunf0TqZv1s8TJr8ysIdzCYPLd2GavVuAT9yZ38
45SYt1ADa2UL61tHfTMkCwvx6Nze2/csJkn/7c0RbnBcpikXdiE6uuX4LlW2JKUe
1RXnP67Fv9MYJeEEzvmvfDf3awL436f9HL6s+alxspemx4ca7VGXMyKyK78Zt6w6
S6x3Rx6oOU69Wrw3gjB3mZ3DiCJX6dnW0MAReNVacZG5ePpRsbQyG39cw0qykxtG
QCiVYpP+oDZXCFOsNCUFsGXi4S1Ij57z/2Rqb2uDioiZHRxO7HnUb9Z9ij8oAfS1
MGhR1E40P0u6U+S5lvo02aMAAss7jWKEn5U0Tw6Spq0AOZNWyF1BqQvD9pU8KwyI
JCLjegosqcNkwKZiAWN6V0pIVlzdOllg4xw05/r98z+A4VK/3N2wlrBoCtF1rNZX
hc9/eiu1hdx2dTcF3NrPYDiTVb2H5h8vpalZrCF5L9GbLyB6POFlTBI0qFvnHJpo
VZBGWNM4QUSE1zERErtj6Sy0yrSX5d6kp6duIDYrf9pRMIILGtiuOx0w+mX8lSvZ
3TPKvKizvuXg8tbG8EriDbKEyLniLF++htdDgxHmY9wmUdGNs9rgY1SgB59KLJBs
HL3S1rhNNZPHlOHHvT1VJpCi1+bcWsp4PCjjfC1+CkrX5Rk8fO9XugCb2gnuG7Gx
vdI+r6fcYBZuh0bTF6n2IarMMBEqJf9fR/+b9XdVUQ0d0ks8eAwkPolTQjZcE0Z6
1UgUFBCR1HFj96SQIhbw1gJHDyXDzWyEHhyU8cWi/fKZDRy9EW2sfgHUfyyQvWsR
9TUSGbF2NYjqO+E+Nq2bHz7a6bc434B5QFoUZneO0RtzPUpq7/CsYttPcOgrauPn
60f47aADO0lHJaVhmKYUOuc/sNrHd4DHfGKkWvLtt03eJrLPVdRRW1d+P+8F4uzW
XLz0P4Dbbfl4ojpkm+N+WF37EWR2SXrojtWotSCTqK4PT3hEXlwuzzVf/OFxcPpu
BQN1yuylHmbMA6WZHYC4XlAfGdZLyfIQF3mber5NwLb2jrUxyM9FjKEirtEsqxSQ
LU9uK0v3ng6aeDB032id9ALuJeSkaLTrcK4k3MGE9nYmgxH9cz4xuxuRHb97QEuX
3MRBj/q/Nf0RHJxrtf+pi2J7bNUp7DHVb4NPKnsEArDqMOS9czBPQbq/Pt8XtSuO
LxjzyO7WToUe18bY8OJN6ubE8az6OaRbQks7mg5UlXiNR9U0MT40irZtwSBUDDaU
lfYI9AeOSxvsXoc3WU3YhxiDuTIl+yfxtvSkp4ROlrekNF26qs5tBv58MdPPVnvD
CzsQvC3FP7xgTV8Hn1sNrbKzQ4VscQV6Lerx748G+BXfOJuZRdBrxTDs/u6qAx86
1uvkBbM4K7YoZo9JXmtGuwAPPBjxH+mBXAz0uYVhvs2PndE7KeoBdltpnPkc1Rfj
BH2V8y8ykdFjXOLcqRWUGoaGpO6QurVUEvBeLOWGYwij5D5u0hskRbiY5Rk+folK
kxxhazW/Msj8Gz9w/XKjnvKqwyEugBcavNOjBaztGlSRrN6mHRUQLyDwh+KAJQpx
QSabo0AJmxjM2oJjs8rt7NixUqTjBikmhYhj4uCLxFRD5VLIrNCwRzOiTh5+w/X3
O1YHWOQ1BVtj7NXGpSzygAVtRWw6n2TW96XHDGwKXOYWn69XEbo2vCMLGpLez024
PckuXGW7ufpSWDU9TPJT12TOHI9FN2Del79U7JJqfloA5PHj6mCPXqTRhSM2v51C
IkWodGIQGZyPkw6A4vg4NMOcO3xxWqgjayLCizCCc5acrNYF4sC4+iAJtm7s72zP
5UWJptlqUkw715+N03GYzWVfoRHQPcArU6eeKTYtocuPkXEklipIjjS2wSvEUU7s
SXCskwJotwesKEjknW/sfxJPv80FsU607GqpTrWan4BaOOYmZjO7GuxZ0OmTUZwt
trsWOXVEIwJacbe0vN0G111FOKhf7t77IuM2d4Nrai3UWJDtmgab2YcCA11XEPO8
IGD7vvYf7boLmSabEw/+BAcxYrsVk5CKlZxJt4kCcC26pOUcX529wnEF/r55mpjZ
7QqYHHZSvghmYwjPIHOmqsf9QhDfgS6Pn2DvofcvmsxCHlxpXLEe7KjqSxffHFWV
vf1YspOzAM3T1m+BK1Ro1crITCGZJiALC4NUuaHRxivYBYSPEbrLlbO+Sm2ofQHd
Ay4qyHuVB+6/K93KHYFy/NrVbcSyMdx4EfQqIyj86qXCQNi/N8ui3CUl6cEke6jE
62MdH1tN+NXLus6a68Lk9hPQ4kaWkki/LzNnBYhNhXyRKWetIjSiITKRCQ5YcY/W
4HP1bwtY18HbbkejD21TV1bXCKiAO9j4ZEHKP3Ejsf5fEgtgXc5QxfNaSySyby9q
w3fTU4DcFJBZ1V3A/vdJUegMRljPfL38nNsgpeQ9d6idKo6oNRQct9TMeO9KUlY9
6ucqsFdBKYa7heHGqvTLeH0bAyjXe/JxcJMdP7xYWw1J5MxR3gWl5ThZQufWNKS8
ljBxe0HWy7w4ur+40YMBsLNkBFNWXuV36+x5HImEfly7Uok+E5q11+thUHFb1mhz
9GfIOpNNTwGDo24jm5AyXw00BzkrgdFHAQ80IB/yswIHUQFnfL7CoJaCSAcDDBSZ
lerbQ8T3Vo4cOJ6xWB2d77aB3VJoW6/xCyyaZrzTtpl3oNCCpvjJawcQwhrXQkYq
hHKJtJZJu7RB/C6qNMOn3zXWuVpF+UUp8yrg8uarzV5FWxcRtsT2df7CLBzKlxJ3
NKTYDRIuA1wT2bpYaiw15OfqecMiuzcN2eShvclnieFJ4v1bgbTTScEkeBJJRpfM
cg/y8JKRPvObOHtpIVuUWMbBHL5CWr/2fpYrpPOKrbpAwKfkrj7vVTgm4mDBS4zd
3XqaJqr3+GL58Py2vO+EBKnpa+OKRKhDTgEUBlUXYcG9KZ9e50PxUeIekC+K9v6x
GxN5FUHNAHIbn9XDAtcFkCKPE5xPJx/TEOCd6QOJTFynSqtkbS1jGhDE4SrC8hMn
8hF94MdxHwz/YXd+soyT0Oq5+GKAzuHWUBx6GsCioQfwASGiAaLY3deD6BAfyrAJ
hQcgQJrKFcfB9r6WjT0KWh9/9e0KvrhAP3KB+8C1XTr0RLpvmUj52zTQA9qWz8j0
N6VJmdVByhoJXmtz0ETxp6o3j3wQSj09D2qY0T+H3IcJGgcBO9serFQUR+J36d1a
WxmbmXNY8OylcAWJe8DxUFUAXI6NDmcsSTu+iEBL3xGTFx+Xcrf1KjaZ44OVwos+
iaKkZuGhMxhfkzB/7X65Pt3WMTdDyNIZRl4oXtGYuxexnoS3h/iWyg+fYYMDXdha
L5/l2dzZYktKlunVsJtNRUMbrus6o6G/eOK/zxbw6An2RXTid+YqckzNq6uw+tXt
sRlssy32P2Ske+KCQHjUBEFrfOvHQuIK8b6ycdu7L8/rrJiyT6y/VI/qUgypGO5S
hbDJMe8iQzWuKoIfkH2rRnpEClgaEytn6HbRzo3NwzRLYYCi5pmZMq84LCan4YcK
lv8Qp1NRlDxgkd9lk5HH98gIC/s4TJ/r8Vj52qcQOygxmCMd22WU304tZBLFyGWn
yD5kIGUEkmblXnw1UcK/TOkP6fLu+QVGwYmTpzwB3kGfB6yFK+F4gkP24x4mOXaO
JAL/z02i0QwUvWWPFd7SQ1lRYXPIAUBErNdnk/xvkjhf101knldkcFqtI4GxIhyK
7aNusG93zy1utTY/+eSANLHyoYez2hm16/yy40qWzCsRk5QhKykTN81cR0JMwIcX
H0Xxl91UJMh22XkhtRg7KeaLDTr9qa1hSKYF5EtX9zkzbBSfzepAEOpGrI7cQOy4
Q1amsVJp8rI1t710m5KLsZ8kbmKNDO8O8ZJwHm2nLryhLhv5FbdG5VzLoYjwhi2T
3rdrOvpiAIc8hfPc1EbgMhivZkEFwKTR7gkmFIdA16bgr+zRuX/7Bnvlt8Gp5U7o
w+oopzRC1f8q2/pEopbFULb/G/GRRsn0wm2JDhZ6lUyx9RL+RemsoYz8OgxhC3Qo
yMCe/aC4hpUHs6KNz3qzUtL9y5ZPsjK7Ar6Frqi44AxrpNQtOR+4OLhFNO3SRzTs
WvS0MYR64vxeqwuw8useHfpJ2whwLfmx5uC7cUbymPHreQOFP7Vr5tD1HVYFw6Tc
9RiyCFnaOeCi1hQKUagE/HbW7Xun9hbtl2bdvaM/aIccm9wEOjjeuMhLyVf2YutK
My7Hajy319Kts6eW+dqAgZd8kjw7qRkwhWNJjfA281p7i+6YOACBFExvUmOSqZq+
ajcml+l8+mat571XKOcc27t8o03FPbGdMHK92ehKSnICzqO42XuGGw+xif474t0d
gVtE4iJlfB9WKJw7sg+P8XFdflMicwxRSN9qfb74GSy5L0y0VMi5Xv4k73pCvBEU
0dkyiJ7Tkc3Wnrz8XrUbMltrtU03Ph1iQgFKv+QuTuSwA6Jycv3nLv3EDQpfHOaX
A/CXtD2rEp3r4zidpGKce+A2WmqTvSpyaVTvIZr5aJt3rxrWUeF7fjOt97EmjjwP
QZDmZj1WXjQJjw+6Canj0bboKi7calCDM+aIZW8E96AJgCq9xKFTxQ552hx6Pm0W
97BRqWMIMOixTgx5UdpRhPVNUlJO4H3p/ysxo4dMBaXDPVRYfXH423M+dPjADLEx
UrEhBkVNr4n9rJsAa9sRTQGMCCvZm2b9rSlnAMJZGI7/IudTXNVTF0Gp46EjAFlg
8louihuQzxc80EOLxEzm0jt3d9Dhvsnor9FcvoMUXwEaNTEM7jtFHKwgRHIuXuYg
nLNGrt4eLnbCRNKdfSf+hB3Z1DX2MW4bgD9hlADge05W6d22cCybkbA82w8gsGil
4Sh1ZHoOAVzWj4OG1hltnEFB+W3hoj5km8wIxIOgd3OL/KFcp6SFSaceMAcg6lFf
KBp80xQO7tOMLjfiGks8VZSMqB5yH1vV+79WYh2Vhkw6rVKi8vHcTz3UewUbsdMf
FzIejGzA6gsZrNC5pAULbwG2RilW2p1kMMrqILbY3V4XjoluXESZhBsXGzknhmu+
y7zmaonfOgcg/9TVz+qTevQ9Jms9LBK2IOzRUVnBpaaUdhhyf0XQoSq+wfzuETtf
1B05Kpwfrvb4vjyay1Sg0F8xj/syT6hq4sArCFybDQ6abKssY2GHssvPkjvy/plY
EwntwkKjff8tCerEU9UcbIer7WjykE6i2fvtsTmCBlFKQ950Mkh4FahOAMJZDa/P
Fiiu2Amx78PgRL35jfr1ZRMaWMz0CJv+yqgKn0agvUocOURk7A8e8ZPwJimkUSh4
/zBa63GlPai3iqeAMeqrp6mJnu93Gq/Nk4lx6F3phTlbtlGtCdeQWE7lRQVkUSPG
ihshrpPc0WgecEqWf9eIH+M9xahckJnw7kKRCMUtgG+NlY5+93rlphk5r0Zjq80m
6lsH63IkrSkubf+32tmA1jESN25YoVWb1N5+R+bx7JUD8MbVpfAtbaXxEV4S/dHo
Gqog6Y6Jk/uv31waY6/TWSLikRb3mAVUIK0/eEonrYEqMWV3mRyYv6/Pocc12bcN
EMLSvSmw2s8X5xmliiTxUOewWYcoFRDgpJylpLGrVdAoKpJzWDWVbP/5CFDknplN
Q9FucPnw8wWA4VNRLyURiCF2cSM32eBw3jYZG/V55lBpJOXnzHMmXRBiy2efjlMK
MTxMJPRBLzRcJkfhrJItRcX5mu/NKKLz+oMYe5p1j4sUe4UBb5/Nt3T8DuzEEOU8
UdtIvn1XxutyCZzdeBfRYTsN1BQEQ0/wMDmG1B1hwoOYwKbBQhsVvwzyJDoa05Ux
GFlIMIQ1/YXCvrINZ13fZfF1lqJfBjDK413lNcSUFBjsmO06ynta/r404WCLBonj
accc4SPs2cf6AJUOrWqUdibZzVY4Vumzs6+levkBfS3gbazc3sAhIT3f9tUG+wVr
Qdv0G7ynDqO4uZMCNgeHCOIY8c+uBHG1SW7ZTM9BJgpWXgpmWT3N+iPgOg0nxX0K
7Fexdgafb/OqDF9gkMwFgR2CkJqcT/AgF6kxbvxCgot7m53As1mVnVPV+RQBrzyz
+6nryjR1Zecanj/lTggZLSWUVYwu3jd8Eh14cfjZfauNxtMoIs5L1/yNJvDnNq+o
gxv5lkV0ekbby+HGyXrgP6G+ON6fcZzz7noxDkyKqZMwVFwyfCGJZyJ5YBaR9ITD
ASlECjAz/SIBM1tHAyIW3f/rC+Dgqvs0wz/PnVAbffj2CiGaNqtVwntWc9z9f7Xh
bZit9z/EfTU4g2AZYKgvv82YHoWEqvCxwkTPnx6pZBj3O2sIiRU6N4H0Pw9Ru24y
nh7rj7X9Aa+Tym38yZPztMrq7RZy7/nUKsP3c5ylwBnSjCNKy2+Zqek9dNXBI4bc
j/o+0pSPwuQPdPPjbXri+JoHaxNGxP5yh3ZRniAvKjA9hftbFses06HyQOcWCWrg
ovJFvV2furS3LYow49mP1JhtNx/cd41zsF9Xo0BZKQ50jhCBSRytRyBkrnKpi4bE
8Vc0Mczle/ibvnWOm0BbqjVDAG8eSlbxxMU9PZMeh5INb5Gw82JY1gSlEqJlE/nz
Zb1DHVLJULnOwN7v23TLq6W/31ZxIGfpzT8VuIIISAQPiGZxMIBDWPOxk5sM3nLK
U4JapmnR+EYGtFZ6QbsAsMpRkin+/6FdKxSlXsgbIj/XPcXYMStU1tpk7ZO5IfbT
QSKQUTAjhNBRy5ogoX1pT9hiEVzoUOlOgPSyydKpbmCTrrr32fbIH4C5lrcrwtxs
O1l8ISQmDUVHIpWXh95tCw1a5RiteEVOjJDZWHTVOfvQ83aXf/0UJ5d4KIEip9th
Lvo7v16srJlp5Wvh51GR4PI+U8oswhpyu6u7/IpSUQuT8ZbyOdpMJy41r/zrE1nS
YTe0wSE0z8ZSIw42UIqh6Bj06UCktqeHC0GHzGyWHJa4h+KvAIVrz0Qgy7/OsVDA
8JAZp60yYo4zTkfO8JXYd0FeggvL2Y/8kzcXM4TpdVHXZsTMU8JCTmAaU3wlUJ9e
nZetHb6be+cBrURq8u2lmdtc/7XtuymAcdchXDsjUuSnBnSxwYxtgZ778MAknccv
jqA0Q3H2zQAznWj7BwudDm6yCLZ62XQjmxkCA5cn6hbGUAuPO8vSapGNcynwUlT3
kqR4JMLoqCCstlSTtrR5Jkqttj2dlAS3Fye+U3bJpiW/VvQiI8BJBGZeKrgFKHtR
QFItvzCVKUAf5KhLSKC7GjcG2FOSVO4hH03Bsk10UGhxj6StgYmbrpJRiNJ2BmLM
918xjt3fZ8qaLsidKhhEO2zWhT2HQhyHowRulOjGL5oiiPjwi2J/46nALLSUsLG5
aC22uNoiayL5p6xoeJVlZcQ6rX+VgQa/z03YO2XtG4bqJ+zp92EXJRBHOS4pbOTn
l81baDk1k9t/ZSY5cYJLFN4NqGme6ZRVfD1cdVEZi511Ps7HL1y9K8d5oMj65fzZ
oFEPxnUyEQ5ZIEthA1/md9KVop+sKZE29g8/NWTRjWJ1plapuxdD1A9M84ACj4WL
W9sV3DN4f9/7hNbUB4U8EFKQ5aS82tJQ0KzxX29Vy1mvCSo2lyx3OZHlBlitB1gl
f9lQm8MzUgIWMwjWT36JLR9zop6hBuvrttJLw/LGi/UjF37HvLK6eU+oVUykdvBu
S2utQXW18nfwkVPA1frnqFrmea7zZ2JbY/LidQ0kJoVhONb/Iog0rpBxRPP/Ik0v
IHxtVPFcj8a//DfY/4WscKPY70CzvO3nzhsQ29oNuTO1ohaGjZiYkSXLtG7HIrvN
XEIrSv1R8TkxG7SU0Fa86XhYkvbUe0ld91mmtK1H6kxMiJpv35jySJNF+F5xVM0H
0+XzRjElgLvq2DC3nqpo6vHcQAUIy2QOd9v9eTJPHzH2u/BHtdc0S04FQH4zsVof
k/Qrga/88VJTgPX0UZG71XdYcGWClA/KBi+jiRnroj93fHWmobhSPwekjJiYhKKW
Uv0WrzM52TlJvo2leEWQAlucHBGsYpIA8MFWPaj6VNofU/BgwTFYg3MQOKEs8Fo0
fuLupHiXSd6ldgm5W9srHrSN0ThH2rl+ulCc0ArIkvTWzWUura62gfQ5689MnYgA
KwFsqaqeS2H3BHLDu1a5ZRjao8jNLI2gvQlMJtnZyo/XgDT6PQJGHTZyvI8MxFeV
CgGMIRFkCv2S0cX+noJqPV0ou5q3RpTDjh+zuxOIJsl49N24OosGu77nMW20DsfD
MCC/MQQD4ReKhDVuCQI/QLxOZb0II4M7OYEt03M8u3fP2pU/TkSLZoZ23IXemAZ5
BK5xMOSwcWXhkMWOwsu0x2yyeLYb4WbYW+ohZ3l+9zCsGOWoF27+qxMmd5dfkyBn
nZ1nBOgTgCc0d5Wae9gqj0+3DrifwWqAqO/8Xc9MnPKJETIBrZs9ZWREODzDMqC+
TRN2kDL+pZrCK6bYEFSe+0v1Kvi8UQ1psEZ4V9BMu/SwU3RfKkaqupDUQ68Ye1EK
EoCqH2ecvdCtsNlQPP9vk+vq0FJlORpxycSNSEAuT+0b85JWxt7drZEFeF4q8R0j
BSXy6Zl9UC2Cg/styW0YqoVPWFn77SBj4Maz/YlVGyiBT8jDvMfbSDzSNP0E0Mfq
fEMWi3OPQ0Q6wq2ab9o7pX7scpn6JI9+VIPL9Jd9jekSlJ6b5cifpKSsmQxCiM+O
wuJXSvCmwAzdWHLfFNpGUFJZJHXxS2yHzGXr3FQW4nh4zHysio32mMIiyLWnxCQS
s17IheeMSkXqrPcqeNfVGfVwQHWbS1JrpBUoYa0kL4pVSPExiZcb5ywk9hU6IurF
hX7PLMHnKljQB+3VBwXLo1ri64uB3k6Nc4ukRwoHcjQcc18ArPSNK2MbArALrhhh
/iC8ma7GtXuhmMCxpa2KIqdYaplUffYOjfzTUWuQceOnIJzicigY6/89QVnQoQhX
4KN+uSQU1icEoO2e5hYodmsMSCpJ4gxLFp4dE7eKaqbBWgLhchioYx0hj3bE7tJS
Dat3ljXT8vtmgoHFp1sTBJF1388qVcpRiUKtPzO1exhIwLW/RKA74jI2kS/sIo1k
X7o0S7sEVpYtL4EOA3+2+W2sVcrCajG8blR5Y8QT0kxgtHRMeFN11sNEpGpVnlmH
qNYseyiWmfKmKSkBZwNFmZ6NjZvuNIvhJLMmNYVfDYO2BEWaRndsXAOEPLyHp3aR
icwZ00qeuhOadTFwxwAHQcpmSTgZQKz6TEqNqtOCxKD2CEvs7SA2yBEdABmODW+2
uleiQO5hZPhNEIZShRFk5fzdCkVu95R9qDdm0lnK37jCjZjPIPVPY2YpcU/zgkNY
bjtIjXPfIxXmIzLfVsPV9mBvPdC/02RCpRNBiE48k6ORqoZbyTwl8KQzgI1DFuDC
YhPWesxh9L9nPg+rEpdMc6lmR0ppKNCUXiqgmVSW3gsd4Asq9PdcRBVv6Bo0FCbE
e17PPwqjF24zT+2r0024ffR5PhPrC2ZyGLh3nvX0vRl5LBK5WS40MyMuemp+EjM7
xjLW2jfnmc+wl0qFt1alGa+amp5fLI3imnQZUaN36LKwEmEk4J5Wy3UnIoaQlNzi
OpDWvw/F5c03854lQNSH6hZhRLK3Hbpl0B+SgVWv74dK11KgXRhNRhOVlTp6E32l
198uJDf3vr7qHiUTmM83gvLR+hWf7kNJISxB1yhGwMWLtI36b60savJcN8t8fH96
CjAsYAGtAOOYksDoywRXHMGUwP3SUYvAx4n8AWkBjNv8dfHShJMyNr7iKSL+53QF
MTlz3nFvmlTCnWvO+AzzEIdC+Q/hcGQ0A2HH5G4K+IJksfsBj+ypexiaHxo8QjOg
Zp8HUdTnBfZuQ0z708pxnLeNytnnyrRDPekzogPnbBWhc5zok94Sj75fuaQwu5+/
Yh8K6T3R4R0oFOyr2vcEdijuCxSHxy6/1x+Fmt7fTOvOzufm7JoGfOLuzJq0j4WM
6Rm5IIy+T3TVOhKqCO5sorccPy6VRaz9xliI0dpwbeWzRruhlI6DeCdGN76rgTta
nchEaTnDMk9ZEEAOTijagHdmH0bxLmc8YHFB01sd3DgKFzoRuwxzQeLuaMgShKh8
/woFTOj/szL3oJivQkSwDlLMpqxy117iOfYroBJ8DwXbEqOpNMZohk568M6Xj7LF
+IDuL+NoqCPKfqsHC6UyJ9iU6lqiVwxXRTMucByeXZ2VlLBmueTo6jgHxfkqffWR
2qjdrkNettXqt12P1M2LzmLVflA3SqHWgd0wTsJt4RjrzCyyTwTPRSp+NphXYRpx
C7TX+SFLHuAqPztNHIoz/aGFZaaYXYGtqgMsYaPDa6rdQIBdGiCdlDorOZOxq5rN
xaLUWX9vsmvBO9p4OeJNJNIbhFIOQDgezxwsYglg5cTDU1XBE+6XQTzrpNqX7YRW
oNrQT2om/Rl09BaqDEPkCh9LZegbUDRlSdeyCJpyPluswUGHE6Jon0YYiZPc5b6G
sydeSz1uMWE24/gdnR/0CeOHVo5D3VbeoBavPyXgpxXC2D++87kI+XpkQzNhQ3L0
voK9jMSfaTVrnAopBPQkjlGRDR7Eeuk4YVFC4UgnYAkl1EHRR0C24F2AW7Novx9m
Bzw88qZGsn0ncv4Sgg/HxoTNFyqHUaFiv6dnXT6m02nF954nfxcID4vFc0Ar7Lg/
hlZMJJaUiLKVJF8OXjvcSBkJPOAE4URt9cGyXlUeUr2+njmr/47EVw7RZ0Q7dC1O
3ojknpTithMc2DJM2OTOPUR4hu5QHW+qlUONANI2+VpiTEgyP8ZkN9i702bp+1+R
3cDw8B7abzMs/aLLaa1DqGKqcxgcTOctRkrGkYgTEH68uZguboQ0x/0tf07EwCor
8JLA2+Y0DNadXYScVIH/sCNK2ABEWpO3uHDqkibwy8zgvMN+nbBlZuGrlBpuXfLS
vpOpQBm0hRhuG92RLdFHpCfarMcW4ubWPxLjpceVZXU/cNvlGeuaurj+Mw8xR+BV
rqvr6aPvcEGuFoytAWKcfO7CQZIl7jG5kiarjBr5nSwzhFJJ3VQzi9LQ2l26W9Tp
HXyK+KrK3nxVJs9yJvacuAkDcTXU85cyDkAPda66w0joDDIl98gLj/pJFdEsXm9i
Utnhcp+0qcmwiyZFX54tNjIL+g0CU8ZbZIVf5Txis1UgpzOZ+NgMjQV9XR4xcZWB
fV6kUUEveZiFmUvXADbENTUZGV+UjcfBTlOuSjq8vhsRN6NcBIcdm+kPyv2JgjLO
PEezCOLDxULQPXSgRexx78+6ZH1VJuKKA4sDoQ5YsQbMU5Polj2DaM7/HkyeTtX5
jGsFlGUaHp38GMN9XGDojDufpG+xE8WX/QuFNwVDhwD4f9gmhbQHOZ/t+BQXnktr
K4e5fMkSgLqJ4sAFjIkT6GdIVSqxUnWS/w3d8JGK/c5ynBgS6f5wvjToEZHaO8vL
WaVSJEo5f+TFufvcdJuT9xp/b44NQHyNUAK7sN+OPrRjhnnmOuA+eoqPYcIohKr6
/MYgAnUa1q7MvySpoR0GS2uWrU08Ikr266j1KtwYGSZEjxpMvTt8SxuzFas/CZbp
5pjw80OMIZKOc/lXBmBQZvwH+l7SBCUCSrGVxhAd97DOWmaxk6KPJuMOkIDQqdoz
ZHgACHPlwTZYnk36LKtJoovM7wcW5tRfbtgz2CKPlfBv6cGSqa5yM/FW7UTaOzIW
BoP7WQ4iGzFKeCIc45w9p1hfXEYZMhGJRfHPh3thN+rTjSRIZGZPgUwROAgZ2Sw+
MauBJnHzLl6Esw3tSp2dglGXrjDPTKWAaPZT77HH2zEK5ehL0AW+O2tC2YLen4w4
YNbf3rqb96xE8a4svU7UO3/v5OmJhRb4dqtCKoPLwmoi6QYuDjpM91O8t08g7kcd
nXA6zM34TIVjubCG6qTGbbL7ukcqazltj54sIBhWjNxC3xKccZGf34Wf4TwoVrnv
BVj94b8w+U+dQIchtnRIUn5aHF2jVRUNdji345UNQQwepiyT+UG3R6evU3inzbT4
RKOQIS+HML1pYq+cUtq+YJA0ILf/k0l0ft78HvT0gfHkhC/PNDFgWOT4V8ehYGPx
0ZzDcgqUByxywH3iRyh31CZSk9bK2IulLxQjR5s1zZZYlLKcPW7O1RunW8/GdlyA
6is+Yw+XaCQ3zjh1ctXcfxRc0l+v+mWIRr6Ft8VAm2PkJjuuL48sHRCkRPcdBkGd
Nil2W4xo/R5/+DB3Ri7nCw2pWoVJPpPYbSbSynMqmwAGFhXK2s5a07ad/fYHchV7
4Y4LqC7229EXQLzxOez0XToG/3anvgUS0eAPps1PBSCRHuM2+CZPIyvsB+rIWEJR
5aMoNVQac5WQXxgc93JFx9/TX+JWHCyvdy9zPDDGNEbObbey0h3Ngg78c1Wr7kBg
NsgkmlaCgJUZJGj10R/MxDJNOxDViGWAPNLKeX5TTalk+9BJTrECCYKrC8GBgrbr
YgWljWPteJMMoJ3iTpek+MpXTPjr4e46JjeKx8XM3UTwxAsgDSyYT6JYh68ZOYh5
6fxtwrqYQpOX4D9OLt00LB2/67bqmHD8F/GHhlyfgEP1C4oCGPj24yNaI6m2sdjE
wjzGdoz1NdKdT0eywI95cu3LwPjiKtMkHFxGwgUwTvsL3f7zf4Ou2EY1xCLsJUIh
gMSQBgYVr3qlGU5snMtn2zJFwllorKG4Lz/nG0hVIKAUkII+QNBDlWPVfhDQfvkA
ffIS7kaCVDvWegMtZEGu164r4TnoPqmQtzN9LCFzWk8m8v6MYwF4iLpNyZ5LPzcN
bsfun71G5vawbZ7roC6OxQ1yVM/2ldIpFlAD6RInKNhaGzwy44uHSLTSrKixvXBB
azPUhcvdB67R5T9hnzH6Nfu3EWlTjMfCVGrXxIdYpyJBRE63Rd6eN/BQb5QRTGLd
gtCvhNTGCoctIsXZ0gfISuxZBIqlWokB+QancU+LUdExataAjomghR3DcWEQ9Bad
KEujdZaxlTh/RKxtpx2+dmOxL/fru5h4I6vu6zcE3NLw8TP37VeEkvEFVJ2/6YnQ
XvxzE5YRY5BsT4inNXqA/R1LMoxymF2lZoUFBZqxWNcr4RtiW9biZO7YpoJRLE8H
3X7qyRD32A6YTSBmQBDBS1aRweES1YL2qFIa9qm2W/cFF01enFyiDGYKF/XOqNbi
vcwr2m9dNRtRlbDvYh23zChuTMN9r7+FKLAYBRFJ1dmHEEJLkgiOsqcwfEdkV9t9
nbxr+u8XGZuNky1ONr6SB+h7vPYhI5tHrVRLHfwk1SQEiHgfHf8Le4KffHfRdak+
Cy6fpxjCpLIDHmq3TWPdWWvRu2BentvpcE9Ye4B/KDoLgxusIzYVkH5aezOx9z2v
EhQ7G4wwrBr+ZdwDfQDA2/2UkDaMfS4uKPRzL8tqy4m4zxQcIJgyIhawbkv9RD7q
NSJqwBL5JwWaBJmDajLD+YJrkFb6Vm/fumcPhisznYXjapjO08ROFcEvqdqLLR1g
cbLPW1dbnGzF9dR33yQ4OMVQ5Vn7XVNQ4zsSW1d/YXoxwr7Md1g3Sod/Jau562cC
qZ7s0E++6E8HcIf9G17DW/Ey7n2k+qGcE/Eb1p0XJfGRkeLZtcXG8k10Q+C2BpXC
Ch9mOWxIptHphO5e2YkKu/qATVm1lUHclls9y8sxkKU9ERh4fPG2YrvSCoUkg0bF
JcBdqjy+rSGKQTZgmLzPCIVMwPo9uCwbX/Bj9gCWBdzen3Mr7fPrvFGQeBpLIAgk
cbdSIhqnhh5bNvSV4RCDEHlr9FTQVUkyKFBvFPsfCTgue6AgBmzO9Fpuhsq3b8EN
1ZyN+jrEz7EyFIUatiQp/oZiDF9rx/4gYSMas/+4bw9XL7XIMRIFCX0MQjPJTG6I
yvjtBeV7dvdcw1uZdMA1narUvGXLy1cbPS63FMRZ66udrvJASXgDiHQpG9czWo0c
xCgirr2AeUJeVn3dyakdg7paE5cwG35xu68vA6EHGZoAMfAr3TVnNZegzQwwuMkZ
PbDN2aYD/LRwOPzX/FnBTtgNKZZ8rjgAfdh6zY1QI+5dfSBtmVZ3G9ZUBWak8Oc6
vz/sZKb4mwnFwjOa/vLHTEf4wkY1NesNCMKthHfrd0+fID+LPSw2VMCSAC3r2Ebj
8xXEMZ8iZsfzXcSQm/vxrm1eMv+5+2+erBNMlSEjqlRvI9Zi34Yk9qMjaAb5RlbF
ogtCqLMvE2epd2G8JFZxYHvq3E1rVcjE/VJN+KNc8Y9mQpHB+86IjnVm9ezSNSO6
8EreEx0Th9p/j7hbec45uAYb2hJN8yeqba0zC4fA7GHCwm9OpwSwJAbAbUd98WJb
XOUKx9eXGBs+8wYng+rPcH8wdqPcE8C+AWIHn1P4R/xWP2S1342GhRk9miutgFY+
WHR6sJuYIae4RWOcCuSloP+uqcqA2Wifc7f2+whn8q+YBlZVVQ/A8Fwtn8nPj9Ce
GSYJM9Z1ew7ON9v5WnpRYjnKKOuvsvyrFiTg5QHVJ5ohbINktqoFQUJEjohxFyJ5
nqzphYCcpX52VosP33lzSo1plPSDwKf6xUHH2zEWYJwioAtPywhkrYYKwi5MDsZW
xMYQ6aT7P0CpqgajsqPziyNJOLqFZr8QqUwt3qQ685Q4cQf7nhD2hmkVIYnDYBzs
fGfbuZgiMALe7txHglEWkS93VLxozN3jNHgaZSt3/gpVOZOI1GaXhsSlnIy+GJYD
H045OrSWwGcgsfOlHjupu53TziZHaw7zKhERb1ZYQPuXXcBuqETgE6KLnbHcAY3r
WHwdIqk4Y9XTNqRS6yUk/cLdAFWPEMTny5M5/KmS7kPVFryoUYs0JhogdTb8vLzU
CbGJpaAT2Qa/j/tmNFyKjUckehmk0rGWgrPJZzM39OmcMM20B1Vwo/R5FM+HAF9a
8YKk/aOTQ/P8OT1VSpESm+4C+ftsyiDsfE/gFI76dufB/jM3Qsrmjayve9D7RbeL
VPHBI1FYRgkgnM1Es6weI8BD1VJL43xEaP3DoXceqDUAnUsz1Ao96PVgYIBSJk1r
ACKJikOgmpG84mziQcWIUTUnG8w2znjZEQE1JKP37uCnv+Nh6rm9aB+rKeMBkDHh
TbouzOAj6NzplEQhcp+fNL8G6uvBMvn4XTn8jII6NEHKkw3Rw1/bVRCbxctXIsd7
Uq8uU4hMwLzkHNl2zpEAz2pUkz67pUJjj4o0K8f3wF1ljonuZBNv5gsQj4/t60HI
OLBqRTDja5inGr3lNUBs/uHDK5cFJxuUiNbpSdvfJ3BqdqcDz9OvK+nzJ5lC7cSo
7Q8soWU7mVVtWGjlYYLKEcZ+TLU1EQWPHlA+M5JWRca0Lat67dIBhaygYJPVAIoT
QX7PLBqAxOBv2x1MapA9fOqF2tq0KwK++OGbnRrBPSC9mEn+Nx4LxsX7pMSynrV8
+K/Fgs5Gcxe87SGw1GTKkdBXK/wlsUgXcPXRnIJyJqTcnwXytQ/UKWDe5OGzzGaY
E8mcq+Be8DAreJJU9Nih9cnnbZrhZWf8n2+5IXEEH4MiPDrFERbTp5zxzWHURz+m
QO+vbdsMNql6QW5e/7LB24CNCSSYFKcXXrDygkzohRs+HdCMElJuXyo8FKzW9UC0
SgK7aJIuIDwRPDsVFHF7boZlbOlMrWu3lOMUSpwg2Vn6ZTGcWqNKcvmEOvql4oyr
lGboAUmhVfl8wrh9CU3qsYvto/a7Bhm9/V7bwwAigzwddF7YBrj+rmt3YOltM3h7
57tgWd5vU5M2o60zrB892zqzuWzDsNBT/Ck5N3lWWPwDE8tiJ4Y5NDkTzXj/C0gg
d7+RjhqblqViiHaQzxN4td9Ni9wQu0OHL6Cyabi6jYN2JNbdSiGf9zDlzj2vC+xs
cCVN66GQdp+OePo6Xff3uOHw8tpgytu3sFXEavnnmizFyKyqYug8tKMNEljCY5OC
Bohsm6reyzMCt9yOh+Jtwa6Pujbg+/sY4cePVSUu5Qq1UIpiokehRg5o+tNAPSjg
uWGT0ejcp8Dap+c8NeZDrfhrTt2pYWDssE1Z2PAILn1M5FmKtgLWvwxQ98UcNkva
CDq+AZG7lDqNc+b+9hcI2wWQrZmcHN8E5fYJDRyvPr063JKrufNEXlC03qyLRVQE
MdRdQuLFtNiHW9ciMsYLDDvTkl99hwT0zqnhc1HTzxjU5zBCrD1ZE3Ao5Mq17/hs
FY/pnNp9PWR8FoPpjxpa2sby8MJK/EGzt/oWS7buAR3/NSxIC88YX4ZJ9Hx7BLVn
a5u3KiePLxnTbhyOEBUag9/X24VXhmsdS+plBIcj6fzKBSkgq3diJJ/pQ7Re8bx8
A76BsDm5cYHEBiR++uPKxVi9xkVg1CH/7czFCkLQA19j7F8A4XIQ/S/ciYMVDKu/
k2TTxaru2l6q3IvtAZL0FW5TwDHqCo1kE2RCXVXCfF7qsotH00VV7e/pKkFMcvzj
yt1EgK6peZ66kugZes5178Hq3wt5YWEwl9B5EoMueDn5373m1jVOmIKJC5+DhiyS
hw1RoMe/G6zEGAbna2WMmOpbfLEDEO2xmPhltzgvzybW3wI6Zf5eg8napd00cb34
CGhu5bou+tYt9jNVTXNiaednn4BIZPqywlZnPaJSl3nCyqIY/ei+pTDK7ysaaT3z
yu4z0yzDaonCwtLGPh58RAzE+M0p2XMUpYYA7OpwrIyZeGwuJxbaKG+Xjg9X0pqx
MQntdwsrIeVOEKjqNra0oG6s0noYJPv1Q90rlU6XbkntvGlvgOu8Pw4wOSDvXA9d
V27WQgJyIWxah1v48st1hCPkZwvtEoW3MMkZLc8j2XeNL3WTs8u2nSba1+bMJ8R4
hKGkC8E/8IpBj8ba/Y7OKau+I2MpnAVnHDrPAgT5KowB1rPA70fSDz5gSGeqOQSO
1MjlaUK4YQMUwWj39BHr5aQ+pE/ZGheAelUm9E3hBVYKAeCtEuggzHA3KOrfU6ty
CSMBh9Y3sBE3tqh0kMnYMLbiKdY4D7EcKoCXglDPMw0WnCsSWXXeAE3fA0NMRK/t
JxM+SZoRn3wQVpQH7zOacy8H1gg3JmD2SOlkgW+hLq476jNDoZhv4Axr56X/T6QO
QNdUiXPuPSZRUiNHrHkJd+kSaK4Q+GfspHn3TpcxN4VPf+7VwK91qcJ2Qu5y+uA3
7HOU6O1aUrvkXxdWBWQolp/hE6pxhjjUWW+C0cCv7tu7n6NQr2KbYsLQXpgGZ4Qn
f3KU5Uu97VT7GqKoNQCzAtpMdu+l6Dz6s1kUhRrJAr6SORMGyA+7t3Gn5Pyt+em3
7vD5X8BMyes9rwb7s6LR9Ujm9z+nevLRhRtZ0FlcSpXUW84Rnwqf096NUUxIOtAP
wf2zqiqDZpCC6LZEOXrBnpzgA/w1qi8IMKS5/zw1ZJJwjNtM0IOdPfzi22kMNUf6
nLQLx3JgOXLKQiqkdadY2BTldd7ul5wtNXJ0vogqmPOFZSALlRkWIYExeIGKmRIa
2RqXlwad4aadNS86Dvu3vpa7TTLEyB6OGMkisScrJdzt2+Ag7bC2pVst90K5JPDj
2Qg0oIzXnk4lwmdm7vtiXxGpPLB2zxfYJ8q2MQxcI+csdxCxEDAOqjt8hxAxYlDy
hjUOFDYmN06KQdcabW1EZXTH2f14VZ4JXMSfGtgSEfa4GQ14qiic4rj30bW3htOY
tG3TnHoHOSJ57ysqVak59f08ii5rZNIFbZjs767usc6g3f/AF6HL7XC3la0wRWKe
mLygxNyygDSaELiJJ6ZIYUx284MPNa01IixNL7wcBPIkOgCWNjMJ4kKO4s/lXy0j
1WHtPTK2PzrFg/55AYHo2ruLKNPcxjy1m7n4d3WqZkR9Kaa9D2vgsAzOm7AMPqYQ
Po3w0gklVLklWsO2Lmu4zp0Int7AvAOgxHfCMMr97zSoReJityqFltHbDy+aA0fH
NpdupOPDI6Q8UO9epWzkqazfKi92OG6iK8SOaLBIzN45fFSmUEUYx3Syiryvy2tu
dLMIXM/vukD8e9oPENgVvr2wBjML7nPbBweEIV7ANfxtNfQrC4uPh/B+S+5zRmXn
hZW/HOhr/WonSSViu6QST30SKgLq1VjQthV5bIVaN426pHFPsAhzhjJAHHq5lJHV
uvuhvVlxFLE7IxautdkO17aHhOs9peEm5TheX4P6xAh2s8m7ceFv+WJySg0zRxYg
ZG3nT5swj25N0ibd43v1dGqVs0L8yLBDoleNgtMN6BMq2amWpw1RNe3cZW2TqIqD
HDOCLl3TNQHMpLDW8anoAbPqdnaQF/MQvnA0D7lbXNpsYmWD/8pq+j3IVuUCowff
B48oSbppnuHFicZC35cEcBXU/QMszJ0bfn6pxKdvy4KtAcfoeELQlv/HZfCSmlma
1JBJdaJ6DQwptC1eFihq5Rk7KV/WOugB6bvqaiMnITRTgxhxjrjP83mZRmZiz91C
ZiB8Qwwx7jR9PxOLPh1KznrW4GiCA7ydKJ8DP1s2RPaoPQTwYxGj4/eT+C6vVZQO
vR+QfxzdpHKpls6hpRl10wvUOxcWP8jlYVsFCoxho4+Gv5XxNrcac11rx6AMS4CI
WN8U3IJ9ar1fpXa8FNxKAa1tmbS9Nbs2ZM9MMzbohP+xEGu3WYMOpGiH46w6aZKr
/3yb6Jf+q/O/T7yXQ3zHu3/fly2vTBkQWWMFtypCLmjxGSfW0YeVMebjRqr1fVsH
iBQc5ALraJoo1HSBh5Hv4o/P9dfgwWuDwOl2JUwNJarFzY2UfzGFs3GLU4iKKjDi
bYso/FCnBrS3vh5xydSWK9/wmyn2e+4hRtMpVonG46dHU/nRUM49pL565xNMLK8R
4fmLBb2x2HY5pOkFqKWTo8Gcf2Ryl7/DDlg2L9TVbW47vmFppgA1wCJ/dhVihzya
cZKn2yBMH0sWG/pSSA1QCfViqefP+XzOJ7+J9LKhOZggTGBC1MG4jT+QYr9/a8sf
kSi8Nvn3oEq9LFqV2086CXf3+CHCvy4dE1qqMslReTYuEcXyyJpmZoq2fxjM/fL3
bPoxpDmb1LJjaX8sQu2dRiqW2UNcK4E0OK6mhoNQQN2P0DSUYnAjcCxgKuYntYyd
McIQyt/WSWpRGi70eMbrEomHxlID+8jnIpqT53OHhVJLdEFYlzLBciSl7YTBJ21Z
uM74szcBk10OwYNiiQMepX/d/xhawpB9nT91LfDIi9MOw1qCcXG63ASnAbrnbzvo
Lvy2JgUtUhImgFsQ89W6Ii3vQM7tbXJvGoSlDxKm8ksSEYFEgBR1mTlM+h4jEuIs
xnGe6879wxhIgFQe+RMecWY61Ugfy/Ot0tO7NKj1ME2IBMHm0guuCXVo5AIkjc7I
nS3iPRTMkeWTx4C/QSdKG378NNSsnHVJeNzv2Vjy7ontgapLL+cDznlp1uvnvFyi
lOeV3Q9UAn2C6qImRZhRxzyuB9RpXwEC2kMwdDCi7j23lHKWBSk9eyxPH4iRDXuY
hNZI7FftZJ60Kd/5X+OR7/bgxcN4ZrnppKgHsTgFcj6Wtoco7bVjiXE9YgvlL0e6
sM5XICa/wP2NEd02tTZjwa50ibAnYY0bn/GaUkAmOvKeOhvo/0kqnFZMFM5ckNCk
pfe/eHgQbVBvk1y78nlxmGLmwBu0Ae+aTLhhmi2NR0Fvnq+jbTJeQxSvUd2zyAcA
DszuCLm3bHjws8SOAX9mFcb67/fuWR37hYA5KZThBN0YE0myf/bO+MPvbNqEVoJd
NjWVDL24eELwpi/bn0jsvq3d2HJu/LMQzXA5d06Ms7dcnF5rhH9UPxfyO+Tnhi54
x1dr5ukv+NpeELD1CmhDM91MaJRA2l6nEDp5lBfkHLfKoE65+I4Uo7pEbw5PQaoE
QEA/mvst11KIo1f4dihq+Tih6cqQR54WVRFE/DgYCzmxkp5FE5uTcrbpZPtMTUwN
RZxaL1hgy5p4Jqp+64smy4SLgQMlq6BnvHfzXJ5TAHXKMdwlhiUX17ekzj+0dwU9
AMoEoCxn0sajVxYkKBXVCBiqPG/LEkHIMMxOc7Rr6NBospMxQ1VLcdLrgHyAqXmT
VYUKj9FK01ORqMa11nOb8Wpji2PdTmG+bbqWoE3mppY8xMczkXq19RhTNgdHG9Qx
2n75WeS5zsQpSnNaRHM3jbFe6o0J1ljqSIv6PnrdUQmRThNBQYiyDeiA2HeQ/FNN
N/Zg8CHv9A/zMkCJUAXFyadW2WjC7vKeLXS1YSN/1fyughj8rqRJprgD3OHgWSxT
HDnnjwy7wzcO2GkaQpip4cLTSyv/4yw2N0Es+IRLMhA9Nz3VpvW3/J+ASExEcGR+
fCKBBjGxZ42pH2+K1rG/7hZM6uL61I4moMXFE7O/00ZO1MZEwzPAfmd7qlgZl58i
uJOExnE17ZGHizl4eGcOuGxY/VHfaJFt0N+KihD3BDgMDUqO9Pp7JML1S2Kdd9LP
ZRikLJRl3mgUoUzcUdAfW051z0Cl/FQeUKKPOF6A2S6+wBKt6xniKhxika8oZlNG
ASJE2pVU7sidEAJl/H31bE7pd8nwvkVG0QhnXqnqy3RLY7pgQgY/JSwvfjXSj1lv
LGaYcM31bEPL8Zg0hh/IVUHoJPmcTgHTMuZOeEIRBegqxJfctn94A4/X5Kb6Thlq
oeS0WY18bPLaddOfUPnFmJs7DswVnj7car9TW+Fm4FnK+EjasWVHh2h4gCZZlQmG
qjHzMDaeutZEalw7SACLfaTbzKBfb1Ps/UgfsouOPiAfaoT6OiUpsuEzZ5ZmNwG3
fIizvtA3qo9Yt9/DILqfpXy10SiDdZtN14YzCIb+xG6Lz3ABcmqo2POaj8WD8Ovc
Qreoqc7VNqfrpzexovc46gpdAVWNssk8S2qfv6dvSZ3FMEnmPMuMzkjZgNrfiR6T
deeRk508QsRiQs2Nt6PgAPI7V/jM7Mb3V50KlnYbHnl6KtMu2vIYwC/Iw7wBA/Y3
aIp+o4TLjdefXIbQZdf+e5dt9y1PyjOYQIs6BcAtNISlUoHxE+3IiaPMNaG4zyhQ
Tk5i8IcsA/um25y0kXhIQF7M2xun3VT49KJzqfGjzLBYT5de7GtJPP1I0u15bCHH
YaT994G8VCSZl8taElf5x2MxZp9m5bf1aplsrpDIaxLUaE9LqLTk2mmVo1Kyeanp
JK45ew5XuTvif28iduwiePtplXW5Hxeqfyr6XZeamAKD26sGoo7AsfjnfmaNlTV5
3mWHXEKT6FblrsQewL1WeYeyFU4m9iTWtRH69wdPle+sORBk84Yon/fCW+8saUUe
nivDtEGNUqDrnX/CCqTGB+9+2+DHZ9mK089kLh1L/eywTMD9HjoP/vOZWof3VRo7
6xGS9HbwNLe1XbQ/MHUDocH3yNpzWZ48ESCh2fDs4oyDdge8VLrauTR1hR3h8t4+
FOQm+0MNtGv3dutb0pbE7PcoGEGY1K7iFVYEnrsGmtocM32mq2rdzHDT6CUBjqJH
/1hBoXz3hhgZ9bPTmEDx6tVZF1DnovqOR1xWbo19bQj7xSKWAk9S3CIJAyn4rg66
yOoMxgl0ClV6ECoijczEXmHgYKJX2olU504bAyd9y6H0zDTkJ+sLcAWmeyi4SBVn
zLRUZkrBVUF8y03RV1+DBZQlT5RiVx8wBOPmo6bqhvXLovWjghim2XsSSNUex5Kn
rZfyAyZjXO1vAVFL309FvhsRAN0YspDGyXAsq3EEfpAQDagxgzvGtyIFm1GWmrJH
IFWBhfrnFw6f9KS5Xmu5fEj1xcsAP2JUyVXKCChxyW2rAIwuYbjgiuRVnlG6mDFj
ZEsnJHvJxsPdYP+QuQ1MjI6wKy/m+JU0UYtgbeG6vk0DE3hgM1b2vCd7VDLTH+QG
XCI84VNg5DkNkGLNhPW5l2r/jEpF6/b4dCFNCWao08CCIQ2PvWLbPK2g/P74EQXw
0amHmp/GYXy6UUaE6oMsRZbSNmocI90oTrdvMy8KKzmzgNGSmGxNFDiQ3UIifFRb
j/Hb95gbgrfMMhGfOYIAVHGgG2ssKF+burOaS2S2P+kjnax3A2B+s2x98O3o910a
AEGic4fS1zda+tYpKbTDT+5lOssv7zRcvv0K39CJ0ne9neaPDVny6xwvZg8vfA3J
BHVVv7mNzKmGwfmNP9ZggprgHjgBsjdX08TWS7uH8SgtlOon3aRlvIdXc8o+9XKh
hQsuWNKoSgl1tpv6vgwzFx9jbE+OssDxljigVR+rFLqUkr+aq2F8EUc5cORobqO+
l6/H2tDzHY6C+VC/BARhDoup9jDqcSFTXWDrB9oEZtjHYiBys2/DztgQJKApViVI
e2RmwAh55AlfT2a5OqJCJsJCLUyn1aG62IPiadl6mslCCp39aBhZ5ayxCVtjX41q
PiCJKJYKejnR7R6mO/7rZsGwkADbrje11kTtj+Athi0tvLbt6Zwgai1V8LcEM2+i
l8N83UNb6FN1zGTXHNrsBmiAX5FBegUrjLAwtt8q7KE/BPEbDBf7Lq4bs8k+yzn7
S1TXz+uneWVF92nH/FD/uwD9vaP2t/4z67yrGPXiGu+O0sHtoqPDZuq848Cy+KfD
DvIAW3podMGxLphL+jKw4ZXdtt1j6ji5J8VZ5yodSnxbCAy+Iij+R5vUflPZBfrO
fKSGnGcRiz+aji0xbq5PKJIsuqBEgeX+vLUbCVFC0WNsy3dtFFnNvlqaq6NvjV9b
sQSAi8ARL53d7zYGQ477dYCc2NrBHrrvhE0eT6Fey1QxFgybRtUXL5poSn2ErJxz
SxDVyIVBiyHvtB8CWmxaLFmvh1qzzI0fkxwYpun256u1mrGvOYE5xlK2fDaaiaup
hu9+cLcqn4fI9Mx2M80/yzHrZaz2ID1vlo7v0llzBZoHnDw1ckJvUtUtV0Dw+7kI
idnlBa64UGcj58CdzjwppwjTww564zT933/b3dCD0xfZCojs2f+W6zSTfue7GluS
av/rvNjEFf2z+gfPwTd6Xal1aiWPqfOTXqENxHKByUNuF7/ZS3hmLk0o3rEjxnRV
Vi0NLd8d9LrFGS4X6k8dcq30IdjejavNE09YHODF16Expk5jUFy8+9K2nAVsfx2d
SymmlglmaSp8YzhCzKeRXOV28eV6pn194PwT1PwbzJ6lS2uP6Io5z9iXra2anxnz
hHjvHpW44ocO5f8HuC8GzELNhQG2pmlXp+zqhXFxXSzvC7qd1d6X86RlT10/RJ/S
tWPYnMxPkVbzwCxGvIR5c3YE43Dvr4GECOGhkWv1imMmA+bp9FGfgoq9VNOPyw1S
E8Q9QoGbymlZnzvQKYuOeMnxSH+xwDpywgy7l1hL7LNX9Smi8cZU2iur76ST+UrO
3hltkVBeoLwruFiuW4fieWPHsizEzMDnMbmzwTxxysCcF0Hqi7S60N8cSfpT7IaP
RizkKr2Ff1OZISEVg4T4zIAlrcAPNZ+Cu/Ko9Vdi+jesIU9mp2U5wpGwZc7V2H/i
p03+wboZbNhXpEiWQ+PXfiFC4jDK+AXaPDV9yrH7kukG10vB+G0YH4A55K6kMsYW
60zwqVRKHVISQ83ptTYHXiisCeAvUytkGKOilMB7F+JeYjChHKh0DJIbh0cdtu0C
w0+g5ApHGc0H0wo/uPwahWyVw0BRHzbXNQkuT6hsl+jM9utbfiWjiFvFtgsw3pvi
8ActHeW1UCoH81VGEbap9MohGD2QIZrSUf3/h7Rc0mON+ZiPv11WuDFlh/mpvqEK
q3NhRl9OMjFfE1htjvfNUxTtXFQOX9gOl2JZNMCRjHu5fl+ksavqtUZxD5dquPQ7
3iiKmRWlQRsFNzWgjK11wOJ4qik4tHH0w5CLyocihMi0+sqc06gFWNl3tNqp2iQ7
xafSs749l3hCzWjwnEwsI7AxTuw6WvH98LNBXnY5iQy36rVTYMrPdH+Jakavmg6B
M+bk4iizbWVKruv1PHUnpPj5DLaDuhRsN+FuDbQ0zlwuB9ajQofAr3AyyLLR+V3s
zLAN1JwvyvzpCdao6v9iIlOlexPJR92/QcvRp6c9OyJpyNvRnIC/xhDe3SvpJbDU
tSB7O9+kb0HkZFL/BmqX7Cqf9Xp3JeFgkcSM5NRKlZlyeWeY1iCsk6GT6/Wg6EPv
QuwT/ycFZUh+FGiO/xvds4dUULzKOk4TEPhAsntJjxbfygXuRcBbX3otrmmqW0rU
0VPR9PKNvLy+QR/cARjz7wzVv98dYNLSYb2EY8uEPnnZd6xC4YeggRqej+yOjPNB
ezTUuBBwcFI0JtpQryGews+8k5o8MeKqID451HekmWYTclBQyICUcXyH705GL+Kv
g7gZocchG6dghA4lLbR55bBlmZ4kILqkLepQPQ2J/H/sI1sDXajMsmheXKN+F2gc
XyEDebO6CDymdGqJht4f3SO7/xWxKk+80SsS+kNrN8vhuC5Z5PbE2l2fUfUhYAyb
nGKzKcpDEaQryg9YJlK203qi72NSXt2HnJHVPvJ/PYiJ6k7rSbXBhH7SrU1Ag6ly
i7yaXvlbhkxnKZDnINHy4Qs5LMlOaoDfRiGP3sr7qg5w4zkDlUZmEycCnvJnBi6k
zPupYCmPgUeoe4NmMev9yJ3vHXX+NWUgOW3tpWLWiRGRxbrZzv5/et+gpiLSBBbC
Rpb0nxgYxIOSD1VElbtTFhI/Z1VV07BqpmZg9uHkkvo9HWoWjTOD4Bdk9YyegYHn
WtmPThAwTcOQsk0ydKod7VU/3mG84IEoGMNZEZqeL7puAq/rRGHduZhP5jsgKHTl
iOgvsBGiqS2pkBAui/5ZerjntTWUnkuCUe/aZnfCNdzXmen87UP6Fnr7bgwUXjDe
ObZC5X6JW/wDvoLJb6gAN1bRh2OYRszf/3UwoZrTifG1OAlvBxStAtOFtMLeKp5s
6PP5daZ7ScAaP+KenBqSBLnSIStJuU0ZjOJX/TwBtWDU8/IdtDxmtfTYnVyaPIbn
q010fl/gAQqXZ0SJzha1Upvd1YdWLaH9+wLXZIFlddNDFxCA5OmfWJ5Isq5GBFFg
7h9E071KCRkwuPI+0fPDmENMAny34Ni/cpiAVKcNKjo6WND7TDN00AWmeqofbqjh
mMCIsFpLjB+llTnh7MtqC5E+9Ym5XTQF7rQPmkDcWuaTH9nqzgeb/vlAYV+RBDUS
SiUQe/rxZvR1SiPOMYsrwQ7I5/SJ0fUJPFSntCYwqCpDThEn053QHubxlndl7IKn
W54Unn5VETKJE6DBamB82ABi/504aZ7YAlAM78O3pZUriMZVsZ0PV4D0RNTsbm7S
bBa/wtHLe/yBZDu1g+NuUqCfVMOUc71qTIelzUlAcd2tdZ/R4YM5NMDXSnJ2W7lw
czloz8M84+RHKa/0WPW+0btRJBmWyTPyZwP8M1ZmnCD2MdNhQwHwGz490s5mjAtI
6dKO3AKvOtjWAiGbMz93lj7L9/GjUfT55wrWI9j97iNAwRwwWCem95yW/Q/tFn/6
DMxyTDbCx4yDRhzzVOEQAm2oQMtEMZyk9bzWd1HHsxmb5NAI5BpA/780KQrmGvY+
nTtNtMvdGhDAofCfbX1r2Bqqa4SLso6JGaYHSHuedM8yKRgXHPPNWoMJgG2amC1+
FqxG6+OM57X/kHBiCsAozyA08m44dmgIGpFtUq9l4w6A8kBjPhulUe9zRAUPoPh+
53Cc4GDNNsA0vc3KJBLveZcfxlHTNpRWmRijkacM9SkK3aMAkbv/4BElLQi6ZgpH
czEkP3ts7M8vCKAIqTc0cYwyv3sieDYH/aJ8h75ZZBuHH8s8EOAv80MwqEOPnER+
auvYTlHdT4IgvVSNrbmqJHr/Htg/XfjIiWIAYw7xBKQ6tmzzY3fnosY00W+yszak
3B7o8/7Xwh44sqqSGrTxgBx2wYV1tFHUNKt3wP10EI8M8/BTgDnn3oBr8kMLttTQ
FfJQ9rybxzpVWmb5xQ/ge21sh+HSL3HRdTP5K0mw+47ZpanY/KeCqKWFV7Gp4LWx
uh5gpygDce7+PsVQISzpneSxlYhTd9p6qydVo5JPbCAbPwxxYSDLajkAQ2OiqsR+
bK6Uj4y08YLxaFCVibxsWXGopmHBfvMjdCSxvDWphvo53V62Pyap1PyhBNcrtuen
uiyuT24pFSqp8K/hoB+x4UByaIXox9mb9h5reEw7NtFENe8mI5A18NRn1PjSHxWr
ZWLSS3dlvJhxYWG/ZO47+q6OZeJ8R+5AYAc0R/8nZug6tVloup/r7aHLpl9TJDAS
lNaV0LUm9bbyk0r/2nCJ/WaU97Ge85QTUoA9ihqOukiTG8trscUDeuhdGzzLkVCn
GnZvvE0ygg3EU2X1YpLunDFl5dTCQdsqvQeGUQjAyhl4xl5/obtluaMKP5I4R83/
+t/KavQcL/uK6Fb7hsS4poDeysrsJ9g3hFrXCUAlClXwHchAGrl+N68Sv+fsFltc
7uDkYF3tFjrCOQBEunVlUVE+bSso7/otX/7OZ78P2XkWL7F4qzmwG/tPMVQzUEXt
yQid3AALvr5vCDzFoDHv5hBdhHlHVHcEOp1xIEcGX7lK2wRVGHMOd/mdYhSB9X8F
vM7b99b+cUuSq3UgMvd7VQkvdD1+EUTFHO+u4wICw1nZWJBBWqIE/jcwlM+4E7Ge
j7W4xhrlKaj5kgDCRDA1oS8pEq3eCCDVXYNAvRrY3a7jxVdBEWJKQDaIFLJbnyWG
jmTNjlVb6B81NwiY0C+L0309lDsKEIwhALgmE9VMbIcCbWqN+5VMo8bmMwCRY36w
npGcOZfO5Jx283I9zQcvqPOtjrta/oQzxQctmnkg5rHuqxsV6d63RGp2UY7iNDZJ
wTqCygnIuDMzgdwXxibgi/eZQSBsVwK+4kuFnnCbyUyl8fnqG6S2YH+niLTo4k7J
pJ28g8X+5h/g2GXs13z3eexM3VZ8LbIslhhfQjWYaDuqFf1TibKjCGJJrGE1Do6C
O3QzxFvXtdKH1GRbL+z074ELA85tQpsl0+854jjd617VFOU4Uv45up2PCrxlNuy+
jiYS/lRRBxVJpeZwm233oEwUi66AgMvoc0SXNXz+vAqk+AGxAdDtZkBGIJ7Cyo/i
V+4y8OixIr7fJ7lfVhSfZAU8OeW2qd0sPX4e4eqDjR/W0u073BX+e9d1xBI//Jp+
h+hwoZk2AOd7KP9uEDK4KCLcUAv3boWBH1R2jc5/+L2WgphZ8DGlX2SPXxUjo0+H
1ksE2p1eSwLKP6fXW1G51eAcISfWenVPH3nNMcjUCk/6hFoeZhgryIAj2e6bi+CU
fbxhE0unCwYiIZSYCdrsQ1FgGMbnMC7hUBeJ3rAYoiV5jsP3t2TKJQj17Ympkfsg
df3UBApyVnSbcZGdD5QfKzSJiMVst+i5Lb8q/edTapOVLMti+z0xRi7M2H74hvnp
pCaD5+PPiWpZvGdhO2iMN84urhW2mIS7y7U2xWYqpEjOXnHdMxvXE+BcwqJTtNGg
kE3p6475Ek7Ap1VBn82D9m4cUQCRGa4icyuBj8eyq7x5AD07rAAozZhed29+xm9q
V+KyFFoV7OZVnac5QMrSQAWMLtF6zE2MrGIh2gJz6o+1iwvKdX2PiQkbmIlaEBAS
qZgsViEiMgNfEEBgwNMM9O/Mw07WzPF8C4ulBIpFr9NivUL4nYlZPtOY2yR7KH2S
jyp92oWjEgl1uA7rCk7T72KeyVRXcUXL0b9Jkozycns1BYwPf0CJYfL7fRWr9MjD
iaUT8ul+OfhbduNs/gqKmyvyzudLp0juizthugJmOOxAFUwNoCFFypUGEJMdPHbt
vvCQh6ZKhP/Gv0dzWHUfJ2IFtrlgrziWBCm7VCI6su55UcRpypmm/pN2MBtZnW6r
GJb+p1yzmQnTPN1UG8CWDpq3Xo4QIGpFXNQUoU8AxM441aClOAzor2xq0Ttvx5zc
Rurf2/sh/BBFxI5/QdYzJgn6Z7VTVYwWq1QwoSaGcY239pGamaAV7403i4YZXHnQ
zV8BI+kvMYZHmEOHVJB69ijAdkzOv3ZvVeNF+2mwJjxchPr7/X+e6DwgmqWEKG6m
/FDiyejhW4vPuyYq8JF75ES8L49f+8dEsQ8U5KCwGeDjFpqhRWcWq6ZnsTB9p0le
moSwL55CNg/7IiUnMK39IkaWXOmMoKsw0U2mw4+aG0+W0LG5WAgHye8kHsnZ7gMf
TXNb5VAGvwEiGLnF562aYH/a08LI5h3HNN61YR/nkKC86wVqkTVR8i5rO9qB7AQb
bs8tkAhRvU4rLo0r8NA1MWcsxxqYdMYbrBFqdA9/cQnVotL1DYuohGXcwFIQSpsr
9QmF2y1K3pbfxCTbUWZ2gZ2eWbRZ5zAIbTKCppHcOQ1w4M47AewmsLwhxPg7fHy4
4mfRbyi1OW65qto1C1O6hE9JyRW+fquENtbEP6ox3qzjNpWHsc7JDY0QbWJjxYyQ
eaAyj7ddeOGx7nnRY8KqT3ZCY5y4DTENZoZevwDnweegJIFwmbPPhiGUbKS99+QZ
hM8rg0TlgJlQV27e1VhmKNXRJDJajWcS8kRH9dP5nGCdzg0hGcr45W4ceyUsQdDv
AmbId8PCvGrEd3a8o8kYSOC/wYPpUNHDGCCSUmrOCCkpLVgbCEAp6euO5jC+Y7f6
A5n6FMT1bo0FdIB0iXaNE56zPEAoDrkZ12/XXFSJ+EFsqiwuY3zpbbsRwJ+J6lGf
aDLAG1HlakLKvN+2NkFMh3UZSlLlHsihhZFXLnuG3XduuoiJOqDpQB+3zfHxgPNM
UALZ0bpW8oB5JRlMvBRqERvBmUf0riEtsZ1WWKD8hkBr1EDjhVsWbKeiVMhT8+KN
8VXRFHvgRWdkuIPC0IHmgeTKJcAPShNjwWN9tsegpZa1GIrgVbZD7KCg3YTAA2vb
UiiBrIs/EUXPmVMiOn71M4oAJTPJwao1jvWvG4wlgDQEU30CX9lnwM6gZvjJgbpz
2MBZB84lK/DA08JzMORoyaJQhmh6OI4txgENWTGd5jqYD1d0Z+bGmrEWpib7Mr3E
3Az6EccFp5OI5tXmDEQyx7t6yh9WvxbN1WatgwdTQLTrEjHoy9ZulKAuU3SSvyv0
p4oPRn76cSavFDZGF+VkrVeSFMb6aHrWix38Hp9llar68OF1LScLtc/gl6IR4uO8
05m/4f8gV8m/Bw3c5/3cpF/XDWFzDZsEN6YUIp2+UJIZXzuqbC2pUvSVBFHNbhlI
xbjSfYYK31PoHPfw+ugyZ7oAW+jpCUDg0UXtIhP+kSlG0GUaFd0efbeEmCzNCWIv
PbqOIjdOZsOYHzcVYCV6+Rrklubt11tpyorcCjnGFDKWdZYcLFfOsINaCQipJO/2
rGEOuODfpYaZSm6r/EMltXf6qY8TbHG3NEGrqxEvEUTuXvGeE8GGPTMphToShtL5
fgP0OO563cYkZmdNaoRq+vrZoi03XAvt9XXcEOhHq+Zc9itmqC6PrSO7bLINvqLi
o7fCa/dfflsQAwaLwHpX7f7jzZUbtJFrk7v73Iimax+R4FQcRitGXeUmQQU4Eyfx
hvX5GMhxKkKSUUX8fD2HO9Wq44Jy1LHu6mpUdDiDhWmraCcroDjyNZq4dv5xEeAq
ZH1WPREkQRwUnBvLXTXKrS3tKmDgXz0CjiXpXNtJT8AJGuNvYCKy5TDGlOuXN9yB
vPsA7+7p8SUZnlzS5zW6QHR/0+Qp0KNyK21073lbErJY7SvTbGnMmWxNoUYZ/Osw
tVmNKhfkXi0/IKDnxJU9KX/4jzOmm0M+rYqf8UMd0quc7FH1fBoohDsAkz5R3djC
WPo85DT1E/HKD5MEonIb8ACBSG50sHiOL7dPFQ3qvCTHWxBCiCMOvApgD28TasNL
sK1QZTKj+8E3scekSxi779nQjEBLnhEGSuEVmqYNdia9U3E0x0IBGFmvjeYmpTRD
OkzuVWO0zJPD8f1nSCpeYJw2b/K0T/RVPg9qma3Dbdrx7wA32nk5L/uKckbNlXNV
e3Gi9Q3skWUeMqigw2fhNFPfJ2FVfA4jNE9UjaZ08vdFlXwaYIk1RdGfQHiaHY1O
q92EvloFrHzuFVfgrD7CPscJYYYEtpJ3jpixKeOwUALpIsu4EtBK8e6Dj/4bLlFs
dGMpHFdTUKqHLRqKb4c6oQxQQTAfSYZtGfipWC0AByu+cscpgQL1+cYhry4EkSU+
UcSAYxHrzHVMeZc/ZGvZRIuoweve8IMXWS3RPbISM1lVASO/FXuWirA5Yv1RCoZf
37c09rt/dHDlsiaLEO0EH53qTlFW2RP7HlNgQhG0rE9aiRtZeh+p7oUg1rZGds7/
zFXfu29skUG0DjaVOizJ9POG8tUvr2wZMFUMp1gpSdyk/PvQyXXNl1jO4St4UcPO
g7+F+NwrFKYA1YGqVEFfKU7gMC97DbdLnaYUIDeyDcFAZgm8KjXe1jhfIiVL/xIY
4X2jFo8DpkfBKQT2CfrLFLEFv8CsiXpl/NZmDmDt8dmfht1EPTkIwDXJSs2EKqOf
tbRcY8adkamm9dw47D8brtatnuIpyZfniVnvOwnAmm6aTqfbeCu9C7LNLmZK3cXs
pFpTNf8pQsgmq95NDv4fCsgwy5IxnyFaVp8i7OFXuuNHOGfLYh0plCWiwz8fGF6w
NFp8W9sc1xDW17Hmb+jLopNoHooGo5LDIvurz+whkhe6A9J58N6f1rkNMDupC/qS
vu7m6IR8/JoL9RVTtmpn9INeuwcl9NltK7mtTfBLwlL5htATxpuKeATKcAGF2mFb
KRdhk0P3LJC/AyYsBOsya0su4j1kzOeQ6E4s9eWZiXU15ZUsXcFwiVUYYKPEKm+4
pnx8dCBa3G8yIVQYv2wDEN68wT4cvQNO2YcMHMh7/1spoI3E0XS8P6L/79Ou6m6S
JOXOqxcoQiGag+lLdVLpvB6otRhomrzaAHG6fYStVNy83qldSIJAXS59oxsFgdyp
h6ntpHv7wHjI3LCVdJX3f6NyM6qjt711XLr0Ap4dLTuwcVidIpPMGrSZl/SvTaYI
qms536UHlx1AF2vexqMGIscaq5Lmn+ZQgTBEX3rYJt4+Iame7bPII1Y5q2uthmWY
Ciwl6QOAY3TqiUndwtpVHTWr5DUqO67KUCeMsbwZmbPkbus1wlPjM+bvXByFlzXe
m1zAVuXG7J+JhkkiqgLz/wRkqkS7MQISUgp6MM4pRv+QdpxRdrGfOQsczcfmXJnZ
FpmabDeQcdMY9PIkY+qvN063v3ruNMQTeiOv1QhUTghDggcwJDgpHQ2LR/mQFpT4
9CkVkwWMqjCL8MT4IfvZLU2jkVAKutu6ArPWEKxvtS73c2S4f8YYDeO3GoGzvjkG
GmWp3fv1UyA+nCLbFlXSMkg6KQUxaHX02FGcLaIk7mXRwCtyijPHDUJPy/HPXFQ5
oFVDEV7Gkg+8YVPXDhRs39aNZwgIWGJD6h8SculxavusU+KoIMoo7KBMhBf0jxR6
Ik8TJ6BZD2dUgceZ02LnbinPdb+ZDjh2ePQ0zdvZTMDz0nWgVaFcZZ33V7Qgkyp3
gk+P+bJeO+JVtJrapyQOsz+rkqXyYRHW9iTlXIcd+sy3bH4x+5zknMHUtHw5owd9
LTGI0m1PbZLZpvFh2nHnq3UpE++u7fTgPRqGrT95tgaBKaA4oWRUMfGEhiWsBV1M
vd6rodINCJVYSB12XawOO0ojDoaqXFBory1Bvyq3l+nWEFbQjWGcDRvhiIrBEiGC
cOPKAHX1VsfJ8I/vyYoqOLLDlzNQ5biazjWc9GNPHdZpa2Wn1vrJmBIltcNd+mwf
v4E+r57TLSk3XW8kX6ifuKt9vNdldjITch8/tjvowpLZb3BvhLPjsau2xkv28Nm/
8PUs5sny++ZKyEtWpX+F4+I3rVg/zxyIpojH4D9i0TLeQNLVwZ8iMNnkAzNTQI78
ubUUZWPtbDk7MDZmGQG4BPsK0aRCE9/d9es02EwJ4vRZCmGk1Pixp4zSkzFpG16Q
7e9/jU1+/I/aq87et/GDNAEd/jlwo/SJz1582RmhjgiYIdA/xMqimiIVkc3J9qdt
5l8b0K1Dm/3ndQUO/N3zuRlbGJe+JlCJ7vnIgmVMKt5GVjJbIXVuFdq1mzzYGYKG
4fkGeuDgSnEFBxBcRLMEefqlbb4DqI18pzPPUANT/qyk+JpJMlWxL6PAKWrLsitB
kW8/3OgKh1899xLxQUhl2vBVOd68TaiClOBfKDdzdweA8Qa94pyMrOxD4QdwgxYa
Rl0vTztaLLy6/X0DygQ1A+kipvvaOx9uSi8pNxl4+Yc/VkkCUXh9p7FfX8X56p8O
zXb/DIjimcq6hkjdm9p02mfzZFHiBDZyQMifgT5fkFVNSgLQGOAIaRpqtZ6NZyQz
6ut8Pjn+mcLPT+FKgKAH5vVLR4ZJo+q8R0DELgVhtJ5hdIcfjrMBfGUbem0NRWAR
6EC9sFKSOFcvyuRCpf8Cx2LxBQhxZHOwHM2U+pgMZHC2X0hz64t5XgZPpxH9U5a6
FjP6wGBpwS8pUPTWjJfI8YJbKQi6FrIqbSIKj/WoEzfKxLX2uNPwKuuJsB/DqFLT
P9q3yYktOJ+JKRuybI3CVWlnKJ1hVngQiFaJsV7xmRlQ8bGK+JsFTmYOue3tCix1
fDEIRf7sd0fP5CHUOme75UDKHMr1iYbU6t7e1A+7ZRC2kpW9wJXAH/QYnHASDrbt
5L2FzTMW4iKtTjm2FF0ciXHzlBiLokNNwmw79ozoHoIPLk4m8O4Nd2msXKNlAAxz
zcvGkJ/OPKRbL5rS7DGfyeTxMx58mcqM131aUqrDTFwKH2j4DX/9ejjoXTCU9kPL
AZ19JeN7FbMHe9k4aFG+pRXfcUc6ZY56wiHF+6mYtGAGzclliwU8MGaT+ej72lO5
ZU6cqV2rbGenresTph6jGo6eFk7XUTUG7sqQGLB2QLhAbVmg8wA3YrNLFkhp3oL1
MgBLsXSx5DDRmoAQzjpCFbUWasUzmHl4D40bfd6BhLogF9J8RK3E/DKgdvY4A7/X
+lYEOvIhnKo4/VibkJYQpGyR1vCGynPvNtrcI6YNu4+SOb4PckPd3bz9FxuuJf0t
WWutgd7fu7gSz0AWexv1g/w0Ea+x0fP6y3ksmPrZ1PlnGq1SKkwO3F1STq2kOKvr
5jr2qwxJ0zkgjb11bxZMlwPWb8xuk/0z2J32TB9yDeoNF3h1tLRaImPp4NMxMGGo
Bq+WFDBqsEjDmiY7JtOn3Qi4wLvfqnIrMFdf4LgXtbXmy9/jCkDHekxYVLFpNSLl
rhBom3Oycb4t+sSynwm7bdEHaFtow5x64w+eXZatPhpF9l8ASJCr+yh4EdKXfAHA
pEWqswkf/6uQzgBhIXU8EC//ZO64lqR6iNbLJYhsKiiiE4Q7xtnqN6jZVfMVKSri
NZuYQZaIM+SoUJLmkqN1MGMk3uvZRBYlq4PkJ1olGJyRXZv46Y52iypWr+bks1Vp
TOLs8JlUAJa44oXAweRgBQB9v42Xfm8lvTbdAbk0y65Fn0O9hT9nXQrPtR0Oo40J
xovi9ql24geaDK66BMiwXrFtt2+oPz1ThP7QbBfqpqIBZk6qUK+tUgj+av/j5cvq
CprHivwuavTTi7wapja01tO7+Lpmb9J6aQ9zhfWuk35fqka+X4rCLv++6QkHCneH
DEs9LG8290kI9MyDuMiRkUMwtEk5OY8R2fCMtvq+6VLqc4jyf3OPiBiNRh9M5Kx+
F6H5fntxeM/36TRnDPGrvyMFO+UHdBhsLlspUl4/yPqqgtCDmzL92mUSx/e2J8m+
OW/33/QlacVherOuFRXkHWOTsH6yRwJRm0ToJITTiwWxw3v7z4WJtCWWKVkJsi8V
vopdWGoPB0QUsuSfG0excsbBbFZkNHChJGCo8Rjasaphex/9ss8SPMA4NmaRb3vD
agPVrz5pENtESipkAPvfZf7h3pnMIIwXmlQ9OykToKKjFSEEGqMbWPSYuz6UrPab
6TJ2dv866lHsXZ873ehnSSgVXz9ICT4k4jlTXwGAOmHIV0ml+bSGHt4oIJaPlhsr
Wyl4+Ay16hV2mVuRM2f6jhdWXEoRhKyTv4trTE5vE5SOZOcNRSfKe8WtXLxdyoPe
nRb1wEk8nHVYa7orXeTGFHiQyHvzKx/t3vFnPB09EUjNGSZrSgxvVizyp39ZUMuz
otejXGV0qvr40EAYkytXRTdTdssbu3Xw4sI/wp5vxXuFZsxZN/ru8sFrRFHjcG/P
PA9g0QfY0XBybyfwHrdFG7eouR7I5wv8N9OTTlfeTL5W1Spsok+ha/hXlzWnUvhH
NHjtfzz7N3GJ8+ND3bSdbgbWHbEII60w/zqZLneMOfSUCJbNAxxkwO/Pm6rzABpi
KZmbSyWM2jGvzcbQ0mAoh7gqb3hAXSojzf3Nj+pzlXstOmy/reV7dzqVpXawH8K3
DnTwyPGKeNMUrVIFGNkSgck/FlHe47v6EOU9q861H2LhpaFd81UyoNIp/UxFpXIq
nFrA8aB6SWmlCa2ITYTMfhld/1xGT7vGjRJSZdVm9IarLVV3L6fcEIHSX0tkj6+e
u75JvJduWFZ5W9tN5T4BFhwsUHc0drBkb6PdYonTqyearL9jFk8cQpkdZcZJRG0H
lU96Ps711lcobjnyKMh9xi28Q45rQFiUIr/flOy5Vfx7gvJ0lACO7ijIzoEt9zVI
OMweJGZIWUt+GiNTUtt4mufgkBMmjFf5kWbtbfYB+l5RZlNF/IgkbklimUK2jp4a
1qIeZkB8uVL5MZZRIsTQdtvZG63KHQ+rbSeNpsRkMPB4A6Q7G4Sz04dd9iXYimpH
ykehwe+dsVgWdAXNUBnriB/68Nqbnm8yf43k3nvZ4Ze0EplTkHpfy82kxDI9Wlxe
ehzMuqyelBVXOQgpuj6i4tZWgdMPiWNxe8HlGsOEjWSFfJBg4rOlR3+onVTwWvcG
8V9lTlrpgzuHSvT9cbXwzCzqyLim9mkRV+O41jxMLema3SAf6KkXAVm7OyPDKejM
iO6zhoBddtT3OnKBmrAPxZMvHQy8kCxYd4UuRXeR3CWGI5lznYMCzE/6n3/oQWDv
wzOZtAAYJYxAfP+HjdyuMhU0NJACYL/cpCFfls+QEbnb0Fsc3jV6SwZeDCBV0G7M
dpSAO9jXj/NvTMlcyOaUSwJLXVAQ7aOzbhefaAlPTNcPpqzOtaaPvSBho5Q5m+X9
Lb0q76WezK8fVHQhyVZ/9VjKhv3d1gKN7i+4iuDve2XMv/3uZYnaQ+Q5waCalmXf
b4RGuvLjtOD9JWV8gkhJUcogFsiAUp1AqXXvvaOLSfMzl38CDZPNKDPKtalWxL/X
iWwSBxkeTsemwhptNx24Mc9Q8dUso/YE9T9YiAItL8uNWmjEDzpofLW2RpFLXwMu
R8AOHLh6zJnnK5jObhj1/FOjJQBkwxxFzRFCmMlVSdX5/N3zbgd/WSHAJZ75bW3o
QlSh7e/v9ovo188jdywPkNgXIp8H0kCFoy7kW1j6zjz4ax4nocaIsqPQzuucN9RP
fBabxWdBeXfzQ+cN9yTp5H4a55tIr36AdYz6MvrWYFoh8hwhm0c/gbABsNEwRoJf
EPVc3X209UV1SlKaX6TPGj+fYI2zxjmUyHR/EqJXXI6gL8pqL8h4lc1+RR3A4Lvj
P25B0RL+GmzxHGLVHO8gnViJzf4DoO3XP9N/lWm2C/3BVwVfBaxsF6+9mvPc0gqh
JLMPuytzr6T/lpHIvngcqqY43yuyVM2gDgqxd68Dndtf7ETqxsa1Vt2hyvO56z2Q
ZVUE1euKaHhtzArm67g+tOE5+HaVXejlqlEh7ga7uXBcGBrRuHTRRgG9NDtVciT2
HO8EFbsU7h+EAjLumFQR4snkcG9JCqmqnVwFCzaNeK/ekGLqpSY+8+7MYd+Z5PGL
zlr9VqwnAKnIq01IxJpYemeHD6i9a6IJgX5z4SxOKQAGjd+WTAHJCGKc3Ud+G8NJ
OIeYwyX4HUtRb+JSDvNE3DVuesNVl6Y2qn8teDGh1FUQ9/jLDYicZGRPHgLMLgIH
+5Qc+IIVrPNv5GdkDr2AxAHOl1N+4Uxq38M2EadCQWsO5U7cbN+jWP9cTT8xx6zj
h8y/Y7/blBRUGEORLgpMpGZcTz7L+x/1zrKXK13STLVfeGADdzrmsz0OPzQoHkLS
2BI/tAJiivgCVVOp4lY8Ql2LDia95Fl9wfPvxa/+84PmEes0ZMenjAMYpWmVqCUy
evp8DDexqiFEStUEQeKFD6YfgZnzwbJlnLcA2w0Olo3nC+m8J5ZoVN08C2/t5V4K
LUV1BOPxXdlgTp0rSvcLTN76SzNwSkxI+euap0/+N2iqpCSRR57BvHk6x9wG2KzI
uZEnuDq1ue6c53TI4Yi5FAS9haShCY9oT8LXRrbmFT2QKdR1Eayc5mm8erzj7yQZ
lmhSKjS86nK80Id4pbaH1BdhPmXyChKL8D3Iwymlo7pCKzloympPCwUEBvJ65duS
Gwb9zuEHH6ZfuMsKjfkvvSafj+HO5TBxMu44zLrPpySIpB6ZaPb6HTnZHPHn/rvB
vdX62vSfEMTLmHp8EPORyS+a2lVKBMM3Ek0F/79UFbpyaAIU1bn7wkpYRDLZYuoi
oOehaXMViq499/SgyrsEZBOibw0zywjMx5mjPIgTi9wDEtlhLmzR3sSedn8m38Z6
si1zMIJwtz6RNm24mQPpOS159HGF3hzUKjIXz2dfy7/Yw2nE4iSB17zOWG70x+Qf
GU4gENqvaZDHoDPfLK8WpuAiJimIaqu/6ixJknldaxc4QUPsCYW4hYxYDeuQQSu/
GgcGDqzBOEJASI3Sf4KRZzeYtUxmBDBTZq5knSbHwrGIM2/W517B1d6yJDk3zjzG
Eu269ZOCRhn1QE6SpMhY2rhbjvSKYs6koC3Bk6cFW9azLa45SQvTnGX3sFwxW0Ee
v5SlsBRKXmcvLfULa8KazpOzA8P+Z/mhKj1vWOQe85fOQV1w6dGbbC8D/e/3Mglk
MuEVIHvlGzhbR7njh7s+zvrJCK0xBEp3fIGpTFzQHoFn9+EF0t8u6yxw+WZYopur
Ilg0Ht2psKBYHudL81OASjxHqwRZ2k9r8kUIXFgn+pV/Gm4/VmIDTbtngTI3ADFY
E80iJNFk/38nGT/vJqC2Ua+h7ia+VpCmjQegqF2cWgZ+tSg5uM+4AotuDgy8HX8i
WQWm2OR0L0n3g/c3JZ35nKzd4LQGAmdDhy3u1FXCSkCmY4BdcvnKUosfcn9N3IQ9
ldJu2ugd3XQa7lsIG0rNijeb3h14EHTruOQPwNtogiPQn9jJfEWmm16CWChRGQey
2875Zgl9V8XRyMmCt4yio/wE1I1acdxooDvL/T/ICQVSZHcvIF7pqXl0Q/SWgx3H
dgQdaob0OQuL5yKKyMcZkqZ4cHBDsVSBbJqvG0XF/7pQau5eXjIaEqKUp4qml/un
2tpWgh/wvqTnucItiwrA6jVypbXfPB+jlVLaXDlGlmf64h5yg48yXu0okLqpqGGR
w9lxTNBUtTBQiTD8/TDODqt/+ZZj0wUD5gtoqkCVNgXSGdKX0MVp5YwXDU0nt/V5
4IqqRUmDNqyadHaO1wTusAN8bs8H2T6VWTjkrMt5GeIcP5hPeMcSGaU3E0TSyF3F
U/8bwZIRvrUatmQQq6cHhCRrIxMvyCqMY7V8SvaDh7qhDeCGQt/46xLed3TWaBf8
2NxBJ5Ln+2a/b1wXzH3YXWLtSOVHQG2sxD7sYUOpdeZpxaa//Ukl5qX25Lv7sHWR
wZsZnuYIoAgkSEYK4D4v8l+mKP7UomjCRZKMLD7SlPDZgKfpe5gFLqLnpYfVLDb5
uqGwucWj4W92qdY8hJCOd5awwlvtLaakY0vRFwacnLbvLIL7x/KWVmsiHaS9Hr6Q
0g1ocUyyCTA7sVYihqgm7Qh5hNfgmRKmLFPPzZ/0iz4T04UL/3pii7lL/jBw4l2K
csiTpgh08wWa2JLRJX+kYOgW4iAJno1JXo4ueBw4lA43n2AxaGXR5cJHW0f9ak7X
YD2L22Zyly8fcmdRA3kBYQ+U/4zu7KxZoVLCZU10bBKZPLO0BAshyrudE6tIq733
xkRfAobajSB+31khc4+zqN+E7bigMgbHUZU24bu41d8vtEYd682Cxo0FoAGpsykO
df3TLyN4z5eBCon0p++dJmfxuYI9cP+TLkVphUsvI1qWiql4WHET9GWhVQPENdac
YrTOR9d3Oawbb9kj0BaCi7w4DpuzTWF3ujLNa5+PhNH/rgmmsdMP+D8nTCdr9+tL
wBS4m7BpgzkkvxBViwTkXRAkR+Xckgd5wEcxcGnn5CjrDHaiUz/DwdhYi3Jwwq7w
tImO99jXA5AuBFgTZWWnzGzCdG/zsOD0TzelEnKyTN4OkNaZv9kjJv7/vZCfNhk0
VG6xCJvNQ6d+eb7oj9BZf0J1xyDGiIR+nrR4ejkmPcpMpH4PzGx8L6OcUxBUtqZO
VZKaDcV09LqL/zVfaXZAd1Vq1RW44WYSHz1/zihFc3NVgNmkqJYDkY5yHX9JuJAL
b9RB52vzPMSyEGv3l1dmC9yeADA4YZgH9CYRDcWBjXYpr85bAhbhFgUvYCtT+ghn
Q/jV9LJ/fVNbzAbViMybyyyUN4ehzQrKyQDfSTmMfRAfzN95hMSiy4HrUVTNLIcg
ycfj4om+A/wzGsX7LuQSWzBCCikmvw6grmH9xM3fsTkmdAPd5nOPpjIcF2Wr0iHQ
hXfHnF/bFOVWepHjaIDc/JId8Ygg2o2gQCnzfmeZL4Nkpg8jOibptr6E8SPvAwAC
Gpo8wCQHaEj/nBf7SSCp4k6t1ItXkMDT5Ndh5JL7kKHa4RqaOswOjZ/1IumkQp7Z
oMrXHIMEWxlRNYql4vu+i5rZZVvJE8jIi8WJx6VXdZI+D9paVTcROGAiabFGUS0N
uIm15dIjXsEEaLJJTa6Ik0CE7h3AasRhsUaYZaEz9hYmTmoHdDdATr5zJISkn708
MfyDHcwRxCfgvxZKzeH2tO3bC51ue+vaplcbbMgtrJuPvt6xvoJMH0GZ7e+IChAx
TP8I4XFd4asAd0PoUN2/UmblK0HR3iUjSxVNPyT+vKc+4JoMhH5MWhfdI88DzNG5
N7MbRPKIn3aUMT4ALF1CufaojI81W/mzEZ49luC8MVV1wJ5zupcYlZ94aVrdLd0e
tgxD/u542V1ljH9Oyz7eOWvmKY5Wd/Knt2KUF0tIBbfrP0bAFhwKZtOKgoIYMC0U
z40ZhcFAAcajqUQAmV0iiIzJPeI2kLzcwdvHG2dONPjfPHO84QFp0TPLN9GAubms
nf4y+o+iSW3+mbQ5Rc7t43o6V4hL2rdBFlVZIGZVX0ATBDP61X4hR59E7BI5D0of
P9iiC58gfzFN7v6G+II0U8kB63R2SXyTob2g8A52MZrJzlOt5UPN3ypWidTvukWD
kFN0JbPmsZaTfzM6Y5XD0x7es0TdpK+Ya0zjk+F6UJyH6vyPuOpA6ai1jJJgbU5l
ogqIEH5LhrwyCIggErQM9JIWsNQzIjXjjrXSnvp++9kL44XSARsSssqYaSWr27fX
3TqgpYQbNmoOT4NQpYrpOEoFr2jDiSY5LTqgT9p9dHdlciT7x5t0ugR8qsthKN8C
daqFti/4EFxO9OeFobnLx7BF/lUEvsJAto26JjBdBjTSM+zVYLOBY9JcIUSbwCZ3
WXRPKnWIoEarmGIcnmPlilZrhYugxrTPKjFJU1cn2YL83je64RXXMxZQTEWAa22y
iBItgT3EmnIbeO2tdo4D2/WyUyp3OVNvdpU5546G3HLFifQY0zwHL8TGy0N+W4++
s/ndBGgZQujZEpJb3Hi6kqcdxnmXikT3P+fXfHL0/kbUxPR4wLu1uZgLDJkbGaDv
ZMf7iOoBkcE5iC6oCmwPOZLO05KYDG6pHf72+mqcKuhYf328cpCMTIguZIw389kI
/Q0efUTSPO85ap5VRXtaCPzHytB6buOtvDFAruhfh1rSlDs/M+M4R4EazYhXZP8E
NSz2tnE89FZTFOL9JJyxDClUUnUUMqmjCLaz6nT+6p+oYJiPFY2edOKvO46bReG3
7hyLcPjP5WjF9GDHH0PZUIB9Z9V01a4WIVkjkOjm+ykXj1BsYmwt+WDM6T39uYy1
Me75exeOLm6Ws6nkLphqHPF8CfQjAleALhxPmdxLYO5axy9qHIbLZENsYSvNTaNc
ep3z+A3FqvVy2oV6pfbJDS6ItiaFUoDOZcKmWUqDCvYv1xePRowyZ8tJcOO9pa/9
+FUg9CZgh1QCeTXRVQFJ8z5zGXcZE0rp3ueUCCgTAeKLrnFC59xyikfs4114NUKi
q1XgVogcuBxtKmkeQeuYlTL75lMpwrY51DL+G+bI2CmrjdrlDxsMkNCep0aHIP0I
+FfY2ruZIPdZemd8okNNjIL9eI2KN/wVdvKDrkFtVyxQs24gsrGb94m/K6nGBhHb
uEYHzdxStwk3ejVjnTNiYEUgB2T/ZbYnBHlsJc51tYbwj3ATaED8c9K307a9nXzR
fsPC0Y5L3g3Tbj8J8AZMvQWCxNhZgRFwoIdhGaFl1V5As1TxDuTpUqSFjvTmmYyB
H7MmgGEs9zINrNKGROVZIv6XbzH/vxeFnoUHmiLjvnF8m/6QvRbSElOecskqlZdS
AGchdxE33kC0MSBW4LLzbR8H2EWKoBlKCuwssMuZi3YsSMzxa9Egvi5KsczppxAN
NHEivo3sphAkivPh2fPcAsm7r5yWBdaIvrjPQ3tXsb9TkuokjWnWoWIib+XpaLxO
wGAj4ZNNP7aM/Hp4LuS4CDFD1Y6QbVbF0OLsae6V7kqF5c8UsSCT375OSaNzTQIf
YomHAxRtBsG8qrkdOyfLk5W8sAua2s/K97Bm6fOo93IQVY4SBWhtqFUuajlQS9xY
MK2vFDVR4Rfysp8TtGxO90WVJO+C/vSnVNqC6NFRciR3C3nVyBPOWZyUZHPqUszz
5NGtuR1QE+VO2Weo9K/oCAWHn1lP55l5xjWhvSo517SK47CnOKz6pT+c87whekfb
wtEZVp8IJMqVZwCBejI9uMIktvdQKyEnXDjhv7dVR05qr9ZNArBXhxyPw+A76l70
lTT5YkSwrugNdxG873cvsAnB2aD5RbcpbvX5rZ18/ARPntX67DQcHPHlL2HWMbyY
+OzVrq8KRlIWKBvXmt5LhLfd/GJb9b7AdXtxXTpuvbZU2VRSOQx+J0ej3VrjIdru
n7hzvB0o11RDsLv8OTI9gmn+vs+UeUKydp7yJLXWjWQG+PsPQ1iekWGf5x8S7gk4
gH5+QP2Jb/V0KvQ5Y2mx45LR0Is0IGusFyk8ErD5Y6XeGGMV7ONcMu62vmKZnflD
Jz5Rc0YlklKq2FiNnvO55QWWTzLmC6iGCLR9MDU5Z7AqEfHcWsbYSSX89vPH9lzZ
2avDRH8eZgCq6sIETCtcfm1L5tAamVakyxJ8mhgIbwuypI7+mPqhqGq75r7G/0YW
FJJRaDHktgGtvTVtHqV4QlnaZ+/c6MG96zYYcBo2RrIZwcZDjG88NGiSgAojP0Ow
q2/J5y/L+hCLk8Rcg2i6MY9iXHBW+/1YTzJLy5XG0xBxlBElXpXk2CxJJDvm0dwh
9AZRttpbEY+j0gRz2KRUuUW4sg7LyS248Obc+z1mjzHXzhHNUiXnR9QmCcYBROkR
hkb0Kf3UWJcUDsUqLu75+EiJRoAlRWIhduPpVXaC7Z2NqD2yl1v1rZ/BH4L8ve1L
ZpG2ZYWpO41qeMNHxHgFvpU1O8hNI6w7wRQe6RT0rFARG9yZCwftgWQrIEVe0VTb
hvJfZnXRNm/FWde576USG3eAjDLC2/Q8hpfT6mryM/DQVie2AtyZJZhgeaoJam8g
QxQ+1EgxBz4Hoq3Gyje6sEHNsFH3VvCQpPQMJfyt8Y8H+TPDRcveKQvCQpJ/QLO1
Qxt9587eGbdQ3Mtm5yrcR22IpqtYRkgmHV6MubzrgnnuAbCxFEay6cY31kTqwKrv
XId7vqNlOWRUaz4oXRaHd9dDKlCNNjvM97PX2Ft/ieojLQ23SbbovhjbCetYIxtO
S2m44m7J/UUwZrVabAzwVEzh8b2ni9Ogz7cATsa2dSkH1Kuaj1k2weF2WThuqQBK
X54wuPEjePkc7ovuPjYBOrgMN6tVCDau/j/q6IKXXbxgVhQFnJMmb6IP74F74NUe
fGKkvr6cO+xq3XmdAKDu5+qp4M6owoMU61M1SL4jG1bNtj1GA05TzTMrNVvdSsyi
3HOVQVXd1ASWgoNNzTClkjyIkN/wbq25Yi+BYw99DlCw0135/FfYqaIg+q21oDTB
BSq78Vp7FDCbalzqgRZ2epKfnJwLHAYvG90nK5TtXQyKXzJl1Z4s2XcMuAAsuX7d
QyXQMTkcrVRbvoU4ayyfFwUFnWZjHLc+OMfYiuVqlVUByWQXcRqKojqZYUS3RMgN
bWnBbUXqtD5f/lAO3ZqXQUUNORxfVzJ5yhblPUfXT7e4fMJnvIiL7/X4NI+WXMAI
rLZL/3I5GuUutrPt89QLJIWk2GR/5SyvrLXp0gfkUhpLrdIWBsObyTI1ixCuDdjS
XK0e/8r4YKIWFzovA6QpqsXOOXZapHJq8dFqQJljWHEjFkxKTokTVinq0hsN/o9k
Kq6VmNRWssA4TkrzkUI6F5FeFoiJfwKFScs9VFTKZ16LZZ8HWNVbTeRCAdFUQSus
1ad31rR7z3ZlySPHT+UYZMxILH7wNbB5udcR73dfF9DYOMShfhjrsi/9a1VBB0fF
aep5qg6XpNW2h4yc640/lj+Btv09yB/x4pP3Ro7A7JdzsliO37DsmdYlp9n0bhJs
g+wKV7N6Ol+1D1sS+57Qfc2aMTJ0Ci8gODZfG2yUnK4QxQ9xqY3AFDuuCnaRCYAT
3WhA5bOIHuOYZwhaVEUGSzVIcr2lHd/GVUUJb7lgYYs8SNw0uZAI27/VLHDd7W+i
7+v3IbhqkNsQZ1n8Si3G53vxfoUgqc7wqRQTePyc/TnA7tPqicYlk71uFACS9C4C
TUeqWM9TCZNzQcOrl3VSGYbwNAVQZ8/q2gCMEdQsGdnGvnkGfGq4fLBiOIhae0GN
euxAidn9trjgQKMIY8yZ6OIZ58PUmbCkWM70AimeNhjpQS7nP5RZ45/ehuw6uH/T
XPlmTmw/5TCuq3kqyYtW3K/dQoj63NI/35Ni2g4fP3A7VOXf078ZZ0t8dRWPyuFY
ax7kLnjdXMp9YA5yjRFj+PPr0D1BqQq6FkXJ53HGiYiApYsZWfw5+gld6gH27xMN
SM4DFuAbH1x7f7xpIpWvSCTrFkfTIDuKieBhhhzes1iPprLiCo60g7Yy5TR1HJL4
3/WUy4rDmi2ZQ95ggZY6zmwOswtwTh2/URqJApgd4MrhdUfnnjjY0TLgsq8roKCN
DsatwGdjXYLRrnhNgv9KIMSHTlBKvaoTfFHmN849MzxKGFtqkJMOEUqBXSDTmmRb
8/74kEd5kbm8c3MrzPwqUo2xZcwuhYnB8OJI/muRkVjU4qElGpl+G1wOUs5uzYKQ
Yr7H0NfqLE64qhxest+Xf8Z5CKRMCPU3wyZEg/Jowq4e0d0aSpjFS1YxqL6GqkAS
W5AB23f5TpKvLF5ETRQ/vLW0sV/OXCJQzbDH6+hP4PnNUON7D771lsVuUuho4aGm
ID/CRUowWDncMyL41FP3WsXOjgYuvDAg8SNk9W1fvl0Hfu3iXs/5jjlPl19joL8z
2BQBHq7RqOsli74wqV4R9iI7/ZZ83Tg7Kwns4TmmcafzcDWi/6OnhrB21KO5CSEt
YmiAxWgr+++BXpIPuvOQKI5QwdDZFMY0GxJSatFQIDDpuxxzKvLoZXaM93vhT1nn
OCcJoVQ5SC4hGUwCwWWQ7nQXfy2nBPcRNFKt0ay6D7AA16f02nYnLL5kvXSHAxR4
857TZk2H0tg7Z2735VexjEJNZvawpemQUknKE+0upUwoSWBKZodQE8Htcsx1afUK
X8zOleD6tIm406AIdXBT+ITmcbFjV8SO/xfU2xEWvBbBAmxRnpf6MgOC4izkYt3R
F1OTx0pur+QEud8Mfz0kLY7eI51CCkyTFbG0diF8aETlaYQPLGFUKN/O65+kg5mq
d65DSxOU7P29f+BlZt2yEFNnmzwVTeeT6/Uo+qDijTv7LH8GMHu2m4r/zdZ7e5zQ
37BB2yaAd8mpM33tZxqPi7Sf4lggrsHFHVDT9zVTKZAstUJZWRUd939EeNSVo2Y+
aEF8nfJuSe37OJ5MaS9lk4l7aDTJn8M2i4dW1gzfZWWkCNWX0UnWzJ1eTr++uZKB
8UcvANJCfSnfuobYFq6dWu/kXFSuCvFofNlGWsbQ8y5jrxSviSIJkQyR2DSZnoED
V/AJ3qEKd3GkWY8mH7knEwSfyrMyEo9aCFM1iv4LuU2gLHhi887DVDoeMsDE896g
K//jG2dpOEa6uGo+xwUL5hxkrECawBDumEV+YQPmzWvXzQqFVd40NZV48HTWMnwC
ddYR/nvrV7pEbn9oFfnm26JKNdCneJzcjzNvN4euuB77+osjo/AQ7fVwz83Xu9yk
mOxkDJR3YfPnsF+kNb2DPUio1d4vlfIfTxZNpQ+Y6o+NbYd1xUafm95C+x9Q5xXJ
pK3ZD82S7GOpQucVl9nkX6a6AdMWbjQagS5YkScfD0IbU29Kyn4jEu8REbOWe6yN
8PkUnqql/c0tYWedf7rNt34itBELV6UWlzGuEErZnNFKCv+5njWjSTuzVQvXDhXr
lxyjSY2lg7KgX3gjhYLdBrLqF1aYmCwp2VgfNc2Kmb9WEcFXa3xSY8kubisOetPx
wl5Q8OubtLRzOTaen+PRGDHYvRNOT9ruMD10qPR42p8JjPMlbEAUFSe5RtoCB3qk
bXq9qFzB5C8AG0yTRwClSkhmmVtpwAZzhLmM9jSaFddX5pqQ59cOtqVEmDI6K7+u
SQU5VzkllXPN9xmS5kLLGX3+QCY79laL7D5aLKaaWNFWiAfErP2ZBiDZSoCdmmlF
r/zKNzNQw50UVw5pmN+9kPVAXCG12QnbaqkKkUhZfZqlVVhZhcNxChh3L5G6ShPY
b/4BsittNWG7FaVlbJclJFEF2gK1vJSzRiMcvB/naxY0ohKvd3EUIU8cZ+aF/kt0
uI5bSo5X6Zs/69Rc4Byr3QSasfgFZnvJoy8MvfAIQIRLi0wN9QJqaDFM0Lx3zhR9
UH/Bo7P6fcgAlu5zV1NKQsayPmQF3H1bpsrWtX4cabpzCXqHnP+e6eXrNlw2bBV2
e1W/ltkhYFAu0cPe4+ezFWR5eDRzBWrTfnuB6omA/lOMMCzB75AA4+yOh6iwPl+n
R3tFbNKconuUciUJ9iLqSd5z9Bz1sRfaFDG8U2Hiqxu89JoUY8HE+UJUXia2F80a
LPGaAecoHEPPlh+6Mfyo3G18riJFySrTpo9QrtIr9Zh0ECcKuO+1S6zlMr7hgnlb
Tu2RTBqMlHCnPDajDZPvsbIRpDLpFFRA228Mj8yNfmoedBLfYxFLwmH+zefsGi15
fOFbut62J7sBRHPWgs5HbDPLrOgnDWSd3VG8E+3yzcoEuIYUqaPkuPtwfhqrTNCw
vDz42aW+mid4YSO/zkB7Hz7h0tGeCxfIeXHFZOVWAkhEaw8cy3IGP2MHe4n2gA0j
ARRlJ04/eKsaQUOaIpzaFfQRJLxkdhQb3CGWU3JHZjuZRn6WypsoSnDjc4LuRdHN
cYaVf3X4L7hz0BNzSFHRM5BDG2K51At50yFYN9PYtxcWxT+rWwn9iG1M2LlFpRvu
IjgMgEXu4x/kTCsDKkEF4rlrmEDkBMU7wdqAvBkQN5Z4QVYqaymBYKt/t82YDOsj
Bics59CyJMqY3GGyq5JOrQeSwI29P2gfdpnl0MZcJtPv7RlveP9c7rZj8TjxdYkG
L4ODKEAQ57oGjFcpnJGckgG12RIs8mvWB98UJB2ps92NkJ8nNUGJ+p+oaZN23SaN
7qFaXlkHZwVi1SFy2SiqFAab6NAwGXC1SmycmwYi62yzch+DZuSO6ghaimOU9DWe
V3V0XvQw4DJowI39/4RGNuLamNTzxvUnSoKymS5EFevhfWtvJpqxeEbQRIK9p9uK
Lb+BXpG9Uf3K/fvdip1nUyWaQHrF646yG2G0MO1UoQU9+bj4WX3FBTiigZB6i11M
vTZnaweiTzTAme6CNbey/qGhJC6MocW1arSzmB86RdulSM3fHGr0nqcv41ox72bO
0ewAArj7kepqQGzgrrpm94m5X1MZivz/ULNj3a/8WTj5DUaKZJDRQLs+DEW/wJtg
Lie+YvxFOpTRqCZAOl7Ae9YPJMWy6CjkMl/85XKTypdpyTMZRiVBCRPz0dSrAIVS
YejzfINWrQDKNr7G3yRRHVdADnaD7bdeX4UT/2K479DCbAThOyYfKVXVx+wEchop
i+TtAodLP6Zii2u7bNK3fFP6mbwbNoqdKWPrWhLru/nRAjjHY3EqOWKluo6G9X7H
ssh5nOb2bNexQtyGuaQBul7mUyVx/DcfYJDPsK6XOxfWxey/KI4Q7H1wYObkd16K
BJ8kny4Ij6yARuZ0ZUI6PiENbvParte76NcH0W5iIhQwAXSmtt1o45GG/WmQQzc/
dM6HilkBKY16+eIC6IKAbiIqWUp3CwzeofeLJXb4n82SdwRpB71zLRsbW0ns7PmX
XhzG6u6Z9/QPo8U7DFMI7ANHjPtIS6N7V6i6Kqb/Bv+i2cWp+tGiZeB73jx1nih7
LbcDXcE2cOheWgmD5HZ4HsXP1ELMLT4n99hwabjj88Ou9NCrGw+dabNulzQ9tMTR
0IyL+jyuyxY5OIq6kSuMXABjEQDyN/FJrqZ9U3VT9UsUyf+1JB2LkYsv30XZJ0YP
6J2NC/ybTEh2+EswuHGiV8XXyYkdOVtABqJ0bWaMzhh+5dVRcoMC/CvFai9JAjfP
SF6kTJS3L5rtZ5j0DfdOIJSn3sXe8aNtXgZClBEjCYS2Yqc6ys48DO6Xayn8vlMQ
L43/Xecy0AVWTepSKAUrZVSCoRP5XFtH4WseKIiykIYxA44VAppwMqXqMRBxCChK
eEfvUQJ3MQXR9ZUQW2IQOcsaku8GYPY4pZ+Mgt4mOBl+rrR6ME5KNh3xiNerUBFh
kNjel15QD10Vs2Tzk4VQpbXuHOs2tpb32LsUnHSPtVJcbZ9/Ut8Xzf9SKzn8TENi
3X6NfU9ndzmAIGBydhihJLEiy3kcOJW55OqzYhOnZGBVNAfs5LV3K7FnGjTjL+rw
Sgvj9W/yLqaQIFy5G8hNi/OQjSH7LDxNtUOpgjjMT3je/qOYlCzfP4KVNnN94559
2aNj6/QeiFmauURU7Y3arU72XvbSquzQXHCxgTWC3gmAhwpX3tjs7+QCd4zMm6IZ
8y+DshtlUAEhx+8Ewe9vRyyZRsre8fKAI7WNzdo8T7aBCavUGzOsH2cPX+jO7TyK
k7lENfzzRbWAnLJnAj0YND6r526j/JSVQUziGOH1nWE/6iDLZfBJmt72OoC2jY6l
QxtYRZGtyoriX97AJFuOnEdBpNsJSBj5bqV07rd6ELod4cy+2EDRswomB+ruvpw7
Tm5d8z2uaSssKBGFaV+Eqw4+Vdic2xr6EyUCdvgqXEGZkD8kyQ94yucsZ7Jqq1XQ
OemAoGJgDJrSQjOHmy6HnWcm9x54fNNcGYBWlI4Q79Nvxyk5vIP87EZ2Ar9RtetU
uti6VOyXoYRFANsEvx0hfEu2Wd/5BcBLuH4QdraRyMgGb7guj3kCm1DDQibLFK5Q
bMkGt7YurxHJW01DB3hFWyDbzyRPLv14C6K8efSQyS4ZOhIaKvA7fKbUs+8EPE5s
aTWJNEEA7PsxHdA+y3KJp713wiv/TAVRG5YL+UfbV1t4k2QAAGQjf2j1gQTOb7kb
w+zJrey5a68aj51C2X2XcdHxBD3qONNoyFeluVTBg8BGyouwpFPgDTsqIUJqXFz4
RGHTX4oCRs4OYQvmZ/pyq/PSE/nqb+taesVN5qgwmTAf0ag9R0MHLU/KsgMqHm2K
seXReKoeJ/sH/oEdwcgvIM7NyqXuvLDWmjkaSSFJz8dkA0OheWcrpzHksv5qzhwV
DnNyooFINuzMn2c0swjMUM08nzZ7VCp8xPeN7orVfExRECE0Q/7rnb/5wUrRMSVt
SRxo+OvkDq36ijz5A7JwSz35Jq65+CdOlQ5GDQSan1kZJJ5ZWs3+iPj+QOYoa5uk
tjhf+9grK/DnLNmOzP2feRM12kAAELejLfRyFEasRuWUiPCSQTlFbb1HmtVPVKO/
ESuOJ/SKVBAMrmnNNIBRvtk9WJ23ViLYXol8f8lOIcMdn5vpf8DnM0yFSp3F4ttb
tQenO5I3Pbw89qq1tsqvxZ2fdo3aThGyTXPvut2k0mhXcDFhKxlGjp4knOuzDci7
hwZ3rWMzXiPMaMVPSUsg5NQHgFzrsB3NNQA+zkqx8i0CLDLbp//cw242VzVqb7aA
poKmqQSyV/i8VtNxR8ZROVNHzUFJkxY6ruffj7J82RZXddbzuhQfx/YsBbXijkxV
ArtVaDOpz142zTA3rQm6VEl4sKiYT3Sf+5GAvV4YBEpF3jXAjwtiduguf7ZWcrzJ
M3eJg406X7B1j0HHLNxcKyNZvh3hzIHcuWOBqoewokIHYIk+JfrOvOiEyATEjkH0
wcxAxPWBb4P3x1K1YOpdpsEWi1qG9d3tPOsUbz9Cq8Elh+C4oJK9RpOUmobuLirj
bteSAzhBBlNelyV+vlOLuxGhVxktMITjkqwvtauILgp0VsiNRid/OYht5jyUzKdI
+juWf4Z6UoEwXlg3W56s35ogL3/4LEOAUcJIz6eeBSCGL0EvHKJlGq/Uh3xAN1OZ
/6B1HhkvUClZ0lcTPZ++5vP5rmlM7a17trNfbCEKVpJPVPh7aJDABr2rr4aWtdXs
rkzb5ePrKxqpajTLi1d2+l7nbTEOHSmPNLwTINAvIztXHPUylrXdBRsXSxh8wk4/
eIFntnjeMvVnYL9nbWUo3YqnbHkMvxq6qy7msryg94dR0kit9HTb847/5ce+C75H
xRXrSzAr8QNNk6fX0mo72dhz0s7dJgEm93G3Vh8LcR9Lk5LOHwibQnoNGjFrnPN5
1EpeYdlMWeFav8MZl6KOuiVeMpbkYPMGnQZZifziJVJkLWP9hcKDjvVK+Lb8uPeW
xCov3W9182aanTinIgnk6o5XB9VoCb7tekKQ2Iat/ZWCGNEWn0xNjDc+DXeOvLRV
z4jijiLRsix21hF+pHR9dGKBBSSvIcOo+6fw7xtsrDSkouX15My+Ts0OEu70g6ZW
Kl5/TmB0lq/RO4vAekOSnIoeQSJGcq3dRwf8T7PCA7V+korMaO1ciaL/5T90mw7O
Skv4mTS8R4eaMqvJtS+xQypcm+tIOJHUWIV0foF6Y6YEOkB6eYMnUpLuhFzXZlSI
yXHM/fi0VJFAaKl69eL14xZaYY80oPNW8ejxwurRtjoQeHtfEfDJNnnYh4OUU1qt
Ty8ykD1RE7S8it1dQAU+OUo08GI2AvgAREei+9gVYu0cB/uWda7XUKLPEiV/rQzq
bWfuYjgznZp5sVbiYsCWgozRL3NIM17Ir2xgD8V/iKAqnq3Nuds9zwUut+zWrzy6
ONFSK+OgvqChCSdAf7jP/K3HOVx/zOb9hP9ki24/Twdj8CIcMmaT2VrLTyLPAoov
HGBs7geaaS4ElMUuNkj+eziUleeoJepTIqeascSlhDMkc8jBA6KCvA+mpp1TBejn
zwxmIWDvhvoqSm+Yn+T+c/EMqmR3GZ3mQUsIl+lO5on541xK/7DUrPcziwdaTeiq
cF/Y7kUSeEOWEU9T9EU1GV9BaTeMawcIqPkwTaNwBZhbY0L2YHqT/mUfttmXqKLt
7WbDyppc0qfTdDaPT5egb3vZCaIB5yanIrBH6OxXfLFnMfcjEYx4khygfaTgCSYQ
tJlgvIg4Xp1rz7eMWklkGa0Uw79aKnpBbW+0sgPurh0cXmXZfdUz4ogOnsnRM5on
dXq2RBmR7Vk232plPcn4sLK81vdjNj5ppqM1ZgkanYBx1pp8eNDXzGwlkRKzpKNn
bm0Isc5KS9sCLYqKXbOkx8oTD0SKxVhwIpRLEUNWPQfW8V4vPNd8ffKXZyAI8Axz
bsCh3yLi4hOybcM+lAaV/V2/IVHDaS/VVkYr+3oc/FaVdcvEN/JAUz6guU+Qd5QH
7vudA4p5Jh0kwqfMK3aOa+ovP7HwMm0f8XBBAYLuzStWJ+1Z/PS6XMz8sBVsKCk8
hLLMlp34Tg3eSFL6VIcDxEeuOqzlAsqYEJdOEyiSjrTfFogSICPDj8WgFjCkaOFa
lfc4V+X4Ttn95PjYm1z8z5+cCzjXCQzDJqYMuElYP3FkLwo4nXdasV7PJM6xJF5T
Um6Hkim7fzLMzLEP1bRJ3+McDat87Z3dMTjfgpxCl3t1iDI/DEnRkTFlVUYYU4SN
soqtYY4I5Pp2ggO90CKRPaLRLgPY2LpcTFUQ+W4+t/Ir8I5ZS17bkjGw2HxT3Xye
muXMmmkbUYZuMwlY0lrKOMInHgP129t+xnzDebqNU3bE01WqxgoenPFj7L2xbEiK
oLbHKbFHJtm1illKrCf3kFLbhEolucmKBH4/lUd/MHOSRi17KSxKNzwXmAJHfY8o
rWf+Im29bKhqpFOQbHzcZZNQMsEeZokrQkvteAUzLofwy1VjpvYBf6ypEsp5EGt/
lymUBBv/MQuweGspp8nO+rZ5e79rK6C1i/vUEBPfQU9sR/iSsI7m2WXm02PRI8wW
hnBJ6rmL2oxh9R3Gn9XDMJEROkOlSYByzw8QvnEeuGRA6cqDBNBBVrZba2PdSsoQ
O3lEwNNa91IOmm0JsxDhgD+M7MhbVYidZcS9oQLZnQyl/2NaPI/rCZzRpoPjsAhi
57gs8bTaYsjF+ujeihFS3Tl+OvULOOuJWeP5RmzFCOQvbEahJmXLHiP2M/6V8Zdq
4zvilGLnyd0DGp4AXQ+UYZ+uUgeCLvcWHDSh+6h+0uigEEpf4E2Vrz2fVxocmdpz
ywdxIlU4GU+wFZ2DQ+pVwL7CvTclSLvwqMKeo97Yda+v0rvwpAPgSQM0TsFoNfkI
D8ZZDaZwwDzyO7dJo2EnDa3dR4G18va+2EsjoluLzXhTaaC4KF96PxS0cYlQ0orb
6y+zxvWMBNlIg5hzSYEJBMRe0T7HWf9dUAaUBWo9SHXmfdczJffZOI9W+3GQMSrI
JvFnOvp0SzZOSKZzyzdMSvjo61OLxwvki6fbctcbOTS4F17zEM3RlNDF3E2TZQ8U
teO1b5wW3oQj6UHI8NyoLsdMbglXOAwmUCAYmUo9LdHZoS4NmnLL22bJ7sHfpgnG
WiYQ0X4DS4G3RzTwQYtcgh/cId1sfigMkm6OVIrr9oxZZ32xwuOkEWb7mqOvzZ5g
Zky5P7MkNb12mxGy+uyPrAZx/nAaZnay9LiniL/VG80vwrAlSgcK3C4HIYmEaGMi
OdgpWxNvd+vycOVmwjQ1kjeQm4LXRSCG0SbD/oASiU+yuJVxxVVfWxBgwmPXcuZ3
oJrLKIEnnhJkmY0Nw+Nm/3lsq2dtyliv/JGp+I5pM4fKHjoIG9of70RPZ1jsIazf
ZMHuZLqFzjqLe/IxgC8GibXRjmYTBp3P5HlIpnA0S0aGig4nRhzorg4U7UHkaUGv
o8Dso5ENvQU7uGbJdQstFCF3v7agb+sDhBAoq7jtBOkRRMSDQYLJeEu63owLO0id
AFvrFIPCTUh/gP0ikj0xwUyWvNHumifZZzouN+pBPmZ+OAa9J8dSV6C9Bgts9yMZ
lPtQbeq4gOgGKigY1EnKGHSEhV1FmKNHoeFZGyinYoQ2x5J9gSBzSmDXdUhboX/X
DkTrRvhS4ozHIzfW691yo/MGkP1hPoZDr1HoUGyCA6dIJ2hRZN6TGP6uCt9HTWiu
SRoOw00/zloJzND7QrQGuy2ajFpwSZmpwSYTF4kcvJRqTHdeC789WDFLia7t6c2Q
3rePIpvJUYdnJTssX7J+JnCSZZLt0LCx9mx1mdAWc1hm2l0U5GRkUgPIAPDCCjln
s9T14eluIBs3o0OK7u80BZXLu9u+odD3Qbwu+p1Mp707IT+NvG5tLjtdSTF6hR3M
09BhZUNKhcfeOuGCJ60TwEdg1QS04ZaWfIaXpblfJ+YuloN6IXcQKuYYyNOsdv7g
HYhXDoZCEp469/l4XtILaqAG4U0k9OGj38GN9v9Xd97pCusIeW1ntBLxgkqsXHQc
jQbGaQETTQpF4t/XvdfV2beLDweo5xfeXYJ7XAeWspoUbZGrzBkl0+hBBYhkzZfL
YnErR7c7fcN8N1xcsr+N3UnG80j9pO+TvvLKvhO/MV7/4MvtgIHPtpMAbILlQ679
V7bL10yC555N4zuTsLbO93pJ4uscKk0Cwgh4GQ3Tku8RwCRB9u1MHKD0CtqiCJJ7
1ggM7LBCe6A75GVb7hC6kgU+lu9XSYrneVkUuvjLJ6HIKBQaNTw+AVqMkeOwz/il
nqL1KWPbNr63Ph6lt1UfmOXYE5M/nrJRm4tzb8725QXkKAbXDV98g+cZuc4iZfW/
Zi+wUc5HdYLS+bwfa8OebSQAPQ+u1fx2/RHtaSayNSBoKdmELveTBZ2CDQ2MUarh
2+FNlWqgiUOvtlx8It92d7waFT6/XZ5tVKmeVrkiuXdEcUjLqyU8P3W3/6KM23j2
j76ZKtg0hs7dLUsUKhUPYf48a9FDX5P+/pCoH1+bm4d2SST4gq0YBqVJ5qL3mzD3
qLrusoSo9qo00ZcwOb2v3VH8Q+UX76zuviNJB8vDCuHHhFOCMznjgwPtZgJvgN+L
lNaefBpotjv61ci9b0oTK5pXlSsCo0vliFylQo2EeZJHmKu12iH92WESZwWonJBN
0Ln9x8XKhUUOM/7Og95FP4ZD0mCJWujDdQ7w8s6+30uxNR+xJ0a/fkiAN9Yg6CjK
AaykND/+ze7v8w3jH8CcB8bqhIi1kqvYlQCvMotd+wuWliziuPc5I6T9XPb/WeUU
zm0FeD1SOYpsiQ/OpZS2q3HsGjBClkasmXBGbiLUsNEUuavx1zLM7JLz2uYXlzkE
Bb73UoSkZMa2TwaAfSHQFUrJeb9xJ2xZ8J0hJ5wCsMaYfwz2O5sLxHnqbXT7H7eN
fwOvhHAbmz7fmjzqEWRTPckFaF5M02H3PXXZV41MTUg8wNoNq2Q0X+61EAzmIDuW
CI/kXWxrksJd83sVFXVYAfzDVL7Jj33x6LvjEyFc8BdQlskMdnvudUrLiz5ZTK+s
nBTkiaVOXbQShGaARZuWZKmLdJJOfcYJIlKLfGxtRIRx5WsWqib4F19FYr5dy614
JBVALlc6qtL516RldGNZG00y8o99bv7u70aiykyJiTyCwPKIuPYNZ+mr49css66n
9znHV2wlGoX+VUhhRdRagla7gkET1wXwblyBlZLGoC0QWjXzqtN0EEPkf6q9DdDb
1AmSNKsXUJFqiYMftX1PbyGwlV4K6TcMzTflgStF8zFhXyCHTEqonAxyhhOI26gH
qa871d1sIMn13Ahra1XjSq9IG0WhgLFDlsjQ2iXbLl0qXM7ZjLvhQqrWFZH9EXPk
zzCkVgamnXCJfePLOe1bjHUXaOjXe71BZg9WbAIGtMEZkpxkQgUTYNA0PvHfdllZ
0sGnfHOcLCuCJR7PVMZ9WEbSBM0Jj+nwO3tR35AqCDtbP+Kfu29nUl3gyjItfFoX
sh9gXElEgcACCjQrdyXBPJihP6LDFNNxsx35PPc9lJDTs84WULQcte2P3qUNlRzE
KDFbWS5RNt5a38pYSDj4qh+zGbFZbJrEkP4MpJfxIkO4we6TtG3Bm/jsMt/v9ZsM
PxyJpfcbti31matXkgSssNJEP/5EEs+UNRlEQ7OCerfv2EYaETraX0ynluD0Rw/p
tZGkFR6vDsSq51ZDx7TWbdJCywvL45Fe5rF6E/9r8BjpyOtNAb5rkS2Sk2N76sbG
HGBqLQjPL8se9KHL7JlN4/uF9/K+XDKQOBNR4Di/E4jqd4OB0GIqGdZW8u3i9GIi
qnJw4g9y9Uy0HGLIGLUOz8EI+kn1AVW/k+sHKoG2rwUOWrxT92sjp7znfjKTuRoz
lMvGtD9tZ8S62TH0fZSzaJ4UcDm9pDaj4yshmpMNrpu9EuEWFRcvIS8gjThjjLs3
/fR0jUZZvBuoaz3R5hxTk7z+VjCG6i5w9KMdh2/8Xm1X2e04ibv9ypmTK+qdiSBA
9zELLVpgxPCS4incUrUy4B42mMjbxhKinft20fZPvLIlFCgvfU8IhOuYyy2QFIlS
Xy2Qhnr2SIX+X0DWkFH9+Mwky6oxc9rcoH3ucQ5P5YptCc4SPfWgG5MMBnEyCg4E
eKHKF2zFAPCordMRChuEtUDvMpf5SZ6QFCfKGNoZyFtN+RmaVycy1dThyWdnlBHP
k5WwNCJtEpviY4RKAY0HrSN00qES5siXfapvsRTX1dYxLh45WMfOWpSpSwyOYeey
/tsymu0hKfK+GKDy7YVTsPqCYBSOqTo9691v/hORuLoS0HyD4jVhL0Zq9qZGAkyO
K+XGvSMKuWpi7iNvJlhRFS6MUMJPjgsPVM/y0dF1cr/W/7h+ULSF4iwBqwyGn9+z
pCTxMpgo0UbN3jtx04c8yXBBRECHn4NFr5XOygY96fx+pMFBGfryT7wvIrIH3sPW
93Z/adcPt2t/GoZTzJjYlrGh9pyPNM064zW3yg0BPRmSoqoX61kWU7b+trlKRGrS
g8WKNfvL4oiF/iwSrXB91J2aAYRdGGI7v2iwhzM2OREW2clePr/o6mTG9St258Lj
e90c18h1vpcuiL9k+w7UHxy6P1Lnn3cu4EMNTQdqsCUy6Wl88j72heBxQSUZealP
LEosnDun+5ZwY29DQyQM2dxxAS7NMud8bPac2O4Bv2aXBXWOhRlO6AN5e9mB5LAQ
0cjkylv/+vFCjZccI/6Z9KXIszjEKUUvSlQGw+z+HdbjG1bpJ5noSiEdobcgVWGm
hG44257rdCmdEee9kRMNb+Lsgf1O8nE1G9SKMLJIeGvh4Icqgq0n4qkkddz7pLuS
WQbxFEEYu7YJYvyjoqiTHqudAAn5+ZQacCjHN9yVh3KOL1ZaBKBry4lH0NfPoWYd
al+TGfw6CuH7wBNapnt/TacB9Yi9TXyY52iaBo82f+Q/cdUcdi28l5ksUurbQkbt
QAG1Ccy9efams5w5EzhmX4zd7F9eq48U9ONWzn+B/+jp6AsvN7rsUKf+ypa1unMk
Q1fzaXtGgOWqAtpUMqVwZQ4UbN+Gm7t6WKmb08vFBkPl5AqIxKagCdhKwUjykRDG
qRC5ypBicSifBvWgX5K7SUWHM1Z+mu/+EQp8pZb6p3UaMyMZ4Up5ByrDATrgLPax
nIoX+tTacShT353NCPYcca+r2yUDRPzim9UdYzDYzHXM/Qf5K+b7wDHYwvrDzgJC
4bDX+0zoJrGQaAJtLFqwSrvCDZYNwe4rapdy0ODeLRM/1jFcwb9ssXcEhsNOYyZg
QOmAW/6C5+LYeD7QtDflQdGjmUKzsifb9RUwE2ZQ4DT9trmABf6Lmv7iD6opCuTA
+Bwae/PDfXLabxxgMl/rP8QVuh4F8EwDrhKhRATNX4PerEl0evoxmZksiYG5+yzb
LocAhIY+kJgxyxYJzuxAbHlYuSee0UrHY9pxaJbzRwByCIhtiA8mwfSL5HYqxz46
6W3UuW7LaP5IPDGZxbYSltv/fAfY/2MDvDoRnNkrXo1FcjOlpXDewEkHnkzOr13A
dbMM3TZnq/67msj8LUSwFhCLCIzMFVoXz7JhykwiOSv1a16pEhG8jcKogIX6/4cP
B2oq0vDxZv1sSIxEn+ryzgSQ6cwU3v+EhizspQSypjDYxIVbJqFxpzhigOYc1qMP
uY+GPsb1qhki8nW3yvKLZ0ldwsMxdDCgVATCVCjENLVxQpWpKzDlzBYi1PBqOUHz
Rkx4ctCtIy+35Xc2q1J/TCp2s3qIKg9UvqPWjFfBCrfFG1e3OE6bvzK6Z5FrJ1BA
Sp5TaUiERuRUZASz1BwlDoPNJCAZqUxwgJLte6so4qzkd+PP7Q6TpBeOB26k5Ohe
uNq7b+CT/jfv6obZ1k+o3YzhK9iKRSBBV+zCWyh1u7Fpda8IZ0bbqqMEzqfn4bI/
HjdHGCLmiZi6tX/+vbchxBIWxc+mwUGR9F4K2ymQcs+fcB5lx+FKU+MVG+wk/i8b
5ElP4/WxxfgyN0Xbf9g9CTy8ZRO7j4mPJxtMERQFZq4LjYx8quy6QlrrHVfFIQ+P
wqGWJ9Ia+ew0l5TSsGXHqtvFv04nvd0fcvfR8tAEmu8zUE84zUIXxsgwPE1UmXIo
kX2HwZzTDIGI4U1gbpb0/6+rVp2sYb17aJ7PI3AgTzfTnnD/tX66coCzEhfwRY4S
JWuU5ZAFbBTVLp2thqTCa9XJ0DsAjL/nlpRJN5GpQJVW5ACYJ3cR+KGpWWdqg1eH
2LTvbfuhdgYoQrt06CrvPXz4/+oOdtc/VWCXa/l08ujPAMYGXr2xNhxPhRdaqmm9
T3ZjIxnBNa+WW+LE0pKsQeeAfcNui5ZppeSyPv+KKs+ZTXaUkXhhtfxSfvf+9Fe7
fCV3yLTcyzPgba127BzFYQJcu/8gWvrNAJ771ytM1yk25WLHIbWHbP6C2eWKcdzd
nHn79n+oMR0Ex6NtAaB6ydSSya0oweMRZIh3K8iMO/maJToL2gmDEG2RfMpg0vuT
UxqmrbCB6QXvdkq8ZMKPbxpLvslIdJItH5Fm2J6fKicynhDojFcCqf/6Qr9fLfp/
QQ7KnMgJ/rj4T7TTydiV0WJ83EbRbeWqlQzhJDJet7PjiWjPSWsZDKVZSyCCkUN3
SuweEx5WqSfYtmwA2rrOzSFNBioPMgRafNeay4PvljYsORLqQgfSqmN3YCCdWg9+
923OTjOVzR+27GyXrVRxwqo8MeeKIQ2rgOn24wVQs3wQeZzveUj4YhLuV8CxF4ln
4CckOK8uk6i9v/CKuNMTShtgui8qqh+2zgyce9oRx06LsMqoFm0YPQQZhAKkMah3
LgjUnja9m0O7h61RGBf1k1/IVjPV09MwtmY2S7YGw9MesKO8ipznrFdkj8Hm1sR9
Nu+8lPxUeTlu+9wUFrDflKv2TVf9BE6p/0qJvyTeFNz0xGV41TMfzSrb6mBYuVvZ
36JQAXKlR/djz96AK50wiTptuJjAchJMbHYAeCTtrZLJPDhNsVFdPtZ3CZRWPWxH
KZotSTTRhz09wGxaVxuud+ehjp/SI8aavwqFv7uqcUd1Yngw2LParVOIClf2F7Nr
j5leGG55yM5kMXXkIptacJJptX4TbLkSgciAj0zFw3Fo0H51gUvionO0hz2nxw89
P1s+urbup+vwKWQyFsSgDNhQrgAaU1QlK3ERNpq/R7lTCZViJfgZTHWbNOhNDNCg
S0cvPMN8GcBr8FDHZ9l0BDpxspThlFPLY2urKWMrOPCMCA8woCKqMYnXyjJI3l6A
PUzIBbGJns/jAotaJMFpPwb5glLP1qqjojaGty7VLM72xKdUAZfYNce45csprprW
wskVQSykiNbynBBLWQht8GYgMePIWw8MqzzwfU8J+fzCymCxMCB5XhFEmzwT0vKx
BgfvmnTknhyHDBPbIxdDD2COxEMYKBDmOXxt5aRpzYuMrdIBL36ZmlOEAOHNe7EO
N6gzPIbeIxA+YxSeEc+W7inqNbUHlcmzFsmwMAmMxLtD8xiVEmNCTsEGQT7i3EGl
k+Ss/bVvoHqw+jovQgswFgKU8oidFKBK409MEhiJ8yiOd3sC560LuoznDO+Aik35
T9ZwwLaGCteLZwb9TVPv3uU9YKPL2bjF8lYsE8ghxzZDJ2Vgho5lctYHTN7vu2gw
m/O0KioGoKqd85wIpsxerJ4Tl29itIr1lAn7EGo6DaOm7SMfQBF2rH3S42C6lpY/
Frw9NnC+MYFytftwuxA13OqYns8p6N/hc+67OiLXHjEKSnylLh7kkb8+qrZuF1nA
MDZKvmBQTlHcSZvmt2Hgx00z8FJmWhuzVsr5AHHr+hyUlRxf8uZB8nOUJY8CIzHc
lrDaxu0CaPqPEHQIE6Xve75p2AxydZGTzr1tij2ELOYGkZp0V9Q4NpDasHcPGza1
GuuZFShmKs2a2BopEUum06/FbgC1sWrWpwgar8q068GrgAwwYT4gkpW37FJk7M0m
m2JUywNNsARJHBPmuwop2DA9FUuOKJvnmHJL+uO0WJlR4gnwTvXTMbNCLaS0D8oj
qkrxOJu7048lTp+rMfNrwP8F2uW0YhhV1QYiwVzYMLfRaH/ehCooWRW6PzjXP+qX
90ebZrr6V97b2zCwxYeyvyj3jQyaAfosdGYYCrGIf1iYBx3d/83V3iU4GzAp2lZ+
kTegYA9JwC4oazfU17Xab55dV5gpiKzJU1bnr6N1YqkWIuAvD94iR0Y866eymjc3
tqQ+cqHEy1hSyyBOlw1Y74+XL4rhkwtAKGabdNFzPO9vpS/tThYgNM1OFFP924LS
fqXp7nMtemyOvQkUsLtHYNrUEjyZft9DvygKQLRHhKX9qk5TwYyQUBE3PU5efd9m
0ZfBIfrS2BnfUEcdIn7uyUjQZciRe0Cdm5vxdGP99yxKvmyJ13+NEYgWsCoW1Vv5
qTecpq+yGKe7AtxCuwVKaMdyMDyQykWIVuylJbhFPIUD9PY1WreOBG/c3sjZPsyz
GBgmZbR9bGufZkTht8MbcX/z657Ua38H+IsMMFBUilA1Q3wsSVa74j23IUns1vKW
Ok9Ix6/4T07FPzjMQitxqOjM6ni8ybquu7qPS8STYycJN7jwirgwKk5gRFGVYW4f
xHfDduogmRRU2NXJMIgBKGNUbdROkvw2SqjdBSb3d57woIBME4vBP1W6hygGgOmH
78MTEIyeO0tuH0AkyuLydDjCmswlrnGHexZyuuNsywje8bqyjwr17T2i57fUYUmt
p3BU1JhPSy1HrSVBOFdesbx4Vg6Ti5Tfz1pea7gz+lmCF2AiKKhAZG1cOWD9TVx8
giK5r5cx0Gz8d1xLRM1b6axNcPoQbNxQelafp0zkUjAq9V1izqbGUBq1xRh1RcIi
JZnJdyu0TR0paZu8cK79u4ums8W2rucZzPgTm7J00PFIhlANGOAzvRGv1vX1txps
AssK3Edw/nYFrO/miOrsg+Qy9hoPsv6ldrl5/TsBJrl4RpElY8D7q4V3AIFR1dXE
iXr0gR99qEu+hWSU7cKaCPkp1k9bu4o1GiGj06bEGJip4NoSaffqWWUK5CY+gDCh
FYkmC4oeGiMvbpFd2Rxqfdx19Q3tHxJsvY5OOwxw0WXbrAHZavHBtS2qLDdbPmYo
lLi+jXxtRva7d2nyBSFfDLT+GQFXmGwRJlb7nO5P+x+hU+GacR1hUeqnyntx8qq8
6guGhBWAV+JZUcI+w5onT9oYVcr7jFZ6WbXZ77/vYgW/Ko+z8vqAv1wRwHJ/cBHR
dc6k8sZBBCglFIABCs24VxGA8zmioXHhnYsMCl9eYBSU65cIy6v7ZhR7YOcbD+LO
ILnBxRggdr6CkPuAVPxUuu1O4vZJzZ3eW32q61HDE9M7x0TKPfk+NBEDCghzJv8t
XcD1dSSwCoi8lGYvAqKzs++5Khor9QjlsoYS2/j+NtOFER5cm2rtRQhawrkAzC4f
weE/G+tUsy2UAeJlfy1bTdc1Cwk4QAenOMSueBPb8oPahJ/5uObNlO+NDXO46xAn
FV2pqwBaCA5/tdibZqGbesHBXJG365n5XmI1K5+9bzD3g8iCOkg/pfiqtz+4RyFK
Lss86fNEtiGehZXjciDX93s1r9yTxt85xb+YImXodtiCND1S9c60BzEuWCEagfil
Sog8DKC1H4K6PLcLWV7MLbiPzDgAx6DMn/GcgkE1pV9wpaG4xPCtRsaaMEc4HSIM
aUxNtWjby7a09V9kMHb+t8x/C79PGpFp8Tpjj7OCJm920faisxVhdarZyJ2rN1uu
H93+VKrUz3tgSGk3eWUs8scoIAO5Bse/zvva9sdyoOa0/uhWh17Um5gbkXLIMx57
SycpYEB2pPpsIoI6buOinzNeg34h/wD2zt4QyG85nKmG0EYze1o3Ypsy0x+MKTg+
8mzHyNITNh+rlx9TfW896nqH7z3yRCDEs35diIbJ4JhrOTyeM64wNayRsqFJsqv2
Z/qsgxqyuiM3raqxtE1ceocdZ5K3NnUbEsiTLM3lzQ9cL6gECYi3NiRzz7K2k96b
+EB95WcLYAWZpDNWtpdgr9ihDX0YVrhsztwfa9QgNgxWUdjRZvx4hsJNJuKVSFgN
G0p8JT/flW0ZiqwfY0auP+WY0Q4B7+74VCHtJFe0vtEtSDXuBrkGy8KFj/6SlSpx
CzmIFYlNf8u1++yIW8cY3AmrU3lh1rbJH19WlLK1OlLMjdwYS34Q27QXSj+tQkQU
Ufp8ZYqdXABR7OZUdI2dU5NepNMd/CrrpGMDGq9f94NbQg4FZ0PLNO9cSxORQVSK
HRWoEGejrhDxX+9HJeg3763UkUIWTkzMESvs9rzqrHWNNsK1tzExBEQfDN65kaS4
qUAlof9r6/dJkeg5+9l9zlGwzICam5K/j5rR5s2wsqKkVeEGURVNjtyFL/H2rPKz
6VYtYCkOylWgzd7BB2oOSkoON5hZAAs1Z5mHvL01WPdsXeo+IlqHC6XgI5R9bgxc
5blGXlQwkXXaqKpauT5K7kcPrwDs81EQOwMa6UYi3du6LeO9pC1BHCrT6Syg9tH2
4hWI0fdFAWtYYev7yMUDh2CoaJXadr5OcR02IL0Nfu5ye6JM5gWJagPy3muOeMoH
3fAdAbi6cE1PerxBqvH8pkc2YuxYuEWo0MWRT5kphThcXQGSpQFoDz/Q+pEoMRWH
LHTb/YBcL1nQ0JaAqJDBodfjFAQ8fSvb0xK0PHGhPchQkySOAKfeo1krKGAb/fqu
JIzH05NyMyWRzFjTMXTE0kuPFeIxz2+KMkMlHWPTnE/RwsV5XnzWZoKagR7/12X5
8sCtu/6mWH+xRjalodN6HTbQjQskFd7AyTzK/obv22PdrYrB6CC2pIERaJIGoWPY
3Pt0K0GvbNFYxV6GkW0aD9FyxaY80NdEYvk6FYpI/a+oB0pwcPrPyjfTyZ0HjvnX
y6RITw1Tnn470xRUBvoH28j+j3OnHIyo60uz4soUv4vV1SJ2//PJA0uVZzEuUKm1
g6NTvg4pC/WudDNZdOlRU2+xS+VqPO1ZzHGRQ2SwDEAyphZ4fBYo3oOYV+lILVi0
oDqKkmauI8qczAhDDUy/W38wss5Qg5kJR640ZQui0EeyjI20n+nnX+BDuEincMEq
o1gwhx9gbQA0tB6p7ovKQU6bp0ahYFKa45IaNNJRVM9QnPL1YzB9hYQofswY2ZQ/
gDxXwPD1DqRp0+T58eDQvC6xlzqa/rzUln1/czMpCpADJYH7mcjwwejZQflXEuqA
s66R3pS2Mwp3+iJeUwCLdWwKJC3jg+FgVlIwonidroCEEejUMYHO/yjTeoibXlzD
H2Z4+cO0XTLZ9lratSnVH+r0Bo8W0MVScWe5pitfWAKRQsedIvxmssg/yn+AckDC
RQtK0BKa4KXcN5u5so5GFB7MFrrzH5f9URAgRoe75OG0cTUjgbZG4PhJS1Cw++vK
0xg6lGtgTmKPNR4m3+ishTcURiek+0SzBZkZLPDvPQmPMnsogmcMwn/wKpT4TmIZ
kFESEWkPgR/shVj/4tgBMsN5ZgJIcZpLSYzJc+B/2+27psaZj9oJDmbZJatl8/ze
QatoWANGBnqft5w7Ds0+0cNaB5zNKtg82zacIeB2RRxzIZgglaGcIXuFsO37R/FI
MOiAFVwUY6ojqy45BUjXMHxaPWci/2YD6EBuhvWtIrutDuLcP8RCBUkxYRt2uTdo
wjkMUhbRWDItbeCjjnmU9nW8tHK1WMoYaW2JD62IWbXjqO3GE07Kb+cJR0Dw+wrC
zfKkrlieTxJMcZK8pdR2ZXmT/SOVRZ8bD4DfodvBuLaUCX7dfX6fuQLB4aFcYpyD
w/cdhaB1vWUAxaCjMKq1o2DW422JyZZKoG80yjoOzti4XXcrsu3pGyhvCIyAQXOf
1s6FLcmfSqcAHIfzeb9AQDUOOL5xfpZuTZuiSo/v3b9HLAihrcub5LpQZ04vGauS
k+Uzr5cquepaCoKen8eJLpY6lqkbJndz3nXDqjgqxDSMgJ7JmknoJZjqzIObXNwc
aR5Rh/EENUUYHjhlFBbaG9/ebFy+uArtNVra8+Jhtfd4PtDmCMx86NUOynTC53Jb
GZtxXT+lcsQxZGzbymTesn5A0wl+stor/MonEoIZhzk0E8ig1ihlmVY3vg8r6HZt
fu41wkOmsklv7yTuSoMHldqFeP+zvQZmc7Ha0zz2NfNet8bVblBKy/rNApaVKdMf
eno27ExYfXcHr5R44fRoUEjnWV+zIhOFDjgl+0IVyi9yQk46sLJyn4zqYjsIQf4a
aD+JbMrEQGFlpERbLaofSAKNmSijunDnNYFPQGMkVPFWB5Q+0BEyJLU0T/wTFEIL
Fqr7vZ+KRKCg4VM61vMO2lYAmw5cJ3GV7lHUUHXEv/EcCPEm/n9sRvw1gJ8sBBrA
iyKwsuWpaRrULYWIBxIWm0+fjfG4OpWn1gzb5mGrzIumy00JhbC5ElyAq+nnuIv/
/ikbz0DRnbk3YFbQshEA0yVpMIQZQ68nQiOCNTuF9MfI3vCiSwX3Nz9gbONqAvjA
IndxiawyAgx+Fm++hjr71JraUHE7oCC0kqlw1+/deOuwnvZVpV0D3LPWr/BHpBg7
2ci0RUsyMH8NSFhF2Jd5/t456u2OuuZ/p0kK4NIcWoVrmbB4SYCPV4GJgPexG9zq
cJaZO9vtbTWa7/9IQVgrTyEjOvbceCoYov3/TmB12fz9wdmjfnh6KjNCW5ahkYTU
IuT4xAlaahCV3o0f6wKd0W3L6VTQgR4TLQn2mDOZhW0hMYNCJfiqH+0AAVGLBn26
m7FZKz64XDLJLH/qa1x0c7DVzPHfRXgpV8dsBNYAPOCOKk8zk61iyyOK1PRcoZaI
B27FpBVN4C23fkXVeKJW7l1ixVZT/RSXqgF9v3cFjU4yVRyAfTnenQRJ+A4dWKiY
uk7xXUrx6E3XW1iOY4sG5N5MD9oQa7gh6zirr8jfV5U7ODWul3WN2KyIGDy3ksvK
9AvwNwEtZyTMtX25ymAmrlRl+WiyJm/oXpoUzQhz4kQduhsjapBCfqp1DG11s+ER
wx3P7QHBD208wkjPMURpHQQtVCBMW/zVAk9IKED6Mh28i8JagLfyK177XogVkTp6
dt7Np4cgWYALm3qgenZExKgfDS/btfafK/012DnPH1h5jafjjOTx0VDdQzYin4X3
fOJ8QYvfQMBqV7/6uLufvAAkaVhb5Bzdjftt8n37iGX4MYajZA978ZmFIx/rRy1k
PcH9Vg393+o/nT1ki+dp17IqxFXyLVWLSup174wlMdufqJw3BsGNvXMFLT6vHwNG
IBC1C/TlOLyZnSpPkJFRPHK40Bbify4tS6fGZn66SIjGVxyrS3bv3xyCvsw483kc
RiMOkZheLny7ekZEwp0CdmAAfC/SfyqMTciRxwR6Y1aGfDV5QUNXW9SOmbdJ+IlW
N9coNs8JsP5DKWdcxLbMyP5MLyOP3j2Yt+HARwj4iWiefpL81S4LJwnxjaF0G8dN
JbkgNP2zXfIdcg/WsOeyXF2Zt0xiqWETxNdnQsJ4tfDDH75MDwYEdC8A8Ms6P7TH
hiQO4QLzl3B3FEud5qcODPjTq5UJz6JEAx51/MJZ6A0qEtg7z9yQMWCfVMWBPcgB
W52BoOYQpwZ4HaUPlM6AsoCgcT3zOohR8iayqSfD+VoUzLn0Krwf0GiC4dTRhLxj
8c0WIXD7HpN0DqW3yOwrr5GMNnWkoVZyrVoSJtF9ukUR5eiF8F4eWwSbnAW5BZxH
6c+zRAoFIuuVnj6cr6tsNCuRkNP2NmazLN7TbmJNe68dgrXitMbJIcrPsr3FL755
Dih3frTfXo+ZdgVDkOdDfAVNvvspD2aY8hfdCdXRnkVYJtDu/jMQ7SEJ8iGHfTv2
nntYLRbzoMPVm5SewUyisvfc9ofiFi0Nj0pDY8QW41sGsuzmut/hYRg+RRh02kHG
RvWF9x5YK1OaaJLwGZROvZ3vuyxUSLX+MShh6GHObSHaIuNrMx+Mjgn+AODU9tNX
Ma4niU2olqyr1Uos7bIhmDKoqlxBZr+eOAuc2BqeEbNqOzvvvmWUeRDprNCu+SrV
ot0+dVv3mff8TK9KFsQfyg7Y2KlcnmiV200G46h8+9f18Ef6/velShP97K3ZX3Lw
82BlpyZErY6cLtg8c+UQq1PF25JpwvDcBpCEbjUMKuWbhoW+19STWVzq/CRRAA7K
HQZGquZAa4mtBwvRxDALoWLW8LsrKGoLovzO5Sd06FF39t8uZPSBiSdpAFvnmhZr
p+M8lLF3/Vdbm7Dffk8MwM1TE+xNPpETxQAqODBWPXsHCkIBoM9G9Af3dwuJ1T4G
YdnYBAVl/hD1QvrNjSo4E6xOahhZQXeShRRN0RVt9Ohf+30KKkHLEbndevEhHmzk
BooIItdgnqEUDktPhUlJ7/tW4ASczPv1Yuvs0wk/BbqrqhWTMmMn6ni/3QtLtZPU
RxHYT4dVwY1zPl5rU84DkDgT5QItZl98Pcfikf63ZX9GKazjzRY1iKRpGyD836DW
ek2e84Vcp/xna4n7h6MlJ45xCi1VcJoyb8dBBxA8zM3VLPPL02CpURoQNcWC4C90
ryNNrMQhzROwB/u1dOW/Nr1wOk8KoX23TDFl2ROZhK/DrtYYU4O7xSr/pa5Jq66E
ZhxFnH3DR1UDgKADQqta1R8Ul4q4PiCcEbTze+4Daf177eNGn47b/ZKjw2g2kJMb
QwBkRQYHsF2NOLpwPkQOZBgWgUPFFuLaeDxERnaHQlW64zThOzYDmOYVMwUarVRe
hzdb+SrnAkW9FkeLDpZVLCPIjA8x2uYZMR5LAIYu6mvjqkiyUg7IwiOLDUMF5Pzp
VMpFWTDFBDmNX7RKJYYpmONS4JqW7AJMkLh7xjD25EowqJh4OOzBbczj7H/mg0jT
RrfQmXrElyuDfmhbFGMx04xuQZqN+RLEMFDiLwfDYrEZYaFfXP1GhoXLyGvBzK/S
RnIC0uXNHv0AvgCl2BgMp2SFgeQ/g0VGctcpHMBFIWPfXdlVWqgBQSFjRJ9jIEHl
HcrW2ADcA7cr8l+OxTeLXn87LZHkzpfdS0AinZNwFgHtCsoGTqWc0Rc99M5itWNK
k6iI0eD8mnd8AA3/v0nQ5n3BbGgD3caIxEiJFX7EqC8s3kSHkYFuQlod7mW/SlpJ
20hADiKdU8ejoIFOtinQZXCEwjRcPxnOvm8HbzYsoUlgr4XXBSnyv5P6cb5UJXwb
BhdKeq2FAfVxhcI/h3T9evGEoFGxrHOpnTEXZ1a9zTTxtmq6lTkwZHzPtUeeow2v
aThMfYtUXhER6ccYxwbuyhv9XS2qaNxYLwN+Z2HReCxWNR1ylRst1qU/pyShLdkc
JsoAxYUWrHlqMGmewMM2eO+PVZ0ZU4VzgxnlIgQ0WNoa1JuV56kO5ojB0qjkWE+S
qeZtIYrG0bR5W2LwJl0oNInqmq0edmkljGhuAhLLjNUMQwMBl/fLLx/Z0dwxXlwc
Q3fI5kdNV3Tu9FK1UpnmI2ufU6yS4zbZRwMRL6CMh9TFqIqKVkfVLWrQ01i9QZTt
8WpPJyOCie1hks8O0E9SHz67hzm3Gc1rUy9zXpB/0IAxegOISRrq1laI82+dVOZU
AOd46xE2iSptRm0Us83ylZnw/7YBZHzt5oQHHyix61VR6kAERNAmoJ+sfnyVqfI4
JALuLWiwruTRrG9OFgM5tWW84VkEnOAl4KzRzYJszPEWtYVnuAgyutXzOAPA+53u
5Q31lSyjOTX01LjSyeqUMcipr0krb2oXg83hOqgUh13vMLf2XshuNxzu93SYb8WK
brvwireYWL73Pcx0w88ojA4ajwTykwpjwWocEGh/YNhI2ypytvNqOqmN1niVpzzi
h60LzaHDwa8hf95lzDs5JH6W1H6xCGSWgDU6R6ry8yQOkfQaFQUt7DwSb7ObhTCV
ht+za29d+wpyU0eJl+lemZmGVZkzlTWjxCOHZ+BD3wseKujgjEjUTEptVAMn0vvR
t57FJkKU50zasjyGiwFePtVsZ4MoBg5jPlDanM99GX4IDAJJai0W7aeUd+Crqn3H
lOX8tu+oa/twQ2tYtArcwW8EJ2NTHMNGGA/m8zam1dyK+oHa79ziMLoVFFkUthe9
/SVeXxG9O4LKP44JaEPd4x7K8oTk4Wf3Y5twF7dyqjVngkYh0i3Yi/EmCIvqB2Dy
3PEfyL7Wx9kCUTwS9ctnB2OArmK/wle9J32Zymk4xm4xwUi1UvKCkhWbL7tpeWPi
FUB8+sDEZe3XTldBykahZxJZfM935ek9wXK5igRiFlrmwO1eXkTBlM3IsojEINLf
72MeNOgduufGXLQQ/6YfWtV1ONcqddWNx5xMvU0LjDRgptS+mpYAZ+awvhDcBW7Q
+k5NdtUb3Of8q9tEJmJMMtpiEOYz23S5dXetFerD6c6S9SB6vHSuyhWcHkJEBfQF
EY+eMzd6HrRDSk/uDm+8VRcC0MzPIFythO7cjvTiHFb48b0NsgDokmSRb7layK9U
1e7skjWFrTotFSvt7GVmEkE+MGjQVPiBXNFllaEh5IA=
`pragma protect end_protected

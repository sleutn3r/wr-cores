// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tY/JCFJc8AZgS1/w7s9j2v/adL/JMW5IAYR4hR6+5MgzWusn/z6H3z9UiwtmFS6C
wxFXhwNWGOpllxcoQnLJk3PIbK+7SOx20qR5K4rZL+I39vQMLQznl9y2nC7g6NTX
aOD57nFPGQ2cvISFvxqsyukI1eRlce6/R8AOT7qHNU0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15888)
XwNwXddYhyNi4nA4rfaGt42gPK6vWQoAE+D01GWR40cEJ5sdYccjSGoZz6w3Y9qZ
Ib6MySH4oO83SzbMp/SVk031Lc9Byk3NeMlacgTkkfGX1OhGcaQ5nFlnUdpi4F6l
aUm9Kng+cVCtpb/oyCXptAs2gWJ5ek77O9p7vvmEufLD6S5l7XPhJ2W2cIT2qRf5
UG4NGBEpdJiiO50cGl6oN/8KVEmIGf2gsgXscwXxPWEEf0uvGf6yX9WlPzAkL9u2
Az+8Uqj7hhhvgsTc8ResbA5opzC8W9P6m6jzCqot3tvIO5/coYgyahPL61K4icka
6vKLbVIerLLt8H7cPO1QRM7zDpOZnjs04uqmhZFvcFk5cbS+pWVrOnfp420/j7bi
yvJ58dlm3kgJX+zjXmltXnHXTrPbBYhwgFPRjOSJGPs5ifMcZ5aIw5Fy5zxy6r/k
NF1mZ6C10bN5U9L3AGfvY2LSjsWbg0R8rAPaqhLsE63hXlroQK2A1qbVFDQyOvY6
FgulV6mgeOMpf/nMo9EeZjieklXxuiDpJuJ9c8eZ1+hV7+x40r1B5IQJ/UIhnUBW
e/IcUodCUgnqsAI/IoaaSEH8Kz3kZQus7vw3gCrePHsKNVMXhhRBvrH6+L+Xb5ml
HqAfc6xu+4jNmVC/C2L/5X+bLhlV+vbPubBhD+s//gOrEUMDZ+K6ZR+snY7y7Auq
NaCxDM8Wmu1pMPTlDaOZtt7eFf1tPzekvqTR4xGXiTdsqQz/J3GOtBc0oIJq69Ku
3LAcy+8G4xQZVoTknUy9I8LfbSW1Gw7tHteuQpjzmulYpes9LDQX6vpqENFVlLc4
E0omK1P305dogU47/5u1DnuKxZC+22p1a0IFiULKiouW+U2iDg52Ca1nzWWZUJFq
8L9zTLZU7iY8lh90fTZ0p2XW+vz9DUKYHn8VTXHJsAKaArzYk5ahQ+S66HOoiSCN
n/rFSOJpVPgnUPwrhNILh6B2SIrnX46pqHRKCQUpth6zwkBNgf5EeXBp/G7LxmDE
w7qnbNA66YulQUrLkMGU+jWEGr72SHSKVVj6vLMpsmjeR3lBGNZYZf4HmMUrk303
6hqlmosB8eMwS7luq9SfGoAn9DouGHp3XsdgViUIoFtzpAbssY6InmGmtjf2SRpn
2L2RF/ltRlvR63x+q9vZHjyNarTHsOwOnZL3OtIKmrYLDbR+eL7jb6NC/MQgv/Nm
fBWTAwZSKJbGU0MYaVL34QIl8oeCdQBsxXlBjIvwYycaGuhQDDsWnI2LIOvjiSfx
ktZFaHhXARrfSZglLGO9hIcPmSgGpZYEvzPK/53H5lsjAxJJSaxDhhmoKzxbjftG
EirVo0/+nYhzoMNnTSftjkj5xWEJEFntHSW9oBkIrMV4fEbcROEfr2af/04CQ4AJ
4PwIO86tQ12IsgnWUOkpvQyz4RwXz4z0uqBxIRXDuFZ69zWbOQraaGU/e5Q8rhAT
zVPDtbw3n7CHrmUyWFpuZ+HYywDKVyGja1I58YzFMHFs0vdRCveHEPQozBeC1Dzq
8mnLCUstgaoecLStF6SXPrOoKlHUGsEI6+hwDHYGC+MKcdxVVsTDNfcxSlZWcYhf
ZLykyt76jjcmnDrmsjYPzNAaACr/tDDxOBqqb01HZIhVuWywvlKXNAkGgmLUMfQc
0ryM8YyNNmicGCXhfmX4tnhZGO022CR9BBYT6mQO5bVBiuNCAFRyhPqL8ypHFD1V
rMpTudzRnl68U2eu3qKAAxVngcaGhyrQXRlefV5SmRDrww081XAqcqJ9NtAnM2Y0
K0xzwh/EXpEDpzcthAVFjBUbn1CO7BSpfhmRc3j7wyT+ZDTQuRe6ls9qSdUHXpwC
AAN6PfKK4uCYuCTo+WgDmvVaNg4V0hvO7z0CmHmhBOMF63WfepOdeZsrOz5SIsos
+x0aK6UnebqCwKK3ib2hRdUM714SeVXP0PGEtIXl6rja0mvYBAIy/pFRvfa5rg1d
XB0vqhGn55ttheArFr4dbbW1jVmnC2W1VvYBIBEI+uBfFKzfhcsfv2YD+ti8g58v
pPBAna6BI9A/nlCeV0FoMlwthfq4ADGj/45D+/Lg/bWU+Od8JSOU1GLaAWrPr7uA
FVWkV8+MzpyebE7VDGX+ZPp02VswE05xUH0edSOVUW0XzbGT+bCsbCqhUKYztpqM
x6Xwem4fEJm0txfXEvs8icN1YxWhDvaWvLeiquzpFKsefDbxeLDG6QBeASDysktF
dQNIVlW7Ou1ypukD4sG7sua6VkGgbKKDwI2wP54J1Cw+g06HahnTbHEG8AbnYI1a
jU0ByepECzLWwQdoVGZGZwKhS4TuoQqRPZUp9rZNhg5Q5LYZBOHPAKJft4ex39oT
Q9tNMlH+zx6k0TS8mC2QuGRfPCHC9GFJ9m/2yfTL3tZ4u7BYKHHzxpC3FwrRXAHw
xAEcM6Ls3t2/lFoefdu7CZHTVnrCkBzzd/LYTiai1LyLiFbakmIlRLWsp69K8gpP
2oXBPArr+tVb6lhopgUce2diqOPEaO3Qc1V5T0rMOQCBljng26IWY1TFyi1m8xyQ
CTK1qkL/xIu9x8gdSwAz308N9orvZtznQfdKtOJmkeqIH6uW1FN4UpYZX9TeoHhN
0723N+8Qeq6u1QjUUCOd1qN1ir2VwsfGu3oTk1b888vlYDiXLiDGjTXVUkUKQqjJ
kMgoMAVGeyXRy0nwJTyoj5MMSC4XmWn7IXG/pot/T1V4XbOYFxdYoASLT7DuLBQi
LLCMsuDxvqu/4fjamghKsiwfl1sCnIv0NwvlpaFzDp2Fsymk1OSWJxzF+woZTzu8
dn+HOUyCK7rwL4az+84xPpte08PxrD1M/jDiIlPZXJUgPMbJybCn4nnDgSA8yqf8
SemsBNoZaaJ8JsmkpgNc91+R28k5iFuLhBSVH0Q2pOmqKHLFiw7z2vsWp75XGC6Y
I83Q3c0+JV/Zxc07gOGAr9n0J6kYJIVdSoqyWRC1r6dC2GsEgFutCiGR3WK39xCm
K5v1JRdlc22fRuklyWvw9LghCndpeYXPaKTVMROrjDc3gV3K4SiQr0vw2spPunCs
CKpDl5Oma6k2yZ3113+O621qIxAFzWW0VF9gBLLZG0ArcX3J5Z+tx1kwgvfbOWun
AWn9thgtHfuJlijVgr2r3wv1I3LjTkAoJkywtHPw13r4hcmNp/YTEZhjryEsWyCt
X/1/g3f61a2dlLhsQ8GGT6gSlRnNB09Y/ox+s68l1jVQfojKbRjE4I1CIs8pjX3C
AiUMqCq+c/5Pz3VIFbCuyZ7ird+YQ/6wqgzQ6EguXAlG6tOvH93dD2sIbAT+hTz1
euUTdBvuBGmDry4vKVw1q3TZ9ZCb3Q22NPSmWg0w1uxEg/k/Ddxy/Tl4NbeYsDNu
ME/OrMJTeT7YOHRjEwACgN9FKATS5ybmMTH5UJddRwX4r+mX+LBQRXJ+zmZMEDdR
b9Fsg4i22YUhDINwso//4PDoZAqzTYd8GJFUpM5OgKevvln4hHRtTt3bwkPbRAnP
yxlX3PSTx3832KfqcnnW0m+xTEB+aGYFOZTqLXCglsE07k2rT/2/17FFU1ix0ilI
bFK0F4BCbStK+oZHhMI2/XVUQ89fGT73zucpd7p3yDZiQwjLtwgg9aA9hrVmKmBI
yBsLPgPAt6ZYtFhXSldAW+19yjGscQUV9X4rQ/GlGiii6IDH5PaKPqq4ZnzymLa8
06P59XGnlhAlug8+2UvD6TRTTmgmBOmbR3vGuWBUnWuG0jALliyIQ0kNMifrSGgZ
FH42iEH8bu5qwvPVbl6LJ27s/EJyTYqYlFaDVy4Ehk7BOHZw9pwN6yQpoWJLTLcS
g57/h18D5WcbmcKEJ2/3L1Xv1XkaIrVG8XaGPPeeUOdhXfUwgWQsSutrdb6iBArl
PJaNJD5qH0Gk0RpnTToW6d6Ui1ta5GWb+7se2estslUhqR48iru1B79L3v2l2j7A
YF42BnI56j39Zfb7k4f0Qp2O/i2/D9VC39VOIO2RCVFDrQ+jZGrY4+byTKvgFJDl
Bo/nYW4E7UMV6FZN4LKFtAnUTO38R2lyl5SDvjG+dGCrLqGYJKXhrZ5NW/U/97TV
fB/NslMKVwYYlItDq4ZJFCA73Arm4BQcO4osgWVTr45qdnTQSns0AjNBGeIEwgs7
RYpXeOK3RWW83V3AvShCFXbpPnarriaEWo0MdLxdkEbgTZVecOxeIvDim2zqPyfd
7M+HSdwldmKCv+HNKMB6nRV6dq/MSmxYq+2MlzbcW7qCo1IK6v9kaDibDyVD0D6B
8eccuzJoqpXrYJC+I13dUh5BRAtc+AZrQlsdzciol3vlh1GyY3z4B8/uh1tq1R2K
Vx9+JZ76kog7ubRKXSozNCbREt3zgDyDGOk7E3KzXPHYnDcybRk4FPhg0dYZ811P
rH6gDdTAL1bSzZZTcMA57phUqObdHnTZRPThrK0yF+ZAgUlQwVGfjm+Ha/T+OFRC
Yv8Y5w33MqbMeIquaLCbHoY1O98Peu4abK4baQjqmhVrABQqIHaGJmWZgMuQoAq1
nh0PK8yb8NYZi3EWSfFFYaeT71gGffv8JRAdT94IKZRFegNzs0KBh8CmiJ7wURm9
qMLjKASygR3mL00zuhQyvyAJ4NKQzkPUBGuinNoh5t5L59PdsI64q6cI40a7R44d
M+qvEL74alY65g9Jyt2puBDbL1IXHTZoy1pVCYp2hE3hxtv209wTTJdVyRfFbtR8
Enurcf6TjizVYHpDk7qnHAcgbXwxAPtV+AnjznQqn0CocPiTq2zdkD7Laar/yxVC
6nvYYFU7+i6IUd4Dp9toxq3u6avQ85pzhizD/DXuEGdD4+/btvzYNxNkWphQxr6u
PaTblOcqwpZhFXjPf9uBxWf5pRJ6wnlXhqmlw5U9jDCokWufSYYVSrifs2LgU+Zi
gtymV5a3pNxB3uvbUlxI8DOCzxDWKt1KKqTTUd5eKnzCoVb7ey18pHBToEFtU8oc
JcCFEqwlimM8Mh7Xy/jLIbiadclWwtGGfA1UJ9md8/tXqoLyyFdgWfJ2/cRdwfH7
rauohXq+9ro/df4MFk/CX8yAY8bjFDNhjX1ZiahPX8vmUoGebS1AfEOHe1bmZV3W
RKarJGtay7iKWJSKq7BPmIzKA74jcHzmEFiqyMJ/j1cMOFCa8HwZeIsEx+9aCKjW
IPvdFgC28LFJR/BTNNDN/YP9qJ7vbS55MPtgAavlNQN26JidmfjFoVpkDTVi7bqA
masBxnOSA0/RZV/gLzMxd8YltNO8TSE4Gdwu/PCZc1BRQTAuy9tD3cBoDsCIFxSa
/ZPDBjRKXIRcLDi25y0EhhZMQmaj83gmtYuZwe66OpNwj51EbTV8BwAsCM9RpMYo
WQSZdLWcu3/MIkbE/hKexJDnEN0iJanag7EjZj9gyGLz5W5XCAn677JbUydFW6ZM
lluIqQ8OKmxSg0C16q+khMWbJZJieRATOrISNCIqz+8+FUl2Wz6LDPN9IiHox2J7
DWYixswpyv0dTPaAwUwp06W4csnkAsop4/Eh0a690sDFdjiGRmx2WaGEhbnF034b
O2FH1FjnvDqY8U5eLMm080Tp8G/Q2t4F/hwsk0OrCIq+6GGN8mf9S38pniTER/x0
bINjohqoip0ou6XMFIeChDHGtmOAJ1VaSTDJyPertNlNK3FbAzrgcBYJ4epAoS9v
i0b67Hu+vbmnd/l4ro8C7hPIfduMb9LQcitenW2o+Cx0wzuabMM1ftRO44dKMF5K
2o6063UtBAAxJPmA+212CR1vx9B0KwJ3z3jAL2hwZDbgP96dFh4M9pRKW7beeLz+
+GebhKDwK4tDV5bsD7iAQtCxkAgcAgGOFdt2fWAS2uEjBzctBVyEqtzcwBEOlr8O
qjp3G669XJG9kf8j3RFt0sCp3no93zY9Tl2SEQJL4GAHevh8kPGsfuJm3zzpuRTu
5LcXT4xjq0yEvq/l1oL8NoCSnXpHRLvy0OnrEfOFjRAMVZ40BF6esBJyfwQY1iWF
XwvRXtG467LpVTsvtmZ1EgYUw6TEgY9bhU+GHBsHTlMxcDe9VhUzQtt7cFNgT461
FnGFroKIxg8xEMMe0aUpUC54YU1dVStftHn2vixV/G3ABc+SnbRvMpLgPcLaHSwE
NuqBecla8XBIWoAtkBlqQk49FqKuRfw6LtUimdlqd5zUKaWrT2+burxSAVQtfp6b
waYakFpck0sBju7OwKWEDgO8HQyxXhLJTnc8KjNIHWz9MDMDBKLbumrJ6fjJkF9y
/KsTAApsouo9/nBM7HTao1o+Wl1ZRDweA8aEU91tpvNAbSpxhL/Mss0+cO+mEZhj
bC9WB9hFqBcaXMbVpx09LcrbSST0fQDsafC9KdM5cpWIPauMKFfOFjU/kH5gBaSB
y58YnLUmPgotI3e1f8rIK0eF9I+lTrvbGfF57NnajbrsO2yARZurn8m3grGUFT6w
0YWVcqa6d1hcNKIGGySRepmw4hAFRozdJiifm4ibWSakvBXSoca2C2Kov2ifIy6g
wK4dBVbPGxaKrObCTtmXj7uw7r0Yi193ITb8k72/FpTL+1Ejd0tXAcJNIOwXvgq/
s9Dn2wlbvyodKZi6WY2uwiwunYzv+2Wc9+lBY5HjNuKbz9pJtAUIG9C6+vlnFJ2q
eoVA6oR6uTATn9jJsS+AfCtmLuojkqEOJVnQ7oyVyhw8mRhdC/QZLkUTbXYPvZzc
pI5WVaSixG0ORX5IfIAgRFjx+1PE+dbZtsGmjiMFBxVghKjjcC2tx9ziZ2UDFbav
3OU0dfhIqmEakJLowZ3mwlHBUG/OT5vmVr6aFJZaeYUAFVyKviK6XQ7coNEI/YrA
uCvCA6S5LLDGjjN/D0ZbF0FrcgmHRponnbxtCZVA/uCSxdZBnrZodIBMyif1TQiw
ZjNIGriojhMh67cPB+2oSrkN+Y23OvUpqxBnmVzj2vnlPQPsS+KDn0PWxBTbUZdB
lv1ipnPxk+azlEwi5AEaQMPkdFFQqruSnsx8zB4w5ZOk2GELR6f4bslOXBDIRPVm
wcckVx0RQlqx2uctszEGL1bhfu0dskBHOQKiEryswX/ZuJibxZrfS3qGi35qF5a4
7WibZSIkkc3lJjNJ8O/FPMjD9UAgrP1M34L7+bnhn7goa7YM4zV/2PFi9zlwtSHz
0MKEul/nXRhpIObJfpNBOMyHN6FKn8EbU6M4dhSAi+uKY0stfdBzWPhJwEkkit4D
4Yj12izJYl1h9UpAVbri5T9N7Ie5jtFDLVvcFtZggY/QiTcGrWyrEX5TJ0XmFeGj
p9AFcHFvrtJBiVbMHy6SzHxKEMZmKgx78yAlysE8EYfQViuwgnIyHPQoB8LnrLOJ
nYdcx+5f6UYb+nxiBfV++MKDZT2NJJlz1NU9qCtGUBZTzdDgqcMZ2iq1m9Ov6AKU
FFKVtI6g/Hqr1+x787i0oHMSjpaH5aChHFoHQkjBu+9D760z+tsv8iOryFh64E8A
RT147xv8t/v87o/Y2Q9emlGagKM/7f0smJ/q4m/+LzAaVUgd7oJRXn5OaxVAUXti
p5VX5NgOZ7YaDP45OSnIDjdRBqPXDvT8IjqzqjReGTGpJfNNSXEiUDGYjZrns32M
fb2chfB6PFyC80DZYNj+JSFknm4HCA0VvVhG3tijzk2xylUF4xv9C5sVk5mkr3RN
Xc/kO8qT47bBIwWgT0aunBdz2LS9ezUvrbZASOIqAn4E8VVHf2qgivgl6yTpzW6M
nH6ZKP5FtSPdV13bHvTDwu0B8Ib2mKwG2A9ayFT61yni5Svn9rzwvvWmb+Umx1kT
3VrHWHr//w2vfGVaE0bbp96+AHel3QvAbmIHnGh3gjvmZx2xbi0hWkccskws4rvz
qg8Q9oc9w6qZ5UnUNE66mm9D5YHXRJyXL5p9F4k++eSohYRmhDitiy830+x/C9bz
51pv9dObM57t9QooRd3xVPIJYn7/jkUMiNYhhy8j1GYoNTCCo+b3CG+9/D2SP5xs
fRtb7xrQYxW933pgztCfctf0Tdkk3LCU4g0rZBx6IXqzrU3HmDYreVVGmZFlgT3+
QoAOWgPt1TTiZa1FAPhePU2Kl3/ZiMbA165xAcbFywFHYW1yfM5e2Q5tNffDWuHr
SClzlP6xYBPAPB7GDdTb4zjcysfPvWd8MM5ZPhsXFWOrgurX0qpm9PveMBxr1feP
xPGVlGbpNtBWbaTF+zQEx8YGjpNo660jX1c2I7Sv2OoQuqDAnFer/cplC8R3Like
Nl7WJvmBIVvvuho9zs6PIA2gx66+a3UOpAWIx7GHLv08xLaoXnYv92V0jD8kqizZ
VxnNMurHi4B/Qoo+vtCL0cePbULlHJh654rSaKj4Lezr5hPuhdHY0Gz+efHfa73W
Gw2kfIhfdC1sK7ya+JPiGu0+f6Qxsm0gBSfIbQsq/FuF4sBeHJbkH0b7oU6XqwmR
7hwjf4RkLcIQsBaMgi2aSmv+AqkQnuF09v97GK0g8tf6UiZKe0vWCTUqcY4A3ffR
l5oQse+Tj8pAz9tdv+iNUe6kZzri62tUwuBt+wJ50kWnom98ImhpbgEzgVBolerV
ojhqtjUdlQmM2JQz80CQSvuycCFlYjOYHS0ei0mwTrgJHqGhPhL+DPgln4c5i2G7
eFJyTKKE47JHyROKvy+a5QofUwNaG5LE1BWDpNLOCwuBYvLm3L2Wdgz8qFGsIMM9
95Zp+QDnW3+qAMbVuRKINpXyj5bxi6uomHIEr9JPsEKp2Ca5E9ld2GObcFxcL7Ib
JxSomJC9KOU+NbIeVkyQ+IlvECHGCqaqq3LBVDnV6xXKKDXayxz+KCk0pVZzuRc0
65utY6WtOkHdEveZPh8VDhFvnv6wdH/90oHRfvexUE+qOXBvF6lzUYz66BfwyHvD
hzt9HhVWoyXDH3xMd2uxRIYNXZneW0mOwAJ1HLBbl9XOKyD++HKaTKDsPHQaaWPD
FU6wXrOX0o67URyGXegtONdYCDyVtHO1V+IgEPx1cypeq4aGTaWeZZYAxWkfdoB4
4aoSx+v6+OTVKX7JdvN0cUaBgkdUHqFgimH6xD7vVE9vOpiqqV+fHNB8SNcnsfjk
+fR1C1Qe6uXdYNuQD8STwQAiMS9Ajxy0AY32hyA+WwNh5AVPYJrhLPrBPACwcAG+
NxFm24HJm/x7yM331nNdRRVJay05ulLUL9p2fePxN5pSrvcYYNtCoWRr+ueFWYfx
iSXi/aBxsVCFQ8a4fDrUTrb2Dv3r50wSlS86WareJdFZc8ECnDvNJzIFMA0BbQ5j
KqwXhSh9qR9jG6Bmrb9UmK1cgKcYOM2ELHcRTA3QD6ZmdYZBMcaUyJ6p4DAUpZ0J
rQC2jJYJksi3CvSWWwPsvgEnccr6DixmXMOlCMQRZQpMY9x1CdSmHGPZFLW4UJ7a
qPt1E8bOOj/pacpCGtS/SwcRqdFmflh96ba7P+MyraQN8+SRL5x1eWx5ZTa+XICp
1vlETMI9XPY/QsKtOySIu0A3HhmergVXfHfqujVRkOo2tAp9ygq7+BOdb4SbzypV
A5dXkxPj8gFJ4BaeT0ciwLVCJ8B41ZGKukbVfrCSP80hscplHUrGfMWVMZi3ASGE
Pp8HDTo93go0Q6+TykgNl6bKBFh4TeuwSQRg5kA1GOkpoBvX5mkY/QX6UzwXtGDC
CV65rzfOeeiYL0CHUBHI8PidfFr8cukntDn9OXQzxx/3a+n08sCFplf+DWLwKhYN
S/gQqLpLt/3A4dlWm5cWb1W6v6N5BEo3mkmLFxljs4MwEMfySh7kkQsAx4/k/FRI
kpNaM/VH0YUqMJJ46pywnXq4zr9KeWj/YQvKyvxqvyOrRkAWhyFqT2eDcGPIyQgY
urbTKj2L5HSCyncej+DHr3WKvtNKXXhmnk7dcmyS6PzWPXkysjco/8apsONe5ZKv
pOlCOqorfVp3GgpA5HEk/KmWbCRVa6mi0o1YNPHS7G96K5tIlp9XRkW9ab6Y2JBT
PBPm7HiY+Ou6c9GE2sSMjLlNrlkh9C/g+DSunTFko55JHYp2gzWGg+Hwtt/SxANg
GQe0UdvigdqOBAousg/rFeBhBWsqmjcEOTuNp7v+AOmS//9xGoSTW8x+p7BM0kzR
K9Ebp0GSWj7VI0kc+cnGu1UNPfNEHbVGwbAiOh6YWQn1v/16clLJXO3Xa050da1z
sYAyxhz3tL7Ac0wPn0z4vHm6jeAeQXbGUjpN8sUeYaV78J3bFkak3fEBKGmPCZkw
LpcA4A64lPKakHdY1Zp7AUBgtQzXDxQt5DShykfCZpbz/QsvMyT3S4suik5vuPac
z6Bc4RzMy3akW6eYIDP/fmIxLrL75AJIhR+mcv/f5AtYq4JbrT96r/p6aGEENNXd
AuF43ChsWCMujl2ewRTmtmu4U3crpgMq6atjYhFHWYxbtPn4yg7CraJppCskij2b
P+XibJ8+T3zdKXEKwyybuVheyR61XsOg69zr/dmRU/H1RY1RirvDdoZ0/FfnaW/7
blTJnOtF7odnHrvf58072wxX4at42uRikPg5BvIZmAUUCbu8aGfW7IyA1bcRK8iU
aXGa0Isz3lU4Sm1AjiCfUUPtUfjNL/PilQXWGUK7I0yENPxeO6oB5o/nQmY6zw7x
0PUFJHtOkcFrTy3Q/qCkyCCAL2CGosdPsYoUsuMWbToilld6QoovT10id/y269Uh
qpIi5ZGw+dQrlL7NCTpMQkQdJ2AHz4Mt6mu9tGSEsYxoK35CoKTDES0tacxxbTra
yGscxEXSHtsmhxIVICesYFPzsMB7guqWzs16COvrspL+DaVNvrEMdTW0nv9K8n2n
6bnzzNd7fDAcTEBCRk0GiyhTCT9X6Cx8cks7TyXMCS66+xMhQNCTm86eNJ3gFoWh
fF1LQ3Fn5Q5u3TyzCu1IH6vQRSL3oY/5UZp/t/hN5yaqkCEn3VrfNDzcfR3WRqn+
4sZC6bhH6ibX4WeQNIFDrW21DcNoJdQqBX3jbpDaVEPLNxOhD/9Zi2IRTzFLyAeJ
Ly8twMhMQjpu60KxStAzHTtN+EBwsb79Tj22e01RgxRR4schtvmcL6Ms6WBnlQ2c
DqLhfQRtF9hhH/SDr9fXhfd6DkPAGEcvFVBTV3vDu399GAswxDPNVmCDk21uP6t6
/Vp0E7PGYYVvDXlTDRsKtYSMFpWV0NsuOYrQHHa/XEN9DH90ZpxTl1x6k4Nr+VY1
mRRJaNLJ0sqhc9shVdqeIWBa0sO8Gnausihj64ryko/u5DwfaRp5JGxUXCVRuS4Z
kwMT+3iIU7n3nEYkuNf15Z1uRf8k7LYoD4R1V4j4Qoh984oZ+n7tc2A9yHsxxm4n
0+RlN+31g7C7rJoph9IYEsWyfS2FULU6UAqnfjguvl2xyExoFMijfOf6mVVziqAB
WhWgkQzGM/xXDe5ziXJJnK2IvoWQqUc/9l1hxT0gfWNWVgk4fiK0smETXmrYTN9R
TiX39bNolIRXMaiMTfFWtcinzJaCoYq5qB6JOZdwXhu3whEP7BJbb0hHy1pmeeqo
3YKJUbA7H7xvOayEfNdy8lPUCZuXwuEtG9WiBEyuepscOcTE7kXawZT/wGYiElWH
AGXk4RqkqKoSKu7MOKrVvNS5NS9ycfXHaT1UjBOtyUelquOFDUEjNy5/yzdFP9o/
DguYbd8rJvE6WYnkyJgojpEQ1w9Crt3CKVzmlsdnUPxIfWlgLcH8VVLKdn6kFw1q
LhmH8ZzslOYR4fHuQLkg6PrpiMcICYeHBXCSSG7+8cb3Aun6G7lnB5F3sjJ+Frpp
ypEOs3eN58pPvJqAU/b8JZ6yPz0dSD71U96tIdRqd6TTwyT1F52fuhpVz+tUfX4t
DyAG6dF7WNTVKGTEhEByxoMn7JqDvtm+7rDJScHRt0joywwNnB8cmyQjpjCiqIL7
Cz7Xe6Lutwme4eUW91Y8MpTBL1qEfS9yZ39GjLDfr1vMcDzCn26pKGibE0LaxdqH
FjY7l26tb+qxlfyOdxGubzktV3KkhNCTweVe/H++024KJPPGKme4SOqjpGWEgTfc
zFC9wc/7zdbDqYpQIgLBz1jHj0XozMxSRhoIB7VEFOwFGxUjPB7bRHENZG6bVTjs
uMoj9S/HVwva1pA61U2AQFrn75SA6YS5WKjdwHxoJwa2dLpUrarHZOBIx9b1QwMh
mAH+2ODPBoJtjuQLi23mHZ+2af2BWx25EQsRsY6om89k79vAeSCX5ExzYMp/YRoo
W2yWuqvIeL8GsXu6zy2YyYd7yCJJDmXUGAuxPwzc3j8nHLscSttJNVGxL/+WNYqS
1LNNmi8AfgOgIhrxFR20HziflHFJjY7JtUrd0BxOrFvRd53i2Rg3jH7cJQx4DnO9
qmdNwljklQTaw/mi15wVhLVspwYA/fSkj+uOCHRqRPof9ozzNWuwXjmUb/fS4UoA
K4kUmjheSgSQrWf6DWEMKrCMA3h/goqzm/7oMIQdBIpPViIxC8+VOL6l5OYZ97a0
sZ7VJIVXeNFerrYKPdYMVjjFnERzKnIul45vvWo1m2NnPjTi1lTz/ogVGb2Li0kB
o3ZLzeRNLSXRoykfWhnNBVGIUdJpsZkrLguM5zOlw+mI38ICKtw/XONiQIoOrcqZ
nqNh3bXPQP0ZzT4pKN1YwNglctF5yppeOuAUBRQoB02igsxfKjkcMBL4JIMQYR0h
6ISF59izKPYZZ0n/t0aq9xn4syBi97JjMXESaePm+dDvGU0rEHE19J4ba9sZG4os
hDZrYnEvfKXor/ATra9ZSfQcDmhyXG50cqNY/ks5GxoAAowkjOOahobyDfm53eZ9
PrqOjAtTdny1mUj217IbhM6aOaSG3sw7la0ecCPttaLhIrRU5KPb15cgFieuaoXw
bSDhsq8a/rPE5CMSw72Sph4uzPTJAquML5D7LY/pw2yPB9zizuE0LmY3CKtKqz/8
MG/FbDaxg+2I6uotPl/cyHh9+g96A6CXiF5hZSN9Qz2z0d2W4l0d2+W9p5K2jiLm
Qkj44aOBoSMtSGXk2EgLe2QD5/RVhQbzb9ViM6j8yYVuyX5wuio01F6wto6BbxRa
RQSTJn4O0x52DysaaHXnprC/0qB9VAAUd2Xvn22QyrTw+dfnzlsPaeHxvCYhHVLE
gwR+SoV9uXCKX/G8J5g0Gsme64dPPfzZ+oKqzGqhdkWqofdysQQWmZxocZ8EkdN8
rkIyTL1G0pAj+BzPLLkThqP7/iExS7iKiWtZBLXoPmv2mugM0uAJEJFl+ZIFJSWO
/9eXJGcPVXsd7Y99cP63QL5Cr3DiEhtu+L6d2MHILFDiWLTGZNkE6lG+DRywKZ+S
yOaHfXKw5PE454hoeuMaMsruphOPeyiGa3nTMbZ6jjUVzKQmWQnM2hKkDdPTLUfF
lly05aB1q/4zK/PbVkWEb4rFE9podMaQSGjj+rxRyEtpO4NgsGtQbuGepo0m9DOv
zohyksObZI6YBpxpBB9HeWpuJWJEWBJ2kQvh/UJ8jfrpvys/38FP5i9fbdIITYWa
g4zgPYLzsgLlCcVvSVg34FQ1GrZRvlz5d3qbcWdMirzsscSIj4XrUJVi/r5FR7Fw
N6S5keXz7VF9RVKE216fdZYznubx7WbyUTqtlgivrusPFtB22j72Z+FXLmmd0XvM
ipoCRIL/0MWgrivWUBgaR7R7EerFh6s78o8TJ2CcOt1i2dJS1KPJcpiwsx1NK/en
MP11mcyQlfIH2RxMZaAlYhyJBW9pdaoB9tb9B2/4Vz+Ls5lEq83hveeWoQr15h5q
PvK/hgftLdabwddWt9/bQO3DJuS024TcBh0E3Ik9StZ4EScnwUxVjC0zec0um9Ov
Hyr1gjyhVl39LveRgAb4WsVr9t2mIpZ4NI4MRy1SrHRRZsHmNZFLgQU7+2op+N2j
caSZp7U87h3zh0SkBcf1eudhwv1pbVoOHTg/tpUCQkPBB+vq3kzjY4Q7myXcttvf
Y6nqdiAUJ5VNx5m9zb++tNenFnleTyiPAnFrOfdh6tQBkAPHFN57IQ43glL1OdSz
fMkXjQGP7gJDxGsuRcgtzghG8PPVZhWC6wXKreTqxV4t2+s5tWJE5MNzq9RL0CuZ
QHqUr+T/F551joO3WyCDzvHLPqpSP6aI1WycZ4NoaYYkVYNRH9nAHZwzd09Ciufq
Yo4b2A1Cfsw6DrRhkmKY3OTK1Ak9J31GGcX5c9OcdSialdMWBBXdO088ElrjXVVH
9UM12Q1jsL1NCUwsyQLbQf4rCr+LozoCZVoX1mgviQSqrysr8GnDPsBLqJ2zNWQr
x7Q4mGD2EFN5GLbqjrTOS19Ad4IMhLW25O5l//Db6M1AOP2cBdgMcsKKvJNe+6HF
+kMTIqc4zuvM7DpGrJzmU10TqZ+ASegRvoSlIj8dCojnIi5+PDIHtOKYaKjHefZY
jryO6hzJXkCFrAloKg4aklwcZsqLtr1qOmdAlGfbS+WJYbWgkg9sdmShxXa0YJaw
nDoGzeBHJlW22Rdoh8eU8gw0ZRJ4EOz30uaUeuuXKgQwJTHw+R0Ja68vcZR4lq1z
tHlNMqRTwD0XeVB0jptax4kF3pPDPop6rSltDvZhjAi2eSD9eCkcqzK5IGpqY8RE
WpPNpnxrFhZRf82Q/cptOr2oJQ2u8wK+qmoLqvErlkXc7Lp6hJZdM7IWfuWrIdKl
wVmbOxVvshSXhx4XSLhLdaq1tjDBKg7diDiuJ0DLbQxsHaiCDPOOJWUhjig38JQ3
uTAU6J+l7INn6fcYlycEOf0xqn49zpDRSe2IgetQjB9iORNXmoH1JOORD/gJvIZm
8zL1mnlFcJ+yzmLG9bd1c5SjcxBj5tmN6V5vL2JdkpjoirQVR/VJykeQFr4T34Dj
gF6uxyx1fCpbWks7bo8qSQK3zHeG9YGWzYBY2m4awNoFvrUNHpiC1vlEbRKJMOma
yZ+ivb58HazFl0whEViJPy7Xz7ahiohNgc7T8Oc+MZoKG2+XFbUNwf2QbkJdr6kK
GEwb0ONVcQnLm+8hpuBG2H02Gqt/jZ6yRzfm1xcBDJZvTccYZ6FVi1SgMjXw4e5e
IPyEEkkITeEpEuWQusD+xvtQgger+GPHAa6mxSiZnWQLP8Wa9/pO9sh27psAPFrW
H6ORajQNYWKIur8k6bsE02f7nTbmEJzRIhA2+jfdIgAvkCfiuV5+S8vd6Siog48A
TWI99kiT2fAZ2Trllh3tkfel/6VyWETgyPEFk34M35f/z/fizTASZnUiPOXBVL0h
f5cGKE9hTS5dYEAfjI18k/4XJa3/eELAZHzMJdFGaFkzscL9mXk6XWbBQnRqJLIS
sktsIK6x0jC1GOY3oiJX6Fi9tLYygVPRjFhN3RoayWC4J+2pKqAjp6zS+KV9fQPK
FG6mqPYgjcLFmpoS5znHruMZxLqv2PPX+3bS+Hb9BLudWA275ZvVnrWe7o9tlHf/
FWWWsIJxGwckc0ejlzt+3wWhnTaW3rdR1vNpS3NDVG7qZvgShRn7MII+gRB5l6UT
F6JOnqDVx/8HZHqofqxWQqu8ufyxp6LS0YgsvMjBoGriFZNxGmGvkRHCDEXIPush
9LrcTGRCF14fHNFuccQ9hHVpDz2o9OWdC0XgoV0EXuAjvC3CnXuDIjJu5i1tMJK3
Drvx4ajJQmFNJrnxC5VmoSqeD8ohetX5gT/W+A3D+dNu7CbeXhGJnJLFSQ9m0nWl
WKxuKa7JdbzuSV2a2VN6tvE8gg2RTLpaBYxCNUbVK+A4j7S9k2Mn3d3/Ov4ANJYb
/5p9zGGLIR5Fd5mtVe8R/4/0a6h3ZVTGONLtZRitFoIH5U41Xl6rHiZ/Dh1FhGuY
MKkLTYTbTmgsEIMRP0BCssUuavjVYR8l/ARFg/90leUIkSACO2/wMZ/TmBN+hfp1
gmdqM0SXA9m2eVkDRLu7fSvFt7PVIP8vEJK0YrtcfDM6An0crKXhi8B/4jrKV52k
ICJXE5nvCV182jm4VwtsG1JGDgs10wCqJrZpCn8dbFo6Zqla/XllUi1vwU86jaPQ
UAXXpkfWgH65gVIuzWCcsU4MJ3eO3lRnN2I+Dv8RLwouEKftflb3UK5z1DQkkJXe
gkxU7QCxB12mFMaXy5merQRVJe/qFQNTk3tHW7178dpJgO+44kUfliK4hV5M0wTL
ne3wQBSyp7qXI4cVCrihfAu2AVELGjRP8hILMA4O1h9VsRVKJB3u1JClJOOQEQI0
AZTh6HFMi0e8/G/k3xwDVu9g4xzHBk1Q+pJq/yvzgbfI3bmI9R64QRs9r/Y98KRn
NjgpuK2Ji0IgocxbXhLDFO4kT8uK636iMY6T0zAe7wjDXGHMa/WvuW8n6lHWXknq
pAsSx1ywGDR7rJu0y1zVF/SsUc3Ady7AOjK0MOrRNP5L6HvpNbBGL4OgXfgl74XH
W6/v0dIIgc+djE99pR1WRxOn8G4ZxFmOYmDP0rXEeYOzW1HGxErijs3frhEZTpNu
6KmuB/TnB9BB3VJRyUTQbbYHtsvEZvKe8kHGiW6XSkSNYgl9W/Pv2WGhfiAuc+ur
2o+Di/k3sAYp4llfV3K187cPhhbTQX/yNnp2j2qgxL+3n71LvYjpo0HzViTFsZrK
CEer5qqxWifVC82bgu5jRib3dmTAnrc7vrP9vZg/q778BqbUuME9KTNnCiisnTZX
6L0Sol4KmAtdr+bz2DPUzz+5SmDGwMzPtXICllkt0nM2WS0OI3oemdFkLyU9OHGD
ELx/2tqp7DUoi3vueRMpesdflImiUTcHeCW2WJVaAzz2MtXRReagbyfIYc3HlCte
22+NQqxxT+xICBGBaz4B/U4q+VnIvehsMxsHhK2zBooh0B9ytT4ztmCoYjjZFEJw
t4OqZPfV+chE4SdAGIQ6HPSfRI/GX2RF+odkrc6Pj10ujhZhi/neeuzJgpzFtghi
BXlghvPJcKh0X8XDqLzWRchFE3NPcaLN/Y6ewUT3IqaC1MT0rpYaLtbdxpmXQGrk
BWcE69VRvTtaTkY0iMjVgGnbX/+Oq6gzPyztK5p3iftQdiuruBmURUFLAcKqbF+Z
H6Yib0vNzvSGO1/DRkMGr9ntFijqDaPax7hnK1jZxh/DKQozN4mbl1VQC4loRdz7
x2H5f6eHt1bSG+itfygFHbb15h+bai+MMlA0pTcj2qKneEkIxNatOE84OP9VbNcb
4Hb9HDAU5IfLfxzgDLOKrqiuzIW9wg2KQPPLuJdPcdo3/NMkyocHaOSsGWV/Tqyc
eP+xlRvpG8N0qUfypMmlkAepQ9uKrRIBDbqIZ0ZmmkF+aEV0D6OWcFaYN8UIbziV
6EI1l5SwJWfH8fbdvScL+LNhc4fBZbZWUGB7dkaDcStQeehr6UpQUASl17hVwKEl
OJ8zf8sN5+0hJhHuv9MY7AYjcEMbZLmPml1+yLcLTJ+9hMsCwT3GfO1QZiuJDJHt
PBBlXiDMLVwjZId66aO0+76nKWzvNfygL1rJD+M4FQd69MpwW1BqOT95D/2uvU7y
1ILUTYCXLjlfH4kVgDmBrKzb4QhpCxJ4sxaZtnOWV0Ph5tKatGb/ePCsVQ7JHSK2
nBCD2mnDxTtUuPZ/Cp7by+KvO2x0v6xI3e3dM2oIweR7Ha6hhXeRbSnioMZyl4b3
PAPIpFJcoDsofg/OMExTWJOYl+ALLksRaABMUR+E7HHZC16jGxAamd2BTo2uLTZX
4cdlcMyYLyRC/1BWOs0lGSm28JF3RQ2fUI9uXKeqEgdxfW6hDrKgCHbbvVHcqM/j
mDluS2mVaV01CwNmGMEL5TqlOnlJNLCnfFVh98Ao1Zhp4sDbwDUZXQOjW8U/872+
HxZZjws1Kem66YXRr/x6VOgYVJofquFKUTzHEiIHmzPO/xtC2Hc9k2Db28Ze33Bz
CXNlO3KZILuMPhvQQ0VUxF0Ss9g09JzDrw7Fp8DD+SSs4MTQoiMoTNciET71jINo
34PvC8P4Q44S0KmySovExIRmppLpZ7QaLh6C5Hg9UymQnFUrznYfcwAWvYEuy3c7
qDSm2ypXggUiqJKZ5Qmm16LBYoFIigjMHiP0E+c37FJK+u7hWYOfEy8/TeztpENH
FZVrtQYYz8AT5xKPrft4gcXvqv30NqP3qKoLtF1grMAmRW0x8OWthAbTxnbp4UQy
GdRRPdfwvU6MLxWpnzGvKvzPCSKMhU+iJk11omE0oSi3f1ybJ+aWn9upYiXqJSIQ
gjesIs7ubP0dda4NJ2NA+dXM9ZToIyaVzzuSjG21F2G91nJHvTVHwCtOjVX9ZVFy
zc8hZonpESF8kFqi11Wpd1By/I3EDWlTfsLZa13SdNlUdpgZ5UmLD5Tr4sGc8xXd
R4kwCm6PJwHR8MhQ9evPFTRbD93W3IfxKkYROKMZ17ld4dH7036pnlGR5C5f31bA
oQwM4/ZK6cgRy3Glc4egw9s/wkcDlJ57zrFeBVnjuMMREFbrsr9iHS5So9Ssw6Cu
EuneCG8gs14ezW69QFP+07uAumaRWEfoWC10aoAcnZnpdiekA/9WcvBuzWKI3cIi
tT4OuYGSdZqxZF+yW/VtyaeOlVrXspwnGE/XV7phTvVV6hIFF6vgmCrzM/i1ilk/
ta7a286OtoI/yYNP7ALg9XfD4rOiO7/dENrjnM70G9Fg4GaSRxXgmp1DxyKloJPR
vMZCjdw3Abkh5QPV8s4TE64zR8P7YnwU7e912j9bInTTXsihnd4zNt+WsU7rpuOh
p+yMkql9NSGI1IU60lMhL1hirtLMfOwn5Hpo0NxqlZ7MTx0gkLiVzgeYBomYfaWT
jxOUWBwm/CNef8D3Uyi1tS349+7UyiXP2/COqv4S/wrPCWnH+7gbPwwePkBHTmie
RxACgnRuIybVmyjk4C3fz8H3EMXiL0FL9Yh4cUtiJEYSgCXS5oLfr3YlTCrC3lDd
R07apdRwGbkK+hHEhhkGSa1WJ2frqEWS7tt7s4+UXnKbrCZDhSowy1MNE2B21osM
NXMHQkhjWaJSkAA1H7A5LHKvdXHwGhlBFGIMQSmRFt26i+JmDeQy6Tc81p/zUmYK
BvF6R063xkPuZlR3UlhKCWQR1OFHBxHy2bBCtocO3a3XCp0OX+Puo4zpVkWW+Fme
G1RlZUIxZQWc32KciBSzblvbeI6zy2+7T3oQ6vuG4wuHfqw4LksKxJqHn+tA58Cg
n6KLCAOI1wuofSEt5V2w6Zdopse3y5LelBZEFgFzRTBxAWZb0MIy9KL0bNztJE4V
NcmYrfjOC1obzWyYaN7ZNBu/+f/01Eq8ZFdop4UvXFySqTe2LzN0eTZr9hkhuGxa
7E+D2L72iDhZj+8zz/Xe64Gpzk6uUuzOQhfZcwgnBQSovVetFN4MpzXlKre4M93E
eiEVoCNOLKb0BIEPctOoJPuc5sXB/At/OvAjOT0fGYBp1FtfEYVCrcNxX9EsWEUh
+IORWAZBx2NBt+sNnGOoHfdjJzkQebxDEQmR15TuRafahu6SDyI9iS6o6XKinisT
/UYfySVbjN8Hz8DCJPn+lxXpWKNnHThrqd4AfPEt3JQkv34qrLbk+zHiyKWFfrSR
XaoITFbKf4u3wGyv9nVUH3sy1EaOzCrx5JDRws1u78EMyDjUtmJzFYHiRwb/xajx
PZ8zh0m9KBCG6inl6/AFbQzs3lb+jYF6ql86CZgF1zHOGwh6x6rdjiBmhdXOmGYf
fVT0Ist3+ACQf1SCf+9OgR/0uI+j9ueY6F3xZyfCXM5WZKe1OW63Xu1KmADh5A7V
7g63WFhPj+SbZRzwl8A4XyPn189+M6WSsI5hkysblcS6J9AC894GGKAfE+pAfCmQ
zKyqsSdVNZqS73nuyq2QX6A7jp5InTS+coqPLfFibK6rf5vgUNl/TTLdKqXwr4nc
XL1J57sJucHFlwIoFcEGBylHYv1x5zVPXxvBe7toKgYblJVn5CSLWYN8i5Fn+Obo
rIBIVkG6yS9rqLImeGYgRPF2fuGbiskauAvkg9LMynYomIQRe1XOKX7PCp7l02Y8
gs4KdDmt6/Cne3JRAHdP5juRBteEP0O9hqBwZdO48i7Q1mW9Cox5cIvzkfek3Gjo
uRZLzX+1yiZnJ7oI0moF+WH5p2ENv3GFRZHzIl4Xh2C8SAPiubS0WMWEPeNVhwbY
4HKj7ZCrvYhE3Rw/CjSduMYijMQD5BzA2M6SM0qbkdH3d3QjF2Yh9yAg2TCtyOcr
wSP0pYtLe7z2/xlwAFpA1IVM8vt+sIsHu0fq2kCrH5uH0N0wNIaenxkGM+/BeGSe
GmpbY6gWMsEW0Q8jujeDjfZ3g296YIbsX9K0YzYND+zw1MuQHPY000PhUJR73wvE
/vqCmFQlyeV7pXgIxd9eHqWyUs4GbYjI/BgW06egjbq29BAgBRtkTP6rmMq5a4Xv
UwNFILZSTjQ9d9dkcL7eMJbZv0m2hcrGkON8K2xws3WA7k9tjhDwpWqF3adkR0vT
WPk93Kwy0nEoQnF49gAnR3N3zbEc83xdlJzixsL03QC8jko8Tg/aJwXUUqhSWGNS
ZO4sRInGmdZTr+JZiNlHxF5XwgMPuvv0z/EklD/vuPxKjyn4jq4M9PUxRnBF/0zY
tVtTsxApOmCxPUwF+pXM2yWgoGnKFceQwNt19H69lypUXR+CEAGZSRVWu1H7NerF
+xKaCcMujdVZ0lTj4uRmukQYFqVQROMCyZcs2WhuwubxAG+uB5lqZeclr74HtSoW
hZooRhH71RsocghrliUlLKXZ2zwJOx5h3+dFpHwseN8Ecv3nPqea/2JwoBoK1LYb
4UOByjx9ZnsWdZ0zrM2Eh7FepkiUChcdYkncytIAGEXowA1aH85X5gSI08aHr6Xn
Bk8OBFg9vC4NlazWQjqCpqP/KE5cUWGSk/nMozmOVal6njmoR9UMA1DkY0BeLPVS
5wOWhcl1CjqyqvNiVHSvSnFAWpZmNVYKkjmFWvcnb+Dung6kf7DvrsqYzeHgjXnc
WYTY70Or/kED9hXcbBxMaBJAJ2a7K49V9bcB1SDHAzjzngMVih4d5yPzDIm2/0au
O/i/vcN4nxEImWcKSCtB42lfA5znRc22hYdKNbe/iOPDuxcwmknbcnkcP/XGRKTy
mWFm4M56Kx4EvQSpX/lAmQFN2jEs7ogk+a4QYoOuCPJEGW60IoJQhh4CVal2nDU/
2jo62z6xTX1+4lEmX2q0ayMEqPDYcg46eV8BiEHvjTQt692MoxTRvM0xkJkSb7OQ
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pBsqC8RVwJHrH86kcUcvKGDBzEnHX8gKEjJ4Ra5arV3tL+VALuA1BDzFFR5SQ+L6
lWwopW1N60I/tTUKbaxuIRmDiWYc07kj4X0yhCK+H/sqZrNHv7yHIjv+CdkDPrNO
zNTR1d3ZsTcOl7fIXnhzI6q4fexMXQPndp2dhnYol+4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21920)
5K1MmHyFClSJtQFx9s3x7eGkvz5RWFRfG1RY2croTl+3q4qzxhPApnXAT7mC0Qzg
vWsIGER1vXvfe0lE1gBvUZIt223qDIAVyeUhchk6Vx58U15ewzabeijyLm9rvAyo
q/vz6lWX50DJP2C7r+WqmdrJp35FnoOUOd508SgJD2QQsMv27NveDOZK6ThrrtXv
aejfW/xPodtOFg6n1u9ccv5JWCahazhuWl+9RLFE+ZvXJ6lD7k8CT+cF3+k1JQjf
e3b4F6bmrfyyRriYQeI9o3FpSFqIC/MED4jOFb5rjA0CR0ayChpiKwKZlNRHFy3b
EvBAmkN8qBFv0dIn8CVhcZPwzh+Knahek9NY2DMGK/aMu3/OrnijiDe3qEmGtRLa
+qW3Vtp5ab/ow3dMfZmONlNIT8YrjGY0Hacp+3WONPtWwrAy+NxqRalwDUurHaMk
O+UarnoaxgJSzYKDGPPWLomqBjA/G4N6K195yWkesA5C9KOG+WKGZVkQzp8vSFRg
Xw46Zb3DeFSWQT5lm2hm0KJSWOCgGQcZKway01L6TESxvzpH3i7sVxvaQqm9F0sG
vo8TiUkj3ZtieVkqpEE1ZNZITmuUldxSSXp2iMZkaDSw2gaCVoitgoCHElFbOIGk
BFRX76+I+2eUjQvHMtJ7+tONtwbtw0brLiczV+Dnqny9ivha9+qhLdcvoFaTOI5q
1dqzfxx+M7CRnFXOsuKYeWhbhRROtDZqKhKa4LUOJT5vOVQDEq55CcBo8f7eFQOu
O2FAjBekKVgmNQE9ZMCfzGn3pYK9Lptubu+8xlK+JM4fcllICaMjsMF+gTwvHlR8
zY2Sj33l7rwPWVF0HYghXqogGeZOAlNqcsqO2yET9zzPcdWBHswwKKb9B1VtcsKm
xesZhbtds8dg7lLc034T8jqDM5dAJ9O+azM8X99tbOxjzuOyWXHQ0hIsWLYtO3A3
redUbyGxqYmrIBmXP7yRvtl+SabncTjwW3ih2F66OAg0ny0eU0h6dj6h6JExeKLU
aZ0eb+HuFWa7vw4i8wQshOKMxLaW1jJR9E84y0Tu6SPVyNia4CHAkYJw5pliixej
GWEukmdYXZGL4KJ8sFODVN9yY1heCa8+1rXDhgKNtQcf5vmCQ1kV4Nr/EmG9v820
SFMMR4pqkuGkpAZW30laUgfUZpGVNXb0+48TiqdyINcY645KE80yBOnCGPyFYKSv
lMD7ByxTbIeOtGWYT7DwXiuwUITRA7sJFFwRaNE9Ut9B1WBji/vCG8vRhjvOEDaY
SbyuUI+9wqTZB8ylzyZDWLhSIUr5buOG8dBLKkE3Zp3EJ2CBF6Y3FH2AbvGBwMB2
sKrUBM5aPFI4OSgIIeeKmlXfpcWubBOSOWDlE1hPK1vQ28jgvNLi/OoJhhYAOdtv
sj0h+HxPuZ7u9r4Lt9EVmP9VSLg/SIoQZUoBoLuuHEB8dtnake20Elj6DMoGxqWn
5o2KWsMBMOzeS08NM99eEwZCCiEb6zinnHXa2zo6oHh2OVCYPo48gFtGExtu70p8
Y/2riJQhOChwECgR7e9FOaGyeFprlJmDIkAR+muHtmcR+wooV2bZ4zGQacRgvDIC
EQLECdQbsHgtBn8eZ39+x26wY00Lg+QrcOpaq6W+sbnmxUAgZi7IvfdRPBMTOdSE
0oOjivhlKRG2/lx+Uy6MwiWm+OjVURcJ3MfPU4pcET7AC6rHQDiwZ8OHJsLVi0xM
8WOvUyOuCnHl/DfVKauSOvQmlogFJIDayxOGM3cKkWr2w6zEAn6F41Ep6KHfnOVC
U0IFY4rlKhrO4zQ9EI5ei8X6mEKA9r6DUywMWYFEG9wR/9bLwx4TEEPXyOHScoGa
euRQYy4BW5xuEZpa8uXv4IucmELyOSyE8iw4fUDHW4LQXzfeMalxdsDtT3mheIHC
5l+FkIpL3satldmCDE5mYvRDGlDOWWbOhOYQeJ5sQyNRKOsrqYZj5GXnSUXdYE7l
eWBknQnkpQRZJKNGUXLcPA24FBDakQKsUQ5/edM6I5XaKSG3bqett+Zl5wIXwnOI
n5laMYWq/EXmCxnrMfTHSnnuBHTD+nmEDcHHT6BZ3DGLLtgnGV89nw/YXlKmlAj3
5Jmc155jUkejCTezhdGSLqPoLXlWKoQFzzlrjvojbAsS721q6Z4ifjB2Rbt11X1j
enBlDeJ1jym06DVRLlJd48XQFxd7PfJAoai7C/x/bamctYo6OV15FOTkMUDejBCM
yCyRSjhfYD8QTgFrpDyFtFuiUR3z5q1b0NOEJsHRyU3NVIAf5oCrl3O+fT0BfOaN
eFEdxKEUb4QuwfGdoUZxZA/cy25AbdNkBzMoadMEgl5AKIhvO6U+nH7RHChz4AXe
fiKAV/i6VRtipWJuSGSFTNLKQAQEOxF9P6x6LVEIA7gatjmk6Zf1kRbYC4ejTTA3
1/XaP7tGXUKiWednQG985PeQcnuIrDY+bFWqIJnENkfHdyQmjYjaaG37ZgW2P0vQ
be1TljLxv6MsxMv9guEq1HV/9gZJzG7KcB+/8zr+I+RSi00u9FX09/MxVbL5Cg3y
HNMpP85YwC+Cl0CXdfFIjC3yiMoR0G8t6VAe7Dcak/11phBU2QSgvzSJtLiPhEJY
WBmY/3LBhZZMgA2LV+6O4jokR8XDt57/91nlTfdVmhv35UBliBb0fP9tuX6XQj6u
KPQVjLwZhqazLei9ir5crbvsdBoC+vcy9oSB2W5B314A7gcq9bvI7sst/GTSbFOH
cO4PbomX11ts8+Pi1OPzAhMmnuLAWhS4vD1UC/kVpsdwF6ohvwGL90hrnpDjf4Ns
62eiMl7hKiD8+he018IuioHjbknha6Pyper9y5LqWVzZD/EFlSo2i/yUwdiyC5kP
NZOy72Q7LlzBa+VtwHjsP9bllPyErtrP1fjgy2fFrsHnBiidaYMTQUc8m/mipuj1
UD8PiSyCZRuNQfcDI5cvOML944ow7+sCq3lko+m43PEgRppnsq0mWdmAF0fKXPX3
87biXhlEjTgW30qpJ8IICo3EXYLwTf84C9kR4HfP4pKeFNhFcFuo4pXiIkomp6S0
Tn3VXOpItXL+ytVyt2u4ri7Pj93SnA1s7XCIPhjQVgQXt7UY269UZw06MQcO/zjW
v34A0RHrqUYu+t0D4wVrgogBtyaccPiIlh/RauYw10HQc/w60OuZX28ab4PCaKOu
VepbLrhkpFuWdXL7WKjpPUUpnH/JiRCUi1ODEeRWgVXGa8OVAn6ge5AqPrD+zWzR
G4qUKD9+hACnMkcS/G5/xuvJUbC0saPL+PCxdfWhNUY90utK2o1cHvLNzAKb6rMR
jJtFZ2vIdWMCKDXf6+BDPOq/0GTi0/zsLngvo+MnmGhYFWDsd/9gOqHrjkH28TW7
Lt9hjD+z9V5GZRejLaBDzM1pMXsE6atx9wyNHr6aU/v9WLA/ZwjKytodrahXC7ZF
gk9/+aQsbeeB8uInFRyHeUM79V7kZXIpXX7lMAodQK9/tKxJO2Nja2h3Y2WQqxxn
QaUE+N68GnMhiN0oc6xoXl8AjXz9eL0NYALh3vRCaQz1bm2+vbm5iZtzX2+FamLp
v4W2TWaRuLVFn2ATEVuIOLesqWxG1yw4l9UonQ9xJMv2dO+UMTKkQXNOiry8U+OX
eLIT+v9Fs9+Mp7tvV8WqOxXr8vsVg6gxWKNkI963drjrnYj1nCT7QpT15nHwmT3+
3+xi8lebNWhC8d8iVC1YEUWCU/LzTR6I5OeqMLzl1PI0vKdo9pJQxtYjCtcBW3Jv
FzcAHe5TOzyvfPhvVVvSzOcuyEK2YD9rl2Ub8jdxhh6JSkvI21iGUVCJ5phld8C9
Jp9aXCUBhA51JqVHntVnekbnkXQBSGaVXKS6m14Rt5paNnGha7BJ8h4vyYljLIkC
DmeLiO+qQLMaWOGwqSAqW/pDm0bhyMdyo4zPVKPhfO1y5vcNvQMuLWBQ7fmgJTl+
R64xyYb/NLEaJvnCYje/XNxwqYmab+YzH7KFjDZJ5ku4a9gVzwXi2a5Z/kp00gNA
2WELoT2FPYV819JO9/q1SGcSHqw421+0iotYqdA3Y94ULT6QB6B7ctaKjB6XUOwb
HDcitDe0sq/iQM5qIH1Yx2xhc6Lg7IaEN1qO4qLLkS2gwNNk9PT0rEA0Y1aiN6o5
LZ2anhfVYxhJiWGaecJvN2zjQm88rf+Z3/FNPslCiePR9duTpmPc2NvAvG0bXIAe
krt2KlC5oYrIK9UDR3FsY3RWzmAfYU3MhZ+xkbAbZ14MM9B/WxVSBvN/ghrwDJvV
xVfYsI+OCOPGQwL0eycWCLFELbtuDPh+G2KUEBcCbLQzjjSzpDl5g0VzCWUO92VZ
DJ9gUvjZr7teQglFHt5aOV4ZmCZU7W6E/65DTgRguBSwbau5SbuvcCrPDhEQjA7/
YpZGIV9lIbKNhjp9R9Qa8P/Rr8b44lt4EmLrSd78sYzxVsplBTMDnEGwgn4h6vRJ
nyjoANeatCC4Np9f368hT2inKi7vOYb5CzoaE2g0SD+/F3tRcCRHhO4nO2S0x3po
okh5ykgEFyTNjcGdKfZBTrepQazhPxk43wPKlYYocmwjJR7Wn+ZDw/1nMSTeM/es
vjheABEbSbNKELtLF6NzG5VF2VVH0qR1ETkrk7UXIKPRRHr0QoKLgcDzl2YO5slM
xP2FpuoygPPS6vT1iR3/Njhxr3FVYUZ8DLiPGgxTQZFfczxihz3ZiyZJX0If7HQD
39TKiDYa0SLOw4teQCeaaWsSUSjc3cJOaZ8RS6kHMiZMlAqukXfoCndvo59tX60+
9NX2W3tkw1OILokDGbozEF2y0c9MHrwaM7eYboShiU3DQcYSeSdjs2QdO9lV4xQe
AoBZJPVUi4dAdSHHloTN4hL4CwQ39/+qnX0jMnFUZlT7UzV/MBOFjHBPpCq43zb8
RkiF87VBE3N1gtJ3909SZ9agVFHWXqqpvnbll6ImmgIdOW01SfiD2crcnCPDU9/3
hOsW8xjCSi90H4maVYyAp4/DHANHUFBjtgiIDNXDZHRy4+pW/MCHErTCRLEbS1kQ
O086a9+KIgpFktcrguoHiQ0e9pC5HmIIZuoSSwh7A5rX7/stj2l40BSbZmNjalIH
Rv775cVregc50G4glULjvmEdivvNB0pGN23hGJ6jY09CTH1pI60WIcCQnXWzUA1f
2/0Dp4+ikzCNqoX9QlsskVju1KzrX4TqXWin/W64vHiLyVWas9JNXUv2amzGehVc
vDdtWD2wkamkMALIwxPJ1o62UYAFAVFc7elTj6amv2a2acZoVcQ9KYxAXIAa6k/x
r+xALtJ7/uw2J8ZgOoJCH2Nju+018TCR+wE4iDe+jSBG522rekIjhHXyrVh9Q6Rt
f5cIy84B216lrCs9mark01EFLIoAteDHVxMn5Z3Q76H9jrmbLbJdwtG7d1t7lkPg
ofAbq7YqXzICfFct6EZz05kgbx0RckM+mGTphpEBnPvsR3+TBL3EdN/pQgX3R3DG
xLLkA+ltVBubGsVWTwh9cIpFIb1/77a/qt6f4N47mz2q8IMFCHWktKE7gHJpnpFg
a+if39EvDsFlr4tccwZ2bpsi/hksGVOVeh5hPh5CbBiS+4pBuE1aOdoALjaVrSjh
bEJg8l/hdoytiB62Fkn44wmu/P0Z29OOHnQbcWt4ER9cJfoWDZQiVFCphlQdu48g
HfuHnrYtd9a7zNqpmzjCS8Y6nhJ+nzg8ZeYCWs/5ZM4J6eB6LSSb06Vj2aq3y8t0
/jrSybYr4Q7y9T7en5HJnGILox8nTRjPOGvdVQDiStImPSekjzY7cV/xUlH2TdLO
0HdlDvn3uzI7TK2B9myqWBUK6enFORYcC7zA5U+GLety9nekJqWN5N51eiWwxPbK
JJl8aTzXGXgSM7JLtcZlvbRYXZBEPvLtzc/XoL4U/fsYzNOsz2/0Ce+7DMzRocyr
clQZQ3sOk3Hdmw8rn6baStgoL+8TR5u9rNIavFE9n/Fl7fRCT25qk+xgh8VoPYRR
BOiCicKuiks3FCtN5Duib/YjprnpMirr3xrEnfGfSverwKXvPRjxWxYnlaaHyZkP
Pduf/yaC+yZ7pQ1Xx/wZv50iMFbcQrT71sW2TzO049nSPUPUZX+GRugPnTGfSaVH
oLyjBVML9fDkQau3VFeApogteVd2K0pilgA7CHdcoey0t4lTsWScyBDBROU1ZBU3
S06u2OIU2noUPlY5P+hCFVPYfc2iVhYyKIc2iIQQCfz4gMJMREgMYKnO/7AxOSM0
8EcHCAy/050b4QL558A01M2nlWaD2IVh2YHMhQ1vfCxF37xQtJgg7mjEIGkZpsGA
Eig4yAd49L0pjpabffMaO329fZh868SG74N7fWj7Esvyk0rl0rvp10NMMd/IA+l4
Gcmyna/SLFJyImOiT1fWvfbdaHKsaqnOLlaeFjPaeo3tGMkLUketp0moKuk1wPRv
Et2LI27unUCTz2KhmflnHFDTHjOiL8DN0vCuQXNKwVcaYuXtjlkF6zI9JjGfh7bE
5m119M+X/HqOl5LTMVRs6gDT68vJ5b8asp2QQA2FWdSzwu9Rr/lAtBvl/PTqkzvU
RURapBC9XB8mPhRYc/upiy58v2buAf/z44IKBgwhQEl17zF8AduDl8lZayWyERmZ
/HJjBUF2mq3hcIlsiwtO92JQo9KPIS0/8JiVcF0Hh3rs32uRT2fOL1D2IjK7tdDL
xzuh0Q5P7PhRzZE2fGa2QuFuqWz7xrleii7V+6AhDXpQj1BQvmeSZbYnJItQzgmI
UY8rzbd7+IdF1DR8LLa5ahJKf9gpF0JONhOjobknL4LEZ5Qi7o3bKkEsYmnRKorD
ScW3APqfcZ+OJx9eJyW/mHXF8k5ETh9ajqYwL9dqwff85f5ukZizBxNXF77eIWR1
Y19fylJ6+Iw8OtXJLn38qOrpW4L4SKS42AYl2hYQDRYFwoENpSlWsD8GglOAPx5i
jZqG/uC7NUhtwlosUeFzWZGsqd9dyL6zSoyTEb65nSmWBCcyal79egs4CfZhwWWd
95DPxBht06tOz+GsWfe8IV41ww7cpwwLXeTI5Az608q+v/plhKbpRGPqPtlLJPnt
kG5UvaZJbAntvyI+5lFhMXetJHnSNUsBqsBKfCyLUjGPw1n+pvRmm9iWn3piDc9O
TgzNdnrS0lII+EGcrRp7G2uUkF2Tg0tco+pgzSEtQflcGAf9kclct6DPCaOgzlVP
FPsT2N0K24Xi43yd8XKCFGz6B3F+knINnpZ/lR8erKE6tJ+ocHeWMwTzTLBJU1X5
/tEhFreud4nzXKtJye7Ju08nbKu5Y5PdEVu6ErqIH5NOdMPh+crdKlR5csWv5xbT
VCuwPBLz3YRJtKxTNSVHzBSbMnhpi+gI+OzFZCzbq2OQiMFhnUPU9fQAaPzTBo02
C+6KB5ADOQKcVkG+2TPYQFUMLpSenpowxbzbLMt2N1FLj9NW0QYJaZOq9yuN9fdg
QFbbYR5N151t5e/1TV1sA4CgJAUOVdzun11OlSjk85jc2e7ZMHx3fWi9S2cUVxrj
2vJfg0K+64SMVCtnls1WNuZt39znLCmhczwJFmXrH+TL3ERmsjBqx6ZNPTbrP64y
nVARQ3JhhiZbAtSNUlfS5B6r/1fbnEtQOOW3Y3jl8KVrYgCIBpn3zpztNtvAsIWI
pNGl/Ft8AC7zc/xsDgkurfpxdXXEVff8i3M1JGwmckrERCcw2o/ZszYPDHq/Fx+m
5vE3IEUCKCv9TrmebtJ/Jd4gIO0g19teLKMD8JpBtAsBxW2LShYCmFCzOK5cfPW2
+m0xpz+rCTLRPB59hNAJlA+i5rD5fT5nnnskn9z4O/8Q+WQpbydjNcHWwaeHuUgy
s9UXiYV4V0O8J+SiXX+4cCl6Cm+S/O9cpjX9jeoE+lq05oUma34JAb2KUMxW5kyI
uFKVnWkMJ6DitSrA+o8Tzo4OOvgvkQj+FtQmzqM837eLt6A+G0QO/axXBmpIq4tk
xxOEFenbRMPLwe7c/Z3MMXtQ14FDUAagXmFnOAQvSSTdLox0YdR2/K7eWjiotIyx
4ZpBm88jKQlwP8uraUuvPHpvXwXDJ6WR+NvKQnxBtTYos4bypMHrB9GBWumBytrF
hTbxYy2icuQb8I99a5YTKHe4GFKBPGDzZWQmjGa+PXD6LmQWlY4q3+AFnUGdX3zR
8+AtQtPzuNhIKbwji3yHO3h3cXh9HhLDTImMwm6hCFUdfpebfEko6dsKTIU/w+mY
veuomLDExJA+vkTBVKOROMEfxlnbdbxKQWPsG6DQMG/jMdKF74eRUeQb1Ulp1RO1
LcBYeTkdXk7JC8FWhv/rcFO0EPJt06Ps3c9Ok22929DqYMaRXpwcQ3FN/UjvrqAm
XDdwEce1I4EawBjSPdvaFYpk/8A4EyYPkfhsdIipVJqgzMbTJXc+8wymbPdZUuuC
sIHoYLoOvSk8UBPRnWhMPymi6y/tyYzrMIVebY7WuVa68+p92/xLGqOHanyKth/N
EIxws5XpxZ4ax++G0Wpc7LXO4x9u5eg6yRwliiQRAlpFPF1MmXq8xRqIiEuaEdij
rm4Ao6yZe64i9R+cLb423ZX3wFLQCPN68//qHX4XBjCvbPNb5B4G3IPapZv1x197
GYFb+mLUVr0lHWz1YKFFcPnQO731bWhxXE+K0GqhhuVnPqqxIJhqNCAR3Vbv5Qxm
mvFSRyHhs6Cm8G+GCMZ9JRJSUmQKg5J0fNwpNPPxFEaCxSxHXQeaWLLQvoKEOdoi
EDe8cm0H/emIqwJqCbb43Nv5U4qv2I4jl/UQATYTRv3gZDvMFnoaKkm5AJsj6zmq
J4IV4/eWwPxZNqUHE5TbhH306JhLy8g0SAdgDvzaJ/eBX/01OX3PeniL31SGYgm3
+OfYP3upZbi9azBWG0mTrPKAeqE60jdjUxh2CTvyoV86p5d3kwTry4zesNRe1yQa
azsHdPUhWQcuIMC4jNH7Hfi+F7fC4ZYxN08Lz6cvRE3aB9NIMCWSBcbqi3I3Y1us
nxV04LEI9BwicHpXKXTOiy6mf+0ZI3AE5YLOglfWEgWwkP0TCFBo57yg37Yc971Q
d5W7UMo+TH4xGj1sz/XEzul/jpYOofHajxkb+MmezVl1LZGD8DApQEWX5fsftIkR
N5/Hu5SHo2XKayaPU5ztdYOG+peuCrG25Mj9ZzIOq3yNFGkS9G7W4PSQJMZEZ+nt
aAi2rLKBCZWxUScKgh5aDXpyVQpdUhkJaw+gRkRKQbHdeOQ8aEPxWh7ohmjYNNEc
d4kZuCYMT1/RcwO9c1LlA4a9ZRbce0lB7TRxI/l3VKMIB55VPZgX5EKp+DxVH5yY
6lsALZtjXvnLcwJAYGCaP3S9vGQOqRyiPOLKRKwFTDHCZ2IjU+Jhi2v8hZmPCkG0
kdkgX7X4Alm7gI0goCkPoVoUWeoLTB8eJWgBRw8z/7iv8qD6CiBG6BnGsPvFhuVL
Kvrp5G9Tt1q2v342wEwkJjH0z/L5IzzLK/MvmGjtYEfFVMxH3+l4kK70zaNcqh/I
TXSLVaMbHjvyVW7MaaYw3Oy3MPUP0ykybhBQAgFLCOrLm3dB0MAjL8LkTkl+zAm3
+mPZ2TqH2UM9mWnx51btUr3Y8ESs6V/4lNylf7H795iiRBzpkol4ET6Dw+e7GSSQ
pnk2Gj7Ijxz/tBM/6a//XyEiQ6cxAFQzVAErPnQItTtfBYe44ctQs3j7K+yduSaY
hMlArOEeVMTx4S8fKx+PltNAUs5oc6UmA3MCbWB2I0WTjeMBGcpHQM009NWJSA2M
S4YQueQ4HWFxVZXVthwUDXviAytZ32TxVLxJEuM0Ros6gNsaG7eCTMAnu6nY4mKN
0y6jkqWOlqYpX+9NDGlRu9nbWlPFXJT3znU445ri5q6p6Td8r03zVUCjD3YtzFfP
EKRMaBwa81wMhaEdCIqN+yWrkAZ2L7rKildluRVLei6mhD3Nsxa09s8+bbAJV9iJ
RkqfIUThN3fiRTznN1ic79zkmzY6GDkW5+Jexgp9C1DLpAyOypuBqMRae8h/K2Lg
YDqyS3naIlUV6+ohrqwxNHuDu38JtC9HgQAMK5ocbS6uPYhR6aGw5P21EJITkFHU
UHd7GlgrWhZAH5wyPSXC2lvAY4BAOlDQO2jNCob9Jahv22K+bg4DX0qScCMe4IC1
1cDCbUt4gy/zMobM0sBD46zEbQKFuupk3SwJmTIA0tII9pY3+2jgdXfNDBwcaW0m
36Ds++bVzmbhYodZ6X4HgfCtg14pCnCqJwURjP+eMrMgbruQ0kK/4yXg44+y8Fr+
jk8R+pszaTk4FoD8EhIAV4v7owucKFwTlQQHxsUZ6hUnMxMqBNAVhkSwR4W68k5L
I3FTL7oaFINQ41QUmaHSxdMh+4CHyKH3hisqcZqgcDr1pqouHUug1nrKBvd82Fyb
yfWG4lzp6msR1b88pdfgeaN5Rvr1l19Y2Ry5u6fOjM6Dg2PvtnVm+fUeXHasjecY
vp4LovQ2rBvfZaFnUGPj6VY2KgA2qk2wKZ4e/s0JJxATzz1Tcqf2O5fKSxCxcSed
n8XzxuYdcmrZ8AWGJGr8EkMvxUK6JxAvrR8EdnjO3Vp/BIR7TkCj6cB0mYbHIGC4
OkGdY0Gd8hfiT7O3NhoXz6seI5NkYSafWd6bMv+MIES5R1ObNq3iGpat+1+CDRA2
IZCZy2LdDoafAJ9UKxTOMQWSpm6WONOrPFddwFC5WWEKcDhxZ/ui4hV8WUy9Ank0
fyZwNt0euDhEQEzqna2jlifY+/GUVq0O82CEQWcmKSPmq8Al5ohHtnarFaaOyVP9
u47Xh1MTNLQnAb5JrXgO9KEy4p9GPmYissZw3jKyCsfdkpaTokLWR4qBB7LIt0ux
aRJteq86fVvxkgM50jduLAS355/deistZuKYIx02f47/0S7yjrxd5gK4PQ82gpFE
o+Q58oNXw5+4jPA2nHLBk1TGmBZrBnHNDnd+u2mbQJ/0E/AuZe5ejtcckzfCiOwt
QMVrdmZH/8oZy4QsBT6gTxTZm12bHihQ3+PbmD6rfvBKWSvMmuTMv9A+3lSw8FWV
PTinr9UJsvSeFs5uwpCtObSA/gnEPY2GVCWICKp+usp9ZRqx61iHTvA1xo5BmCly
dH7nUoZL40T7WzA/0ZYHorikaZi4J+qSEgQ1TUrdl76VJy8qIFCEDf2J+Px8kBrh
UpwygpWgJFjzQjS4g40m/LC+JUy5BdimJoUcIDXwXughDLHCXt3fPeDWXlWj7PFB
z0PA2ler8xagY0+IVUVXPiQkT0hqK5sklcuxa529HEHJ3Knnbc/3ZnCHnpWyguh5
QMlAtrlLFt80ZmoCv7kUaOOHeKB5kgTfMv97q82Rh61fAfByYHwuROMjU98OJck6
+kRg8H1+mJdFzVESyxrDTUyZ3Qw+L7TQXb2KynxGNBmDEwnuMbF0LADDqyImVeNu
CAOmuwBQ+vHd9X8esiKfbNbbWSmHsrFF9a1/YGXPqHxhLa29nB2Cf8wX8/wUuUOh
oOgtvninORZmxKsbDot9J3t+7ksfrGkRAC8CLjV/Pa9oyC0o+f8LLM9DMiT0Nfii
trdI7YRQK4nT6eICbLAWP8OSN9jJs/m+aJit57hIHiFHIEjN0jh2lAfHfwPJT11W
AdHiyBJfyPJJhJlr0REz/g35cN4nuWTdXJbC3+OFWKg+r3qNdy5px1KbQ/Zmn18m
hhn6D6yXPJjZ3TnfeEIMqdsFOgR49WlNG29elWWVKcBCcyWFKDRfA4RjJhlEjKZK
PNkUWsMdXUTp6mwHSrPGAaM69qGUGRZfxpFnM4V0WfOtBPbmzLXHEAvW3e/sDV2S
06fLCcWvtKbEWJ0B8TDiAtS6vcHmHvOjFrD8rs0UiRxDddQ27y8EPHWKpYVSOWaP
eUgfpORILzAmPjeccdKHqXcuUuJQfjpm44FRcJPjp1cENB9RVhjyJCR6fYNyXtfR
VEy08+Y0+dprXlyHjRgyt6v0JQ0olDOnOXAD4jpFXBNnyC0uDjdq4wuWSVtwHeGb
ylskQuydrIsuizx0Cn4BDgG+YSzkmk//waotmsdStw8lzBfLtfRYDuySQ0DxwBEW
IWOvWvUSthwx8+8nsklPgupZiUJ+yh3dYf7K+oW1eQFyvEbmtf2eaVgoTx4GLpZ4
bwLf7KAgeINSo0Fqc34DXhZXQlKkTN1r3mT898NvjbaPUlxD5Ei0O6tfeL1iQPfV
panqNSTi2kOAWylSBGMymhgXhSs3X8oivDODQsAvhTMQuJIH4kNF7a6hwJbZBTKD
54v2RqtHGSJBkrFI9OXVmc+UbzKKlhYNLcSm3Xh7/bbBrXX0/e5qaGdt12hr5QxX
zhbdTz30q/+L9nJDblwIt4cuDRJjvhLCns0zfWFcmqHZfuFTKdOnKD71ydLBCTMS
Zok2LWJBDB0IGUJozTupLtyiW+XqkoWdZTT4NUZBeBY5sRcPwqgLnLqiNga8A14p
/2YHKqq14w7gIOCwaiilKTZp5khVsHoWLKHcd2xHXU3uPKAgPjzo0vecbSJbZUCt
RrQeKi7KmFe3jwzfE8f8EOXcnwcdxgDlTWbMb9TygDIRr7YwszTKAbo4azHO17SV
s97+ULTwMVbKn1Fm0574FFbhDilN4M9k3C/fawF5LnlSTyjBhbNyuBaefubZ5m6Z
u98pkDTjKE2o7QoSuBoJL9P7fi7Zmmz4VpdLdyPXiUONwz6p8RU60g19oL7ImMDY
bF/zgY7ItecKiVQerx3J3xAOf2oCfwYJYDBirDvXK3R6PHXqymNVqGpoIguaSxzn
r/qv8BR5+cbsp2UCJ0WHUqWD1WAOywmltyPpVpV4I9IX4S8ZMkgsPgkaJ2QjYQ48
f/oOfxZJlPX4dNG9vL30mibhp7I4fVmzL1nnRomjnf2MTmwuwOt9HU7FmLS2m4tY
kNIOLv5AdniLxXz0g7MKkdg8MQhpETF99cP7UWsnJRC7ozB74osHxzpqJ8ucAk5L
PBMOXmASLSPljNwtLuDujQXsgvulpPeokGjQ3Vjt2MkXXlVQYud1uWRCsp+/kmNj
REuDr065yEPVaMLNcUNY6elwAkixrc/VguiRgw4A9DafwBKROplDlneBY9CoNYQi
zpcYRXBXEKSjvNEj9M5gC2p2hY37990OvWYb0s7SdRH09ZmzCe7+NAXX0Gv1S7vp
fgYvrTjmnRy9HTFKvJEk2k71tzh1s8bJG0sDaIEMDiFkOzaRAFme1I8OMAvF6JPs
aeyNKiIt4VscXMrsVNn+/BkUrzfOqXqZHZ9mLbSU3AryRhU7CFqmK5rQzske3LXK
qEZvyCaItpp3GQFJf5VE7HkLi5sOjYk0ggTU8xIcKyom9jOpXLFRzrsLuZxRyZJZ
3l4QfNXRq3IkzzFeTt2XW8KmHrX8+dogm9pQXnaM/5zvkIDAx/5nllSlyJ0gPlm5
Pm4aWyOe4vydmuxbRRQpw5vL8o8JNZaQfcjNzgDkSlgVdDXAw+E2QjbjTqyiPJEG
Wo+AHSvGa84/rDC9oD54shNCmTi0VtL45dl5cQYCyZUM5yhk2e/GM3NDXjOOSQM1
bRcb1jOwqw2xgvPLgR/TXlY4Nbz6BJLWKHMaFdx90U654ZWW2s4E9Xx+KrAEYz4I
VwnAdc01qa/QAC2KZ3ZdF7UfPmwz/IyZyvufSOPeKeLdyGUIaebO8WS4YgZMrT0G
DGXqaYDgwZGot4ERfWEdstqQR3/6ZDOtOyBF5LwqftP68SJ9LwkhPgOTKu99cInd
0VQJUFui2LwOe+HrAfcsOWNSxjTSJXQHtdSk+vx1Vlwn6uzeHACOBAolVbO0pN14
E3kZ2tCpKUt3dakFC9cUWOo7RHm3+B+aKIaj0apaIQMh2sZlGmvSK8E7ZqnK9xgO
A/UEFDqvvgVThCZCSOXIuzRnxmSCJhnXGA3X//NfnYQbtfkO+D3Y1zDpqTtbgn9C
CzTF0AbbEI3qvOocF1n/6/LNet4czj/2Ml6SMKeavSjfVhwItXQOGPG+l90u2SaM
zn9QCcHaJagO7p2gbYwRMqiTbyQkMJ9vNxq0eBn8dD8IJ+YULemm3Y1aVkkimB+S
8M6Tcb456o9S0uooOTEf1IrVh5aM54CIeq5S+UlkApnFMNCKpJMgI7ZQfHnxrAdW
nSEni2kmalPe6QtG3Yr3ZR/P/zIGzPGGyhwJbmXW/4kFHWiOt4PkWEMPwk2F8GAd
uA9f40G8U4DJrdh4KiajFP5Aon/XPSi0YWZ63Nu13joqoj40Q8nrTiHgkhQ7zuZI
zU9aYcOKYFvXT/abl1Z/cviDK7hTph7XjTDlO6OaubnTARBcdnANjTDm2Xx8cryT
6hNQB5aOj7eM3loWFBCsDkmfIdR6xmA47LHx5dGu2/VTgCujmxUANRw1D/G7HL2t
V7o5/F7XynBZLXBQkiFTRVBRG/kCb1CEHgSK0EEt/gvfX4XED8RgCtaJX4zjjcbW
SPpQSeqSj0plzdkeUdcjAa8u2kVPcqIxGVAnOuUPwVuqxqmW8mBYB4Q9JK167mhh
L69Ap9iCE1qUFFeRriVPZs2IctZsVkZYB1CUwk9Ln/Cm12Rax6t3YY/L2wh4xICz
6xIYE8xhW4vJXAujNmgxd36Wm6DtibrmjrxK4XFAo/33uUBAKRM7NYEgIaU4LeLS
hlwodG7qM7EhVf1veZaQ9VvkZPj0EUkNBW1U3qcgXFNSsoVBLh9640/DM3RZBFDQ
AkHzGNw1QtihfdiR81Kxtfa5n4QWO20x7t2VnL/6klApcg8WlXUnipPNHSCTn2rq
AMCp8/NNkXWscdldM5Kb97QWrO3nBJMH9v2nS7G32qasmoAeF18yOKLBmvEmwQeU
Djji9hFqgqOXrdCx52R01agkcufYD20cG8qRpGxeEsPPshFJjnMOVxnkd+KnhXS4
XBcbC8q/eRb+lxhtk/xO9MCoJMSlLejRbqi5l8BiKezr4vaUIdxIIBTmeZUHOJ2z
Sg8sstbUi35J0SEFGlZzxgOLOEhVr6yr4yLEIp3zRmd9H8WDy6UehNrPg4pDq3n9
9WfhsgBlYczLJMygWcVbTq5nms9V6dXetK28F5mPmXRC9JhN2XBSRiqFC6TCCCAK
po0D8BJjdT6iegaKWn7OqtbNoenqJrEMSbtW2S+WQpoZCO61Y4bPEGV1t5hZBkyV
3g4JkbcYTGWDcP2uLLchc9EvxPCYEeK5gUjAZo9BvdyiSa2hyEuFa+uHsbvXm04C
erFRzMscJS8nDyUazwqhMVyGGItqPqpTjJ9dXA4ivOeMiAa/nPVaImseXYNXGBQ/
v8WyzMdj/fLLGDh1QX3JuzM9p8KSyq5QHCa1iJyAbmSSBvO7zNLekkW1dh4JvGUp
kT2K6Uj+GsN52U4MIe9/SIGNIpxEL+zb/tjZIi0rGc/FoFpMILfYoutjNW+FcYzP
jtYQx8Xr68CM19u6OaLywgWonR18sjFGSwlkd0G5UpsrfevDs0I4jD4vxnIQfEii
boeGGZ2411mgP7CWrMm4pPJF150xeR4Ka+VCBbBPkGiAdNLghxQcQMqA8x/EBYZn
IwluzbrTyuTjWKhsrnFBbQe8vWso5Yp5KwLR7IsjVBbSJx4CMwnEaS5XwvxHim+8
EqIP/MEhH85JAPepu1DiW0GD4iRzRoMV4gOqfL2svjppLJs410ykaUsoxAp+rrS4
q57ysB8I5HYM3UuneVD1T7TMIAxKonQr/Xx3vSTSHOOexTmxeGiR4ctf76VPjJ7k
aAPiv8JkelkbnxQtekYoJOQtkVioKlHvo4kwVe1Gi04/rH5etj/IDny/StbIUk7h
b4s0XLC56b9TAMhRAdK27kymXiTUzgdXHxDRc/sqBAJPpb4JJ9beWe0x1zBCzWJE
bVXKEHPLJ8UaDTwIbd3SFBVLqF5Netg6e/fQdY+awwP09pj9MmhcvL21yxfZY7mm
f3Xm+M8XJxwx/4QvKiFx1Q68KP4Np8vPZCw3Y5cLsMYbXlxAsf1YBeXCFMRM1Nu/
WTDTQG5/qHauo0tc+yeRQom/puvRPo4KiU30K0sSocqWXm5+bQaA2qBCm2eoV27h
HMI8OVwI/kEKztGwX435++7jXzVncIcp5etVlTRsaNDNK57FS8k/XzguNKzSGC5d
KdwgAYHsaNouejVuNuhNCigSxPoWGcbRHn522uphk1JE544Iz3rKbZTjWChdarmR
5Eywo9hQrGaldRWMFlBKz4i0M0mcP6AKHPEeboKxOt7sIoMOUksoG7/JWg25MPhD
a1bgeQdRWaQNnzMciJOoVRPJSOcsG+T2nFLDLOmI3V/WhN3SJ6FpnLJEZF3zAMPF
mKLhO0UoTG3BrotNVHuoUEmaO5TjwJHArz0hTOMAeSgOKLYA5ByvXLCYALNMKlVi
oVj/8Ey5XeJzShP9D254QgIqshayk7BRp3dQPPFw20X3h9bk1IZjdcekHzKbQ3Kd
EoeMg6NYSMPfFzMs8L6afcHfLHh7WDSSdW3BKsKl9CxovsGReNRuXZDFUyDrWJHV
MZbAU/bSX2V+1isFpnVs9z37i2l5cAbGPSEU0UuO3PBCEdIaX3kyrOJtAAxmFIhM
T1CbLwHN1DvIl3R1RmMg2PI7SXjM4+/MM031uH5hEWc3U7UvGnWBEJnKTzO/p1rh
IX7nZWgmEIZQMQk4W18xt6Xu0nA03CAvQNdxQAVXKvyE6PQ0+Dv3rK1zdt6Uod5L
+ta/RGypLCGhHON9EYdLYsokZrckYNlINOQo7/AvmoSBUJDxmbuIrllRlBWAQCK6
VZQi071RSCOuPOnhh7aQEw3PawTSTLmQ/rLWh/Qas2BC0VdjADpVQ9ddt8CaDuoV
6Pn+RAMb/lSrksiPCxT4YlLKk38ZQZSDL1to+ezQULxCavq/eKHKvITuPAIHit0C
IMsBAgjlIW4TcW+Gy6X7JNtrWTejsGpwbu7/4x4zQDB+KYrKHPWdZA1j5k3AGLRM
ky6gvG6aGxpq57x6xUpu3ecEOQgfx46PN6+qkezyr92wogxjOE9ChpkS/Md7fdMz
D4EktO7YDPF7IFJIdYWobmN6Q/KLm+xUo8jknp29LYW124HCBj6we9S2NA9pDmgi
sv5b9/C3GAtS7u2gyuT26B0ivMPzlMcbeLiWr5ybTSfOsgtWTf9uSbASobioTVMU
1JBWQSHSu8KnjNnVTSmyo3eGwTOO6neGF1QUojV7Jc98JhEGyOcudb2rh7Ipy9S7
2nQ6xuuMTyh/ffxiZfep+PmOEJL+rKJ2QEpVQ5QGQUFFtCTsLXaWbdi0yke5skSf
lQcCh3dIqg1aBm6v2c9Ha3O2s1f7Jf+0NtwNVGFuP1ji/Xz5RatTcPb+ZlUrJE1Q
Mu7MeZgjmmt4zj9JFrEoKuQiScbFKWjiA1dFf+zkN3Kp69W7aMyfKO9Vk6vNx1WG
Jp4vDxQkJuVgRM3SfVQiQeCnMFtp9JIFt/EdNIhQinW0jTGuAzlJD8oB+n0cBlvO
wmdEEc25WNEub6M0FvV7D+p1mST+9Y6yr3/5tOjkX4nsavEm3oM5Td0wWCSF53Bl
JFTcZHsTQsBp9DQJ50U33l1yxuAG2THaI8SanKqgjm2BcZbrKmLacvXr1ViHOozk
fbZev0uUa+N1mDMPJrwsCyRx2D0/fk+KlTL62u67Nvh82wPEgpOf/HfvJGmBLvO8
d8Siu7kLryFrMqXmoY06lnVd3dlXxjytB0yP6SP/UltcSX9hrDwxAj/B7XhuM+Cz
7odZ8jNmDGlij/iaQf4v+2+bR+/NqIk8i61k6Kv6ffFbdpRmPpGT2ljqa7bp5tWA
AKRK3QPwdnHxkTCP9w/1hnUmHeMROjVvFYmoQknxR5fTENHNTDkx1vaJ7+NoWoZy
gdvXsA8Zw+QR66nXGyHUPymLoAD7w3XlaGAWKsG9XDCwY+GZqRpG3Vijr/CVmvs6
2ool6NjfgHIiuKj0vB83ki6KJBjA5LzF9NvvmgQFQ/huJjMOlahEScrEuhn/duRq
cz80NJ7TVtK8TgbbhD9ykv44+2ag/4QJV/bmnfryqzLdqAliGJcCECCk2V9AmwB9
ifm4bcyrTAa6Q58IMXwZbBk0ZR14jlpJm+A0CF04xK/1Qsi5t0VRD2gQ5tkwBKts
VTINLG2JV16PI1+eTbo70N+QYrIiCCEi+WickAdKBZ0uYywpv/rVVxnb3ofzfln3
/I8tDYb77ArNLcRi0FU/Mj1ZMzajUfuVWvfU6OfxAhMDoy9x0zZ91wTAUyGtGK0B
nRJtsdbkKGQmIKfSVgAebLVPYJM3Fy3HxG9Moy/65Ev2mw4xZKw+qsCyRQZL8D8E
7sfeapMzb+YZWOWLK5wQA8ZACHrwXjonS6KuzJ2lP9Bf3sBW7GrbCZ4QWQsz6iyH
nlBCxNnwraeuoN3PVpRSsptmtKccD/QXqhKRqg3iLX4YRHFk6tpaUhsEg2DnnndP
aOCGi/rgzqDHkAtLNZwBJNihNK/Mri1U0XGG2+BYBDEWFn7OzGSc8DRLafeRxoZH
lfUJdcvVTiK8CELGUCQpqiShEoiOjSgBaShpDz9lOXCjP1ka3+Ssdtn1LaUUiFC8
OFvm2+sV4Me7swFevn0A8UpIpIALS1M9jShYzqeIJiP6GT1ReTiApkuvZxm90Sh4
5Q429M9FI2DwD1daWCsyJp+kK2K93gv6W1Bhv0GapdpMy54w5b3crL37ZPfS9lAZ
rdolrcFbgBNkrdi3N0t7dEUmoGn6b034P4GqFMWyYUVXEodtHk98bMNnNB02zDDW
vxnv5O/kZo3AazulqKGoUBQaOCSwWAefbwooxEbOjExEJXIyuRVrQg5Q8uciLVGj
bAD1JM/VCECO+cPAxx4+0rxn7m1o4s4Z6PWjNwN2z1EH802DhaMCtClx4tOWWwG7
ni5lGRPvNKC/+5zWK/ZrIFVpgAC6EAe1iTaJwi7pVCXbMRaBEiP7rB3PV4urXkcU
JLUUqfGC6KpL8dU5JzSd4YLWbP0IvZzVs5DYzGDTmQiP4AtT2yGGroEQWxVpmaUA
HjxpxsjSCF9jx4e2/OKEfUKFiuCkq2FABmEsJ7SNEixP4rsFNOl0IeiIMc7fsEoV
Orp/vOuvG3zVbQ4xK2Ps4EV5BZmxUwJZPis0RoxA2zGzf49AxvjkLqQ+mG+N7lfT
UY4SiocCVouJ+rMct837vW2uK8zLNneZX1R7IIVJVGm9Da4ZhwZeiqohWQ4xukGL
vPdF4ZbGw36lUnJKSNhN/10RlSEyQq/OcdEtOZVA9GtZHBxZJ+yFBHeLsNdG15yp
VsGc9l3gxUt1Nhd7zfUb+1FD8lmPaBdtj5/Idy9fzWIV/u7EPEsQ19mvuzk585+d
Eqa5eAtptsZZvczDTc9Rl2YhRcHlN9kb7YvB529Lcoe7JyLtWSzfRs7og4NKE8q4
Ou29lshn+CBpQPVOCcKRAw2GB4Z0KjZ7a7c9lleCtoDv8PhD8GqlBhuG1UMoyQQp
yhllmRLtXcYdsrxNnW/ojbepWgmMrsTO6EqBFDCiwVAoKZyJHP0IWEcHxju5PZa5
VIgZHYLPUUEoI8vSrrzDEmI3lsv6eTZ2aWinNERS/mP4Hgwg0PBItnped60SJ3Ys
yNFkSLZEPlmY+uXqYYfK2poS0BK1IdZoTS1A9goj9asdbhOc29WcwEr4vsXbHMM2
Oij2jOfJA953RASLxYHVO+2ZiLUsBBlWFCZDxOtHrBjje1T2tmYqaBl/Oejnli84
tK9n6fgOA+MSiaGHyLtEC0XVim3CwEO0BmvmzzR7F2b8wfBHZwAvRqeD2I7z9eWD
KtCq+cVfzUImhIJAD5c/GOq22kl/vOVY4d9vyY1dzdgZBg4XV88gi8Fku6/u0quo
RVggNhXC07DwkIBjHkwqlW3dPegTu9X2byStnGzkTXuBMykkZiPCX0DWepA/dQIV
ChLUrmDewCGJSXyn1TOT1+IpEUMpz/g5T4n7NuoXaV+jwVRVtvd7Q9e4azDvb5lo
hUGFXXbO1Pf5+SzANXpPoIk4+0TS3OA7i3RLvCbpcwyF7xeZVGFVN2X6aAwmiQtr
9Vr+CcSAElrr9CqsQfDvCI25XhAk0Ny9VU581PYORspBEQTcv/D3awWpEE6lLymA
9o+r5MrYy2T2AaDzC5opOrNZGbckz/JrjFcHYxaAlTc72QNE2R5CvugQwXbnc5AE
PLOCjK3vFMcYQinIqp9BroVHzMe26jV4wTltpR0jmtfHy842CuRMz4kizPk+GUGS
5O4djWJ4AEIMeXJyK7LzDjmj6wwL8v9WNrxPvB3/eFB5OMCHpLM0djjGnKEzVGCn
beQIXL04Y5xnWI64nHvczrByvQ+q7KBaN+JCu9FuBaHSEryspw4ozCb548ZOYyFh
zXYYZjQ8Vsw5sCZ2N08tQlS13bbeV2UAMJ0flsSzTqpeoZVD2YfxyQbGOnMuSJ9U
liSgN19mm3D8S1aBntA8gFWS/C8m+RXR86GNBYqXXM3/LFsrX5azXVZEe8XX+t0i
lokhJfaqC45H42Ge0ZK/G6EYw1cwOStic/JNwgeMVI7Sh3RgI7nnpFzk7HDombFi
KF9C/f/RoUK4ZwDYrehwswEceKVS0GFLNGH4UzBRnVjovSK5Rq/pShCZpEAoTPbZ
WZvaClzjtq6YczzhWLj2dr8VTEBwgcsGLoxtcxfO+oQ9F8z7GbjJJpFCen/DSsDv
EdBbYFc55+1mWpPGN5mtfOemCJYIStHXdX+4ESwlnINf1vHMxXVSeA501Hs7j7rb
0kax+a5UclJIgeHZAM2/TdzQ+CW8m5pjjT/3t4qF1YS5cvhUKkPKje+h3yYhmjfM
0Qjb01Qum1B/IXFlS+35AXxprRud3GRPDEOVVeCQyXDvXQrvyFGmsytjaPIZUUAn
hv+0R1hIB76PESeKl/66sojTAIjKx6OH4+DZ8IAX/K+005GrfN6ZFRjmAY2nZuNv
gzzDdbBYEVNpSQVoC6w050CDWGIECSBCat9yqlKr/Cf/I84QrF99MDOrCO6rTwtB
+0+Y8+LtfX0Qpt0xY+ILyEK4S7/JAOCvP6LVI7NJmVJ6k2xg/pLyYz8V8JaW018Y
WcF4dnPNCnWMpJVCKLT05l8ZpKV6WY+hgFsFsdQFdw6ZUZHEEMww92ykq0gS+Fop
Csb9hOYW16pqkVTFNdg9WtMiRVsqoj6w44jEi52B83vp3fu7/BWQUumE6P7TlJm/
JMd3GR9UFIR6XuNzBV8l0lZ7RhdZl9fEedumwVgM7gRncrwZ3A6cfNGrZJsGroXz
Ij2jFEuPD2xKvd8uUu8SIj8TlTpEVxtwAiVIyY9ZQjXjl1fglNGH6hn94tYnVtn8
nNNxBmzb7qaf8LRFVdpJeHQnZCu7Ed4pRw5ZWxdMSK9XDq4p9Y/O4YCwFq1abXuh
83MxyWtEGHjYXVAjJ+H0HcZ0xFQ1yaitxtE71iNxltqnHBu+Eni0P98MD8z3pkMp
of8AH7sIzwJCZEt3zhID/ZKekTyB4EbH0gNuqwSOc/meDDrL8yd6voS6uAMQLGDn
yTp9gYbTu8vVF7xzKRdO+0ypzmADog8XzD5DpcgelGB2zjIqWGoHDNwa7U6NL1on
pa8WGZ7UQEZzREs5Lob4FNirC/jfnBN5+4tBFg31EFvL2Qknhq/c3I4cRTLIYDQJ
Z16G2gJnA8gDRYFk5JTOtI7p3H4VYUOynxjT6CKOAa/cLTEC0sbjnWUQxELd1J7C
Pwor9Ho7zlMdhAnw3xt7i+6s3BCgQG1sUUdGlkrJbRqGophRIQJUzt3MvyJKeJUs
jGQ3zxuySRMnY/79QtbJAwdTEHUdt4Ffi6KXXlnqtO+64dOH9btyuSKhM2hlxsk9
KgmmbG6XRD8dKX7MMxdu5WVXOCk9WoNm8rzYB4vwA2g9SEshkHiQHPbZ2cbdjV3N
DLCodoLMCb6WUAzA5iF6DGvIVoYtR2yMftW5acDbKKYPaCBS3gRFEdQMG7Z9dht4
ELqQfcvLnsd5NUuN38UETD3nYsh1msn1F8ZX+bJ6WVDAZU2tPqCPW6ecS/4HrPfn
XobX5L9jBJXM69oaeDvaGhAN2ZGn8ZtM7wuLDgaBxn41/vn6ImAPWkvjZKdaBQ80
7BNHC7vr8Q3yWQDRoiiUphBfVKyDZq96SNrYoex9+Rq8rrmeejeQoLKR9CYbBRN5
Bd7E6Q5l8vbqmJDqLnhPieJevSSfbOwdIMBU/ZfYb0k0QE2KmPjm0HJFU4imlK7Y
UQjo57Vnm+ZVPEkpk832sa6N7N/00k2yg7rzSvpH7KtxTLpZbtvsvOTd1ISEvaUf
2C3/qhfWSu8irhpjOzw+h7oPf+MXgVRcYxV0MdYtcpUrhFiOS4Kkj6UT2yYpxi/y
b2qdumqCc7z4YMXIRvS5y0uNgMlTl7dolaWOql//OdWO5T4lBXAuf8tbEkUeFzoX
yLg2pvaSQtsrv7PpDCVBKjzpd56GZHCevGiC7RDXIZG7QvmYnUqTXhmxOqfFbkpE
Fpq9nIs63I+l5WKk/xR+siy0vhE8GMzY2NnhyNZIfp1+5x3u9Uje0d/z7XyZRfn7
r5uS+CBliC26QUeMiJzwCKlUNhTC9kvPsb1MKI7sQjaIK+ryFwa/9uXNrtGQ0oZQ
ulEcxkyGy2QJ5ZToNm4DQMUCpdmPER3FcsYHN0pE2T4MB/kOoU2ax8KvBhm4wjed
mvxPz22jAb5m9iv9pcNOCWsOO5QLaYRearJtDAg3Z8P1RloZM1ZAJRWJUBDRswmY
/arzaQmKiiE9+j5vIJinz1xFBnrc1kt/GBoPdGEWMBqUpYud0QmeeDdQnmZNI8xy
ZfIAHYUP/null2/xrqk0hgAhlhM2JzRMflODO1iD1nLsVBiqiejKIU+r+lo4DpG3
RkBC9AKb6ZUXU7W+38wv3tgaB7a6KapoKyVtbhIbgxIjftGFpHCmCPXRIIZxIr91
1aPSrn+36HoML8asG4A6rn0XiFEFQxiyCgsIrv0NuEgK+z6tl2mzHVh1PACJHuPf
PtobEoQJ8W9yFEm7k3K1DL6Bd6PddNBjklhPxTZAeHX7p9SObv4J99eM6Rq5mcu6
jiOu6SjKbDcsl3MaQtuf/XuDT798bAYxlAWmpdcofPxwlyxIGqGzVYy8fBpYx8wQ
hqzCZjPBSMMnf7FDtXrm3dkgr+3BJNLJtZpKiPMvLF0spDVtC54MKbJPoLVlN08f
3Gq6xuGExkdQJ6t2futOIWfrkTA/IcvLzHBbElDLJHzIeA0QJKSsEnsS1mm+0/zG
VY1I64n26RUA0NozrJJJHlBaWrMcacE2rto8CMRGEbGNHR5mvACgSYQQMhhbl4Lw
+oE+zev2opWcD4Ocd/zZjpWgBhLzaoj2JQ1frzG5TKTU8bddHWD7uD0H1eMgwQBS
IB0YHoxC1lfZw4JN7ecD951ZhfL2j7XkpeamH04Qqq4SOM+AZl+RAA60cjJph+XJ
jzh8A9fdJtG86qx5rw8RH+cNYZVyP9acrWs/4Yknxd5SsEU5iJZ6/6s38AzAEvTY
YU2NOsVg+6xpJ68xnOw3Cnj4RuRWXJYZp9YFjWmN70U1l4Q5cCKmzBZnBPfaEFtS
XmL5r1Rr925Wk8okBGddHTrhnEKYbvm74UMTpHDyeRTQAKc01AR5C/wGMNwtMbrH
G+GCifY7dcQSVMnt33TDobgFtxxO7vLika1iJr7CyCXZvRSUuUpJu8Hcq6P/okXy
hZxvH3Tg4Xjt5TnXtUVgktRVSZ7XEqfsynLe64k5t0k2Uqt7e+5GN0uI2uLUhDHo
MbtzCotVlDRvXNP2bU3QHI2aw8MyFNftFxgfiui+AonIChZG6aupwiGxHAvgoIxn
Bj8z4UgyOPNc+nLMp06ZOnhDw8OEprrMt46v0Q1lmS7lVUuPnoxlqz+7lErm9YDA
9s+eAoCAGEadaL4WXquAJYhQnAsEWoQ6+gdOT6QsCzlBX+0uACw+Y/BtGQx7J9B5
SPfui10mcCPaC6nPdxNLnifdMdURaWaZPS5z4xERw55HMlXnL+9NzeFWS0YCTdIs
QjCIuVYqznRcsvyzbHKVqjV6fWM8U/x/OnrVip0Ru6E2TZ5yiatF8etSrwwOuT0O
Y8dnsCPp4gzp/TG+U+eDuJGX2A0rSASDyeoKYaG5Ymder9X23EIICfJdKyvdwxo2
KkwUz343vaEc02xGkHmHNgXDKpj+iL0vRQRiZ/svykvRXNGy1HYx4iyW8AymtcyD
aOjDi6FPS/iAgsxlFRxFO7jNxlOcD7Lkl4c3VbJvOUbqkrZfTRixV8ibQ0tdl5ca
q0Xen+p+4DU6oH64dZ/fJRMr6Wbg8UI7T2WQACBditKpLrx9TQ6N8i31SQemYUE0
tVjiQUsrUq6J5BU5rBOSvFF4i/WBAFPlWFuoqur1MfF4q/CGqbleG+zD6Bqach/t
eX5Q/k7YMt00Nz3cV60j5nysk2i6LMF8/k2jcQi6PjclZJSWBwqqST1TR7hjEyKr
uAQMeXwVSTBM0p1y2vVur/1TNgvTLbjA+KQWPaRDZT5r4j+gXoOemnO3ByFVvr4v
EsxBwz4Q9EpJHvgkDzk37b3rVAVkdLQvN65tgzRqnUDOGfDbuEbvKdaLTwIGzMnQ
B4Tsr3gKz537TOUtyG025abiMWEfuJd3hxpWtk3sbD09vks4iMS3BzTnZtcDkOZr
A3od7M//ud/Xbe/xZashrL4C7dDM1WVk+9BupvxCmVezU+Er2Xpo4Ltn6s1sOAtf
2i4YpYn9/3sZFwa/ftoGTlTRAFmXj+T4JJgKUuAWM2QO4yRjfcYZXBWZcKtIQEzY
Cp4tP0vSl230bdTpLrfCieyYrgxgZxJgctj54ZULwvf15AtAWHLWNT0Sa4Zpt2J6
ZJlTKPZBjXJ7bz1zfFAui0sZXzHWoSoyEWKHYZ2ZdJOkNDkjCvLU5WS0odhEa3+z
mwFunpWtgSPEc7+bf5wL8PZP3cxhCICls4st8NH68mkDKWuLTpkL5HONqZRwlO5r
DIDCnHcuuOydsuXYq8BuHBq3BC/YdybpTM693Nhh3aGLlATGeUauelDH7y0UAzZp
3QwKzeHmSVV/LbMwopnGssfeNFD75Rzjp5ejOEpZ3PsLJRQ2kCvTu3PgUFDkJg/N
F3BeIMSluvYwODmlkAG/JyfnzGwGrQhKBImGtXGIedzogKRagPNAwue7MGk5KWhX
AVcNeL2eMZgSBBebm4N34SnUxRsgUCzxNi448KZT2nka3c6tm2lF2daKjkq6HyFU
KFo30MZI/FYdkMKBhoLP95+Nlp4rKWk8IZHww90KDFGS+jCqP1Rt3E2O/8XVJblL
5CIolnrmVieCavr+BdSHE/XHU+EdtYH/5DB6miKXByHPM1MgbluwO5XSxQeLbATX
Y0Y8ovZtJzb3P87QNQNAyGaHTtRS9ZoQ5bzr3P8i9AJGGAfa2tTZGtoU6tmLl/d9
nu5hh1S6+tisQVsfEGLAT6xsdzDenOTqddFIPTUvtvLj2GXw/jl0PRFv68MIlgr0
ftshO7wlKOTgLhKBt+UZcDK9PZcld9F4Oz5l8LYanUOdD6lmIqnlkhcZ7H5GHAr3
O63KjpiSZs8UIkU3g6jL/UXZMoQ2McIzSv7NBgmpDDTaUZOG/olcHLL5QSjWFeep
HAgDLN6tvfij2c/oZq55vda3r0XIv2+pKTXHV0KXTAgdmRQP8XQj/9U1FnDUeO6B
8qazINnBs6R1SNi5ylc4ccIx0PiQYKC/bhsMYjWZWb5b287Vy8MQNYPE7xFv5a7H
wCAgXDVTptyqQDEFsBGClEp8AXEBEuaak15UWLgr2pvcv3fKSr8xRA0rNm4px7RF
DC8K9w4m81Vt51uPJGiputs8NGA4HfU4mz3himCXHoZkuL+i3q60WA4sl5FnbS1c
ik/Fvjy4ruRNDVQY6P4OUBZyCBDTFj1NVz4tAnK4+wKsRTfKBgp5gNxsFshItOhd
ViqBRnkdIro2HhUR83jTrYA/vHSOEqs1VDmHyr38X41twzboAD4RkFB2/mCCUByr
0ajR+q2MR+O/X0jvgRUVLuImU4omhmetqYBW2L1MgzptF+luo1fBpY6k/t17gGlY
OrkqpmFYlZq4IZ4HD7QoqG8VilgMjVywrlhH63bey+6wrDjKBOjmeCudibcUvwX7
keBYpEdeSfk+y4rkD40mKmaaTOFN7e1qytg2juBvIeRYAiqKPt/hBEdFiwwnx2x3
/qmNSCxPb+TYm18Gvvyutv1w8tuM/uixj2st7v2loDha4F4EGzO4/FQpfcwHwwce
EE0lsjVOKJxpkiUpW3AnmCewBxo/Y+du+2OeiUCabXlI4XFp9QtHaTF4mSzVgkbE
TW6++7ZgMg9uazaVb6AMIgBAT700wi4ZjW2lvfhChvP6LF52gMuH7zK4pbWKU5kC
l7delkTxywHhK8L9wB8RNzB2CNUZbSEubVsPvul1bvYYA5f7stEsM5tAWZM0v0Ul
5f8UTCJp0d9CD7of9LGv+X9DRF8SXMFXSqA2W3vMC1CYNMWpou3uyLiDEwCHYyn2
tPduO8w+7HNNlPxDm0jmRAoZRPygVO9zhc7QhVG68wzM0FwJ6rZXbptzZBEMV4Ag
qo27QvJRvlpBnLXnKDg82+8X4wWHntitUHXfbtgMU7Z3x8lY5qWtu+YlyRTUY48P
RZVMI8zTqtBLRH2YPgakG3B02vLIrPegM3flFkLzhSr0TspEivUHlu0mAFJ/ScTv
IKMtCRvArGjyib0hPbfgPEdRYU1xckequWw27cgiDhN95ekQL0tltWKI71msLSEM
qP2m98b8e1LczCL6jZVscYqXzcRJPAlpXYWEiv4g97hvz7eKJFImXcL13k+lEYlA
ESeOurxoheGiF26X0zTx/Op60T8PGIAvqBOiVzPKiySNNcArd4Ff9droyv+K0C1R
to7RC5G8K1W1DQNFOxY98wQV89MXNo+durS+6iic5E7OGj1jZ1nSeZevmronlpC8
2GzFNU4R8kQCK4+BfLtZ3vlWCoc7snUduYCbzF4VDqCyem6xmtYNrmmxVi39A72V
Y1FNMrCjskPjCqMmhqAAS54VspE+HylRsfMRyLlqvFab0/GtbSUh0sNCRJESGwg4
i1CiEPpttsMg2uJkhj8dPiL5swdzG9dxdZ12TvtLaIzxox5Z0wP04ywaXLbJmViq
Hpcjcu22ppXTAnqT/PMQlsJfrivk+o+sy3mGDwU6w797d0wpw2e+tjIdO7VzqLdj
/BBNLwTQ2QwLLJSfQOyvKme/HRNtPflRPtscLTPL9RSDV5FfOdc1G3PNVpMbR86b
t05LWZuLNKAok6aYsGAlRaE9vLjqNIH3Byq5HpjFluNHo4IHVA3+VMXVxHwfSHfx
esCzdOyX1Ymt85odUY74BMc4OXHCXScpHW1XzrcB4Q4LPgCDTRuno6EfBCxneDKn
ffw3Dq2ywck3NxI4lD/YJq1DNE8UZQb47RLdOKA+/AALIfxErzn1mlnOqpcOI4f7
lUFVSQl47DXcRmthAHcB7otTNPqvKZj0UNu54a3GCl+OoLb+zul+viEZCai4dnPU
ENT/j/OBC4u6xlSBndtdWcPyOE2G8ecbqDJ///f4cfl6p8OvVwpa20j0/QzdtwLm
ox1Nb/Xprx6et7EPqPHTJeuMxi1n4cw6T7hWKamzWKMGwZmfkzSIhqGJUJny7aU9
3B5lBB6ppLQ6ZV++aD418CbUtn0niTPX6zEfssKc4WJoWUqYcpYq72R9eVln2zCF
0rR4uMniNmADAmiLXqf5/++5K8JPI/G+4TfuZ7SGo8CGlsQNUQZhbeiuKmvGMyIo
ygLpGpDovDJL+E8kHLB3CRVF0Qfh2G+6ZpLrjoq++yqJv8U3zlPYMfMep28Mifjw
BKtuzIgATut8hh6QcvTTxp01RoHlTc0ji2C1jm4FBQl2EbMmdZU+WGg3VC/BolRo
fmdNbEJpamBsanki484COGXHm4e4xMnz/ngSqxXyJtLiEl51rllyXcMqPP5astY/
rENcJMMOUKLaqtlqK+5hAAf8bMiWbXd42m6o90oUCDRRHaicBEEcY2Rro/juiIsR
dyl3QK6hzx/RFQkSWAkvoSFNHQkbjRma2OACr06I2teYAZRI4C0WpTiC7yRxAhFb
O3mU4VgEqfp28wHXcpdl/qfv12HciJ7qxnxZ6vr7EY6lFuttBQft/ED+vVk9q/G4
0NXfS7VQikGZQxSE+H3YOg5CSLOJJZRjV0r5HsDRe9vTyw0tbrjB+wQTutbXgIzU
E3T98fXaWD+30LIz+NujBuKKVVjL8TmrcmiezxzOIituilM49FGUCSmgbLg+9Fpp
P+PqmSjg34gfOygjC6zcKBJpXUf/l84CR/LKINOWQyxvmPUsYJBXCJBiU8OtOre7
LnYSmfdACyoJI6awA3COcDUA8sdloAdGgPj5KuAzdehJwk3SPjE2Qz5vZn0yeDA7
kg/gwncFXHOyEQVR3xxZEY7Dq3LNqIPU6YZBWmrZokMislQxS8QtG1j6R5evcN0X
srDjDevJfAxqZDo1suqu9XEmNkvip0GTQ1VUWIYolAmgrZW+8GMIjLnFVhHXXoCz
+p02JOPcFWGHH41Rz2H5H9W8IgMP5e7JNUhbuLAhw9Qcsx5DP6mLOuP6Lw6lki7G
WHUzNdlmplgBCIKZFXQtANZz43sldM7YFW022WWOCl2PjOOyCTzngsnUlCnxwFWa
wXsOLT3/SECtTwJueMW7dKaRhf4cCs1Qp8RQ5PFo9Q+lf75obCKdPAX2bPaleBCM
u3lXzb7bcWZgZDFrupAkXb8iwx8mGKDdtHNm83qGA3E/Ne2uYW2KQT5Tu1MzNs4/
V/aPnZVPpBr2Vhhax4EnySQ5jjLWvICMBulsIVXGRsd/lHdCW2MH6h8c7h4MJn9M
EA7pC3sseo2F5WVexQkzJcsohp7/vKJQr6J0a8DJH7+IjvZNm4TPSJ5K6CLDHA7c
ePifUNiRVSr50VgDpQ99msgIiPzfBdsXx348yRZ3bVwuIGX1CxpB3HD10AWqHBbs
5IP5+nzJD1ov+LJeLOab47iVA3o95GiB8qY/XznyuHKNG9fRrB6ZY+qWVFN9VWC3
knzayfbqAj5Zvl24L7cSyij6eQKRJkFt2CUo7zpVhrnKWKI8aHiqGE7pvLMHkRJ2
auMp5ylIhnovm5YDzWYkv1XgAzI1we94C8MqUToDt28SoajSDCTs+hIUGuUdvQGx
ti6exg9nwYw5GH82aq9XvXEA1QzzAow2YU/5m1m8U8k=
`pragma protect end_protected

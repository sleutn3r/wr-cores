// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IjF7MvQKQPCqw9W1+L0KEbcyTUPP1z4wmC9UqdCHIm6hG5B+AKN10oTD5iR4J4Jl
X0F9mzPfA6w2ncuQU7kZaDeTtSinwW2/X4/inPrL4zuPNWJk7i+jCWJMGcHClDL8
CfYFXfgtBdPHLSVewZ/7cHCiwoIv/gAFYTPV6Rxi+9o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
71Minq5K3AtxQGAUuUnV/nwCYSi6zL2GhWXetYV6EPRZoNiBuO3ma6FcnqcxPAcz
Vu+cpv5ErVG3oq3n5gJAG+6juCH0/z6b31LuwOVyliEKyq2zQ6yFTDWTRYZSc9Dp
oy9iyHm7VZ0rtq2e2Oy3qXayZV1KCjnnZRK8dxAh4I0ljlbBF2MMsD0HLO67OaKL
6stIT4oGSy63y/JM/u91am8tw0DhNm8oW/DY5zWMX59aj8zr6Izu63VLHaNeIiev
5ZYdou5F6ZiYCf3ERLTCIngqcihmr3DfSj3hAt6S27tTT5+P9JbzRmHABRr+Hoil
K6kl/KQMOkZwgxLfghhjGKFBSKeAJWT001oHK3OIole12T1rsKTBrgDdvzYvbU0H
N0clkiGKy7m9jC/zbcVUZI5iQAJDLhdr/LljVeEMibdYWZaLy1YEtzgikvJIY3nD
/i8AFUIvKDInHvOxZwwd0P8PIAu/y9j3yw0ip8Qrosc1aQiUk2wmcRreG2vuYc+X
uGB454M7xZCuV1sIbUTjC9JZGFt0+8bOwrIwpS/2EdBO2+cRZ/AKlFUXmWkDZLdG
5yoZHlHVtZSTXyi67zCh2tjCD0uKYYY7MmET2/4eoHTuWBnudGcUHeFCLQkLHFEl
t4K0NqQbJ538imq+VzSIBvxTSLdHfweu3wG1eNq5X8AbTzInnWk/fzquDb9mnvYS
WzI2owh6npJ5AQcR+oRW2uMlikXCxydG6LxEz+nlNkKGR06y5hiCzok33fDrIBEi
uTa6fbDse9UNxiK6XVY7jDHyDuA2/v36/VdmolriDkapAtZmBv0H/Jkt4+YNZHMh
VjRhEPuLuQXASWXYS5qH3YRuaX8AoacOZhZE73mlY40VgtNmmzMThS6FoDzB+WHV
9Vte+FS86HRVdqktFiyonC30A8vDpmEYe+E2PdXxJtRTw4KlR/yyKICjm/4alH3Z
5UD5GcFA0+M1PULbZRF4FV396oUpI/1uVBNs0VTAwBW9eBdGYMnokKbvVNB+r6bv
hsQ9q35kdTGBbrLbHWt4GrsfKjvayYNDRE1h5//COT0vhCS5+YwEDu4FMkgv754j
O9bRi5qqsUaiIUTquZC26zWufTclQ+bgeppL7VogglR58yu2KsmGhP8++PuL489e
y04Pf7UNxthh2psjIVEU6brz6WfbbnE1qXVPoVCtYo7MH8U9Hpd6nJ+yxwAtbLk4
/DydNPGQZa+J3M5d31CkGTImL/jIQDddQ1Lh8Ae2Rc18ATkFl6W26jWAwXqXO+zt
2B4kPQSZKXroutmpeKNPSLTPkzGpqWTmOHtTfFyIydTTMWELjREZ+R52udT0uJV2
195zNDxorN0tdPAnFw21STjpbhnHnlOY2nA03MmJsaUVDb1CM6fjNY+wRndUv1hP
9fky6LHbguT7dfStu4Od/OMYFWkeL8PstFxHIhEp0g7tfSyRX6hIm8qUa9bB2CBA
mr5dwgnj8nlElpDWKi2ufnuevAhlLJLz7s2nEZsvbIeRfKjRs5Q14SPoTxUnND52
5mumh3LkLRZbd50+/lqPc5N6uEVPYPj19ZwCfvdNciJm4/CShGUL5Qw2ufAdhvDj
EggO5FAtg0gAd75Ped0lK4UoxcQd+BXAcJYIvsCV5i/Rih4To+oxpIfJJ+mFJ/iT
gT3GN8nSwuRVNGLKATWlc3OGemJ94fDnI538/BnmKOybt7Fg1vnrYXyxIo0WIdql
SUOlbW3C1BFSzFde6Ayvlly51WwydKLbr0+Vebgg8IjH8nVUZyKWdW5EmHIhnTii
O6OxgHM1gv4IQtyHdHsAhCeraTx4anLT01ccHZNOzlFEW68UYeAX7u6vsXKUwgPS
e88R/hE2WWFLa1lZdsybs18GKFPUowUHd+KRc/ofF6nP/c0wTL+5VVDd/oW83Dq7
RxXr3P2/T52uFPKkvRXO2hcHhxSx0aV7FqyMXSvDSONVP6vFHy2PtKyECr3kHv8a
uOrb9qiuWMFRWeSy8g7Dnj5VXfNbl7l1YZJ6AffdxRiDB5GKhzA47XH4m0xsNJtz
yClFtrVXsj08mG/unzz1Rot9UHnZcJpXV3iFcwRshx68MiqXkpc/mBgASxBB8Mut
ROuPnU8gO7/iWdDh3dQfvUmigkk9ZoWmTxeccwy4hx4ww0M8B11ZRVMVMj3pDdPP
e45H4ZaOTH3UO1GxQ4W+sNgeoVN3djcLVhcc/hcbs0HG3a19Yqu7JRkoTKMyrMZG
VVsbY7ePhR9nPnAsPseoR9GMUgsyqf259+g3PWD53BjXAyYB33lYAtpcqftxDo92
FkdRz8FR9WeDhTinyr7PwPgzO2qMLJ4JsEIArKIKwSrShOk8FLInk9uuB+v9cUiP
FvIEjP+5SCDKALC0WMbEk6u6lnt/bLh6JYHeisYHZ/Vc7RtiX1reR02D+AqAa0n5
S1ElnDtMQb7o0oDz1fEQEox5PB1mlznT0WWFdaHAObp8ajLtHVmbnT3aC4Hd2RF7
8MuVojdbPnpHqEmgJx88wd/i3OgE7W4O9Liczl0ZyVlFA1+6bvRmyz/Dq4uuTryL
SNV1laNxJ6zJpDHJnkd4HU/QtxkUE2o9SSk0lD9FyCE8AIzqu3STEB477urcu5Qj
Gh62/59o0tL2/yajK7rYhbbVzILQ5fK5joZxnBPAM8D4tvTt6XqRHo2gKCvhOS2H
3I7rAWeLwyDA1I+x7121ltOgEcGr52fJHxw+8hI/n0iVqZMM/xiuLkLOkViBLa2S
0l/Gg7aUEj08oTr2F7DnsVfgus5pMHDqfpRMJvt5Ud8/aZg/bpVsU1+/nlfxI/vt
KvFwo3G5maLJDhvGJ73u0U0oCwVSwPUfypMJdh873A8Ji+9XHC1wJRKBgnsNZlRM
IzBhDP9ylSMmqkXHMUGVjp0PZhwbzKEujeE2Wg3pnZs5bbZIvmxn0kC7fXqfRf8C
3GalsWuNyTNPmo0qRKWYhiLFkwOSQKpu0LBOxpkYiywR1jK+gKw6q+gHb6AqpJTM
ocCqQJ1GEGu5IZCuAx/1RR7JN2+Fs6r8M9fi7dtj6+bMr2wYg9B2yYdcUA0mBMZb
EHN9UqTXqQjH6c4lQ491FdFepNaimB8g+rednY/dRx86DSzBr0DeoXLAzAqDylr6
w78kQ0C5vs+zKJAxHy35xiWW7jj3wimsc2J80Vaio8ppf2XtZ9CnWpZ5JbJ8SXer
4H/kvty4Qd1D2y7QYvylav4MDPb9GFZGrVER7xCERFFDO6UoiUHa25DgahTKqxN7
b4e+sW6+7qYrTReDJGQcKc0lb/5ZZqfBcqKf7KXwk1O/lxoeEN8/i2srOPgH6fYb
T3rmgZIHqDjirrRU4UMzesWFQumXculdWnDJAIZUWufJyIAihnXoBszIe7oWB2sN
37vM7WnjSFGufxnsHhQp3QbRzMdp9bP1LxtNjmGX8v/dvcAJRV6Kl8hWtyuEz4nF
9ItMZfFkOO05T+Af6GPwGRm7u+XK7LCNBba7EpiJ4jZ0oz0JtShHTbkNGcvpOeXV
NgJGFgsjHzBj+Z8h9OgRvW9YB5oVjJYieu2cXEYHCyRHUV1wrks53TwL6sWt5Ovm
aFfmHdFyBt9hHcij4pZjFT8zc3O11D5kF2nY5P/amoj8+Ng1b3EJH0a5ClDv1ZmC
Hh6TrmW1qUgPF2nVU3rHWjLuY/Q0bIVZw1NCOCoK3ofvkF/5XCLoymdFabSfM7O3
PO3EkLZhYKYiA1Waqv5OgHCz5/Ri0HidfW4XW+axVa5yM7mmgq5JecFU0R1KEE9g
VlGbUk8/6sD1f781A/gypoyYebPF5AnEBdKozF18M1z132WvDsYDFwLycSv27y0i
xV+449MYPvET4g3ArVgb6W1wZr66MFCZ+elIEN1zxFDMvwQv1qdLaetD3RHyTcdL
bP6P1UBNR9Vi4vDqGOtnPqSJDOM7VA/l3fGmjKOCqTwnSVS/GRcZBZ361X37WYi7
xXNt07hLXUv4hHwy8EbTE88C1t3Uiq3s/wMVKzkyNceMx7mjFPtZBvz3kEAf8BHa
DjjhrYwRWrrCl5y5YoxKJtQKSU5BBKSRB3HWFlxBd/h0dFEMT4ydx/GKfdQcKJfz
NpcoFFaAv4m7dwgOzDZahW140KxdnMQRAEEyLGKewyuhOgk08e5bcRzfQ6gMgrEz
04PjYUjrnl88d9gYv7VTRgAvKKN828PtwH/JsXFMYC5IQsljHa9TgDsuSKr4di4x
qF/37cWMvnSbKVyyYCTjumciY5hX0lPAcwfGprOQ0Pk=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VdGNV2/Rs3oMG4Z/5uPBMcAQfyceLMqbtF84lHmZuq1Byso5KuodiClm2U6mH55h
3Wl1YVEwSkxkpVzFLSR1ptkpKGaNEKNouIX6v5wjUQQnxuqHSF2qQ1tmG9NjHh2C
gaLWa961OPHShw3KVc4/LFBqK9X0BusD1p2w7eB0rcE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19344)
Bo9FIZmEtbjqhte7RWx877KtYgAVXcTxXA31/YfZN8tiAx2RHbp3ZPbxxfwI5D5b
dJLTMFBmjzGArgSzhpOnIwMWIn66U5K+Qqa3gOiBoKbSg/oMtwFf8e4JtRsrjqpt
5lK7FopN/kFjdTXbogFIcU66zfVs0aBUYw/dDTAJgMlqBwtvjNhRDdP87fXPaz46
7fDo4UcowJSX3B4XsgUpzeHYlwW/s+EQAOnTZlWtf4AGk0V+rODLRPPe9c24cGeJ
/8k0mp2s+afztzUURPnUqponHVxgJP8XhuqvPJSoAAcEcoRI4Ycg9EuKFxT0sL/m
WnrUDHRjU+tKB2q2Y9kIyBnZj2fI/I6Ly4vZdQEaszDMy3TyiAvEGLBHc2KiJCuc
F/AweZBaFUYNk2ruAMBXzdSWrbw0dPBQ6mFvOhWemu1AXzYgFjuK1bgIG6esz5Qx
DVr69PBtrlqkvTVlnF6GKMJ53JJjpmHpKJDKNm41U/EJsvG1eZKYERQqIfD8SotL
aoahaUxfa1qsY+MbZE9BLqE853/Vz2oarXAE9SE2W2gU49y9SEnnZbv3dwFnNN6J
nXiZtXk6McEiMKwhb4ZwASxxuLI87dE0nEqN7qLFPP3kTdrCcUEBbHUehbrJ9x2Y
hXzDuVmfyddnlrV4FK7wh6vUR8CUsZKUSMBu+wlTbWl/V8I9YwYH/Z3pvlwT1SZd
58eQRVWv4b1+EFaeV8kE6JTE9N3d4QJOUG4YNuYre781r44ogT9fY5pXCbEHtPBw
sBucnII3R56z0f+DagzNvraRHANq71/DaQkL6S8kwp0YZ/z4KUL98RHC4iO8HbEx
2bgXr5zBo5/9TcCg5TeRcwhUP2uONwVgxRLvAsQU5Hy1ZPvE7tPjZe2bSCPreE5E
h0piFCc8cq0kOjnuydhZt5k5E4/c7eW5LxJ/76W4Mfr3HetVFk6kZKVqyLo/Vqff
2e6950pDyshxsiH1Y9s3KKnyj5K+JgZxj3G+9HB8kAHe88maKlf2I82vHOFv2IQB
D4DtHFwG1uor3pWPlMIMT0OGvcGcFy20JyC9paCvnqUFbcPrg6zrdraxhIRWu1e+
mDN4RhddGKfNZOlQEg6+BP+LBVEKTroPWxxpu0o+hz1DdbYiAlVvw4K7hfx6r6CT
W0cEQDN87Gfy4cNm+DYHClekd/YLyLMrbgFZkZPGfVHl4Ia2bNIl17M44tOFLrMv
+dz86nByeV+aA+FdD0sKkvGnZnqww3iwWGs/MCaUudhj1FI38z7k1GnQd2a++Bpu
u5fibtkZfOPbmKEeRik8ZoMB6SoRtcf9Y0s2rxcw6Oz1LvO1wV834G6uy6CFgi56
VkU5ol4p6btOZ0lXZBAmmseWqE9Uu6skeFGnbh1sO1TnfUFc8b9ncgJc8G65+Ys1
entGFo5a7AQhGPxMiouJgo/2zP1LYV41KB2mCylbb45B0lcsPwfO0A6EcnqmieOG
ZNpmkLnZUJ3mkMFeob+0+QLEyqWNJb1/7NAmdKKECqGnM27JcUYUqkWXhRy7OWXx
HkRqb2cNmlwBaYDd6Y92Asj4UX0hIotPBU5sya6eCLeiI+CK8HgeiPlBv3RYigbl
wrjbNrenqcqIACEQ7cXwvdgZymxGscRuaP4SZBLf7m8GjAA9PK/2eaxbGm9PQ4qA
XDE7QF2VZttC18Rc/OEaFtL3JJRUWbFynz2uZecOwZvquvhDhiARs9eWO7jxK5+L
dM5U3B2Qgz2M1BByRJSVbwcN0sU8Yfa7cbkh4m78HolCM2k0gjkLdsag7LUb4qK/
zsZ7i4FgEdCMwTBl4SpS3Wehc7bIqbK9znNRNcOSVAR3ATIBF7kWCGDsKPKbY+5x
2A6N+CrAO+iy/Mmy5bhbYdEyq3G75UJvaOlSi12aqxiDqrZaN3X14aQJtPXVNleN
kuWNCAh6wT+PQbha40qIMdGxp60Yt4PRT7Tw1cKV2dpvE5jefNs0hRw5WYuR+w6i
MHmxwM2RX3QQEOtQq5tVNIO70YsfrB8Nlu9WhP3vDNVwJ1qhLY7Y+lG88kYhgdQ+
F/yrI3UFo99JIMmx9opqHpazmbJhqGv99QWur+P4bqN7uxE9NcyeeL3Wp6Z7CLeo
UbZ1/AHuHBNAIhMGQ3iZDdHiqS2q7KeF5FKrGIUFl1RVhYMhgeA0kAUqdL88Yglm
ZBFazjVp1FG7p6mVgGlbeyQT1pwiXCGyQCkdw2aLeQKuhNwP+sVQxirqRFioXEdE
8uFwv2624HEy4FmwaLQskUEi/de5inCq4sf6eDXySvXCdY/gJQP90QKJn4PaPKUU
noXjduVLHsdQsOr/S69WfvF4KlhlMiH28cdjjNJlBSpjA1BAVZZteEz71xvHGhyf
QEu7svQYIDLJV6Pv1DWiZnq5qYWCVDGGUu2iyzm8YAH1Hmp8hd8zrzhFKCW9ZgR2
gXbJ7hW6Ul2Og1YFycBhmR3XkSiFkhCR78Pgm0GwccL61v7F4z8kU/LLobBsTsqP
N8tMR13GuIIbpsOx33eH0P1sEnDDqxk/fLkIpyE4S08jw0fAd+pyIywWHiEPph7r
C8JFGxJl087fi03lOz6gWJVlIXRMT3XhX2Ytfl3guvett7DDJCds1oOzSkerdQof
wZmgdZxUi0BjzjUkHyKw0bTr4whSV/DK7zGFQlsNZfOUt9UmeNL45NPlTBqzvHf2
Vo9C5fMabV7HUOTxm2pJc7eMdbCdZlQUWeHiXD5NqV/IoqNEm+j+lwzRfsq63sAF
4t8zbzTwK/9inRGeE0UthEHLoTbb4SWgAsF6GgGgcim5Zu7J4IP43uKeWcBU7kF/
2pN87x/uXtiy4sVuUZwFVcK4IXE4x7Ur+hWPhq5XV/GauJRB8/8WO1fJKWrMmBfL
a463WBtsHEcN/Jx+Jn7QgCMxf6/wksr7rb+9h/FD7ZVt6mfviRQVtIJ/D/xhC8D9
f1QwuRGyvETWGkGTlZrsdw/JGxD6/uRGmEWFDB8LjpqxLSXgJbistm5f9lVzbgCD
OzCtRENjDn0FCwE0RJiUkwqsDbb52tZXnlt1mauuIzMiX4fDdsLMF5gpftW3JQEm
m+5gR0vc+ySOYftwdOD5lEHPlheeHoY06ORLMqGqhMsdEcqBHFQ1AkScuiUEsAEx
ho/pQ0olQFTMWh80xOn9mHWIVlH175Hx8zT2Jpc8e2of45NdUWsDaWueo3SWsats
lakXTv4e+F+Ze0hCvJvJSQ878H+uLEVuVOQWAIKr51xPkAV0hYKinkPgWzELA9MZ
lesmpvwPXfiQbO7mLigoGqqO3MIFYVScnOCMMNp8MAW7qO64bl7XQL/oGpKpVIUS
hL0Uu+iCXtq3JefbqzdiUBWFUCg6qDZGZPmiIjFSeoGk0vAkGifzTFLfW8qtKdtT
KAJinFJSAh5xeDO+o+O2QOUyoASMgH+5PUoQHDzLG6PIHuuZxv0PFyjNMiWQisl7
BO3zfSCr9F42aaTXcY6ekGwBkfDm8ocMAEkvTG9M9Br7ovge3qtnagcqg2g/xlb0
PRmeQ9o00w/c6hNvjBmScObrv6ZxdgV64biffKKX6dSS1GkA3dYER5juho7D7f2j
obZVGUh0bsnfqWVwrkMoGzSbmPbb0hWcIjZikd4jvBAydpIa8g4vVhR3DtjjcNaL
7WZLxQOHIoMRMeSsChBCquog72kqIZufvU8+8um8N5kdGpadxf8ZpqULHPJORtOs
0tRm/5CqdmAXuLlnIXzY9aYlkCzHTr+9K8tmBu5rLFXOBuVdcuxFiFmZJMjrNJ84
P8OnFRocooli9acUg3NGXbryrEgMrnG9DXz92aBPEo612xXs9Gk+miMm74SOCytW
2X9gq4TfybIE1CqiQ32Lu40Y8YtXuVqT7xFGSA07XUeo6t6J8vOKhwLN7F9R2Wm8
po6m+J11Hl1Gp7pwRwtI0zrZN/HpGDV9yAf2wXVdXYQpUhSLho8aNWGquu88QM0D
36/TvU4o9xbovPQF9BDATSTihLXXKHG2dGln6qMy6OZEyKv1NbTAjA9cSHcerGiA
wy7wkGgHZOne/YaoyabS7Dw5dui3aZr9ZhVzXx7ZpTGFFN3apDhviCA8KCihCe5L
9uDIbgdtgcDofLb/vlnPB2ktPFntyqoAQVwFBuiFj6+T8jCmBmGKDMqZq6f3wkwQ
Y/rXeLEDax9X6Ny8YsHiU4VuvCjKuERlMldQtZbHEdcCJu94D1wnXPRckykEA78e
Qbs47vjDHP2hA3esOaer6AUNvbhFkxqdSXPySkC6ESUDNBJW9tJiFHhDZJT+DZXn
UDGeloe1Vpsm16UnEzLUt4Kdex49t3JnT+NGnXeuxsSvSahBbusbLxfSjlyFqFoK
PMnHwNmBpxTqaGFk0t6Ij8c93YNjkSSPGpLJgJPADAOqFPrESEwue9UDUo5TQUX4
KaJSaDlpNzKBbsOCtLi/4dV1rQgsEU652J+gkPBhbwgD0gye2WCb7nA0OzdH0hFP
pC0fe62sicUO+HWs8ZNDQG9OZoBHWQjL3fJPiIIQIShlccWZKzinDtBMwEtwTwmx
o4G+g3thPxCl7iYp1sCAvwi2O2dziSMsRRAkCcMwDgQayKlb/g4C+3FiFb8zrEIe
XDKG+FQKCnOrnVwKZSCGB1Pzk3Xawjwuw3xWerHcX1U16MDDbpeTkdwm2oZh6mUB
JuqMHWjfVkr8I+TAWDgA4CdQvfwJ/gMh2QA2OTHqjScBhYp72MkX6pdTYukEgyW/
BcxfX09g8mGrdRi80GrXbr1cTTumX1KdDyZknl5GoY+oFDVSUbyAL2XCcEUyW3dr
riFZgCbW3vn3FZ7iNZAsVYCaq+EP4yTqsVk8wUuoUHscN0okJLtuN0kEDWQXGaS6
JAdGSXGQ7saTN1uzzx+xKM+NyEU/SDJa9jwJFOobLl9hIRcP85q4DrP9mvAKhVib
iBG/8m0vTA6Y3Jq57gqFac4mYjKclPS09T2NhdGn03xLtNvlZjCVvv7kbbHyFNLh
R9b4koxYI+ACcvXT8GfDWDlSoccA6QI0GijyBnf0ABj54u7n9rDvFV3S28dvVT+u
5uMb47iRc40OH7JfEcpETenb/Y5ExMsf1wqnQNkkcGC0v7BdoI0Yfyd/y4XL3E8t
pwt96JzD0Lo5vtmhSVC14yJRajtkgucRE92PFd+vhUuQ1ocwhFw811tVtWQQ/yfV
DTVrQ3Gd5+Kr121l6XSh0GL2hGZYDU84seD8kcOS2ZtE+rc4zmLgSY8GB2gbXD4B
j9pqDOKyq1HLUs+q096nmm18I6XTc08L9O2eSQiF/SDcZfJxzPu8qayf1I6gYMTW
9lvgwa5cX2KaXftfAG4hT41++3RM9ERJSpIYdQqeKnaowaIOnqut+NAu3OmlvFXe
jfUTBedaYcjn975b211h8Yo/pupMe8GjM4rFgQV9rm5dCnd0AAKfWBQXI3mng50m
mIh8WB5ka+5isspeoULh23NDc8hWfUJgPTukXQZhWuWS7frOl22O7FldD8MDPQ13
r9/exDzX8oajuh2XIXnw+l+6yUuYwI6p9RFearn+Mkpnc2j9WeL9scqkwx/eFl0Z
p6cED+LI81+f+Ai60IL17YydUouQjdoJWcdvCMSAgnAyG7zoFb/yAyM+nnu47SLv
ulCwIA+dISxEzZ/c0LoajXcw19Z2Io5V49wu4DnLDcW9NK2HYg8WQjIFM5V0FvTN
KD6ETTkfd4ARJqY5uCW71kQCn/6ee46pixw1dDnthjlGyP0N2pW4Ecs54NHOpido
IDkua3Snq+hQ6AhiDjZ3XFxFYtOnvbJTWP+xU/QqaEdgGfYWEsnnu+BDvAWi0nfr
Ain+OUzrXwVXh3n5AL8EYOa6juuS5hfdGUYH/CTNqYzu7rd2hBuMhgckxYyF0lDF
g9qA9ZmGA0Ar5O0+OCajndgL1yxPPluOcg+rrnH5V1rzH13B35nYjwYHQRhVYEO5
Lo9KPOOL/Ke01mbS3jXyQMdG1p/Vb7zzT8i1VUF9ZCaMOA6O1GXzQJGtvKN84D67
RKe1j6UD1TLHb2sfOgD6GBuZCDfTC7n6YRlM+F76VhYymwVQBI75A0g1D3WUBnoS
cXSgIi18vPlRp1H/brz0ooZH+x2QhMd7izXyF9coGXlXKhD0UV5JtWEj6AQcBR62
NWCfiH1Cck6+OMAYcTLKojEwa2ErgWuy4cavQoP59w2HfxwwgqmG8reQEAxYs3Xf
Y2U+CxZ+Q/cNEAJoRNRYfpxMsJMRmg/jb/iq9rzQ4Iyv5VpgGEshJjXLWM2HUNyl
bvAZWG6nc60ijDoqOf+1TyT5JyqOJWq7JKqR2lYm0BqobDNGDT/KyWbPiOjA9opT
9x57rlmcWWdX+LMUUaJvxILNRJf3Z3ATNhF8GFBHATd/9AWtI8NfuFfrTLK6kujA
IcNjJhHIti3G2XRn2NesyeU5kd1r5nHeLm/XeeOABJnJoTjhN49QRgQxPn6NWKEh
fDlUdWqiaOF809tQTMAq9hGdQuJfepGBOm2SU277dj1GeLSaDeFbZVkMYFLZw8E4
vkgoRIgUwRgXMGxla51R2TZPO5NoHS8CZE4odhqrY+gOc+s0oqzKbgjFo0gHY8WD
iUAuiOoFFWCOxN4CuscbNoMXVljzpjT5ciLlq/I2ZTzd1Bw8SyoV/RlKbAZGbDEC
37cwqHWBRYwLSB7f+c6H0hESydH5/7wOWQwpyTA5qkYpsEEzsF2MfeTxFo94LioU
2+kLOdvJJxbQRUHbgrJX4MTgINPNE1QlHwd9wcCdeTfe64XRKGVTQKrKXRlmTLUs
0tRThr4RZX7JzEhvt7U/OXOfFO6AjWxNkyOEkXXnunaXmXw62zRQRha4BLSSKyOI
Iew+xoa4qCcvyYida16/zqYV0iCh/QtbUPl4hh47Tz4r+IblW+Z10of5+gvxTRdZ
HiHbbVA6WdVuxcHstJFnIbVDNcdWEBICjQQbGaasE8aYEiu5kNw62i3XuCdVfEWW
RrGGxViG2IlQUueGtlAkc8TFrS7gP3k+Gg5k9v7JpjgyMTi3OzW1L0ETzHslPMjd
IE2VlCzIcTxSNJrg6x06yQCyMpyWbXUKMoRrY8FIlKumEmRuPzvatZ74p7NpDLBJ
2de02WWXJyUlI1rfmDM9cLTHx7IBx7vwp1MKLwz+dVjTLJkQGcHcC8ue+ibl8ies
jqmX1uBxF7qnmwxX8p2Ih208PLsOD/Ti7yPKkfW9CbuZKfkw4Gt5GwPtA2HAshDE
pLve5ZZL4Nx98y9g80P3ETsFurqQ+4SH2Z7UrNj8P0ViP4+eyVsxyxfQa7N1RB3U
8/zhdxHmmI/09+PN5Sx7/FM/DugnvFh3Rnb8D/7wFQIzu/wdxGXwbTlRiy1eo0SW
ymVpGPK7puHd/ZAcaZWh/x9ICxHYmjKvA6el1dLVk38BT/V/D36nL7azjAOc30w5
XNjPgK40mZws7ksuh2tPZ+gJwblCox+RDpTBhM60RPE1BBDDTDRUbnImqHppW5UK
8DWxJ0R+dfPXUnPcf+qwbqTP3cgg7Mn+0rTvWcrjhLullD0Wu0gD3zaBJd2rFkMT
mS9Zz1+YEnZ5Q5EHNxEz8gRxUS78EWYjIa9jKmUVwcp+NVzKbEd11XczPECuCILK
LZbNdiYOoGOlsHDm7WnWuml16LEEVW9bmMbhUQmga0rqd3141DCZ/IEmZNX2g6R6
C8MfimRTrWx/7/Y342J8Mf9Jkd04qWW5zxRGsRvihfAiaCDMhxgzWkqDECjuUiUJ
miCpljJxOILyBgnl3ebfaLVFu6x5n3PVLuaGb3teAQ3m2uw6/H3jt5tuw9Bk/yT7
IWX11A3zGFQTaPMGDq+k+L8xHWty3lpDntAaI9PyWmDFew/OhO2FaPuJh7Ook2P5
tf9qx4LjgEttpB1eMeyFFs5qxjB1ojYq5hqz2dHa3fxtKk8DlYeHq6LEBBCqh8Tn
MmJEF/vUHIV7nmCdAoUl7Vwb44rxcgyyQp5QKWAW4q6BfwojWDX//B3rC0lfdXF7
pSqRuSZlXYUqUM/Zj32eG1AcvMhWndNG4x3CjFBf66ZM9CjnVmc0JBzOuO0yNddU
VqP3z517WIsbPLva5vaQ1CLs6kI2wqeFv9jPcSXYmI3awhHkgh26cobFSjJgoe1C
uL5OD1xmEuV1z494nA4PRz9byjnF9cD3tmCRj+P/cjcp/3sMyw2CwvD3S3x4vumQ
lUxbQ9gxUWwwcHILiUlWmia9DssvPG0m1XYwoCRmNSmADatioHnZr3zwO0GVKxFG
Flz2univ4hOKlywSK6jIpzEaeOTNjpPoTCg+M8mnp0VTs5fBhAdGROSPUXnBFcoW
nqZkh+N+soWSdii41TZxF0GjeUUWFDV3LDroyWYe/y5D4zkNk/O1E4O6Gztf3tKV
cpqBwb30KEpz/kwZEikddtuyDwzEJI4nEQqk2sfRx4zm24G3Z18OhRKQIfSXi2+B
/Ry2KxWaYmf+swogoyAbZ/My4VQuxGr7n4A/E07Xu3wrnHFQhfFurOPGZDZnWJa0
ZJDwvPA0evCyGtT/fzL8tAP5N+s/9tjyHvy5IKbzFi0LkzlkIQfx5NmO8juoOsMb
kHia3IFjek++frNqoqqDyjVGHTy6t/BMRnyK4RO2lSHiyo2n3aUDjehENr9L6htG
EtyzMBoSbw53Bycuo0eqzBSvwpM3Hpf4GPNE0p4Dt7tuU/kbBmTWa09o6VHWc2nv
qO1N1rDRJX3Q7eCdujDbaWmv7aai3/+3WPWAVIeClvg46ouLZGU/H5oiA7Cxj8qp
q4lWUrM1OPtW+n8JIaBH9f4YVUDn6yGaIt9zue63MkRLhJjTAJEXbXbSN3HNapRC
nQAsl3ITQzh2n9Is2k/CzWByolOKtJrbNHniHf3Tlcr+hSCAHKQNErVuhwGIXtWs
Eu5TEDmOrtgP33NdJ/aTvra1lzrIz9burdNn5jBt5KD8UpidY5XDuBk9RkQnXx3F
6oDHdo15oR6tpWGFRRGbj092Bq4ADSJMDM6qL5YeBlcciBZDsY72/jj6PXbqoXJx
5+S/FK70Fc7RnGy4Ay16AM7m7cjJL0CQuhiE/HTCZieONbLboNZjCvCYSFprqE7M
i6n2bfpkw1ZF/4ckBwmAgnOhkUlNLLGSejunKL6wx3iFYusBzXVwyKur//ie+TmJ
8crZsZQ3HF5JtDwAm2qCf6IKQ5Ef3BZkbMnjSQ8vC3uTahjZhIamRq+Psj3ZrV0W
FWXkD3+hq+ItJdFltCazbG5UT6eJZD2OOjEIHlN8qM+f2TkRWjnPNJlCbv2kSxso
1raNglO4G+4SiKLdeYgqKKoEAa+yaC9q2iOBJIMDTlZH+Qk++Gi3wA8DzZqR+AJk
W1zZshtGhCJkV+64D1DV5+FpeqEzHUoFV33C1K7r9YCo57OMHRiVhjbAeQcsAjtJ
8hFqpZ2nyXcQO7ceIs/+jByl7iQLxKIOOwzCPw+05XBMemErcJLUg9gVPCR7NNKx
Z0dwBE9cK7pY2vLVEFlSj8l8wVhIT9EMQvWtrd1NbbFN8OtXKvKv3zHV6k0DQGyx
2tGXCSqunHhMIq8d7JQCGB7VI5pMDfDn5yds6nfW3zQQSCBVRJkUIhfOeaLhmwmd
PczrU+TJVv6hVhDXM8cpvagOsMDvV8mnxVhUQBfFbk9ikUnlLOs7yVZV+0Uqss96
U3WrWohGrUxsext8a99BnlOYa90BJ3yDU7lL5ZQgdFei1TIXhOB7Z3+X1HMEkCvu
0TTw+6EfHzTML/L9gc3xIJY86RyEwK9VmXoR4vUFyu465ezAjj0mgasCkLId/Z/k
Ig3sVKzspjkYa+3qui+/u6xIjpX5xcmJVY3nfgUNuQYTXmxVbOQ2hLZBcHq8KZS7
4xUQEDYMH9yx1YL48CYb7PmHVJEJK54PbwVMepEIqdGeRgizlHz7hbqXytdvsn6W
oN2cC0Kn3nGHO/jgaCvRrYv0DdwaxIORlps/Jgt2LAbGzfEpYYU3BBWWjgT0By+R
hgTAwI1gE7sMlOSJp00MmXfEt6kGsKZEZvxUbZmldZJdbmNH/Eh/aTFfbZEMGmmD
xWJZr7+xAs7rEWk65wWjXFCpmcSfCZtrMMXVE999X3bk9xV36nnuLoWSbfhCsWmk
tPaW1ECGRD4HYZzhi/+wYgsuTnzcRMQBxwRPLlpcghbTGHV5O0GZvLrcOXajIXxX
K0TxtlgKgVRX/hDh1YMc2VYgQERpyar+qt+jpe8n0d4f0llYoi9qgRwEle4D3Wwi
WEQpI9rAeg7ENLMiwaZe4eRURBA54HQS6w8E0p3UWSY+yz+qhyBCSte8ijLGbalP
zXxPE3UllA+yCAKIv77ourqWRmOkaO9yenY5LvqjgPFd1vAgcYR3FlYphDNVPCyY
Wuu/1Psxb4742f4kiu3bRA9kl8OHa55mKzOSlF36zKNkB2dOt9aP45a3HdTXZ9N+
ZMhVZKjgEnvYkrbyYIAzv9fjXROl8kNslyG6FUDBwijXl1F9nKvMNy/pO8Pb6gO8
d1bHam4jCvWgmbYpRZBkRdiHcB13kggwVEjr3nIg7bxpTQctJRt6TXaE1q0kL2z3
g1h+uKeiuqjbZ0ypgl3D8QBtbjI0CTFyS6jbRGBRHFM7rUXlF9sz2o7FQZ89wmD/
zMWoox35LvwiDO9ZSvTF9G5vjli/r3sAw/mZuPgky2ijBXesUShc5hdIFI9rKf+2
Pj0w3JN8iW2PIOXFbIu1aOOjWRPzliGnlhLPpc3ugPW+l46YnuRpWoKF0HwhLezt
UU6jzIrmRR+8omYpiFUxlZA20C/uz7n8BQBgEKSfqgdvkZekcNadODdbVbzKJo4N
BMzXTMMPYjrAsxtlnBgA/++4hplnafGX6stZAx1x9T//FtTXkOmM/SeA09k4gwWv
WYt33i4HtAMjzlWP8PcJreYh3rnLB9jffNY95lcXN4ECRaI3EEE4Y4B0sPOzdrXc
DEiZKOLUD+yDsfPlIYF3j/g9nXJwjhoZQcxfhZlShCC64seADpumGPXTZ3jRG8Hf
lvc4bxyoyyIsOyXNcYS2ryOzlyu4xl+wUuln/VJXjx3sejZXg41L62zRsfDRxvF4
mv2GdI4teca3rlBcaeOXHbJ+ABONqqY8jHcpQDQ5Z3u2u1IkF5JgHAWU3m2TYVpm
28+ZZX5unK/LBdTr7M49TJcc5yb5LVNflKrc4s3TBbNhhZBUAfmi7GcvPK8WS2D9
DTxfwDlvI9VgJBdeFVc1IOOO5mkC8iAYgFXuqv781mWjGewbCBKBnJXPTj4N4SCK
B7FP8fOQUIqg0qHMWWlinWX0yhcQlpE3z7Bfu20YTOFfx9SyzyfsYbEJ0GlfsnUg
NzE4qDlaYNN7jrIAV4usNiIKZMQqLrrQFawp1A2uGfevO2E97dkbi5X6sYhvTQXu
WdzOGTaWLWxAOQfcJcosPDo9FXys+3BhXg6eIA7TP3eSfr5MbDngaeSRkUAaWuYd
f6WBXs5K8zcuFrsjX4ucsmVZiAFd5K+WOs4eAQA37XDLEQ++cCjv+t2gLRgeKyc6
RWZS8AVDNAq9dZ7HFExqsOhHIXluqLhee7aFBjkZHMUpsOgua8clAJe57u3dEOJ9
tJ3uXLBl6FcYq77lm1tI6EalS78Sk2Or1Vjofk/mWPGQwmsu3vlBy3YTa0cDU1l/
g1oW6+h4Oz4xgJcHPJzOewFHynuaTf2ahG+kUKZSiTJe4MSzLnlOTT7xcmjGXTBC
Nz6TYBvRHZGKkB68EBPioBRt4NfQsjm9j++xXTW8W6fXJz6Vh2u5+tJsYod5nztJ
sAkFoQW+rfCGOIGkUV/HLPpG9Imz7g8atbsdDPmGOoFxWXWLB3k8xhTgEnLwdH6H
GxTMZHcX5NGrW4V4103KqIXDo3cTgv9/y4LR3779xOnoZ5SaEHWh7nayt3QVI4ZD
cAuUOL636qKMRC0VpkyQQTzZIClID1VHr+HVmGA136V5R0uRWsXHkH7y753d+Bkh
hchkXgKbAH61+C3TWoo+go6wUmuJbEdjaiVmN5GMQR/SXO+VBqkAlPPjKExhjX/2
K0T0vuPoOiC5qVEkOmvVB8imkVirRDbmekohz21Oi0+/P5H869R0YjK3HcTw7UF+
e8u9gXR0gbF5BEOMw32sNJljxQDSLA5JGfTudN33+H79qfXEwrzJ4Mpy8GEC9sYM
i8GU5JcKT1BYbSYocmy9m9A40R+2iNveNBk7AhM9d53Vn4n9Bfdr/laGwmzz0CIe
PCLPuO2RVjTey0yKg9tOJ7y5oIsnItkF0ArYXb962O/nBq9913TT8wDFfXrSIYsW
1YoFl3VitcrzT28jX1k6kWhUg/u3BEV+XBlsJVF7Xc3P1ruzvVciXldzj0i1djc5
fPtdtOLR8XfiVbSfg7x8Sb4Yng6tNTBiHIUE6mhh0Q2zJ8WtvdCpCKbv4gyx/sWB
OSMPVsW7qmJWbEcuRZj3sLZPqkrLUbWIoagUY877Nl1HySIZgQBdRbdzxhlRCS5T
t9UBOPx48S9I9PcJK1J1gfJ7hOEpRSK3U4Mcc9rG33sAS3iW/KDF+f83iq3cayU3
rGAjrPIUN+flmYUG9TBv5KOyU2VwGY4i6ZNO41aXaMmzkth3Pr6FYWdUNjN3maDe
50CUlCpTPmbIaQ54fAAftBnaWpGRsa+a8QaJUfKS7dzOrUFFcJpaHXZYZN/1hDmq
Mh8jQpED4yLgS1yFkfNAcaEUylDjyJMIrDBh8nJ/1JoqOrdirwxMldpiJ2pwmo7m
Rfja3PB/2dWxCb5ISzZihVxDPhjd36zjuqyD99Z7CFgNMhI45xGuoAIw4kKgUZTa
ojzp5LeEvliIEQhssEa6ZO8Gzh07k210kh7Xdbx6iZrMRbVa4NIp3GXksDljwjBr
nsrmilYc/loQE16dWthVFQKyXBznlLXHiixObjpArP6YgQBS3e2mrtyunLIKN4bN
dy7uwJi6vs+uFzW3fLCQ6SN+RDI5P+doKFoOdzBQJ1iatSc4vnNk4sRuRhT4PZ5u
c7wU9oPGVsCeLnoCb+3XbNJ/sIjemhh0yeQ28mblbxtX0nqvhxWeBh9JwtxyijcV
nYEjJO5A6IajvmTThnEI7zWIfTOEqj4cDwkUWqHHkwQeQ4LYu4gC0hITT+iVG9Ge
OxI7tEzb/Bw4yW2kUa0sYObCgmZWK9rCGZPiKoKARossyOm1ICWhALA4jsk024cF
japvjLQBjMvQqt5+20yJgOvf7D+0KCpWEMDKrYWVV4p6ZHHKtf5A1T6SGkO2GZYd
G5kRoQsBvJdc5LwkWkIU0Tjo2fvfDSwsBtLAisDudIDI33Uw+zm0o72tI7Ix2ca9
I3DLu46yKRtW2aAntJclVUDaDdFAbr+AYM83+goTqFj+SV2srUKfCoz+aZ/ncW5S
7CVFBdKT9SlK6dqQt+G2v+u3uBSuR3ZdkPWLgAoLwam7VYsoT75fkWhEUt1G77O5
YwbXVpRZzueE9xOOlA2Cq4zjDTkX4k+xLDutmoYLWVcJ0qPeSdk8wqORDDOnEWyQ
siLPoljyXKoBIaJ6AbGuKBe5mSWCcOj2JkHm8zyUVnmtXsN6zq3tHhYC6A9l08ee
lsimNuN/vQUF/Ug1VVu/4F+rvx6xWdgd2nq2gTJ+jIGjbZ3GHasTnb8qE3pmVOh6
JTqzmJQCeV5SXPtBpWNvwOfE+2taq9B5ogAAJ5XuqpGK3+XjUvJYmUuc54KKLLIH
4Z2PSvWGD02oPGDHc2RSoAsLNnHf77h4rczRRBU0AQqEVx2WnXk/S+u8Nh05me5V
FuQfQ2bLWvlAOsSu/YpRR1+Ebw/XL2Kh/0/n1pt3e0tBcDCaXZtVw0ZDEsijySci
CNKydLe9b7YXeCKxs33CtlkfLNXXeaA0gvvY/27MIB+cXkZuIycUkoAHgKz3Q0Ly
6pqhR5dAhI4nh0D+iR2XIFDF+rEEeXJ+b4jJzu44tYdgIBSVASF4wiOPGpoaDNb6
boNvYj7J7Iqz+YPegGIR4NlZi4c1TJB6ZJ9B+YpSIEmBCDKaw+MWUBiYrIAoCxSm
euCaLFwfDnPLBFesWYnclLr2pyXH4mizoaKhrDrb5CRLu5A0B6pf+kBp57ZQ8wia
Tvz2Sp/Zr4u/Vve/3Z/UEpAD6+/vmZRL60rSjgW1hoPRsSdFm23K1sJibydrfVgd
3IkqPM7Dz49iZJUZ8qTxnjBtDfbTtqwjMWImzfjM5xfI+TXYmH3yMFtQKZlDwSam
2OJOFtE0188BSLGBOlLdFV4d0Sf6V21NPxD3HDlxUubVPZEl/GkaQJJESYN9JBpC
K9mrGcTtXCmzee0yWeQwPKlym42dZghcoUUAkg1PHQ4RyMmH7ektzG09V+c/Sn4D
zAmR/u50vuyXQB2gzvyxAdjiEs5zSZ9mpHBCumDejPB40bw9hC1ddRx2PV9/PRKq
HF2qFgL7tSGdEZL43aKXAGzfu9iR6qn/YL5QSYA24MRntAXaI2X7ekg6vZMpNq1G
OOUBLwxSbLNbzD8wpULQoOSD7Hm6qkpAKUMsG1TM9IILR5AOvn0HVcpMJNHANCIa
GMVF2s9wZ8ZueVp3W+M/tAAEeU8wsZQWZMAPVM2Sxv1Cevc+g/IKYKUBADCfJCaj
m0lslH1xOisHx5AWT042bK4mgv8VoOLbr/49WFeMQZzB7EwKoHSjHyOp+Lmshf7t
gnTmWw2NiSu6LFoECa7AHt/BmQwILwkzS1kBGnsuCV1VBl8jbmSrqWkO/lccTDNZ
fyHwZq5CruYyPkKZwUR5+8/xjid68bXtEiiykdtYO1usSTManc7xJlUvJ2gPU9wV
/z/NO6XAz0jkXnNdJhPZgehJZxf8bKbK1Gq2190EBjljOisK3op+Pnpc5riUHTv0
Bovrlun+T2MeLnPcI2I082qV9y3XZ+UYEwsjO9aCUzKXOYRA1OW7sLdowWLlmwMK
6443S6WKGWgj+THz2nNEcjDG9m/M9OOJ+pRqhAILzR4dvHysU1uE0/1iLRMTWRiL
KABHGRZVNy9turwKVGMD5YpLqRRnGyZgmhO4rhPyvEIYTkn8xocsv9hAaNmN1Dv/
mbihetCg7WceP06lRdsHyWlOUr4pK9sbEbe+yLg/XXd3hcjObAGzV3IOVZ8rNR5U
jJCBDJ8i8APH4EGmDPTpukFL+bhNkzuNiuF8zSfx1oabaBkYKDPKWyfSbgYjKSDd
E18T92mFuBc55yKIitiR5h0nnQ/KY5tjaLP1lsvHQIytMBgGwyIE5/QIT4fzX3di
A83x6kzAXTmHa0GbeBFuiUm2PAVM0cEEde8j+gzIh4c/HDaMoyWm4BfRKKjxFNzl
MMZOgGIfhc5DjBjTPQvtsrUuPj49i+SDnmFWer7GzCJgDy/AZWPxB2q4m3O9k99u
JKmWGND7P8WfQxClyKik4ACQiYtmVZ/IoYLgdVl0/ivZvfjp8yViZJ6doIfflkrP
+BUrNyJYzyWjcRejf1tFA1i4BY7i5S521uZcrhL8VJYh0B5AititLf8MPiRCtDzL
EyGn990v13HjOz/K5lmUotCeGu7gKmSEgSUH67MrMQ1R6xQ+Gnc5gzWuohsxrQLF
hpKiyc6nGP2iOO3WoMsA9pvkXUPsaTlH4L7+AmVqhwBb57gpGOhetJf+RuDx5aoO
Maoid9lrJBIyCQ0JQgTD/ECAA8JU9j3MO7K6rZgr6KP+nwIOjDHUFMkwvgd7E68y
IVptqROtyvCoBVpeAwgvSczTnb04xHPnBHZaZq/grhOCKTQ4M6LIuSuZUlaiDJJ+
9imFcLg6TjLPgmRXGu5GnQzblQ0g4gsO+qZGpr7fYXSVy2ex/8JRre9l974zYRVv
vOujlVS28hXkghPnAasJ3TLDDOqBREaHX9mKNjncZev815IxZMh8L9V6SMRrGhYw
9MZr1LYB5lapIhv/YoarnjXSr0EqG+FzlZugwdpT1dWqmrCGzcJD3lmmRfxkIdkl
c0hjd6UxWVhNOFg1eLnbfkPqwUwFwTj+lTRaAHqFFtUg9DZIvftQELNbdakwM3PA
uQXwjwOcQTy15qPCZr+9jV82T89FBOrU1LB28qV+R6BVkJ/qvz9ZuxLNnUXqjLrU
x5atsqK3Y/aoEuWl3TDvp7bywfBnMB9rRMkKKJlI/PZRsxpBM7VWdcyphilXJqAZ
s3OR1PI85+4ar4ksuKOTKHbvBkgfWKZg8Vx9Ypza1DPeDOG1HizmlvRiDUXRXlbr
SbMKdzlwR30TUmUxOSHDr9P1cXezwi1DwO9ypmQZeEG1cCkC//jXxOtIJoIfuSvi
ua6+VHT8OqWLfCeLFNgnnfwphaap00GV06bCca48vOS+V1YTU1nWyLe/uNavx63S
Yw8/WUmKzJ0utYvpRApmt5fLtolVi/jt+zWTh3eWAOqThB8zbcwBATNMSG9Jljq+
vmqxweziLGdUdsTMoL6CsBjSEEUyJrREGs4zdtvjGaLWCY7gLICJHE0eqsCtJtYw
veSRZDOI9WbbUjThy6Gzdtucc3fMJk6GXOXkqA78FiG+W5169qTOo+BJ23bX247p
DRdNJO0SrhI7Xd7UJcJZWVSPiajK8f0W1weI4YlW6OosJiwQnjtXDQAhfybJFPhw
dMpFbUpNKEw5FDGl7uMPs6zn7d4HjizyLIXArpvit1U3n7aJlhUkARgfJPesikA2
g1DxMww2Ko/K8psKS9Vdhd42NcmUa5bg0eUWSpQRnyV+vxMZeTpJj+abjlwZ0y/3
X22c79iHuxeCQW6tJdXYuqEGoYeo2B7syRmEd1rWUtUcRIWYAA1qWnMq7AbNuYa7
cflf5GA22y+YgyHbWab1gC2KqtMpq9LJVdj76QHqZPIrjwAgA6XF6ZsIBay5sPHa
4q7AVZ00ML/bKwOHb3iJOo49aV3ajBksLyJCDD2q3gr+T+vENG/2AAmZWzKUxpi9
OXlLisQNEiMshD455INJD8oedxYZ3YyzPmB64p1rE8f3sz8sLbmpTtjVw4MOYlki
1R6CMP2fVb7iqZ1Zk4u9Ed2TsN5l0BAxA4SJt0xajFFiWuKiLJHKIPEi7J2dSsbL
aEX69CbZkATfCfmHnKTL1CbOVRXzxbaDh1YKRRQLv+V78OqowkBg0t7MPAvzwiTT
nMRV0854BiDoI+2cbubN0SfQdGJ2Yq7MNzeYQVO++QngOja9eAISideu9A2heis4
ReQwaoXRVqZSUxyOs3ftgDCoiPRKDxOoWXowfskDPboSX9eFIjyHPJPcahE2cvZW
sswye1BDdOZcg1wItguRnZmas8ma56b859e1zc44a8GiNdpRb0woci5WZnWjXJ0T
/IwIk8i7yIGFGHC+5hpPYo6RlBYgotFXCHJEpY9iw4F4yLIGCl5lMjs07KU9blLp
HhGhN5e08aMKoud4ZW2gvDzcvcK7r+AyqeV/yykZFQ1GeiQTxpLvUZsgLpfonldu
ipmBMjIovWrFwo8LJ5HZpZiRaxbglQcNvJMM+ihHiKf0ad16VNtITIhECILrp0Y+
CemOBV+Ym8dFQrgLh/aNkxqIGxF9r5pPSRjleMVDsESd2v6q9Z22U3Pa3mNWHwlJ
fxlqRhEFGD4s8Y99N8oRLKdLO+WJoiPEOAPq6Qszk+RF73UBx0609sF47Iq87BjT
G3Nh8zrxOHRuL732wV9dvbuelIoB5qWaCY6fjgJaqb+5IHip/JN4dZub9+h0+oK+
1FRrv/+HAQCzVQbHRcI5zRj3xteMhanCV4rEXmultFezTE62oCFyRpPvwrYlHGG8
jFrK3CeysYbPSsuLvIealci/8w8Wia1tPsPNqqBAxOrDjWZYe4g9DPVyNvhR8CyV
Qlg9nOodmv5W8SCh2USBoaRXUlzPubdhUsaUh7xB1dlimDPJyn5UFs31Y59xAFc6
hUaWuxqLR1gQf7IIcyRk3mlmjsF0My8Scv/lDuJZQ5SKdt+Kan+CtTzpQjTudps0
xqJwt9E+/p7C3++kkQZGx8rg8q8NBdqEa2fCf9unG+D++1fI4HgC42rE5Id5WxkL
zZhB+2M7NV/1AhFE6sRpE2RqgVaEOLZwBgftwfyvOORkYYSFu8fXZbcYsgUawKcW
3pezRoJ2NbRFr17EkRR/pgEUFzb3HRCt3slykusWT78be4pzR94nUWMae393Ebhm
KAqJ0GVU2Ez/DcEFeYJqou6az5JoGLWnfPlvw4DawJ7diFqs6EwlPdJ2hz4JxFNo
0RH4uCTTxMXOaln6KpMbSwlzm7ypYRebSy6DrV2S7xIqcYWXhX9WKVAMRtmMOp0K
gAFNXyC/BqDWz/oiVaG37JZI787BXIrYeqJkSBU5P8jZg9RqeelxfY9bUJ+5NsAG
+q5EEo8Yd44XVpW4AGeITsq7fZZ3z20mgp6jcwVepCbGFgwIvv3gvPgJdMMpzT8h
DMUjvDd2zL68oh9XnY1OTjb2im3Aw9n4eB53TaBBA1uVNTXmQEC/VwfgJ/9/FAiE
zM+/UvC4DnaQ/goJg6+YagGwva0tfRE8gd59arTuUd2bODUoW9kRCOkE7D7ohIcc
OTav3uMGFfCFtRhy7RstnE6KBEn+OnbAhoZMRY2gDbZ7gA4UGXjX6m3L/KUfUIvc
C7BNbdS966lhd19/Ui1gvlxAXtGMX+IcFAk5A5HDKua0xxcBDG/Xj9mgpfIe86Rf
7yjhJnl+pW6UEHN5+JXpodWWq/5B/65IbPPvWyTMCe/or7gl2i4TDulALIdHzGyO
WPpt3+UiQX+yeMoxYgFmTtBoWCeeY9qBZiF7YVmj62yFNCLpUj8frUf86qHJEQAw
YEvfosf25OyiRlH4LAEhYcIF4HUO2uZEMlpZiVa467YZMVUF4Ru1zjwMS9RsKpM5
rE3o7UoDbcjv+RlmLghSianW00OUt9eqoGRcgBqV6fUGzI02uFssOvs0Q8ka+9rq
CTtbL8Oha5lt258rDminHpnItQeonQKLF9hUYAavUPxfd1A1Jsmm7Tt8uALK6WLt
tskIMZai6XRm9AaJwsjg3lSOGIfIg4wdKe7ysJknNMnO32k5F2vovt1//y3KXcMb
kE9XUuWkrwyuRFdQFq21l9nhQzWVFyR0dP3gXswsxtmQjkiZJba+lleU9O+PwoBz
hswy98Gb2YyvYEVKpjUWBKvlnVgJwJLskVJ6hf+dI7foZWMQ2/j9r95+uPhu+nYr
Msm85XfKe4AUi5lj04KBFV90LlVjxSHF8yqIfJazuxzUTS2wuMOF6whU8eZ6ptqo
DaahWS/kzGMeKfsErm89cZ5Cn23gmLtNnXf9pUx+YR8JzJrEpTpygwKPN+in/AOr
fQKsL9mpNtBBMPXXZmUPXiI7fajZihMfVJIwB8lGDQnBa6bYy+qNjPQEfB79rqZZ
P8GauMYlq0AZ23qi8Z0bHRUyG5vKjuzysx9xxrUadK6fw4kr0V8iyDL9zv4nT5n6
Sv6ha5qbMDjf095c8lsKc+sAb43ZYsEQPxptatSKiZdLkbcXtQ1qL85z26g6KlM8
ZTUjs/lUFgam+mNuYcO8zj8thLjDxzrvnAG5DynTLEW8rkszpvm8aXz+c5HzCkhf
GQfGKL/qxLtxopvGsviViBpuY4CDQA0SGxMRHmsEHnFM8C6EC6EGF9jH2ItEgeES
CxEX+W+5RejuRF3xhyibjnfF8BO4zUjwi/41zjzYrmXj4ZE8X8Civ58P4gG+/45Y
syUFXp5DY1e6AiL7E9o3MRfvM+11cRscHbShPLOGJcMs1Bid8uYDxFECS4yu8aUv
J64ZDWlDTZ19md/2TqVg6KftLF8AJ+pTzwI61+HZcTqUBOZp6kBOz1pErIFNMUyT
CZtdtE0BapUeem8/xPwzwDgMyyggcnlOECS0B0cfv33JFKievLV9pxRy3PbSLz2a
mFZP0sJLFAbN5YA8ALSPAgbh6yy/XevVSs7Sbk7S5rGo7tWthQmjHIGiwt7piFmV
ixfgzqU4U5A2OHaqB8rvIbddFBa0Q2wCCyAxljTB4K98CRq/014bhsCC2FwCcUtd
isEtBG0kMNDQIp5RWHPy+lYXRKvRVthYoO3fOlL50kWMr+YQbVKO6wpjhoPyoxSz
xFm2Ph7+e44Rz3V20GQMmXGZLF92sS0dJqBhaGchq9wVzXUxD2e8jTgt3yM2aMxZ
vyU8hZDMQIqsEWgyWlMDSJx9Djh/mwzrUo4Q6wqIoX1AN7WbSdSDy840G+7s8C6+
irM48YIuInrH4ggRWEdrM+ngyvwRrgpea3ccOTvXkPxccefRSmGoSxHnMuhIo60A
Pjub6hGrFznOxtx/yC6zQwm7i+31ZrApD70PZ2ULnks1QIyY/7w1skZ1pmdLumjR
MT5ClA1yIjpY10i6JIO4eswUETvByMwrmbgtJwzV3RmW4G871hG0ICQQb10ppIdX
KvultzfcLf2kQ0yi+sjVtpTtYQJY2SGrX97sv59ILQolLaRZDmLyaXlq80Uy3QM0
CmA+ZPZ6tiWKeZPc8nup6sNVLsu5rdAKcc5yFdaPyAQwLXEng1Ij2gNe9UUQ3Cg5
NDUYt7nD0qY45VcpKNVrwAUL7oNupNW694WYPzQKGW/omU5mWXdLaL1kWy9UyVx4
yJne2mAaMLVCYKvGIZOniWCdYVlrLwaM3fc5qvvtd3dsinGwFVvS8XTZoXvzLAQR
SUlPLISFHMaECH3dx3sZ4m53lIRVDHrCgDX3/37WWy9OSJmP70LysHy2hEdnE/Eb
CFs/b+CGDADeIWKnGoMh23F+IWXu4r0BCP3tKysVOQqYjuvwyqZ8AWPkj4+21Qmm
fkg4btin4TZq3vFWtVBOpVZlMQaVUTJ17AqxWRtsrIvA+ajoaU2FU0eQRwvX5N0g
dYML+4Jt0fY+rObWvR3GspLRbTdrN2LO5yEIafPfJFUf5mapXrazAsrO2uC0A+nq
VQU0UX7rpiH5HAwG46kl+UvHCP0xcgIh6bcGhj7Nu+X3zidMbVjx2zHWCbQA2Yxo
TCMf2t97/SoOSxmyTTsHAhTRURiNqQjSWUoYIqnDPBC4WKSK31tuGPzpZXZAm9dN
lImhYh982jmg3PzMl4SrvZ279jr3iOmsmfYk/9W9/CHBP13t3VhrRRu7Mn+u80YT
iCK7xdA40a/huhAIPQuY7XyuSnU5gXlTTXioymiIkbjJSgk2e2dXkhTHUlfrJIJw
BNHw/3NQYiXrT19iknWI6AOXj2klSiOryYg6zFHkHFYxGvUKVFLN2GhD6FZtatj4
zNvchbrHjMNM0qOFNQVxGsW03SlZhWl3J//tcm2Z1bF/PBuUIm6tGBpVEjrqYf8B
vjqiRWIJLp1ag/KYiD2Hj51PCHoABGjxjyNL77+TxhuospmitWZvkjdrYEM/ZETI
ZvQZbBndGCH6r5Rgm0DIgBjCI/DcBWz4EWkZ2R9D4DtGj5HOvzNUM5OntBJy43L+
1ReYGxpmKFZWAbv7EF5eXeCpeX+IEbvZevzd6qwd7PdV7CO+hddsUe0W09jZdFVK
n4pSEWkqmYwH5NEPniqgTKqh4ayp7qWj0Ib3rqeQuAw9ckhK7EzQ58c604lP4R67
o6CFbYqUCbVFlyWCHfpbc3LIKNx5nf5eub/1nDI5Ot80Jnzk9gdDoCGEBr2HbeP/
uaokn4nX8rVGnvWMTsBLstDt2YaU6lgfJUFQQvaww4djwhuKoUL76d4EHz3BPiym
HYABp2XCoN0o/2zHfpHUzHg0gIRgZQSSShP4Dk74vQMYzyxA3gTgRmmZTD/ST/tK
PMKd4z5a2cY5Cf2feuD0ncp+zLhA2lyze5NvXhozsEpMQQMyquVYK83413h7TC5Z
a1+E2QRF2CJwwXJGAOcuKcF/RmONKl8beI1tOvptNyIG1fTP6aO6apgc4uJRASvj
eeivbVHKSAyxohH46XBybtimr938AwS/Qj0+4XJ0Tl6W54DTDB81E00vPhT/5UfA
ljbYc8cu9dG6Ni6wKiodWAHm/MwWaHLRWytwuVI0kweLPM6fTstNCCR/fiWxD/R0
PaOFALfk6Yc3EFBi+JfdXghcNkjJLlJSo7N+AHalcL3I9v1egdZ92Kpy2gAdLdvu
eNsmCoZ6GbpPWNYm+kibcKpQhebREO/g0s3vm6TXv1UpuD6Krte/kIjBzcWvESdJ
kQ7Z3rJmEevIm1Yv2XGAfqlsBjMllVF7iT9+sss8hCGrW1bfx3ALoMRsqry7lNS4
kK3pGzlH/ViF/E2vURdv+zRtlDPYRBetkmKx7+po2vdTsD3zidJDtcbUH9WI0koU
T0+8WsYr/z/Rcmt2YzXlpa2rwvlt5YEmCwrKMq/yHh7gTPJTpcEb2YMq91xpsfPZ
62pNgs9Zmn0YH0T3i/H4F3bmIKXdSsLPcdYPAQ4kBzqO0b5t2gP0Hp1wCMc06o8X
5lX/Mc9i3lgUgVyfZBAxws9tqA9ZiuaRIjI5nJIL+ZTNKEYEOpa8ANASOKop624n
CCQhPrXIBaihWkTygIk560doLtj2nqztSMtn3lAKFg8V4gZnOc45+C/5qBGBl8lm
YIDUF2AeDSqM47F5TXwmk92/dne6VxYrc02AtpqP8Hqlxj+MDB9P+ls6Hl7MVJvx
sr59XGq8w4jRfremLvxftsWUfT4FheV0CnPhiaziFqOSJ2jU66odNoyr+3m/ABJv
wVnmO6ojYod0zlZllb+/Wd5vFIN1aOID23xLzDrc80mfNaARRHlsZ/NvmcdZGAfC
6NshL11I9mtl1R1tSxznVs92Adp/R9+TimmzQCrtxHiq2vRIF90U166Uzd2yq5eg
+Av/A1cJZEy5KHNVVdafZ+YdD8zQ3gEJldzGN8HrT51k3DLkIvKcBw/PWiZoKZOY
oKn/T4QXvFEiYYS+w3fJ+lv/sxcLZQHyMHitljMts6SJ1n56jyI+hBK7AFedimis
YMfv3dxx0WZ3IZe/Gy2/HUrqoKVvWDXbxkWMDAvlYOOnKxxnuXruHA2LkmazCrG9
vv18MR+6XDpCy0I/S7xMLs2I8+2rTxfr71KjnTCnpRuo+B3TZOPWbHPNX2kkSajn
tvA5nxemyPDHmtPipH7QBCQ586HmVha3zRn1Wq4N6DaCK8V4JaValNDeT9iAPIkH
kccdz+hSXgfO42o0ThgvZBGMfUZFqj3kYHyQs+n5lHERWY/0uOXSmRSo+ZbVB3dL
4H9h4b9k2/pM6DbalZG/Y3Y5SR3NgKVliG1WsERZt/35ngi4OKBA6SZydC2imKg4
Oo57jvkWZz7A0vF1VINZ6Myy2fTzMHPCbF/9kT0PMhOohRr2poPsj6/aq3TrHH/U
ODY+nEPkHHbMyamXwvM+/Lcu9jHN0NWHOsBuT/Cq/4/WR/OC4N4FQPbQq1x99OlI
FHfvqJgXQcKxYqldmPTyXaruO/6b1Zy3tI9lXaH6/NH8yuLkHrhP1V4h5PiZwS68
Vcy+futfv3YcTCQ88/4xA72hnIxpuKbdHvq+DtbUsILrx3agzlP/6Gi8WtaMCheb
qX2jkFhAyfWMdXF/DYFx77dPPtVEE6aEVqGoREaZufHsHkZndCQy1efpOnAIAjDG
ELBymthRQuiKwLLzBt6+pN1kPjhR4AoZhZ2EiRvaTObcA9wJHeqGFfR0Ad4+bj68
6fVPtusS2PxYNdFn156zj7l/efxZkbCiZ7tURHgPiZAYIfZWVdzMxEBTWIgVgB7a
w2MAxjDDqE8Vuh0HyIhIa29IRTKcgBS/BCsLg7tWexmp/LSlEvBPclGBEEO67Xp/
tvF5wGE9MDPtm2P9hyEN+NJIZsngFuVhHMVv7/kF8tXgg0gpngBWImDV7+LoVjbM
gS29mTFD6Qv2NDDcrBfd65L5pe3Sg3i23IbsPAy5YCImRR6cCU5ozClXLXrgaxq9
IYq3LqZTQvJ5rWVhIS17YgQp8nbIrrcuuvQZcMsQjxpsfJSTvk7GrLY/yv+SMmVi
Iza7LQL+BllfaNZLtGh17aTYyIxfa0ZpaLYC7SFwQeywen/OztMcZxW7lhoLtrt8
A+KaWChGnSLdpF/ljxNQCRrT3q4bEz7K803sO1XbIeM0/jPXmtWdt+1GNysFPV00
15GbSg4xxTuBmaPv9vdAEgN28RTFtgePW7J6ztoeZjBmCmtMYYL+Fv6p0SBvJc0B
Mxkhh6F+FCkwfjqxKQxoe+3FLiFJnkk7bS6hAfwdFbxzhRNa7aMTIsjdfe+32GRa
NhuitTXc/TJH4AKsNkmiBrXRClkb8KfBKO18QM9E08NXnPigqNYXze3k6sGcGhbM
WVLbsMfSEe+8yWLsIf3TKVGppjcCMSC7izhfIrUmgAK/eAfFX+xxfqCPf1Xpx4jf
yG988u7JJASpr8TXj2jFq2q0kKAX4DdKiM2c/bvofM2w9PxHhkc5utLTUpQIUSsX
xiTNeZ8J+u7i7WR2KKv7lg7b7UXxj8H24S8FimNTT5m7vTjzaLzogKhS2aTZTE3U
2CJJ2jN8kVV9MimC30EkD6VfSgSOaGxoStwvwT+cbgNCsbcHV3dwgaRTDHvEGT7t
NQulAO9UkZLRRzEVHRDE+mN213ZCfSAbIxvDD412WyfDgA9+8aMCPtxFoOoHHUzC
pgbppyjzpNPjP/OFGneWJL64TmsUKFCXP0sdA0C6TEBOryZsEypp3d2GixZKuh2f
ysPBLqig3ZhNqg/LnJUybEFC9T7hmiQzdWSGkw+UXWZZqOXCOskxEdIvQ4zzaJJG
bZSyXrLipMiVboB9hB8Hlxz0j462IVsI096hgaHm+BX4cAYmjnG24X+zV1qCEBfz
VyPIFQsWAPqwHCKPBnBb48lAimX8tjuS/50pOykodiQgTrr7ajbEoLtVC7dBhTuK
yzvn8wn6GgKj4OVHOLTo90VNI4bWYST156m1Gwv/6cT9hxDfS2f8ruUKwYOguP7O
favaAIEKMLqNZOcSfGmvOyIKEIKa4glzJlAgCqoZJcSEA4rkmDi3vKm5ld/1Jikn
uIWmNHfqieibfrs/5oa2wKF3RXXZbowF7xjy8z73OPqI2S+V06+eheQwOhQJ2RRY
fs1+v6ihH+8gbRuZTh0tz2uQS+mk5QjL6M/pfP3HF9taI3j/ov0goITxDDY6Zqdw
GRBC7pENyMjEAZ99vYDkZ+++neT2la01kEZNmsFloF2s/ZjPo9l6JhQKTtji7yjU
ixXEbFteCkYbUF7LgaIR5s2hEZob3EZPVDtmWYEWwG9aK5bJ7hqlv+YvJCaObe17
TWGcJ7CTFJ36UCyUVMB0L3OoElPouIulAm8tc/HX52avzxMdKYMP3FWjRzy+Aj6Y
9WSk3BeSatXLA/FlOm9/sUqLRKMgtjfQfFMn9mlN8BccYG5RUAe+C/1L5agEyEw/
xPsfJgd0AN3SEGg3o9eJBLAComCbjq/AkChrJd0+1bXjwuv2fYbM8y7pqvmK1gPP
Dd6e2CPxGDRkl76mDKHNBpdB9FH+IDuEEriHX/1EUZfk55kAWlDB/XfwgfgB2rFK
vo0PsuI06a4vGFsfVU8/PVrW1vmA6og0WREPf/OgRx/IhSlOCao0Pmx3nbV8Kei2
M3dFbkfOFQvW7Wr4pvxYVwiAuLAiLvBi0/uG0nNBW0a+TW9SM1iNzBRhG6WmjAsV
q6jyteWSd6ZqirHuVG5xqh27z4kjk6aVJINPb6poFZYvv7KEnRhpIHwVZqEIZkFl
FSw0qTHwp4vKvvGzGyE7awbJtf9Qfs7MSYO5+wH0myR09vRZj+SvE6tAJQ0J1PoR
rhNuxknhWwI2tteY9XFSSu2UptkocDyQBshl5M0qCyQm7ERy8DdW8j64QSaugwkV
bZrvw94vUGUuYlgSVe6S1LWZ/+DUpQM3wD6Ra8qN7VE/hsyTAO6MC1XiXz4L0uSz
`pragma protect end_protected

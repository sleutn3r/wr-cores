// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M0Yjsi9bLHt7juXJUeOI7F0+9WmpgFsM/FdZGvxkH49RRlR2fyMjEnccmbznOnu6
NHnNz/WRHghgfNc59pVLuYICWuZ+xxjXP7fXLpuGw5xJdGObINOtQ1j5+owOPp3+
trnAtxWW/WhGSbsuUU5SmMgKVh3HlHTVdXjHCAmL7MY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7088)
Ly//o3VxLSk72bM8C8lt/kxwIvr3qrW7bmJOF+C0Kn4LJC46DlhmPqYDLt/JTQaT
v16LnI9kYRcu9BX7uQ4mYx1GMI1U/QxZR+4hszZJOzRN16uOrCRYks/vYRIXYjfP
36gYrw5s3NJxVNNOtCMUkePj1xo/DsvOOwtnVXKFPOQvpkyZSqDD5xKm/KBIB94J
z47PJSjQKwN8LQdSXYNLv5/f74yvHVULtU4wUt7MDY08MKM6Avc5+rW5FUwccyJK
iOPI5gaZ4A9K2qhiN5yfMT+IQM/nh2VHtnnGCP5gth7uC9taiXsLweAEHlC41kQn
jyRQqjFmgUVM0/JxcncpghQfLA2h4X1VUWi9sJue6ew3ZroAdm7nLbtSg6rR4xSS
IvVENWVeQo4vYyv6NfEHxms5msU5yBfoIqA5W1sF7EVWFj9x7E0CLG72IXdAMRk7
PaGasc9/Sh/EWXzZlExfZlUt/9QvwQkzETk32ynZ6STeZp04C1KxmQKcqIet89MF
I5uMxsnmFaKwaaVhI2qTrM0iLM/Cxyohlu0sbCw3x9UaWjhMhVZ1CAezo59+0QvH
RpOxpVNYpLzko8y3MTOJ57dnNLcwzlB7jtplJ5yulEQIoQppSxhiC0oeCCnDPS+X
BRXmvwRcS3jdIgjJvvOLZSI31+SDQ4J7YOM4Jxob5ffPCh+YKBcQpegeLucYBuy9
Gc0E+ILeZ0Cy7oMhCEm8dHy7KJwuRjhXFBdGiVxTcQ3cVZko8zGiHzBkbxjUzIrg
X7eRD1WwwSic9j7sGNWGSBEhzB6/YTVrPvzwUV8qbyk1uYbZXOF5EFLyYu3oeq7e
kwS/UADXpdPCmrYLkCXAA2kIGk+g56UWt8x2/dkFwsKtuAaM6a9SFYqpf21DcKSM
vZIQj+q1vjkgixqhgGbTPjwnCepKnQFW8gv5QTreSGNWtr+f5twJ/6i/asfphQXC
wQ0VcOoy4ze/KbKmvdQqIgzil4gzlNvXKcYMNJ2LdRvEi51cbfN4R/yNy3oUTmhy
rRVjMcSbW9CSTJ4slEtal33m4apeBYZ6ffbOYvp5NYsRO+qli6qudExRxXrxmXy7
olKZRqOB5loRDxmq/tMocz9IF6LCpvYvQaDlOhLf3qHdLnVM72CWjlIEWDvmwUDw
yqLFa4p3cMdwpVgfXY/IT788cd+xrV7dM+elEi9RmbfjFQPdSijXS+WQ1LDoTdmr
h4tgDWkkJcaov9H4b9OHQhdr7xI2fdEPQIpaI1eQb0FyUWpq6uXlUqnMkIr008eo
vo3gicffzNyeXZfpro737xzYjGwk7dEEDoKd2fbGId0AI7kPAm/oxe64Pv5d/l2w
+n0uepXznLunk5U01TFMv9trLPrmYj4ih9IizQGRTB1T2SJBGhq0U4uXVkufLnn6
UcjqC4auErLsFYO+n8XebXtp1ImNpd3cG2EaYJ4ASnWpHL38HJsfIKz4br5kgrFb
vUAQRq0mixkE7yB8G+uGLKSERRliKCcp9DEU7k86Hsz4nMIrvtIE4VorWdeSj7zt
H/i/9nhVfFHCEcmFHmMqnb3SWVLRzysUzYfElsEnmTSz6Bx5eUDy2CvZ8JnNtYcQ
Dmy1+cDH7O0xOSF0SBzSHBh5gQ4NFb5j+DlsUmrRVOewAXukpaCqisH1ensFxGFd
OQOYGOsbGpmrdzTtGfyi/128eQxqf1PdUNTovl2eAZK0/g2mkw8Qi+OUoU0TKkdA
WaSol5OPDf35+6dzQlOBLK2PxACzc36+2KQElrbFRj4ULh3DeMswrEFlOphq1TBu
UtZjGw9pa1vOCaFvRpeJtM37r2wTW83hAwuqa0wbn171yarEqH9W4Uv9skH2QPW2
5nAxOmpwifYiac5OZrTA5vyse1UBaK1yaANKwNI2RrcffPGdz6VtBklZYeT5GFr4
URF1RMP8cAK7Fz8GElskdLk5GhEwWraZrRCPDdrUGPp3TEkxKfyy2J4tVuZtIaHS
ofZqM91qOLQ2KHVPI3FWagYLhiQ+uCfeVA57dyoLyce9p9gMrDtHjJep6nEmWlUr
7cRzb5CZz4CymdZOD+qBCxSCPvVzdMXnGB3NIufzrCl7yuNCPrL19PkOg8pgL4XS
51aQsRMn3b8vsY7vz0G5mv7QFRjSwGXeSQfj/Yc2BHBeLB2dA3scSE8LQK3eh0pe
kfoQjMuYYe+cC3Z6vCCRNq35Z00OZLBnVCFIsoAFM5er2iaN3oBgsbYAAd+p6dyh
Woh+qFUWQ+ExOd5h0vR0qL0rx/ex5vrExz7T1APjombfTbf0VaIgGYoRmwMIPyLg
JHMNrRrdxtXmvEA5FuoGBwssVZ+tdb3o4ocN3/G55vvpik+HRCdzpCPOGF+tmBu1
PKmsuESlnohuIL5aAPnN8xDJA0lhh1RH8LYlDbm7071qG+CBeIAHSNOgIYEX/+LW
L/nzJSKzuj5fLQ6Oouu/L76xASSc4Fd7sMwyR26/XRPtJudx6pOOSluhHW+VjlOx
9dYDnea5t00DLIR7Ep305YsH35DQ7+bWI2gWxNJZzduOAG8OXNnMV9MIgV5Bf7ai
sHGr+ccDsAhWMWUeqCsyz4FGXgXgq/JCCyjCs87ZDDmmjQ3CasPJFDf3Xs9Zh42Q
8QAOkjY50REKh5L/sMgOB/tzDCs669a3w7NvCV3Dj2gry2lf1iBJTnckUsDkrvzB
RNKwOemyUvZxgy/AWArh67KRnkMsTBtEeVh8hg9Bksm48QWt8XG3X1Y9RbPgL5od
WUczL8VvFQE4ENGmX3budKg8GMo79llbuBwtdifALGfjw549pdC8UMGjuQLoiAUx
w5LAJgTd28mCMWRVnDGWNzO5Z/Sfxy3ITdRMcDl+I5uIdQHGppUNWO5r0lNBX5Gn
kn/JChruFCE87KAsFkQSzCxHOV6OihG8uq1v3KMQiDdBaLryxea42ET2gh7B9FWc
jMVA8hANg2/NLoP9yTrowfwh3X8dSf+2ZcTpcQKVKN9TxyuNn22pm6ATOSgvYv6W
u+OGUnnv3huUwcZT3TOF4XsjuHAgTTQqUNHW/Z1v0MCGH8uYi2x5yKzCRAiQSq8D
v4d7ZgDrZa4EnMKkGANF/2NuLaWFmQQXnu9iIdg+Ksf6pszkX9xq0i94SD9ZEIym
69h8QLHWJkvE0hJWUd2k0I8rrXm2vM8a3LrvqpcbTRxoAIxt4HFoKDOBqgr9UCsy
cKxZrYLa/KpKCIa/enguHwYJf+YZjpkyWLZNi7B1BMmdCjoS3vp3hSqc7GBWlSDZ
HYgce4cEL7EqJdaXVuUwR4Sizm51tjmqQ1HB0yiCYNgNZwuwc/pz9Zo7wq9KshOF
dPyqnc+PVfKADmM2Gpkf7XWgb91nSh13qBomSCjiEoIAsjrhpTJhrV1eatK6KufN
KR7OTqs95vJL4sN5om+fUtvjObkddtPtMlV54bbfHvutxpp8wcNIYhCi5UBkKQuY
fdrYjR5nkyl5pR3a959J0eGwVIwTze5E9UPEf9QbAsewxPlSMd4HfU51MxRqtcAS
Y6mVkSW6OpSMQVczVnxQkecwzevRfvFrqybjwT2Qi20slRVdQjiWhbkbrTKRihQY
8u0t0x/BwiavQAp5pT9I8MX0TYrjD/Izc4S1hCuFJk0pH/xLL9kMGgE/zIAm4RFB
A/6sm0Kx1QgydZOkQBh8CJlyTPJclfFa4EKIJVsXx1Ux2fNtsDwlNEwai8CofP+q
DjfCc2ldZUgcM6OMWFyIM5Wr+ZMVkyAP78b0ghsLCoHIjRnEIgFAHCW8Jkuishje
Z/iE3JD8AV542aMLdO2TxBot7HtXl5rJmX9PCzgb2JGLNUBNXxt9R1Dw4Bg/k9aJ
1p/g0hC5awV7WT+q3tPttKHCyr21QCC9ijXaPRwH7HNNkQ64nkFYC6D9s23fpHOI
R0U+Ulpji0imXRG9fDZ9ml4spGyJ5sJ5bt3VZbDXwKKJxPhU7kUYJFKlM27TS9Nu
6mUZn2M2/EiqIh+mTjm290TMQjAoB0AxbQcqj/pcYaygDHlINhNLAuvIQAEMX1Yu
CidoY2Iqd7ljh5p8cb9Bcmo4ZVWAQUZrJ6tdegSD43NlzB9/9fK5Cauth2boFBjZ
dyns3UAfdwyCOJBWe30PgQYN5FQGOfbKEg/oDbzZlosIi+q0Bqx4un0VfjzNzE85
IEcG/sxs28z4wHEcQlTtaqy7v1muPsw1nTYh5bteyewn6X3qGnxcbHu04YHB0NO1
Z/6FLwBDCAytFPRA2DSvG146WUSsUc11xOfimURb1wEwXibEHLXBWgLueaGG0REC
6OlOW3q3kYG4BSS1Vvc2BEPingajPikRl7d4qD1Kv7v6OtkPoy6yzULTHDY6ufmI
vMWsip2OaN/9CjW6bMhdczH6COrR7fH1wcgIgx+96Tc/gsHD06Gd2g3oYpmp0tba
ZObEiIGY3N/IzRqR9zdoRrHTh3Medi8Vo2kY3I5W+jat5dSLZpF1yFDx9bnwsKhT
D569jhFnMwQJCILdXRxDHzefKhtPSPVF6BkbX4TK2oKoyQEzgSjSj2Gs8O6iZzCj
N2i0yGFDrqYlhw+genpWf7ZUAu1T8xEKZt09ZA8uz8qiIPp5Ngjk/R6KSVQfeYkk
C7gsY48Trinln/8ueihS16jPOQu4ij36YeHv7uY2nHjmQJrA6M1Mi8Y0s7r0lkOs
hFavGc/sVRVGatoj+yZFk47XCf2sua5OU0lT6pw4BVSmy6oaAwsIhvDzOBj9KSKy
maQe9wLu8VzbY1dRmd43OjHafx14v/0ffkOmivB77nHXPC3UPkCBBHkgN2b36Aci
MHcgqGru1hXpw1gumbWZRUt0BaOWOYUwSkwygU9GjL1CzxJYfgwRtJrrus2E8xJg
EzoCmzVPFf0x2GxeW2+SmjxAWy2y5r0y6CthlsXu4F+6vJKQJPfdQ9LjYgIGuw7B
phYiFPfx0y2WTiMzjagE4JjbH5i0yAcakb8YxKMlxdcrEbcP7+sG99sU2beNi1B4
7vBdnoiDxd1SsowMB/SZBSY9sROaqMWAZEykqtzv2sCcNFVTXmaRCT0aDtHg+Px/
nd1RbytkI8IB3YdCPQwxNVOfmaW6GE9FkXezUM17s0oNsq1R2iKWXsBdJIM3JOPk
wMSleU/rylPcuJScKplWqn3AtCBSseKuliPtRn5M6NPL7XbzCJ2SGNC1vziRBy8s
BAHjIBqAdmbndTlq4nyUdLXqMP5fmPTF0yueMvoO3nxKSXBw2VkwxTtlDqKglB+O
SmmCp9ogCi+erwK1/4eq8Q0OY4vgKvH64uBwM/2M2fxX2d3AgdqrGvzXtKc0UDJ5
CLNr5lmXcjfVhcxUKSPTePrFM0dC1nfgsioeIC+2vMxPowVXSKXXJoUeRkmCw72R
h3qCPaf1bsa5Ml5xLWPNfJ38moYH8wi1ME7oSL+HUc3IbJYULNjiVui5TovyyWSQ
Y9hnnOI0VSfpxBxLvyLcdVRnBfPawL2qTO/6jU3gIuoEEiXMxJO1iT4UUqf56IPV
e4pxpQmuKe2NHhFBhCJHL47k3mAJNysE+YgUN0pcIptAO7jjcBPCGX1dkgt6qQMN
KpDuwapAGlhXYWGUKP+h5Xvb9xpmW0N5lfckD2CHfMEQ+4hb+X5E9tZXQypo53Gy
DWS37HJTHdlW7CEBvmPWqDdtiXbMaVsePBFMbqlu2OymtUFWDJdVk4cUuBwF9ggQ
Fb9iCtgZ0SHSLJZu+w5I/+hXlSx6ZU1WtYyRoUgxtteOpZsMr2SGNj8sSqdjI2IS
6kcyB2jHSfekL/gFvJLe5+2tV3Qu/srB0eK0N9+rd/2LMPJ0IiMp8B7wEP5qnYyG
eWLsIbfrTtsKOTSTzvqMBIdtjXkVUa0xS83XpzOgQ2v40b0H8VqcmIRBNvzaZqr0
voBSWzZcVf9Q6rfNLiiZxepFAtKOYn0ovml4xq16P2GKcWTlh+7/RcI8vto1ApRt
rcmJIGjy8nTtSqjl3BZLdyUuctFo0NYY92EXGJxEGnR0/kqV0zQXxCuKwZGQHag+
5Z5j+bt3j5Q1kqkir0k4urfei5S/cQaJYBAvVXuLRwH9T71syCSPARsAvPpbmfpg
+B68DKJGHiFw3BFwED9OTI0TshbEtbBKeStms3Ixax4tRqO+ZFhPL7RDZBy3Unsa
34m6nKrlKs4Xwu4CSZVmAO9+zT/jD4xhnD7VcIfPGU2qGqtpyp4hyTBTv0Tk1RHU
hZE/VVBzhmMV1nyc0U2bszwtj4Iwq6WXRp6w2it8cBODK9Fq3qfO6jx/JXV2tZCk
0Tb3PWv8yoSamXgEP4ugBIgEvjxGec6GUGz1NeOVQ/TsIrReD1phq32zMs6m0Bfh
bFhjkilmAPghv9spNSCSA4UaALYns2YkGxRlAXAAF24lVj6xEpQ8MYqg41u8T1mB
r1WHqqg6A4t/z8oFOO4OIS68qAyeP/pp2ARKrppf0Yu9NkqSi/0I1lNeK9EVaBLP
cmtfLHFG153SpMrafi3aTBOdpi7BBES/Oxh118bj7IKkgKRtXRrqw4xY/MqloDG0
P193VUmaP3ZnVT47Wk0yVoxurHLMoJiaoC0ZWI2sssMwNIscs2GYGtrXqYWJoDwh
sCRPBTlH5DGdWUl4Rgetd8LP8l46ZhoVyO56W6TOM+0znK3MfFJUW0fcHpuZTQm7
MKCSw/q2eDMGlrUkleGXNKFq6LMMd/nJtcLG46W8EMOT6Ft0EE+4VCTvcMGD7CBG
MNgbmEYZK1zWwIBarn+wKIx3V188w/zmdVxnDQO1An8h3HmhxjURlhXq2RbkX8YP
jJlNgzSwdaSdY+hb9WVt0vKW/bQs8FQm16CqfdKrDHV84oHACwf1hKvAyaYZ/ANd
5Efysv5dsMi/zm2UzpdC3Yq9ePLeFcmfy0wywZmdEuxVkX20yqK+V2Xf2Jlh44bc
8SRHW7kLsFm6845OQbB5EzymM+xtBZOPXizvszQHJkp34rQJmoqLWG1wiVTMGs+V
SgB7cW3MtX/Fo1PDayk6OWQiUa2VgBELUdqPw8cDgovJOv/4swWVdBxyqzf95FSZ
IE0gf4wwgDhEr4X4mcAgnqZVDZAszWLDNYwcJIFOVrcyODPM5Q4hAKL1gSJ14IMN
BKbm4ly2IvTPGJqLsjHuQjo1N27zudJ56XPWpjjfYOYnT5e6rXF/RiBlGqyTh6ov
oy1gCR/FPgAXB9WT9vqQFCM2HvYRhQ0NezrgloXre/eCgFqB2zDheyfW5i60jBXB
xFo7GU7GB3ysuhoEYK/xgqv9qf6NaoSjP3E8i4NDNeGX6R5mLmB668OJEsi1EDl+
1ep2EeGYo5hkOCTH07vkCELp317kjzkQ08u3eWWYBWtco3vm1hOckVFdz14QO+6E
To4lnZa3yS4PqKemFcu8/lBurjBdWBMUXeQXo5iFX4RpvrrM5UGywJgXpORp0G9k
4I4M0vCzuLW3DkX4+r9alkDb6KvzvCJ9EOnIixLRtQCLoCULfwoMezTHGwp541qc
DVsJBHCrl1MaAbcYKVPcU4imzIivgEM11EHGpop33QFncgFVUR7m2Mm8A/EC226X
0rzJPpov+fQ5B6H4Ku/V8RjhI94NymoMIUgAxrjTAGxKjpXc0sbfB20QCAA9uoTE
Ncu/3F4SAk60V/hcZMjuzleOlvKe6LHk4s9woU4Fd5Tbh1bDmIG1S+pQ/NisbR2l
+BT5qz5NAHkPs63cMaLuZIsXWk9CsZZuKDhLXy3mQKVzd8nxfldsXcVi6cMclBI0
4CcsB/u14ke91s1+8Xi1llmlHH8riljrSznGL/Nmn4+M6dZwu7odyiHfQz3TsYN8
KJk5Os2+bgB6+r5KyRc8hdLjaF8uiYo8Dy52l4ijOt40ShjY5jUjPyO+Kk+fXs6S
dBAQMA941ByAWaYYN1r3ZIGFH0pr3lvlom95oz/ApKUaq4077aOGXI7+jchQyojI
GguTjf3tSSISA2YKvm9+/XvR8o8eNqpY3Tq6ZHoKye9imBk6eUE6tVM91I7h3j4L
1aLNWVEx4IVROBgpy34xHu0iPlGXB72rfEE6zBHj1Jj7WKR4m31mEn9LulmCRIXG
/A4sceOvbCbnQg6L2EgTziN/Yk8qvMS6tSX1WgYXSyqL8iGaf9CfmSX58kmQ/nxe
tpAAXTZ63APf/gvcyTmuURCh3+JT+Ebm0y1yzVkK7NEDouNUWuvmWEQAQx23lr7n
VSFLaR0DhbWoEmastfp9E9HSypL3RDJFvJ44VDMnYvZG48TesAouNcptRNbansAG
EoUnyMEcItV6pH+9yApl+LNHrxP8BPMv8Q0e/xuSODh49uFLl7Iy+tj2WbOY6C2d
6975jeLySDzBljFdxVRCyd591yNEypM7aLG1iAlXk7f5ViqX+aR5GdggqJ+fIAtP
vqy7sQukMonQmeRE5MQed8LOHc9xC0yx7gmPtkqzFA3T+cop6pQeYNdPeYYfhyi8
F+sH/fIeO7gOYGkUcwBcZDFJ9zd9nZHKsZITxjlRis5Id7D5oWqM4tbqvvUBLtqD
wDy/00aKx2/rMVGqvzAJcGmE36bz/HtY5Va4G+UFIriGq1SeA6IOhxMHaQy8SnwL
hPsBVRzg7T2xir73nWO0asLANDsv3ML61tHvZVgv2lzhJ/ns8tLVfFuJyC1fP0RT
gRwdG0o4sT6osTEtCgOvtGl6jtraq5jKIgRfzHb3Kur4JZ3LQtlv8AxR7qtDhz+5
7SdfyHfH2gPxT8ITR7tlPIhLbQVYylFizZPBfeyk6QUKGLJvysjbtEA/FJmUgk0v
YJOG3u9N4+JOBVJ+E8rSuCHZNO+/VSwaGwNmfYaPS4/1QkmarZIW/oyl40MVD4J0
gXhMc2O9psU+SyfZWK80SlAKKpviIeKcz0MtL3ywngJIQTocXoGWUFTvZjxUGmrg
uLgg+8NqONbSsUHgfaoFPR+MYp0xVA57GsrhV1/bOyURoOMrmXegeoWoy0AP3FlS
2J/SwFcOSDBF8Re7k79yFC6AZ1dED6g/iuDq6NaWXkdOy9wjoY79N3iFA0kBSN5C
kFpppAOEXEcXibfMDwJl6cvDvY9SiApjnPqS+CBahFcd0jVvHc/SNuArFpiRJNIF
JdCpTSv/Dnq8TUfgn0V1L9/zQyy+Zrfor74oOzQ+W94rBKCB7wvuLXxNg/NklW6Y
I1yoLRRp5KPdkNylbW+itpsPN0rP3gaNRuDvEth11W0hilGInZ6ZbZMY2BS00Md/
YdKSal3kJ5Bw+r68/FXHwGZlyjSRRkd9q7qE5nxGYj7lfCtK7rHwSTrAOvmf/GVh
i7TPllj/awru2lHEZjLj+4/CWUWK8jmzfZKxZ22Rhd7com0K1IT1EhIcFahg3hYB
h5zXFy4KbpHDPJjtyFo6iafsBBVULSincxdnShNO/QHqa1tPXOOxB3+tMOPm2rMn
s7RGmR/x8jZuvmhrVyMroSjNRftxqWT74Z3v4EUzBJ8=
`pragma protect end_protected

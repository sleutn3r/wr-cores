// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lfnD4ReyyUAGOej4P//3AQvc4jul7N80oydee8KNs4okgYaPKy5bnkEBg6DRXCNN
698qayX1LXSVCrh89IYpLGn36fhVvGTFuTS14xn+k3sdnbF1XmAHyKqIv9SevHDr
K5HxnzrZ8eCjlpO3SLIvhpmtS8lplz6uje7o6UBJemo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 16704)
nKg/D51UbdzHM5IHvAJb3oo0oWjLhaIBhL26KaAquWZBC+Jzpze8YM5hAhnhIax/
cNibAFdSXGGXVIRwl/fByjRylMNzup3G9BvouqFyrh9WQDU2WoTzZY/Vc1fz3ZNn
G2MEUkm5mt1WjNrt8Q66RkmsEteBDdBEoDbIkyR+p730iM95c41Z/fmMLYONB8ml
z2OiVLupi4rWE6Dlf3DRb+HVAoq17CyVrNvxJkcTjqisswDdyHpEqIaM/4spRCkD
JbS3BtrTZ/O7XyKXlGMN+3mK9FheZZKED4AZVpw0O8AYLK9NDoPYJ+IuRhAI3ytf
ihLYmOUrtIgPYbZg5sKXAGJlfj+R4DFHY8oaM+WmPOIkQxk51ZkA3SHvtTdZ5yLf
vqO8n4zdkH4mjIAUv6W+Y6n8L2lcPcf4Bauds4/MDStGS7ue/ho87Q6zv3Q8/OT9
M2PVhJEhHWKfneFCV3967kpxQevHqxrRIaByyfeL5kIUYRMXB9m5gj7i5LMJ9Dzz
UC1a717vpBYnEfzqVqZ1J8nT//Q1ZvDSstzlpbXQbJCBpiJ5INtxhZVpo3a6yOsO
wAOO5mbqUrQvyRIkcPZAPKlpth+bXvuS4uD7YryPkuvASRXZ6IhM+29ald6rkxvQ
EFnj9BJZy7ADaZpQuw27qYjIsCWxM0sHra11K4heqei3BJHI/llgvcAP888fpfGc
wS0g8njIO0RQ5fAzFZAnyLkp7FYEvJ9xdNIMda7ZFoH0QJh2EfcB/RvVIV+jYcnj
URW7wwtYQeHmL49MLAEpaBG1pMm6eJ6TOzZY0wcCx0DiFMO6y3h4dDtm7UebJmM4
G3f3ZNDx13kkm8yYeWw7+ghLf+2Xf/IRjJ3lQpcFWrSJs5A7qvLq77lxly6edgJs
bnJLldNZ/FOnkE2575p1flT3DxhDiX2SRyyaCZsTq361DmiLCaKDCixyga2XzXi1
fjNZ+0gmypJEIMDbT/jm4dMx9vThifMRVCMHvgvaD8pAGOr+Ro9pB1Eit1i/V7s9
6gT2NMonfJ2yAjzJ+o4TB5cknVPiavBsicMGfrzW2Ncw98vfgjhY4oIQTVGMSPGv
92WgyaTSRKqoY2icqM8PzjD5bSEUk0KsfNrOn+56K8kF7ohgyyGYcaWGtRoMpOyK
Zg4kLMMv6x5yN/MQLfpga6K6sOmUn5ZJwqWdOjC+iXK9DCMnUn80+dTm2WahFB0d
Zo/lPvYZoAS8LF8sAFXgIOFrVMKsCAVLHFo8jvnRO/vPfqKOldQTjOKGFZ5EVRW9
EUPnmGSWgcdb/Se4ckpecRjqG/EQRgd6A6/1Z0pYLHReipIfUQFhUfHKto7IZ4VK
+OGfsKtzCz/RE8bfQcDT7jZMueQPZuQK1iWZvRra02O1Th4b0sUnFmuldaIAW91X
5QqqrMB/UjGJpQF41J9+FdW5weeBB95g3LGDgzFAbHyhGbDv0FnFySJDTBk6Iyk7
S2GcSuu1Y5kKuoDSoEp4rkfg3IbPY0o8Q3nNPZqsMyvjW6BEgz0jjGtCuaVxbqXa
kaSdXAlxJcVHTNEQUtGVt/WOaKlnC6UVKx6qvS8dv39IYP1T6FcpTsnmuCxxJg0X
DDxBtRcG1Issl/hk6LP4S1cvaU2TWYEBna37O3EqhAR9+zLREDiHvi4UGtx4OYzj
2l1ujoWC5Z/uucdDvi9OMnEmuR/kGB24TuWuKA9HdUj7uPp9XHqfTyv9+zGHcqNC
peerXmZg5kGAcd0Oo0gMtCvdMhlbrSSU5Q1/zEDlCzM408n9oaV51RX9141AQQFD
JzD++yVfV+dSfMQtgxmGbFd5+gVf5gBduvKjEVtjRMDJyQUbWcuG+STW2gzJBh0P
ZrJ//l64JHZtjCwgiv5QvyjCVI/+0D1a2ZcQywIafvtZ4Hisqks0rThe5nnHJtuq
7fztPezRbyJ9MBS+gNksDVW2HeUt2tz7mPdlhkJdNLaT6d7JRgZvalILOU6LpuIa
UJLlxtO6f9SNSGroMFPxs2plWnHQf+sMRnOhZmYsicOIGwApP9GE0yI9yLvGxJah
w5h/OjguqNOGLlZdArREVbesCnbUlWcTvKIkiDIRI5KXgWOdRzJFBbSIOZVyzLHf
t9YMAxtaoXoNtPJaPNojnr3nc0tUOotJ/hEthAoW4RRgZJyUFMconEvkHDGRMEid
dzCk1zSXlWI76Q7k6FlB4O7VbIm8EdewUXVcnkIsyVcCtxXsY0zJ6EAFdDH+ZXyz
0u2oXrhQNNBTSdwJ0L2QNCM70VWY42bJ43uW4fID2/4afeS6hbriwRCGoA9+bf48
JqE0oC7EZXLnOuoTdwCj6u0N5vpSQrrZsyn5tSgioVe5w7w7N+iUvQhQBcKzWSSi
79p5BTSqTlku16+GFiGpz0DQDKtexZTh1hvry/uCTXaVqetfSvJs2lODcmkw5aHg
TkEF13XQ1/ispuqappTJxuIHTP/I0dYnnwW7UL+duU4sHwEA2rI4MCWpF40wZQ8S
BtQkLvM9cZzWEToyC4Qy82HrYetfEHWWgYL1kLlSUb9zlB9+pp2inAAF82Puo3a+
qF+FL0wxZZai3xANBBPnX8+0NF7v6KlyPcov73FZOdHK1Ikd5ZEUJ8+X/KOptWJ+
8fQEjMRcBrMHRfJzPHfEMJ/sOHxjYsLrqBNU+iqJUqkVTP4leNTaY9wcwBRjWPIm
CxvttXBg2XHNqIde251mw1tKHQCsJ7VBxD53O/IzCnyI5f14SoY27w0qGQwFcaQu
IAAl0YuC+vi2Vhd4NM0z56jMP+g9L/9sOyvs4KxrfBzWOKKuitkSg01Lk+nQ1snW
74Ld5mMsXU6hrzbFnnNhfFYWSxpYUGPhtJxHOG7kfyZXmjsGRyZTKQMJZ/LWNvWl
YwTC668MvwzNtIlsmzeaO0/D7+CTsyiQpQvZvM20AY61ufuOeAV15EV0axuU9SHg
v3zwQbRNFnbOVmnu/lWTXe905fib6lUa3MNHZad56seJHgQWDkQnZgT59FeHIOY4
qJWaf84Gn/tb6B4D+sKEqWC+wEvEiIur/J8JGQfWrWbmXBpQGeP+xyy+IiEeUh1h
Ex6ujj2JGVr9hzw2PuzSM9z1bJDZOhf7zFodkKcsXMfXHhikXZy8OywWxyoyCZEc
OoGQGLqcq4HjU6MJu/6Wcng44P4cxjEslXyCHU3BmxHNKcAOqlU0zoSf7vnSa0nr
olbO1cX39vfR/JL7qK9QL5br1Qb05qSr+KLe/JWq8Jjz2k4wYWQqAUDdqATNFLuB
jIOyVDnFyhx5EKtmttIt0xSMol8QfUX3hjbdloa7cJ/Lr0IjgROd3esQTd/zFXUy
jMwmsnzClfoWC8HlTDfreYNNkzFnoqOmzSBwQKGWosL4XYzRgY5cZyFvEuY8YINM
Bh9DAi1NFk/N/q3Sdoh72sisFISrfPFV2FaE9gH0jvmBfnpS09ruyb8+6lDf6GBe
hmCH2Ji8wECKo9iT/9iwkLCZHGq+wYPsyHUYcMjjabINaNu8nderdgrUHcOevT7S
GTpp4t3yE4w+ANziTDjLjmx7bT7oYrWB9gC7FcGhptSM1vEVlDBASWShQIEx0d+5
h2ZeEtdWnbx4WjSToZp4W0CMRA3QQcd+BExaaMlx8yqlfjsvTh7H2CE5ck90dI7e
gLPYmbv7sWQVD1jIPXrFgOjAYNHg5iQAJSAv4lC0EUYgolvP/tBUUbyg3r8wwyaL
ATTE05wuncWxCSdRHbgFeZXo6OwopEhGlFMVO5MjYkrtaBf4p/94+fqiNbVDPUd0
o8zbxT5R45oUCkBSinGVhV3Nuoio6xgyRJ4x/9JnVxQWeZCerRKWn+4kxOZ7WOCY
P6ZC4KN2U4GefKDMaH+ZwtneMfj1x/UdzQ1PKl/Vwy+4/nElaUoh9ewNuCO+tlnX
U0/fDAgfRuuMg5XjI+XbATBzjfyE7QzrenBnAOzveWcTPz1b+Lj4mfj+rNkf4PXN
xh4eXIxfDnLxJSga7s64D+rdfJm5h3nOI61IYeNiP50CsmFeM35Y+pF58Utkw42O
wOa++rqZP5dekqH9izJtAkwBaiUF6hQVSkFRs2GlwUMGp7pzdztoSAVtybhxdyPe
PZAPWA5gnnQOYp4DGHt68k7CMoXXOvdVw4IrRGOvlQBQ+Rax7mNLyx/hoQOy2Gim
NPXC9ZwyGNUIspJEHgxh3fOhLIkzYPL/JNQqLxUuyVrPTkTuHjmBTGcswA1W01qB
wRYX+RvImLwnGUvkB0SBjtotPEh0mGWIUdWBxVK9mHzV5RS+sGJ0EyvGaG93Va7p
s13q2poacNLPU2GB7Q9im1DDEe7f2Z50V1D7nVLf/rbUSnA6qVCtz1lAX9O8nAJC
Dl2LSucrbZqwxsXPFRZMyeKoe0hPl+gxqE1JA8FIZm3UQUsA548Bw7sNzVKbYJJH
GhT5OlaqvpRdUtKl9yk69POHRfEEXmSygRXMFxSGPO5SV4eAjzyzIqVCBdTpvlx4
jwxNhF2G/uLUNZ0T0GJ0pI5cbEPEU+i9gSp//MTMf1C1hRniTgyyI6Qsn2i55cxJ
Wo0q6u3FQydMpryy0WGLSWam9M3H4yw4MpxKrN7SqW0VPF+v+k7Wfe2cjPtaAPUK
fzq0IHUSTRjFddwJjGwH8nNvOgTwN96SMTsn8n9W/FvkbUscK101nqLRYJdNqu3d
n43fxrKlj4Gcf9Xmt8ZTL5ui3U2SGBM5P3zjByKRTqQcEsNjAnuT4s7r0O99QerN
4LL9ZlTbVvgr1uwW8yAIN/acX6ujS6zz75IlfPw8utIYcASN/lFl1jsvdJfHYuDR
kyHclT7l/anRcJh3Gralof+R6Nj/Fun5NeRfvMQg+NE83KhL4sVVaIora9yMORwO
lOm8ERyCU74BM2pDQ+RNLTmX5iPTdBIKXNM2eu/owz4KDMHPZCtDQ044wRCrPHtm
E18SQH/6LIeQVzExJujVg9NYKTxU302ag5UU1pD8jsukPyqBu5fdhXor+S1x23fh
/n/imkBHjTRypcTU8xlJqwL3z3Z0OqaILGUam9lhAB/BK0goa+igqLCR0CZbwhWp
9dk4g5a5OCYJbc+qkVu2ppMYRuGOfNhpfz05hAlXMWjTSn2HfKY2SbSrDhAUAkAY
0oBpiHseyX72grRu4K7niTkWbnKComRTDCmeJmvcT6JUkaBhVnvSdr9sQdmNNm0r
6cgS4v43y1y2puBpDo4v1+F6//jgF+nuq1zYyQvE6n1rgpKC7ieofYQWjMjAUik+
uNfxjzXPqbXeOKfdJUkexkenmVdLdHTAYpwEGrb08MVjyGnNi9FwduvzGe3z5lq4
/eUqhc+NjYi+hZhGIJoPtDZftUkgl9RZ/hKV7uCGw6dafzDos7NvNSx/buJCGbRk
W+yX6rXJxGzkthxt75uSzqUNvzk0YC0IggRHi1Fp4OicdG4IE8fmkyqFpg1zjPgw
z0VlO4YsOvdggCcYTRDT2FlxbYXEz+cNqSwhMky/ItuLVDwt3oO81z8XbVpwu/WC
5zB7XMYjNxz37ptlQQSQvEKh+r/8P4uGVMXOzWb4qv3lqqLsrxka+7nqYyK5WzWX
4WX+c9IeUIkEYxNUZjpDOKWgAiUmcw4Fd0z6S8VR5K20+IuIfx9yJm3BpJuYD1F5
HtvHINe+PCcA01HZycr4P5rNfitHcswmvZJSBWAZQr4IpINfmB9HFNITRyUFLCij
B4kx4GHEaKWAMtQBB8ro59vRGfwoHS+Iaa62n5zXFXN9zWSewpfLY4cWVmSyHPim
2F1gmIR3/zKMuKgS6iH0LUD7y1FBfrIyGs2LhAH4De/wbxCLZJq9C1mDnNwjiAZN
6PKbQR+D4p15tTo2lxP2FrbOLMM4J9DReYTZAmCcM5QGSEmaSrUpIi4weZUClhyz
SOrGtd6zgiXcS3AqeMEuwbxN7K0MLBc5GS1OG/Qnpcr2sycwI5GK0wyDGVKW4o0Z
9Hf/xzAxuNDjcYRYgY7qE7tl4xPlTCm7uIqROWaEtu0WMCB4+T7Aw7WwKt1Fqz9X
lsvHlejEkseT5ENDO14uG3pv8pSXiHJ/BuYplkBBbxgZ5/hgPRh7Nw9MvKIzv5sT
Za3T6j0YW5VSUKMZAfSIKoCe3p0/rM01P5Dd6a3ch1O/dssg+w8lTjvWjHo6lqck
buzrAZUeCgt+lklAjgUfJWjB5sFXudt7Q5+AxRwbWE9Tg1McZrUSERl3WZdf9AjF
eV3olTGj2lGCUwFe7VHq+/x4OAXHTLIrcWf3rZ2T6MNS+HpI64luRN1vKKMjAScQ
u/9NrpQIjICuLZz3hcIi84sHOee+bpZqRuRPeVJlZzIIyGDdfnDF4jvJDAOvMm1n
vZtcd/8DKC5Yy4y5Kl4sqROwkcfgAIEJtBh10/C0HzDyDxVD4avBaXfdp+N5knwn
Xlg3s5EWCvwcibLKjPqj5gJWDuyGOv7hPaQql3BE6JdFmUKntMYb9clQnyirwB9+
czH/x6lH4v+t7irF1UNgBDlIbWyCpzDPOlXj5i28zMDY6xyPjarKufO0r0xyeSMR
qeXRhg0pCI6h1zZmUWnjv93qUS/zL1ixbTjqKqGmJfqrPvk68vCe2PPL/8z9dyVJ
/4RBGOBTRe1ukZdq1xvNSm0oJ7UP+QHBkaf1mV1RTrdK4veU0Vz/yNZ4RKTAeXjg
NREeDJHEMQn9ymb/zoA1kQ5unOpDv7GJYz06fWNDyeF/GKPprOtkjuFBsul6uDfl
VQPpxAbLR+P8N6tB0gKH0J+cbAVJ/y/AdiqGgGM/qaW/UKRzPnjSEBMWlbmJnysD
eiv2hOcskSyhQ6PPXoXggpFl4GBluxfkWaaJU+LWEyclV9cJ0Cc5hYXqCVnFt0dl
1pFeY84jflpGSQSF9PK1j1i84cv+xQVYnhV4VMvYpp271a5EiORouMEucO1Y5WVC
CA/zmqRzwWmckvqnmRnu4hUMb0Ph6CkfBpZlL8A5xhfmicaIKEV5wtx4BoL8zJPd
xz9lfIgwcxrfl+M/bfqB1Tflwr0DMiw8W+tvKso7frmDtBjAK43ddpElbDlFvgyE
JQwOTnyHA3EGq6aFeIob0Tks33TeHMZ/b3NYiwa6IS+FYedFpG1TFSzS0grsL/cp
NkXXDxyTFsR43EEOKbv8fkyQVpTU3vdsWl1C8F+Nc2xLQM7tfEpgcVRvHpngzrRU
7ji0CKHCmq9nSR2M+LYod5ihw8cN1aeSBogbuRBzgWypaBA4ju0Sjdd7nt9lB0U9
HcvbGyGiVQJBgkY4dlFIHgq+WnQ914EAvrhrBBLI+S/PoenAjX1jbMW/hzKCcgOi
FcJfItlL61UICA063e9cdL13tNf2afaQul5nUHP5Byeu642bhLWibNKZJPTTBct6
c5N4tPIMCT6Z7DSgX87+MINcGBxG5XtrfvfjcgcLGtDXeAY4vkK28RxfJZPS1uZC
xeC7WWbAopMFkyjtgoe9AcrJ+sf+iPH+u6VGHdqCl+xBRFayV4LMimd2yjkECcaR
sXYpl0Z5YFTReGPlM7G5faJONKY6SYoNhhRLXzV1nZAPy1QY5zWD+sqzeTDe9kI1
2+E7u/8geqPrW7LPZzT0AFMHdvHU0iYJjVNe/J3FaSsCNaP+UooYRMC5WKWxodu3
XBytOPaHt06Y0CjZz7JkJonJRxQZdWyX+PrubickYW7n/ELmyS4h0FZyIPXY2JBi
J4Qpvbh4ZxQULgjE40ZZxV2tlnkB7jThWtI9ioFcZKIzkAYbAXcQpF9L/P08J/K/
4CaeU/y0FBRaqpru2+b0KBYEZRfgUBo8QsZQra1qNVXSg4eXJADvIm3YsBGsx3oL
+UzJs1nqENIKQZizeL4TvNzfI+VF2Z5fmP2P+S41chy3yFo6t1q98i3Yk+pCj6mj
CogruA5P8pK4MAcO6hcp0MrbloD1JgWdFVUootHXnVllkNoUTSkUMUMDFJNJWSgC
vAnAC61e0h0LBgnz4SKLWg1KSTikh6GNYMpduG/RHwT1gCgxEOM/+AThG40LFLMd
BQcPBhI2xANRvygkmV1VnZiDfKcbChb/Ap90OzBRQm7n3S196CmqeqPpyNI35n1T
yRIj6Kz8J6LAgywi+/SAFGLCSseRduz9d3m10PeDT52vFDkuhZQ/GgWbn5Vff8iL
lwf8s2nHlchklCCE58PUJUbIW4fOes++3lsjgmQYbrrwtz8QJGzcVqMpC4Dizdje
vivreVLhgQPEp0KjsAwV+iCYUbP8OBA8vt7vEOOgD1JRnJUbZG8rlL3oPRm07ekX
M9D76ffRtcBUtOadF/YYWHFzjVmxTBP0nMWFZmxRLmPZTCG3F62FyBk0SLMyWx9z
2XkGWPlHgiVHYi9AFCL4GBpvS7bDHnyYIoHkQoy33VXYOF37qb9LXJqHVamenUfu
SUkwUjaxvMtzQvFdIffwCsnmXX71mEExlSlWpdbkp7HKRTdj4jbMmNaIPZ8FxQDS
BfWY9npA7IVA2adh421+PkoCnzC4h++aND80yIPWeIF3iG5H4IwJYxc5TJU679Ll
JDLaiR9TFfMbiEQueFqMHpYtjmMNdft/AAJzvhzOq51b0GH4oT+P6XMadAcp0/1m
mQCiRP+2U789T1y2rf8kHR/9SOD7NAXnMr/OcUdUdkst5VMRzGbVm0QdAAMdKLtl
Mb0YKOxXeFYRDqK2E9ftXgZ2B1hATiZcguKxTQSSBaDt7vrGFB+NKK/W2qbQQZmR
m/nIAd+tDZs+IFC2jvoEFDPfr9kloJ0NxURKDzMTjY8j3/dsXgsnAVPvLo7pF49z
eX26+01Gcn27BV0vfd3maW4Jo4OoFw22H8xhg9tkwfFKGKn67XhYIAyiF9j1eF+6
ZK6UkAls/lOovbqouw3tT9mz2FHeQbnKiGz2yPhotT0K/FHLF6qZHyl+s4U52YN/
xBbIS1h1CpSv26scs9OBNL4OKhYQhNRVXJlqHocSjc7DdckH+uAv3E6CQ3y96T+B
qSbPuICq0aTqAUxlSIpx46H05aN+avaEnFUKN5nar0ZqpmezfquxK0fYEr+qiBZ3
guFDl3Pqu3ktp31WPA4D8jrqvOheQ6LnPlOVN2hNeyPJp49lDOXBZvgNAZOp/8Cy
DW4U9q4e1K5BUYqSDrCgxI6lRbGiNDPYRNC7V+KMF6E9+CQdnUL+CZbsz3lHWdvt
fMrsXeRCojGevt+ID6LwHXrfe52XYu+bm2Dv56JDaJDa2bA9axNN+cIoZVyXDOYM
Ja5Y1nQwfOjSRUKP6bDBN6v7hHkfHfMP6YM92tci1KhTVE8XsgpG3C+Z7FLNX8KS
k3XcSgj/z/mNc+yJ04aTSejbV0DIy/8Heph7rfQJvo3a7BRo0gaWKfAPjVG5Cbc3
lIRmDZpoXdNC5PaktKIRN2GKUiww4O12O+QB7lJkEgpAjSaw7c/M7TH/onMoeI1v
eARP6XwE8kdSKBJMcl65y58+jGZB5ghGjNrZDMdZq7WSxgkPyM1VHLyNBLctsokf
xyBJaMjhrw2mMggiNVWQYuKA4aG5CSgBzf+8kZg3GHwbazmkmWhEqW6petr7Y/bQ
OicXN5giVziadyKSXjvMV9nsgUnwRlR4aOiBa0vH7JyQs7xJTpkvc0NTSiYh49lK
tcAqBY9UDgZLmkkeLcZTu5H2M92roFBcfF+iNmvY+zcHOUkXsHfXV3XoL4HhcYML
BVlzgo5q68oGybHBVMd7cmsWlj6VizT5wvOfEfZyTK6HS8KBAjOqsDaF//Am3sMJ
DSFa2HuGWLlFFUMqhwoE/ozDLA0p99RgILkrYwdGLufMDU0QwrSpWzELP3QGTx0q
9PlBBGw5QgT/8rA0X0orxYqprqSQtzgkaQE3L7GL9cwkNEbOxvoRf5cuW1vXmnWf
/nb89fKv+5aPa5+vjDXdUTHf6NjhQ/fTj/JgMVr/yetOkAYl3WH2ef7iq2QKTV3z
+uj/XR+AY/YFC8ycTdfkyEtNhbOSxHH2pgU6W/l4teHPGB0GGdDwdQU2oFjHx6F7
XPKlSqcLqDIVd5CMAxfUn9GDrYmmfnM7r9FgP0fOPbvYLyD575ec1jRudxgXBDnK
TyXuxbOKQlYoK5FCGj/a0IzKD5VP7Ji5FaK7HEMwXOv1pR7gh9gtRUPobvGnt1cg
SQFyXWX9DwgK/jj6AVi1M+0ZlnCfYNy3cI2CB8aCq5ZwtCnbqhbzc8vjWIDLDNHo
AFSSTlXn7HdDUlg/eeGMRNzk1CILmcsyQXu4+Zk/7DhROxplt4yNILmf8TlmyDqV
Yfvmd67KOser2313A9EI8LE/2Hp8a9c0PZ+xw9OTcdC5XpW79rdH5hEkQTd6US5v
eHcRASEh61OuWwrLDxY+VAJ9LMFnX6BEbvTXoKLQ6rZA/rwrR+wRspzZfosbjZxz
/zsLFJ56kpnXSo1BRH9RimXUsH+s06xf5Qi2V5WeeSMS9LCRNimYC0M0W2krpaeF
Af7WybDTpGW42odEB23GBS5v5udNLScr+xKmRV7HW3yeBbPpCZXHRbxTvT35jsZc
mrQ00RZlgwE00L93IQ0vgSHfHpTLVWLAYGo2eWcUt8X77qExAcCcXT+arbyh0QLQ
CUpn99KyShNt8ObeRjVGb0bN+O4JqFwOCkuH/nmIDE5PnuozloZRXZUh3SIICZ6p
9O3s5s429AO6BXiSkJHUUewL2YOP6YTLVrapWrz93u9fzGLGJBbuJZQUyf5IDmnm
qLr9sWm/00bvMCwIlwGxUje1B7GZqiFuT1nTGuwWjfgbJaDHVUsXmJv6/iVOC6sp
gExL2jbWFJj3q7mdUY0Lq0OW5dNHcaB/7RJdY7CX6cy2HtykNlYoG0yLeocqZAv0
1p9IGv5RaCYccdEpTVpE2ZhYrE2qlSGWexFzNX6HpJX/NKYIsf0nJ1PLRQlfBDeS
8pEPEQ6yd2dAm+d/Cv2d/SqSPdluAgtvQX/vgVUnxTS/jSFXnqvjaFhTDhBmjKYh
QJ8Mx+nNCquiu3x3un7h1UuTtq4Ixg6zZ8PrUp7ba9ORwJgP8YdGedvfPQt581Ys
BhMV4ZG8TgUWXxpC+dtPnEwiJD3s5NjEcTgQg+x8gZ44yb23Dp7LjrF53xT04oEb
Jzo75iFSAquySer0DuuXm6qDRnlR25reopiR7N+TruMta54B2fAWHtjnCFckHD+K
l/UiOOcxJSbGCeBtmSciUycnn223DUmklGhGybRU1IWHmKqe07GyRul44Ve1T1II
NFd4S3NM6VPoK9FTUsdNo790VhQc0MT61Kh6pieRfFGkfgG7RukjIyhDFNciUNGY
vMSidGe1rezcOnrfJ8j69FKKFswV06PaSrZGE0VYmK65BMw/mpZJYqJfSXVKMbsw
kEQZBa8ujjmd4WyxUitdZ43tvUTdjpFgMUoV1Bq6kKq8sFD2VOA18ZChTe2tfQzO
E1uxJuZSAgD9uElHz93NtDtijHKwYkHn5EEgbos/3FYZA7Jv/Vud9yNgSkDxSv6k
FlOsaYpFf8jM/ccITXO+ygmp2Amek/G7qby+1pLDHYum2GTaWAnqkfZ5ImcQq7Qd
cC1LLJ3tiiDKSsWmY6Fc3YaXs87uYF+EpmXvwUCbYlmO5+SZkb7Qg07EEwQwFwBZ
8QxUUEr7WkNL7MtSsBVcBm46PyrS+hWUdDLfafX1n4C1ERrsxbHChmPz6YGlsmgj
o7JOYcKEcq0/JiRPOJP1HZW1L2gHh48X4VqGttk2hgWq1I8VDxV5PhD0DPKVJvKY
9+pTpO+NtZ7Y7+KdicdZeTDJ0xN7s3T88QSeUsVcX9h1r6tcD5s1Q0NNvwPNNICW
fV/phhIaHAGtJKDbjZEh6u9yzPD9njLt6PQfPzdC0O5Jo6WNzRo866ioNjgtgjW/
027pibkul4hLcdNm7q0E+9zObwKZoM/zsbFG0WQXDZgnU/aL5Vi3Caxfg9U/U4OZ
rf+PNegRj763OeNet6kcGhNmrZbpiH/vEiJ9hBtorlusrr8fakdrx8DmwytgcpGN
qSUpQQTnuyY8/kWi8cXQmFDmERmsU3X5Q/0zB9H98TP0Gf3EcwlZWm1HYbCgcDtW
iIfeDBlOvpcTjMB9RSmPGgLZHQLJgwRgHBl6JSbaBMarI30AGfrwaYK3x3T4Y4+W
qnj2P7L564Uduhg7pYDGJ76DiOtKuqdFZogoCjY3ADSPX66QVZn6pNO1jQ4DosF/
OhDNmVRtCTjmu4N+XCo4Rpq/qzjB3ytPylP+FMn6UNUP6NXjB73ySX180G7Y5qtl
XaUtOuOP5ZirLoaRGR4DHgQ6Gjau4ySVQ5oWc1IHNWPzog963QqQzqHedYX8n2Sk
WFgjmpqUSck94hKIcyVtIhgyTApHbrsSnoQKGR5rbv7u6Hx/bZ6JgJzb3yKLGxhk
92X+pyW+QluNx16RveOjPqc+OtrpzjbrydruWt4GRnk+FWPy/yjd8k2neM5HKTel
ZmvD4DB4xUyVq3igDqBCX1yx/J/o7gqz52LDojpiSctOohHdaH3lFbtu70w6Z+A3
7Uq8W9CRDu0Ye/236jCDK4ca3xIIjdNDhnRZpEDJPyBlNRPvbR2TqzRDKcR71uPT
Ln5NpdNol1HtWyy+Ahvkgl9NzXzagJKd8bzum6WM3mtK7eTVushJjc+jQdZXHZmH
FX9CDKkV5i9JHG3B81Qxy4dzQElpGv+fAeoqi7OclFDCUVb00kOF7tXJJ7U6EGYZ
MEfGqu2v7uqExeeS/DW6eKfSmnNQ6ADGOnd8TpVx0OJHaxV2UTlykbp9zZ6X3/1B
adpvDso97tjyBEhswa0k/ldrdWiJ5YS+fS6csptnJ6OY/+04gnRvCG0JbMeQ66Co
mrKYAcQETuMx21LtaRMLtwWIzAD2K0ev4oYPO+3mOEGEbigg1Fa3PUm8jijhXtSR
FTGhIM5w8S4sYToL4HSevqQ1UsXMoPCETiNAdFqhrFRRxUPX3N4Y9eQRkdlavPs4
7hv2YlLB638dkky/ciHWJRW4uSIFWGP6D4P97aUfXQNn3ff7ptZW31xTdiC4srF2
P7jSdeYx0xYRaCH9HK/kpiZxZr5HmMTp5kM1+XcjcS3vrFv0pBUsPSLWk4mASRHl
kfX8gleWeNkacGuEuQuaEknFskoij7F5ZOGaiiwF+fsWwvHKCOQxyQikwHIkc4Ep
sP4MSwYBzg81sMFHeFYU1ttGtuy/mAPI8peoJFCBi5x4t/PW80e4GoT06yUE0ffT
RhmgC8D8zSdEjO8UBlaN9b3SqGEJGNzNwc/w9kICZt+4dhknsQzhKoQ2Goyg5YBw
q1VNBnYXruOPhYvEkXgkpJkm5R/pu5lykotpf0HfnS7/Va7Cb5P+FG2H+MWfZTHW
8s3dp+u0E4EgWI/RV0YwOzdqrNVr0+Y2nzM3V2xQQaHxIZosOpAAFvQi7+r7n+DV
XLlmEwPuXECHgbrNH+QCpn1igQ1cYabLyNzMvsCRR4S6x1bhILN7MWNXQ1lz1GUx
AJYfRLOkoHl7Z8Ky/lBcGbICnnKBMxYLdxS06LapchvnVXuPGkYaCCbmVa6Fy2cT
vdiL974Bl8q/1Q8zS26QG5ft1+qnbV13gJv7BHkaVWyhGy7gpQiu188PDg0bU+NT
ls0q3Nu6afu6Ir4pIS3jXH7pgNgBkm/8hFvIyHmZxx7DxeYX0kJkKIUjZA0baCkz
byEnh/p7RtEcDGSGAcux0PVqXOgNSMHrq5Y2Rc0edzJnx13PmFhklGZzZ80TpYVi
AwcKKGW5/Xs4KLoE7DjOXcT0n8lYnPNTHuFi29PagQ31cW5k1fUa7sJy3mqSQOyu
HFArXzLXz714dSWX4HNWSrgMczOqNc1NtQtzllwwzwqFpp5BRRtmAtNyAXoK3SD+
W2xpP1TaS9i47XO84pPRND7CQUExgOlzbNUZG4fLuVC+gws/WyXM7GghJJQsO66u
RqIwAqXTdZudP0WbE8hvR5STPmoogqpGSgVB+AZ/Bco5B/hkGzQy0tma5DudtICr
KYtzRfnqj7u9KDkmpJ91OsbEQMPoblryh5V4e8EVuwFnH/tl/A899LyYUhYDwhrp
NWlzoBubRMYXscaiNuZloJKhNsil9DgJSWMxZu2w9lC9ccxePITsRzaLf0vD1pBP
BOXBTihtAKRcXp8GHcpYgz5YpiZmWA/nYb4PcPEOVApzKP+tmOqUE14xCBYY37Ka
OFjIghf2BVNhME31SsITz3yNXMKZcaTpvreD4d3kXQJpZeuyG5/Mo2BXxUa7d0x4
0E0PaG6K+/8CG2YVIF2LLhXuDD/vX3iSGcHXwfEI47png7rSx/E0wTFbVcJn+9tT
KOe/ds/+ZpmJR9sccz5eOY1TlF9m2WmGgUTyNTTtMHQrFr03cmyl2y7/QErZFQ5A
odA2dbBgwUec9qrz7vp/o/yjvYB8qyOHP9cY6sZAYCUpJktcWl0P6xWSffPNakWf
7sYvsazy4vNxCBPMlHdc/+xhIeQLKly+dQpN/LN7mkJ9zcW3FtkGAS2pq1P7LGrX
yx7+5KeZD8/Tiog6RZrTQWiVO4Incjl0m12W/ljW6hyxG614NP20atUtMpqXvLsO
yP4BafI/Bu0VfxVAy9/NO977k97navcKXqswE/8xShps1a+6y0KYQNF+XV4dv4+j
cc1gJajZdrmgPfiLBw7YYK17SDjMiAtaJQhLkvczD8ixnYn9zjaHjgML9KAphulF
Evmese9Xavch2uQAaSdm+YmX4gS2i9POSI/2lpp+oTFgJhHPIX6dUcGUpHE6Gl2c
GyrDZ2QwZSgpoptLZvgFnLO/DXgTdQ+QocrGoNINlJ+rwUefrgEFCi8af9bnOYwy
Uxme5uw4X73s9FxSAU596sXZfiHDLSPuKORoDbgQ5oeBUVGTXRdF/2V3GUmlf7Uu
ZRf448K/a/gys7bxXYZ+osvQS08D4u3CjH9B3r8Z2ObIOpPFMwCVDmm65JuatMEy
LKJoqXRn1NsP6J9n18NHfwYoqPm9wH5Ed5r5DCCyLNI689/hYnBd47qqn0Dn65sC
FwXGfWbrV2XEXVs9BBV5Z1T9wRpetQe6W9oL0qVt4lkWcfCLmIDpgmxxdYP5WDzF
iHHiuxOH+TvkHeb3Wl0tcLtjLxdYy4g6rbf2DP5EhJNFzeACTBJ3ZFvCg9WiX2NW
1rhyOKql6rCYsLCKKRtDulp01JI6L/lA5m+otNOkE3K8q4QjUveYu0ucEVi/wW1J
cHiEBoF7FyDTvkifKfrpm4++X0+qIKmuWkA9CBNOLnXF2a1wRLQYGNY8+cEffycd
xqDED+Ml7qN6IvnrCbW2k7ymfe6Jn5xzJJzTwa/3edj7nnk19+iO647/UKqeuRrj
Jl4NDv4CsoBWfaux3iy3hAsyiyiqi6LPvWyBhOIlTjz7WkgjrqzeaWL/EwG9pZNL
SmDMSFL0lDZCi/Lo57ivmLtctii35TaTWUPDicn4XqVZHf8uOdDVcONR6DOk7tPa
M8T2lKxpFZqIXmVaXO+Fmg0ZswzsBPaXpLSuD23ImdrvQ1zBhmR5HUo4bgKnsYEZ
ju7SAci7x5Lmmzzp/locGur3yfHVZT3sZzDjg9SuyXH5Qh8I2FH1gTLexls+SSg5
H/hkQ5l5v2hMn3L2APDLY2IteVRcbgeElWeB4Ln3wcVf89wNT4cL0ANnvvApa2U0
n0Xq1s5IuLbLW+2FAS1IKWE4GoBOv8/VVuLYTRMwmZsfYyIO7gFEYtcdG5lRr7TM
KD0XIoEd4G9SraDQuP8PcnZsfBXcasnigbBqHAtiRE6ADdK6RWQRIR+FHbebhO5N
2ZcJC7gfe//mBdXT0WIWNPGcAiOpieqrBSkOe8VOZ0oLQNjYt4HBd+Ly914AIMlF
IpeP18vipff5bwPWXiHYJ7prRQJgQ/g17LKmKuUtGsaLUV1xHc/J141A8ox472zg
rxNPBWu/567/7DG9HisRiOx1inh8AjRvrY6oQ6fqDa6Xs/Awu+FQbz/1FJoab1hH
VnbIsQmAk0Pev0HD3xFmgmfLCg5Ivpt/o0TVYIkp+8X33iwxp3tkE+kZWHnAgYZZ
7484XwiET0Bru6DsFk4Q7SnjJm3hVoKQa9jBzrFaBQGOYIchGOsBnFgebl+KiuJ3
p+xnTUEpioEZnNrNCAtEI6LkQ+2iKnL33aFuI31LYTIutKyUhdktdkoZKRkAjD0h
zqZgshIWgmOIatV5toid33PiENv1L7naVLn03csmhNfVS/DUZJUa1R9nYJVlumq+
/3txivCe1Iv8L56aUHLUwSOcxMPOlY5WaXQ+ayE8E7s3F/jJuVWjxYniVQXBt7Yi
iwF7uiNnbKgr4iyFxsE5Qof2iudzNub2yAuD3ZRmPkfQSk4Lm3YZ89FtLAwOwuNk
bW3k1xWTnUwPuLCIep8sgooa9W1pdjy5cAkwwZlBBaJWiVYNYP4E2RsmeihRmmYN
NFiz9lbOfUIHmawmwbb2y5gwj/lotZawciluUMaI3dx8xBz1yNVUW8+b8nTAzcjN
f15StV56M5ADiMgCa6AA+iLMj3wqcjVtW1o6vP9iuEvkCGoO6YSXnl/aROTXxJE8
VH4QAeP9J9/qdV2uu8RdYzmefc2tDrIJ0aQzUalVttAoiMuNNd1afTL+9v1VzA3B
iIqtE0SEcFeiGN0Os8f7YjTW4x6v0oY28cDeLIivEwaTvHCCMjonPlDz7aT/wJVh
QUAMmO6+QCZv2g7RW5Ylpfn5J89sCcWCuWdvVoLGuVlOiKfe0GSWsnfZG/RHQ5Xw
HBvTFRsSSunUfIdZ5EfFoVaTKuefQcyLk70t6jFWb0EgZ+Bgfj5ZhxiDczVdTvLM
1O2pP0LOIe3b5vfiokyqNL/oOfGUte7bg/APeESWuFfdKwHmGGEnqK32GrdsSPz6
b0Chv4Gk9Hdjcswvf0L85GVpzsGbbvF6EQanqyMoWTm9qFsgFAX8VQPfn1DoBTe3
zjmDaKtW+dqNBVHMVfFj3qE1X0YICZRpSEPMlP1w8rwAoJMHhFRpbv+4kAyPncgR
2TFkNOm1uoGYokBEIBW97qLcu9wi5UbXWvV4NRILnYPgIvq0vsQgyfXt/LA5uzJZ
XKP8MXhsPTr0BtFZKjS2r4HjpQtguu5QZU4tTurCl4yHQzovo3wMICe5hjuwKPu4
CWR0UceDcFmrujk7oMZYGr39VL36kzMM7nRhYGXYR3OkLrFedS+hGOZbQ5oqPjs0
8YHyyQcelt3ViDN0SIWwVqQ+qrgmLIRGT1Di1w2UL22Wl+ZavZXoVM2wm+Re0Gbd
9UBPWe7PG4ApC/uROvFpLX7iCuQMBpm9Bk8zPjv0hlreEkYcIHuOKKlrp7Ei9sN0
+AHGUaKvp4jgfzu56LE3HOG3tl5BjoNgM0dDIBRS2w4at5vWcshD2OFloScxcrpp
x88Ol4t+BlvykWit87MEabrZBw7cGZiZ7Fyq3yWO0uyBjRB6/GqHS2B2ANshI3go
5ngWiY53Jz0ERowjZrV+Tgb8V9+dy2PVs53JA64vLPHwJZ7po2Qm1GPAhSCs6Mm+
OWBPjpZBHw1FBpoQnLgs8i9t7VdNXW9BXovNeI7dcRBUreaMngIKv3R5qVNhBIZ6
SnIdv0YDF2uIwNx8QpOsYzYI6hi9pXSoPDZGwS3Qm4SuWiZSlSXmJRl7Ad8IDRbr
VtCeCym5s8bJA74LnW2OGWJsPuQZdlUmdsi7ACZLh+yxTc1Wb6qHmKnaGNdgsM0Y
Z00183Kems+mg7AV0YeSsaBGweXBEje2F4t+gx26lNnbjns6XUPyOFymAMSCPLmZ
bo6m9iMvwbRZ47yaPXlQhqk4HCAs+icDj6xTGCjvqQQlnEDLLRY/mthli3ayKsWj
/ndZNtO/pnABWpCAwd6QZ3SLn/uVpcT6EHgtJ9G3M/F5+i/PgBLfIPKbkJZ2WHaP
HVveU5NPXChllKpLCUpJupOAoudbV2KIemAnnSSxccBJY7uTvgjL8+MQ8NF6fS5G
SpJPg/8r9RA0xtUvGFbdDgO/gGRr4SJtMK871uPEJHSOb6yoGkN4kPgbCq6vW5wJ
nhyEfXP2KlakARyy+CSnQLYiYHRbu9zKyKFdwf2oQZ2jKRMHTb3E1rQH3Xo3PIra
m2zuKLQdTzv2rKY7KaAo6V3QgnUKusep/t+QLgjcMCzKJdhLGh/AhEmyVcPZDMjG
Tn0PKyRTvRpyH2l/qsOLO4x/dbbVobZxutJ0B4Ekjws40Z/4rakSMak24yuB3j6W
UrmuSxHIlJQ4PW4VxpcZX3vH2nCJrX38p5Btd3YZJXBha4pPw7HN+VGodWCpgSUS
lqV68+PguYFZyp1+6vJTZ5YbOZpyOx0h14dgFnuxR/cUGCxV/iYu3JqM9vmQGo47
FQlq1H+tRsgum6DaoRLdnbS6Yp0zremzeyQjjgFMXyMJ4P9HdfkB+vAlqxufDOQj
VmSgP03Lw2qvRg6ro1jxTGeyeziAifXPa1M2dbRu3K/mdlXnVgmdsa7TyXDqw3nb
m1mZweT5na1A0ce71rcxH0NBcJBxYr5NSJbgao44aRZA5oQMqXvudp3yrW08gwcl
B5nERCHWADRV0aTNSkC4of2z/jg3wguSvh6lRYM6CJbAQY5gwNJUp6rNoAGg2znC
vEf9qpR6vLHgtr+XKBZjKZ0REQq6GaoMdbn++WsMRdIiiTTt+ecIunrNuPPGx4Qx
aaOxgCGJJKliuxt/SBCPN3nPBuPAwDq4eyceagOckTiOTVCCDA66GCK6sgnzni3v
mS4tT/fYlUwpVEtQJ/l2/8m57N99iK3vIKYVi1YSk/Su+GuipCszvzZlutB0UDQ3
9NrHWUbc9DH7UBRYVUj3ETC9MVwA88TcbjuNGEfJ9AamAxj+RSWuHjKKL3z4YZ37
8OuT2LvCvvBZfuGXdNmWeXzzKSDXuN7nmlqT18n7r1M14P2yVCGmCNPW2RA1IntJ
VoDO+2F8U/iM2tocueut0azGpdPivMv0cGmpaEL8lfD3xYNMyt5Ub085mr+wsQ9A
ea92HXrzoGBUZlaKJsb097V6zTADa3XFPeBiRDseb6arX02BBXM6TkkVtRWDbggU
xG1SGsEdUOsNjkIvMEMEffyLI9hEaoTDKo1GlXclOXk3xeyQgULuC3oqfEK3iNPn
WZCTIAQAvsccIwii3viMCpQ9hvvGEIvXVE083ai16euZYJneU4VKzIv66bVh6b8Q
PryEKrEVGYbiwiUpOevizSmArl1YGBam8ogtbVaDuDqftfW3LjA8PmmtSRqF0FEu
llKIx6L80RMqDFrfZUfLw9flWKnAROXvdM/etq7He3CtehK6YyH9gWrwrYGMYLsA
S7UvPgsAfVQL32Yv8pJgMu8mzXsMlRTY7jqM4Z9NswvD11gjni11mFNMrk3pK44A
8+piAZ6eD3CLR1Zv9ZG4To4C7tawE1qpmAxTXmlKTuYjW5rVzyl+I7FMiF3TyS02
4Q8epWsJGHKp1kY5xf0FZE8KWK/o2/XtcYmF80UmKPbvvOKISTa8h+kDomKpGOqJ
AZzbpF1tGRdc6KtcavyXVMl5Hqj4ZmSmRvOb0VUD+T7iDWXWqbK1qdzzHG8sJtgN
o2fFUxRUrwcWJ++MVpjmnro6R0fY8eqUR/JuNcp0WKeI25G+nUhvvah6FKuuSms4
W7ihtvf/BBGlcOb/c9LmilEjDmQWaWJbAC3Dvs1ZJA3ac42To9+1EwhrXWOAhlQO
0h96LZ1M/effY/2zq7HwyKVqLodADvNwDw8Xs3jNalVn0oUc/UqOkYBFWMDk2hRq
F8P2Z3WgqcwCrWd1K4Oxkvbf2Y9EkXsJug3PSsXXqfB6szg+fQKhHs9hMJNDOFZe
SU9RoBT8oCkzPCS2+TYo/lx2DdT85gPheekB9duoBXnFtO1tNP7d6IeH4pKtssnO
e+5Wg/U/3UTQqRGoH+DSzYfxgLtOxqXIfK3N1OsikUwKFYt0D6TxzMANkSaIaWoC
V+3wwlVqtLQpM0KgrQ7HleBpCvU+IU0JyufPQlmjQel+uShhZFWq1f6e3WvYJ3rM
WqOCQj7jWnLCNgYPn13UIqta+vH+yrOTj+HCGukVlMUjc5WGUTw9nF4T64aKdfge
/kdDQ7FscWv4tK9AzZxgdg5K01C14Fsf1Pto2Et3nkTDwM3mUAcUnRqP9kUfloQW
Og0yOPS8Xu3Mt3o2V3HWM1Bzjw37vMMJyjhM12m4hKnxwKdqXuyZCzEA6Xq/lm6V
G3Fc9NOtRKpibkEZU2f/TO7FSDEGHSKO73wKk7GgMLFX8tG0P77GzkADLQMs/xwO
7UsR954o3y8fbTcuzpfmND3urocJ706Hi88KCBbTlneGKDddCPzJq+liCXYTxonJ
DRrGUFfDAxKLsGZzEPeeZ2Y4wmKC2nNocrDGI4IYJVgLc0XRlgimhMZ64gOnENeR
4X88UFGxf/gQFivxizKvEuDrSbBJQKiV1Z+434NsMbffxULhhsGpm7ay09EnmorB
weTTYPaX9DOIKXlOITLRqnUx9TCl6bdOWzoFTEm2yYnAlkY618v1MVWogFjH1VBT
IFybX2VuOTBVgIPkSs0PIvHrnf0Z9sk5a+BRjITvPrk+r7rZXmHfBS7rEby3IYsy
gXXK9/CK3I0uZukUuP3mNzICPasQnJG37vo2H/PL2PUub7pOiZ/o3BDF3HFEQrBb
cwYfqVqRN5Z7mfUuT6CkYnKnvwrBMrm6NM4k6fSVRtJLidLLz/Lq6w38HujjMZsr
aAIr3LfDIDP2slQUsZhe0umQWgLvkF2G6B/78OdLmJQPykmgZPBGdWlvHXGucxUy
Jp04t4tqOtgapVAzplgy1OHgC4e1w6Do19XFVaGBnjm/vdGw5hLohJPjFDOZVRQe
HTltVHhKZQ5oIqq1ILUfHPqy10KjfIyd3PI5TEoQBqcmKieQxO+IrkL6ChjJndhC
Yc7eQcyXrLtefzJyPnh/SfapC1vd+RDiG0+3re46im90GegfU4X8A48dBmwrcW+v
eMAw2GtzXzkB9TImAddCX8iQ1wAkdxxPf7mYvGN6j+m3lPBKgjJ+zgWZ4LrVsvgR
M3exHJTENPDfbGw8Q/HhLJavvIV4Sy4ka8s69kxts1+bBBQUeFltfoWFlGlG2ILs
SWoJXlgk0F/A7W5Qtt79mdXcJypWOmdwT/sS/zEQI5VKHO5jQ6/ld1ZWec5yxcIy
xmcDz935PhVKOsrj6rZK2niZe+hVN/CWuWA3AQHA/EOOILBppDMIjh7jrS3NGBNy
VzOdRtR+RMuHnDllhfAri1tULVCKa04DHqEcnRIto9yYEfQl+Ppe3x5AQVZwpntP
e3PhrwT0Y/dThcaHra8CZaISglzet4Lx+xy4v1/GQRNnTzgPLyLkSAZmgmcLCdxl
wRZE2zflFeUpYFAGv5s6faTRInvn1/l0dK9/ZRQEp54LQCJd03BpZYLFaxnLVQFo
jqiRY+sOLWLvVmyNbBOY6NzgIUife1n2FlnzOJFsop/K3JZxWV8bkde/9E+1e/g5
hbIuDqOmyvJhyPEIYP/8dU4sVVq0FJOeqDK4ni5mmLYNoL38KpTvATT9qn39Qpz1
xhTAORiEgGha2MxMDb3wqZgc1/gpJKKbbbqMA5UNVESHEzh4KLXY+LSRqVp82kYq
KBu89lGhgtTJUL+wo+KLTRuE9aqT29HlVzdwMc9yi0DIyIR/d2rdioTMQepRLWu0
m5whGg3rCaF44vWY3auaKSIH1wGc1PiVD+Ec5Ywerz8AAtbkRmCMIHYLDZjisdfL
wghqtun6dAvfwcZ5SXJxWO5WRk9EMCx/IlSbEwMiGOoYH/PvQTYK05SMM8nA/2IG
NDMxyFWS/W31fe4Ts6Scy+MSry9eijMwAA1Qt3VcCSId4PKLkOxlX3byXgWKEGsz
t6NVvc0vhRT9RNDjdPmd7kt4LMk4gpngVd1iEDeekDV4MnwaiU3558o3gje23mM7
zZ16lhB2NKKU/KFEzoo+nnUdt+tVwG2wbygdA9rRZjOi7hG7c8jrUqcyIgqWqzDu
fukgakkz4KAcNLFhel7k1hvDxpbwK+feFfZgwWSsvzgILy7s2KE5n3fI40q9udE5
IW4GH1gng1MBIpg4id/QX41zKaMjFEZJDirEld+iGFQfKkURbfBKFzpg8M9S6v4b
j1auP4XJVGxdN65rwbK3zMRBzUtSOUBcpuNXByj+vQR7WoLCyDAwkv3u67P5GFLk
+zu1Cun7EZLOyRsTp8Z0jV3ghnenF8YnnpuNggrSXXAdkyn1j1kqTo+hAsUV1eQv
EwLvovys4k9PbAijDiUegt2jm5I3yGy8g7qClk2mHSMAxXEaj2PKC473Yz7EsLbA
`pragma protect end_protected

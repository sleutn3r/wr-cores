// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aPlxWNv5Tn++K6OlyiZzgFTvVlEDhlmafc60bo0xDOF6x4y16wVodX8ozcFa3SiB
zF+spzJCjp2LVXcGLa77JBwfBUunqxB0pbVCCd30ZM+pSuSXeEByPBuPD6aOjAFD
pbI4pGjkL7i1y5n+8x8+VtidcKWFQpwvnqak5jPQ2DM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
Md+P+qsVnaFZCZWJfUdmN7ES3WD1VfuSK4mmL43puCSrb/3VZfyb7R0uLHu5NPOs
LIPmHgVoOg4TetyLa5isMlXDy12sf9/6fjYv8fd0mMuNxgn225zO/RN6t1ErY9Se
qPW1+fgAr2MRORb1CmFeDDRUiCQ8LV5Yg5fl+GuIpsa58Qbcg4MwkPBUp73vVhyp
M0HcnXRFoYwdJ+pRq/G0hh7ISiMNjp5zekfHVl54vghfc8QmiTWQGXxE+06XKaxc
UGNvfPOEKuM+DL8NTPwYxxmNfs33UJLHkU5pA91dc4by5wdPHuBoBQrUxD2beQYU
3N+vBCrILN28Ch6bo342MdMfMR/RvAdBoZDCo6A0llhSStPjbSVgW2AFhjspSGlA
pR33gerhAp4PrWwPcRl3exGOErlwa10LnWQcjUUP2B0gtjXGSWoMIAAINlfMH5Xk
0BoaCtPS3ggFxayqnvvmNKaqjYa7bXcu5H+kRBKB0jqpd97KUXymG4JCZIEX6opF
9O3m/VJLeSUV22yj9+zs1BEiCt1jNGPcn9zT9EqoSGHPLVegRWu76SbRwThrg7E7
qnNXcgv0sDnKpIM5hXfbvnSx+KItTq77nMSzB4pd+URjmEHsJ5d5TMHQB0PMrgsK
ziv7hyqmBNypnlZH9GIQDLztr06wPG4fNncB0BpA6eKVh4OOCrXfAxr9JZBTvHea
DdC2GVpDBzul8Xzp2SeLtvKj3+u9+0ELRpWGb49O8tIh8rL6HVPogdhacw+Euu6u
5E8rC1Gb7d55lWLTrxThTE4dmYeBPA5unX6ukduzOUYuWJgvzOFbdfbkhTnmMOu1
RZGwPiQB8tstgqalggJGOs3xmheUsYdoJf9aa4vIXU2J/MXXAVOiF1nJzpjoq3Aa
AvK36iHg+oZTvQJSHmwnzjleEhaUpMuP9ehYrLQjqzACfPgFqzzRJZURtbqPcj1k
BXm8KQ7Q1gpz6ggAyPjiMKl03bLDjDhoQWl5W5Oa6IjEiJynPdlMCFkFWgmKP7q1
RPlodSPPQmGKNUUNxX9q4TggOwTmK14tlP0tn07QyV59hX6JHCGYLUusRiQSLrvO
TAr4G1tS5VW2VK+BGHUxWQBCuiCeTKZ5tIjTdS+wmnseCNagmAO/YJr76h8Ri4yL
fSaKrsQoowfxH5BwpVZwingNdCDK+3TM7I9XS2Wq9wv3vtRglw0W45njDYz84di7
MyjQyaMF8Pg0wI+LR/AiOkeRoVJNWtXEjGjglXrTAtEcavqZF9OHYDy3MX4jQT7Z
EPCXhcHFaDN3+MiE31yNGDgANbtgkQTQVNbo1d8aU7QaYuQIxFV7rzFwsw6eLApw
0j9PZtGT2opnnQ9hQsNk3XoLsuxQ43++hUqSezLWxWfO1Yz0/JGI/OO7y0OuKpT8
Tvho5YoqWqq7hKyTYUi8Nc9EVOc1XVmsJFXj/Kpr++F/vb62ejsC6Z6VNFx/xTLi
Emr1zxsvUmuPdspTzkSDuJzua+7GK7j+se/L343SH6r7ent1YWZXDstKMto8Fll1
jQtmroqOLh32YgyfgSu1Kkr8uJFQxVGQPQhmyYjHbxuarnmVxO5uzjNQxFLoMeNm
bnLgpL9PChnx84PjlXW49b3LLz/SSC65DE8qyRuLetFIC4/zkUdqDSUf5EAUe12Z
VI0JEC4jDotct4fWUYJI5XvuYqA5JJsZ1tyFvh/TxET840SezEwk7UT/2TBQUOFL
mAqGD4q0U6AV7IMIoIEsWyoV2Af/z5anAIUEP4PCGoQIa4NxlYh5d1ulHav1AxI3
Wpn325LkOvnHB0HEG0/u+eQzGg+ayZwx9KYVnh+dWX9eY8ClSaQIIKyAsx3AjEx9
WNC5x5hjsPhpNrLVavykgLh5pDKOrcPhxfWxxs6LbXj/stlEmg319mLjkMQCxI3Y
y/LXkPhFYBo2jpN/U6s7niunh0lW4Vp32aOUhOiYLsWIRRbFPNCKtYIhp89dW8Iw
XaN9wHeIW0avSVOzIox6KfbrhdFbo+h3621281L01XRO8zVN+NDiP0l6Tw7e7pE0
eRNFj8DHYW6cN13OGGPEF/bY3c8F9aguuLEToZLF25OLINdyHTz6GCFGkdhDM8d/
SoPGa4rfrdk7i8U9K374ktPaMuq51m4kx6Uvdu5gHkpTBwG7VHg0TqiVVs0SYjLO
f0FBw/0gcpL3xLfPMf65RgjLF5T7gf77OF2ESL0zECRxr5f4K/kkluXa0uvPgoqW
k9ntKqx9ls1cgZ7ZMuLF/IB/witomcLr4sud7Sy1BqHG9vY/qEyYXfPv3l7GsDB1
KwpyAMtWakTEaz6ylG2xsFlTGzbPl5OYNA0OAtQe6NCrCVjKrXtiJx7Tv39oV9hj
Op2zOvcGV4a2km5Ku2YgV819o5bRiAc9PnVDKoMVCz3LS0jerlRvK792WkArU6QU
RNYqhb70MGv1VHc9eUdlqqHeJq3hIiZzN/QKjb/1WtpSAvBI8Mjs9UC3hp4JfSe/
cd9GuJXzKqXzzfOtNNClsHapG+XYLQsSSxWfZq0BLsV5bZG89BQAVdYj9BxRmDi+
Pf59f2QC4bZRGM/Eu4tz/bETw/WjUwoRk37vyxkHGPIbf49KkezUlFvdL2WaOIHU
slEIJIJAtAX67sL+wt97cMCiNjAsAaCcTgXcXTW8DuPUAjY3E9kQ7LCPuYnziWMR
YZ+zp4c2/hIUcmKqYd4BTPBxt6A1aR7cftr0ezsNEC3MtO82AWfinbRiQEpOOtDM
Weh/WEz5L3ELeFIObVqiAxsGPnGHObAfk5M4dwqdVVLefqND40Nxwsrie+zhAVQs
ypXEQCvoUL83D827LPMZzuNYBA6YifXlti/cExvVFDagfNAOBOoyFg7BRMC9hFps
0xMKDJwu3cUDbY//p6OIQBw+daWgEAp6C5wbmfGBvJqq4RzU4YTPVGSsMBclxVOi
3ald+oEqo+5Sop/p3r/5/pwe2F6YMtV6kj6qJDGpuIRpOGx6doYDAylAp3tQ4Nlm
cIQRgcoSAqRzYnmMtlce6InEjopg+Ae+fT99zaAIahrdtLvNdHZGdcdJXpE6yyY7
1kvzSdN4JPWeK181/GRI7RA8moGLAvZLOU0jdGlo8O+rxCrdK1qZusx2hlgArw/c
wSZpUMY3hFMH4IKq/uHokgfB8sHNN+/X70chU9auQBLM/j8iFprD4OCzfOM17mA7
up3CQZzo8uTNj/xaNQpFELqbl0r49nuJ4n0GVe4GzfOE18RbJP2oNWkIQbf8nt/4
3VZPAfh2ZmFVd0gWIxYt9udb5SwNZUGh2/h+Zy3HPMjJ6mMYPAdE0gD0DTOhPtdG
TI0vzXXC0biC9l6+kFhbksil+q7RGkvbIyp0/S7STHgrXlY7i1sOiBGKCv/2lx0w
huFecuX1agZfXjeXzXejwf8Rn8rhkyzNnZ8cGVkZMAvaK19Qbg6nh5VgVTBib20j
5WAYGWkMsP2/CALLpXWc5G9JqA6IYVtGgLfQfVW/v5RJTaX44yL3Ll2oUh1+a1Jk
ZTnGXzyJn+iNcgxagfRnPuXnrP4PAu+rG6nGhU6BvXrHFaN3wZrBGiJwSOVo7om+
rMriPTJQx4k0AT/5LXxMn0FCILLC57Ym6uv0RwwrEVIU/hDpSPccy2hPV6fUGvHZ
HLYTXMwbPSI8ZzClMr2usAO912DR+YX3lCIVghdEWIKGEuLKTA+3bVTiu4dLfPED
UvGhw1Lh8tG5rGK2IrbSLYpdAvs5Bn5qX1BonIEsHwMAzhGBbgT5FxHTrftn346v
6nDvwoswpf85Aql7H2nzi/5DfR1KAVLUhemSHZmJD32dh3KAMpp5Vk2jgR/64edQ
PMtZ+994iylUKtnghjog88IozdpngK2njobdPIBCT3dCD9vtXD/nanLuQsAkDRxZ
4G3ObRKu+cxzIFDLHzb0gD+yG7b35Izdjx0vKDwXdzF+sZBTe/6Oj/KiIoLMNJQD
89JdMkaB8gbYLoqYjiwWyxTdz/i3Hmaf4I/HY1IaA9xUNIrss3Ue6D5yr9Jz3yaY
ga5JgXrybQAdej9Im+4y0xdMaXNBdFbUt8N/zPtZOcoSGRR4BOzxYp75wPCrxVC+
MGr54OhcoW3TQpBxoDemd1ohtCPC+L5wPkRaGnaSssN9y1HEyb5Ig/lHIWFKJQXc
is549kGjt/mp4Of+EktkoSlqw1lXpJZI7IeYEkEfOpSmmWBvtpc3jAs5+V+RfsEw
hkA7LDYgfeRPj1dok7xrRp8E+2BCsCXNoDHdP4kpSo/uGDQTBRQo+/tYerMclUha
Aqse9Z9EvAAvO914xEtg2oI0OL11m0h/ywUmXztIPn42WfMFJTKnflmf23wI5Jnu
Ko7NtaSAN2RMOIzNB0cyjxJFYoYGxgCNsjrFpToZNWTJkrHpJeMMDnaAVYmVQkRF
TQR/brvXqMVPaiosNUZLDFeRNK06DagNNpS2CkNopdO5fP/1asR9UZEpNEMcm/2g
lFNLy5S5qA6rKTVNQyTBg8xyNBGFvyrJWF3HHLPPZn7TVgwJQI1FwIcyISe6AIiB
n6S6QpZqeAAlznVVWyQfJ9lw4c3mfe+g0yVmBWAY91LAPOUa+xd9yYz2e+oFOIBf
93btn0DFv2gt1+kprl9xRnic3XvhXoL/uPnDhANcD8r5kjSbnKQ627uhWdLmdoy2
6I7Fd1JVsJR9OfZL63InDFBTVhN2IVvxQQncDibkt2sqoGZrnyhRbvRZ1Cx62aob
eSSiNvaeOlCEK85Vn/HJanwYlOLwS0hQdd/1B9xzb4lz1D6ERyUKvsBGYSovSsLy
Uyt8CxVpuHar2x7Md8cqpzIrezbLUcijdoYHACTe0Njn6VJMwxkJH/rLOmUmmdKF
hYKpmiuKWsbFSiOnkpi5bHUQFa4XPj6TI4Q5i7SjBZDqtvJulwOhvgXfDuJX1n4y
fvVxlBeRC1fnnw28umxqxdou01FXMGGP2N9NenqHT38sOxK7BdOwYUFrESBMs7Qr
iXofNBFrVGFFWlp3GvBDTmRnAR2JU7BLgBdbopFO2ku+QkhwuOcyddN0g6Cg1FPp
nUR/ZWAer9l/e9PjRJDDEsLk5PXYoHPPfWmi4d7AOBhA/FivG6I0MaW30REaslFK
L4olnNslixAYrDJIxBhHTtXsxeB42eqb6+rcq9CLKJM0FdrWUF/8AD6oeBQtb+KT
u1lPIEkCwtjUWbizkhnoDj/ZKazZybedPkn1r1H7nUYVCW0+BdpXbPrtacrFYfGl
9yiSp4qxtoo7ZKU3N/tlCScfptkXppvWQtT6s6A2wtToX+P0Zi0a7h2KovETzU4m
jbripETWcDu7RcXO+1yy2LHYzzGs3csbmk72vzvWE7ibjSR9Xp5nZCZjIiiE2g5k
kyAqmQiD4CTsgucLYRH1ifIJGFkJ7dZoVFKcSJy1HQ278B2OC9ngY4GjIRqZCvPT
Z/D2reTif4aViyZTidTYsgIKwmlK4ovsrlzaUeaBa1LXPV3QBLGj1K0/bsko2YdF
rv+tlnE71C77IY+oYZ1slSbuIyXcDdnY1NN1s6car47b7RQucPe5CQZ3FcRg3FFu
7tEg3HMVpB90r+5ZbuxsSw1Ofgc7DNVeOUQmwnuiWunpNHXgMQ+UTIEuW/pm6Ick
N/XbPi/ItgCmL8NGsgIGGIgZ3E92+AiTRaLrxKVKSQJ4PPI5QtvxsWWuX9FK+ecj
QkuS7eyPgVIS6CIMzmgL2Kfu3PkqUifdAw8cxlM4gKbOtSvLfVznjQYdYZNS4dip
+/7mrmsDsKldZ0UG79VH367OC42xL3jrGQf2FneiAZHChzi6hsZT2YJEuk/CrNvs
jBwP05fhthdmy1syBTrb37x6pHiMsMiXNwrgfwPZxnBdDJ9a6Js5SqTxy3CnAP01
+s1cG4CTTTjjkjzrKxCbw7hj6mvsZzs11U9gzWfem/Emd/74k+nIpHYW/h0GG7wx
Up3yGVoZ1hLL3mGLUknQBIBhpBUlwi43ZyMx7Z5r+0Z/gIfUPPBSSIGMBZfuSO2x
Dmxnm3jBWsu9m/jUm4MYYSuaR/D8Y7ZsbQzDkxOv50CWerRa4NMwWb6Sz6ZGaeBT
kVli/AJSyUVDFjod5zl9y/CoeUvVeAwikjRFX1sO9E8bnHRMHvHloQSAsRsBfu1K
T9nr4WdrnlZBO2NyI2D7wIyk8Y4+9N9HPEwJwT0TPPXQRXVTdlBcn3EWGV3gpUF8
5OrHEAcxTolGYGSPINjObxuftBR8WeGUrKMmEhjiFKcQ4NelhCKdvnGsZ+fxXbsa
5LHC+0L8dGTa01R+Bt4gdDIJoS4c/k8wIVcCwKGpSjhciTOQpft5s0IAWN7HriJt
d/unMmRzCpefgbIrLFu3QCRliqqoPGsLlkTE2SA2sahvK92RzEAGBuIIZyfSlzYX
ZIB3LVBEL0DZ0rgYxLyfzlBlw56wfmcEE9ykPd0CT+TVGFRvEhVZbJd3KnJ4BaTl
1F0qjJXJ/c/xJ+QbdbsqzNNMVqXGUK1maqPN+V0vD693rBKsCZwfynHeg7z4Dvcl
wNSTVWiz38qF3krCc8GOsQ0NpnYvqUQqNeWm2d2YZHVBVsQ1b2Wq3eb6JLFGRwQA
DY+mzOCj3urNjXSDd1As2ucsZ9F5oKU94UKb8Iob095s5iO0CdE3hGDXmefp3sKZ
mFKfhXDR3h08OySuXpa0G2dVF6gpyikGQeasGQp62Rt7+fo3fVUDnTk61kIeJF38
AQuVq4bVTYSfElrJ72G3DX+RkXI/gibHNAe9Dy/RZsCgS+psR126HdsBc+1XGAKU
6+6zY0DncnmRdHlEYsyOh8S00cCOLwJylH/PlMLB+sk2886mRrd0tq0xcA/uIx6/
A1L9dn/wRMHONHgeupUrnqTEUm1dKeuMnInVNJ8wWdEe0D69sV9Mw2X/plNJPK1Y
RPEXJfa6jfuTXtRIUJru+l/wMwh0R5n363QUuK2Sm8fUbGhOF7yJ9yEFCtcVwbSz
U0LRcH6hiAA0r1U1H9J55+RF3gb9kVvGArTFuvu1MJQFW4zJVNqLPHXb5OVgMPOW
GnP+mxk+PLeY/vy9Mt/Y+ESSfP3KRXNXu2xv18jDhlrYI4fKaCRg83XLALPz2tLN
9WoZrtT+CXb5yr5c5Y2YpbFcYc3vZfz7NuBQeMd3/T4SHNK2NQ9eNNfTB6fS0VKE
5NqPy+oT5JHpUfAAgzZyiIw1Dm3nePqvbACXCCJv1H7sjrGAcosAyWQ2K2hAGUNQ
ZttLQ5BTtaGbziPKyAOXO7vgy0pdNCAWW6+MANX+SHX0oLyE5gTXMdXYyK1NNitK
cM2NccgVKziLtHLoHU/KjJoBHRJRoEXOOZb6YbXdenU=
`pragma protect end_protected

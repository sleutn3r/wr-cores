-------------------------------------------------------------------------------
-- Title      : Single Pulse Generator
-- Project    : White Rabbit generator
-------------------------------------------------------------------------------
-- File       : SinglePulseGeneratorModule.vhd
-- Author     : Peter Schakel
-- Company    : KVI
-- Created    : 2012-08-14
-- Last update: 2012-09-28
-- Platform   : FPGA-generic
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description:
--
-- Outputs a single pulse with adjustable delay and duration on a trigger signal.
-- The settings are written with the Wishbone Bus.
-- The Whishbone Bus addresses are described in the wb_SinglePulseGenerator documentation.
--
-- 
-- Generics
--     g_pulsetimebits : number of bits for the delay and duration of the pulse
--
-- Inputs
--     clk_sys_i : 125MHz Whishbone bus clock
--     rst_n_i : reset: low active
--     gpio_slave_i : Record with Whishbone Bus signals
--     wr_clock_i : White Rabbit 125MHz clock
--     trigger_i : Trigger to start the pulse
--
-- Outputs
--     gpio_slave_o : Record with Whishbone Bus signals
--     pulse_o : Pulse output
--
-- Components
--     wb_SinglePulseGenerator : module with interface to Wishbone bus, generated by wbgen2
--     SinglePulseGenerator : Single pulse generator
--     posedge_to_pulse : Makes one pulse from a rising edge in a different clock domain
--
-- 
--
-------------------------------------------------------------------------------
-- Copyright (c) 2012 KVI / Peter Schakel
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.genram_pkg.all;
use work.wishbone_pkg.all;

entity SinglePulseGeneratorModule is
	generic(
		g_pulsetimebits    : integer := 32
	);
	port(
		clk_sys_i                              : in std_logic;
		rst_n_i                                : in std_logic;
		gpio_slave_i                           : in t_wishbone_slave_in;
		gpio_slave_o                           : out t_wishbone_slave_out;
		wr_clock_i                             : in std_logic;
		trigger_i                              : in std_logic;
		pulse_o                                : out std_logic
    );
end SinglePulseGeneratorModule;

architecture struct of SinglePulseGeneratorModule is

component wb_SinglePulseGenerator is
  port (
-- 
    rst_n_i                                  : in     std_logic;
-- 
    wb_clk_i                                 : in     std_logic;
-- 
    wb_addr_i                                : in     std_logic_vector(1 downto 0);
-- 
    wb_data_i                                : in     std_logic_vector(31 downto 0);
-- 
    wb_data_o                                : out    std_logic_vector(31 downto 0);
-- 
    wb_cyc_i                                 : in     std_logic;
-- 
    wb_sel_i                                 : in     std_logic_vector(3 downto 0);
-- 
    wb_stb_i                                 : in     std_logic;
-- 
    wb_we_i                                  : in     std_logic;
-- 
    wb_ack_o                                 : out    std_logic;
-- Port for std_logic_vector field: 'delay' in reg: 'Delay after trigger'
    wbpulse_delay_o                          : out    std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'duration' in reg: 'Pulse duration'
    wbpulse_duration_o                       : out    std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'enable' in reg: 'Pulse control'
    wbpulse_control_enable_o                 : out    std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Not used' in reg: 'Pulse control'
    wbpulse_control_reserved_o               : out    std_logic_vector(0 downto 0);
-- Ports for PASS_THROUGH field: 'Stop pulse' in reg: 'Pulse control'
    wbpulse_control_stop_o                   : out    std_logic_vector(0 downto 0);
    wbpulse_control_stop_wr_o                : out    std_logic;
-- Ports for PASS_THROUGH field: 'Soft trigger' in reg: 'Pulse control'
    wbpulse_control_softtrigger_o            : out    std_logic_vector(0 downto 0);
    wbpulse_control_softtrigger_wr_o         : out    std_logic;
-- Port for std_logic_vector field: 'Pulse busy' in reg: 'Pulse Status'
    wbpulse_status_pulse_busy_i              : in     std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Pulse active' in reg: 'Pulse Status'
    wbpulse_status_pulse_active_i            : in     std_logic_vector(0 downto 0)
  );
end component;

component SinglePulseGenerator is
  generic(
    g_timebits    : integer := g_pulsetimebits);
  port(
    clock_i                                  : in  std_logic;
    reset_i                                  : in  std_logic;
    delay_i                                  : in  std_logic_vector(g_timebits-1 downto 0);
    duration_i                               : in  std_logic_vector(g_timebits-1 downto 0);
    enable_i                                 : in  std_logic;
    start_i                                  : in  std_logic;
    force_start_i                            : in  std_logic;
    busy_o                                   : out std_logic;
    pulse_o                                  : out std_logic);
end component;

component posedge_to_pulse is
	port (
		clock_in     : in  std_logic;
		clock_out     : in  std_logic;
		en_clk    : in  std_logic;
		signal_in : in  std_logic;
		pulse     : out std_logic
	);
end component;

signal wbpulse_delay_s                     : std_logic_vector(31 downto 0);
signal wbpulse_duration_s                  : std_logic_vector(31 downto 0);
signal wbpulse_control_enable_s            : std_logic_vector(0 downto 0);
signal wbpulse_control_stop_s              : std_logic_vector(0 downto 0);
signal wbpulse_control_stop_wr_s           : std_logic;
signal wbpulse_control_stop0_s             : std_logic;
signal wbpulse_control_stop_sync_s         : std_logic;
signal wbpulse_control_softtrigger_s       : std_logic_vector(0 downto 0);
signal wbpulse_control_softtrigger_wr_s    : std_logic;
signal wbpulse_control_softtrigger0_s      : std_logic;
signal wbpulse_control_softtrigger_sync_s  : std_logic;
signal wbpulse_status_pulse_busy_s         : std_logic_vector(0 downto 0);
signal wbpulse_status_pulse_active_s       : std_logic_vector(0 downto 0);

signal pulsegen_reset_s                    : std_logic;
signal wbpulse_softtrigger_wr_sync_s       : std_logic;
  
  
	
begin

		
		
wb_SinglePulseGenerator1: wb_SinglePulseGenerator port map(
	rst_n_i => rst_n_i,
	wb_clk_i => clk_sys_i,
    wb_addr_i => gpio_slave_i.adr(3 downto 2),
    wb_data_i => gpio_slave_i.dat,
    wb_data_o => gpio_slave_o.dat,
    wb_cyc_i => gpio_slave_i.cyc,
    wb_sel_i => gpio_slave_i.sel,
    wb_stb_i => gpio_slave_i.stb,
    wb_we_i => gpio_slave_i.we,
    wb_ack_o => gpio_slave_o.ack ,
    wbpulse_delay_o => wbpulse_delay_s,
    wbpulse_duration_o => wbpulse_duration_s,
    wbpulse_control_enable_o => wbpulse_control_enable_s,
    wbpulse_control_reserved_o => open,
    wbpulse_control_stop_o => wbpulse_control_stop_s,
    wbpulse_control_stop_wr_o => wbpulse_control_stop_wr_s,
    wbpulse_control_softtrigger_o => wbpulse_control_softtrigger_s,
    wbpulse_control_softtrigger_wr_o => wbpulse_control_softtrigger_wr_s,
    wbpulse_status_pulse_busy_i => wbpulse_status_pulse_busy_s,
    wbpulse_status_pulse_active_i => wbpulse_status_pulse_active_s
  );

wbpulse_control_stop0_s <= '1' when wbpulse_control_stop_s(0)='1' and wbpulse_control_stop_wr_s='1' else '0';
sync_stop: posedge_to_pulse port map(
	clock_in => clk_sys_i,
	clock_out => wr_clock_i,
	en_clk => '1',
	signal_in => wbpulse_control_stop0_s,
	pulse => wbpulse_control_stop_sync_s);
pulsegen_reset_s <= '1' when (rst_n_i='0') or (wbpulse_control_stop_sync_s='1') else '0';
	
wbpulse_control_softtrigger0_s <= '1' when wbpulse_control_softtrigger_s(0)='1' and wbpulse_control_softtrigger_wr_s='1' else '0';
sync_start: posedge_to_pulse port map(
	clock_in => clk_sys_i,
	clock_out => wr_clock_i,
	en_clk => '1',
	signal_in => wbpulse_control_softtrigger0_s,
	pulse => wbpulse_control_softtrigger_sync_s);
	 
SinglePulseGenerator1: SinglePulseGenerator 
  generic map(
    g_timebits => g_pulsetimebits)
  port map(
    clock_i => wr_clock_i,
    reset_i => pulsegen_reset_s,
    delay_i => wbpulse_delay_s,
    duration_i => wbpulse_duration_s,
    enable_i => wbpulse_control_enable_s(0),
    start_i => trigger_i,
	force_start_i => wbpulse_control_softtrigger_sync_s,
    busy_o => wbpulse_status_pulse_busy_s(0),
    pulse_o => wbpulse_status_pulse_active_s(0));
pulse_o <= wbpulse_status_pulse_active_s(0);
  
end struct;


// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KNnX8jSW86gHu/gxmLaOW9+I98qfIhV8YckzqWS3QX/eW/gbf0rkggp/KbHo9Z72
N6FM93q2eobrd8mxSvf5P1iS/EZgTYhIO7+vA8n+6oNhunDv4xS7WM15gDQdiC+a
2s9X8buzwobNRtrSqQfYOm1N0yBKvSq+SqW7IqSYKQE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5200)
PkuKhA5YZONpGaKKDNViDmjYiHfl2jG4DH1DinSBvDp1OEIV7AncYd6L/+1FvEG2
Or6ikr2HM4Npb/R3vItXCEt7AkkQXQPEv88uW0D99xP9/zVZUF1EuC1UdTNo8gpr
nbjNFgwPesUM9M2P/wBJYfUqnr5wGY/aumjJ0P54zVhAZ+FLF3A6R2dYG2LbNg6K
BVL/l0drCyfmuXWBkvUuq32obKTNytCmpLUYUFqLv+COHAXThdLnZls/i050wX7d
wcQvk14qpw37D7nibm9UEWAMaiEuA0gBEiT65rZh8QUFc6vme9tLeBl/HPd/gq0m
K6sQvq/yaiqUV4QuZMvj6lmpZ7oAI4TxvSWgkKouPAica/pmrmmPdvIyvRFigbYO
QtzgmH2+Eq+6tF0JsRroHciPAVafI0l8fNB028RykDR475HrtdnIZMUwK11+Y0Q7
VNWjdSTQSOi7Y3xuUvIerJFAf1B1vtCtt3Ve/lidZPJ104cYKu5Wz4/AQ5fGvMm8
5BwuOekJ/ysy9ttZGFWuAfuett6gJv7JCUYUOSsC/bEPptzYaZHMKAShM61pkAkc
JAFTGBFFNG9S170ZibWrau+wySyDdmN91bnPZInjSC/q1+7IFWL4E3LNN6PIaEC5
n1iiS9Rt3em+gzm3Y90IA3OVZ+LkRtE1rzdlyAbrqa4KdAwgxlcAhnnK86SETDMB
oKLDuOqKnl7Osjv4c/N4RiXOkhZ6V7F9j2vqRrniOuTuaxU4m8rzM6LAKaIfk3Ay
ds5dDmYCdgJUfOXexulRzcepzWTLfC4GwMR5g44lEJ1peCR0t9+7vpvDZSLCcsLS
/oLsUZYNCivzo1KAxptkqgCkmK1itdBzMgDSF66EBiXku3zT5Y3ROQHWtHPqyeqZ
1IpSfJRXbdEcmeyG/Rirg+EZkfkhKl7xc9nzfqLkAtXwFMNnMlkGhDrIDHpXi6HT
RNkjCBcN5N5AlvJI2XgWacq//gdRyM9wSQ5OEETZOfh2YmN48C09Ssw0j3WA5dkg
DxS4OMLPrqkKlNPwZNl1HcTsThtDmhpnhM3vkHXAbTYm7J2BUFRexxMTc3lTXPVC
P3P9x7J9t2Zwmo7QuqfRTWGTXtax1ZeSi2d8Ru0YKzkIovI4ZuVW4KDYbaG87qJn
c3pBw6+XrFELJ5hULzSvCW+/xzVJ0YCxmzSPSceOwUWuJblUEO7FCKgcRg9tMGZZ
0jj1fkLcFJwktuYSZXf6udopYvIQuztNw5tg48y5eWFvg/YROpmKb62l40Mufa+l
Ztmpb3TRNQJyd82mApH1KDrIBDupycPFf3pHlpipqWGEHqOo5Umj9ZX9Wbzt5h3U
2D/o2SIwWt9PE6RvfP1SMlV3Qg2DJ4Yed/9yqcwYbFQClWr5LW8O9XsgYBt/2QdQ
7Vh1jK9lmaeaEXiCj45RQdljbNO5k7ybbO+3usiUVD0ooVVfLAx3tFulMiEVcGHc
a9BNgtnUv/YpWsGpBd5KKoL8L71SrCf1HuFBh0v1zH5Fc1XNz1aeacAGzygZC7VW
g1oxXovaF9srUmdPWLCZWTt/goZSLebJ6otXVctoaVZmTdBJRBURK9Oo8iCoc6QE
frktMuUUmR5Ib0u94FeKm1QHaKQq10Z/RaD0py+nPsp9dXmHjeHkAoAdR3ASPkHH
Km+V/NBcwTGBD+up4wsECAmJiXUU79AhXrOFvdb2B5W5c1Cw3WoF1gXakcuknA/v
2nlv8w6a7fi2cChsCPC0CzYv17b//1a8vs0R/8uOSGYXpoyx2UPg1y2SeRU1icl+
sY2pELmO+ZIcaK+yrYputFSYUBzGJILWV0srMaFwI8B9QAhkEw6kQBpUVntMgvGY
kSTwZyCLgKW3GwwZ9eS8Hm0wGDg6Z2A32wQHLM1wJPIoC54EYnrsF+TmrkrxNDmB
9xqtbsP/5zT/GrrPch0+WIWP3Hb6MJyYo9uM45umxroVOnu9tOqneNcGyx4hOg6+
BuiTookBt5SUkSBr51O3fdwzQcexeA278OyJFkNR6DMifjuIfkohY8cSopIRQWH9
B640yhNLpnaOtzMGudZ/abW20LrzjrNX2/BtvO1HYvqfQi/tBfp0pLlxq39RyXNu
aQxH5hIH3Y1mzqVrWVJsbtqM8cSbmB9L+japjVpjG5UUog3PY/mT5+pJJZIha2Ni
AqvU/Oxh016dkfBtVjRRSPVo8ygSO/c8uv4Tcz0zijLYs/xBfWu00N22tGYiMH6c
XYya3x+lK2zVU0JGqsG9n1EzZvkd84NcOqXpd7NcsGpmB7VVY2j1rFFOJvvlmW6A
VXpd/aup/DJq8QzI0NUZpqPBnM7g2FHdfZ2vkn37pL23ERgBHU8GDza2RUI2aBu9
eToIbWeXM9KbHxqP1GiOlYPVeaxGLw66Ufrw53HEyMgyW5MEDBX40LRXJWInNMGg
2saoyL+BD5O0twS9k7NUIcP4KDU4FJc9NXRmVGAH+la2/TgIm+DFvbmROf3S3TUC
6LenY8pzVpYMV51AC46c17PPZZ68sHFrboRHJTCTTS/v1/j7sItBafZmoDpg2CNU
6RKmEKCxjgVImv+DU37AvY5lJQ6gPntymXYBk+2UqmEGvLKLbZGjggKl2N5ZM7y2
u92X1I06/YtHdl16cJc2ar7Z979U8S3Efd10eQia211XKFx8lsCvPdG9382SVPZL
3GdxTf9WWzdTCNX4YDpiWM44CSTRCTF1BjLYvebQcFE1IgFKbsvAhh1/dE9+HymK
uXO2mS7qdWFm1xl5NAQ675Amjx3/jKpEi/2KtPgAfGD+kXZQu8VIC3jNAkfua3Ze
YdTuCzufcrPLIu+7Ms9P3mjEsojpQ8WYVwvSuACmxWPzJTLF/9n4NyajY2YFmfYr
ryArvYNWvy1xIbGN6knh0oIqdhAPSWQFWXlOLop+gG+YAohoust8wMeWxSfzC4wL
ZBxqbrdobOTEUMgMmq8vH+PFzn2q1x7KHEFzz6Wn3Gs+jnHxuLKcANLpkFNjyV6F
1Dnydcy2Fwp7kkOH+qlz3YxoxBTyamkcJVuAaSxQFu/a2NlfpdnCiTw9FL1PSDNd
9NHMcg+bRKs93ZhFDABWNtwEwRIzuRcxdwFycb4h3aXQau7Kdbz3iNRmd4uL+En9
S/tUtjqcWdIeiKj0N1FqnAUTKSIpPJ0CL2RcGTEAT2t+oM2xhwWrigGE7S9oijcM
6I7eob6igFRFEoFiIKBgvjnyeMsomhcr5iEAsrmVtzyEv5fZtB/qSTIRqn4wyNi+
EHJI73URWEpi20yYpQWIfOs6slTVMdiBAvgHBKHDiuecDlwDWFsYaM+zk1oWN0Y6
vNnytvMgRajvtl0x7TXu5v6nmmMuj2pKIDmQx80TPZm26XyGRIuj/zbx+k0orSma
ommCo5HPHnCyXXNlTmt04t/8gOh66ct76MBlD9UgFwOE931fcWd1ZugQ0oQ41t0S
P7bn4lb+iwLlgo/Y3oSFaODW/ssunPsWmAmUXerAtMJpahL/PhUUN4xi0JrH7BNE
hpvzRJ1mQ5Ax9g/EIEEnlghOTSAduIhNs67gABklx8fhnb5axF/CAVtJkw8JvMV/
uBrLWBKEO8gwCxndUrPPIYeAGDQ2fZIxUhFlytjXS1CMyN+LTTUaOYtvuBfSwlfy
EHnauJ1WA1UMjK3DDfXqJIYQsEOpQji2wuOo+LN6bFEEQ/pk61ip3tiZj7f6g1A4
fzRwiyUq0PW6+SGLa47LrfvExI3WyyWAOVhmViSMAIcbOsGRD8TJZ1PYFo+SB5/D
FDDSlB9poZbg/tWS9aoTKakEWQqKLrPdOA280EO9lxtXPl8aFxSQUWESAmPaHzi4
5uCschP9WfZATROCkKYVrU9oD8Jxxln7MsjqRY21x2wW85435lu2MyEpNBueUzue
cu9TS+b/orgmGWGMCw/N09Hu5AtlSZym4aoUzK+zzDCALLKYQKkc9u/YaSZL+jGT
JALw1A9zSW4QNrL2eFiuPJHG3+97HduI1k+CDPW6pLShwAOPs0kDM2upAyqJrmiR
K4KcwaHb96+9cAnenCl2f+D5z7RK3ZHKJwnwst1fxzTkPYDwxVOsKScCC3b0BREu
ULdayUofUnhthnr3gg7q4CykWQ1DoSjU+myaJEdDvOlVQsTHBJOlSGesnmufwyM1
3RYBnIYJVPojpCNbFkOPlAQE4RCcIK/r3VyFbekQoqJJceguDvr7QkTGfdEx2Uk+
nSKcvZVjkArCuP0c2aMtJtRDvrwk/MqvVt77UZ9fLIPWiIHtADIZDLVOn415zn9i
VV2h2EXD2g5oeIERIpSah7byzk15LYnAtwENNUaOqpUXfahn83nIJlPxjJ0m58Fn
Rw/nQKK1ZqHaaJ9iwv4Q/dqWWsuyfvFUasSV1VJ8zZjBvT8LrsA6x96oaf2kfP/u
gkhRYUMqn/ovZphhVJowyUPi85PWslKs7sdt7vDGGXBYfNSS2dypJncNTlsZ85J0
OchZPRCj08Nb5nuBm7pQK59+4csqfOgDMZFnFFVw+4hK9qMUFvSh0BNNL2oSfnld
SfaAAmeiWVucWhK1giFGkGQF7UO+n6LZHEkfMeiFzowM+QmvzluyBLMCml9jTHO3
hVYAHrJJyrgLpbQ5BDSzPFZXg+ZUlukH0eRi5zJPVfcR1LNWscSSN1zkEil02vGc
qzWy7L538i1wQ1zn6Qoh7VXaJ5KXPok4RKcro8v8Z4ns+YCAw1Qp9td9cs5BsaCI
N+rsS+tlaThJ3v+PDaP18WUNrpeUyU5+8kSwaFZiAPRFOoOOoPtq/VQC2ULeAb9v
XZftpFJ6m348fP7oP9F1VlErPhClS04EzI8X3VL0enuwkfwfHWfYCXSM4lw1IQuI
dHe7rD+oRDpXyO0fRhFjCKpow0OA5lc6Q6nBjUHm1Z5ghe4KSy6+3mcafi1AMfzs
t21NYrVarh1iVeFjV/6/+Fyk3yQJQWyWDC/EyjFwf5QlVWDEEPRA3ioyIKrn0i0Y
HPeYxeisOTQKwQP0162uXJnHwUI3QLniFDggWe1AkDpDky0Pa5NQ6EKm1DMWez87
aBDNIpIbnBnVbgbEa3YdImg7fHiMBluSK/2dGgQxjeZB1oW2fSqO4N7hgX5dzK3p
p1mTmIieHaDN32ip7enJV9BE8d7s8OPgBJmOOHgWWi1/awKjtoIdfU4hIJ+q8C/P
tV1mgLnZWdf6iFDgc6IpG7myx5VRCUvmtDCtL0/OOLQgZDL0eBkFz9qBAIIGPqra
OAhdpNSrmtS1Cgkp15mDAN+1xCodh8IN5Lc7Z6oV65Fi8jZZFoSyqeXuwwffsyrz
WM0H9i1sIBt9tR5Otcu/XWdUbXj5JnX3pErvelPBA1ITgnss4uUDLszphsvfnD4F
EudEULTLQfp8yHe/CE9tzGGyxdnEcfhoLkl8NHUGNcLIUL1FdPsbfrH4LWR9/DL1
hdGRJbhLDMaFtV0ZnmvysVOCq8pr3BaQUgU7KsuJV0hwMKh4VrkdD5338TVQDJW0
5EyeZQIB1mdekkDPLDnRs3N2wZxKiv4tiAwcVl2ftdEa/nBRwt14MzpF/GklJjkY
PafPMeiiq4UTSW7EloNKp4eOtbPkKtcR+OidWjpiax8tG3sUjkdSNSc00orB42Qp
lG5BzqTqALERTS4IxyBZDOEoYDq8qp9BHbzWT/UJGMZP8BQYjjo8Na0A3tCgVWA1
D+CvL58dOkDLD067wEzWk8vAXTQ2xEyBoUzaGFstd+aYf0gIdRHpdJ6RrgNRAUOr
qe0BYk4aoICojylRLxCO2JMiInHeA0jKiYE2/QbQNfEPINe8TPMDJZvwvZAfBqiA
S1DNOcqs34E3t5NgbQ0/+t2FMnVXPnbLZhtrNzI3OkziYXQE4vwPMLhBgT6HaiwD
t5f/1hsOVgYaHE+AsFL0chopszg+fgz3/OASvAAPTOJZrX2UvmtLHnJPav3yYXtr
59ANm4a9j+jURGoPkhSlmTqBNZ/azksEsvXadTHu9iUjeneZ2CIrsugndY3nZ4zk
T6q21gPVlTOhkbACTiKPVpXJr2LNzd5k7QKQviV2i9PJtoFfvglrcEg/rhYZl0sc
svIFB70Q6t5uizK7T7hWuRMvQj4HhOIQOWazYavLEtqtnUPGKe/E/JDrYbbIJweT
X3sJtP4WSOZU1EvoJ0M64KhJO2bGnaZn1vBRCnFXDO7vRvThjNwB5KL+VuycTO1q
VhJlEswvCP3TElofAIljMWPBWxjSGxP7DI4MU3CUc7MBFWiNEi8ATt0z7/oi4a2H
sHqGji3vowr1dk/hFX+QGZHzugyMI30kGAa9YNUQx+rZx6L7a1fdz/G3Ylps9+dy
AbkfBChx7YDp9W5Cs90LYRsvH8OpLxNI13lAu5ORvUz1mAk3aXef6uw/BxO80MkC
mGpCLTk/vWXpBU/VoJoCrWu54bbP409Z89+b1a+mhKXio7thKAai/GNWTorhCLCb
joivjvzQf+GKJ6EF0N5B82elLhNOZD/OdmXTBPDEQpg2+b7R6VY4otpi9YyqNJeO
qJpXa3ZjXLOzLau1gpFUD9q57ZyFePX0CjqpwpTVsWHiMmWtkKoNy8mhbEpTrk4y
TrQD7fR6jQ6K71fvTtgfjpE5DT4lxo4gDoCxC/zbrOcs1jIZflrVTVCCWiZjYVZ4
b+kd+sJwPyESxqcZZryjaqzBiacbirosDg/57I+aY/JmGBlwS1XYx2t8lcUyAgGr
P5zUoBvTlWyCQ2r/HRtOV9iMytekRnzkGzY8aixSYQTYGR3iybjXcoOvJRD94qhP
7wo0DugjIu1BjQjew9NymQzWGsmIJdIK769ciYqyA6f0QHI8qo/M22qMh1GD3d7T
F7A3R5Wt6kt3/2ia3+XqJaxn3MntsWnHO8g0F5+4uN6K07SySgEaB5KokzAtJXtS
NyAbE16IRDErdzEfs7F9ZA==
`pragma protect end_protected

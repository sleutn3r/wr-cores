// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
heRDTR298Danq5cabwe+ADyTO0KScNc/dyNrtXu/7UauhUe5XqEyvdeBcX3+Fm6h
XHRe4tSAEOADI2x3wEO0mj4AG9h/AYBU91Z8LwoMFIR6Yvc4GUsb3TOy2U6mus9z
q+O7Ngh/DtQDjQInnDk7mAfPF8YgGf877cwLySMAAK8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22000)
ryCVXpungAn6VUeFq2+OmzADjX39RVm549lOrNomWpujdSTckS5IDi4hPNFWlClK
ttBzDV+t72YEMX/Mwo3orVjCc3BMvjtZ2VDWStUGe9UbUCiGeRdLSJIWeyuGie3G
rZQkLtiTv027pjGlx/Cl7u3rAkk5d2RpAS0Qf29oEh10OkWWHeZCSzzy8Lbs1t8i
j8p46mpyK68IY2fFjQHr97uPN6dZwsMh0Z5Ygi6vm+OPH5MmYBzPhVEDWq7aRmU9
CgUGYXGAIC87FF8cnvhVDBiFw/ystxxzQd4gF3JcslDWZvvx/MdjgNjRQ2zLe02/
ABmTRZ9RpJIvKIdHpGzGoUTPVKV8ljWwu/vRUZRGKtNWDqMgJQr3D0+vJQ5JPM8W
/PAgV4eDhtq9cdgzzKz6itbm0nimuqFAGY+YA6xB7c4j5UqTcQVx6cOm4PlJ1lic
V7EAxJgWifBHJYVpYg1FiQ6KKxyPnXw2/T2v66vP/1qlB5VE33iXKySpeB/7l0Gu
YdYohlTy+0tnnNz4ImIvt9raoFDknFx5DKhvJBcn+Q91oG75eZ3D04Kq09paZe+q
lWmMzb2+jmXgUmN47puPa65OQV5vMLcB5ZBGnGSP60t2v463uPNHzDH3+wPh74pF
CdjK1347ekzr2XFMCX7alvhrEFM62yeq/EbTZC4CwVj7R9dmmWu9SBqtMMlNffe4
oiT71PWjxX/G/jibRNm1QfpKhcMTbnewJk/lMHGrdzbYefxoi6hYzKZZgmDKnIBN
dWNqGgt3LdPE9ErMSfthhm3sPil0ynlLavlgFikcBA6CBGuC4xNH+RasMuvz8eMc
fkHvwvr21I31wfHdFas2Q+zJAT87SBxRGNqcLcoGMxDz66SIdBUp6/LZ+p7amfiq
ux52eftphUf7yHRowoRNq0md84/s6w18GEHv3GYojDWN9Dqyjnm/72pUzkQebmAx
MlPNNuMU89TcxT3mHUF+NaVRMmWFcy70YWNV2T0FQ1a9YwPCTZN8Jgh8RWSupVab
tRUtTiydJLGCXKUSinWvcZBayCozHxwyuoubSTVsRi+m5WMH+FhxY2Q1cc+uSDB5
yCj45z1TeDKlPSvHZnLsUvxeSRw+laoajXOuCirO3ApoBO/hXdap1LXPG79818lK
ErGhsp/FUXI86/KltymNsNfy6DwQI2qn2TErT+AMF+bDdAi0urlJ5xzaSXIDAYtt
IN0BSEmR0ePBLNFDKORezVFKOwePIwkye19IdDkHuqHW3OJWGCS1eXLy1zN6Nxo3
5Q8JAK5uoG1/dAZU+Dyg5Q5a0S5ZaQWOOozq7BUs6SD22cu04Op5fgmzRtr4QEtN
QbRrpPdRtHSTNajN2Y0SQLDsvCvwZxL+ouEA6YTVitlECA4ia+qsxrCdhKldjr3F
VFAS3X25ldfGdm++Ary+trGC9cjvebap9fhAeLc7QjF3t0VzcDROD6JxuE43TVU3
6jSJjGcDLo4YDB4rejBTY+fpZuNPQXUdEBAY03r8MiK69PSa0wg+4S6QMTqoFfwY
h2qyTMYezK56Po5SjP2YITnfrKZ35INiUdLoYVt7nH5kThYT6KcUpnwgd+3Pu328
FsdlVEBe+QS2VOcWIJiwObH+yTOOqoQwQKayZnCMMt1K+bUM9CyodRH8TgKdD7VW
vxwCOqw2xlhcyQ9wZyC1C/Sh+Jlo1e9ng4WnVQi+zgUPmmxkCsEFnGiumMQiNwGD
wtECi/r5V0PTmLNV/o4rXCvXM2AN0sQXZfGfOS0Ko30YMeDStR+WIMBWihIuoEE8
rINzip+e/ntZwFGVQQ+V4cfM06JKLH6QJSwgHNfLC1nTHeB3nVjfqeyGooNlXjj2
uhcUs79kJoGtR4FFJ/uxC0n78fdm2Mi9vVR5dk2dI79b4eShPGDRWAeAhpJl2wQV
A/nVGSTWg+tFWELVEoSHSelgMacOevPNAj/A8xxtchRgIh+zG7bZyXyrIVkQCJDi
Ii80+4Yv30rTAMSmxzBMWw6Xc5rc55K71p0Uab5jJRY8WJ8T5Ags9r3oeMtWE30a
eTL4Z5aTJKoing2tQoW0UCDMGcjUySsNP/NTLDVAwkJLoZSffUiOlDJmcAWcTxp+
nrrmCBGYFcVBojPcSthxThPxXnLxLogKRzYqLlkoNt6Xe6yctQFCBd7pU3QqAgD6
CzjXgF+qco4Rol2SYsi7RmZ7VVJOdHejvGoBDD5mR6CnzD77O/rrb4QDk8qArn+n
R17FoDZZmhNcKr8qDV8/dE1A+AyHs0oC9CW1+YVZ+kby5jbeh2NevsA8L7Bhg4rK
sbxB88J3k9+iqsbglUxbt+LajJJq61bWLvzp1He00NpaRzGifCgFIIdHST4zmxI8
mz0Kw8Z8x8o0Yh5EmzSwhC+eL/dxpTsaR38CTt+lpA9kAJ82RtTLn/XYjb1dKSB/
6FZc7M0AwkFUFgGS/gCpZ7t2jpueiMHul5UIKIBnmseIt014HCIwtRPEIx+VFlci
/fBRyUJjCijpCe4syXcc6IHPqpFjyA04JjAyPRyEwPpzSZaQ4FMc260BrVwn3o7j
gAb3K6BjvipMKF4DwHCQwtQum4wRXQ2NckEpJT32Ncnq+r8Fpbm0d84/1Vt8Lccn
4KjR4kQIEJNfLrNgbPmPz7NpV3XlPZDylkrC1rs9UZbORQEeeQv2eBQEkIfXuBPI
g3uXaDKy8ISBVygjYf2jTppY2edz/18U3LS5wWdHOvBv1a+LHQosqt0pDiXF96gL
JbB7MK3OZ8kXOTM2bhTQWECF61vJcRO6m2ZaacogzSP0oA/qr5AuQvZSc5Sr/fDg
MvIVGkpz3Q8moDvQ9HFCDF8gFucU7XHyOCt4pwfwHzE3wsfiHY9vaogeUkOyK3Oz
4BgBYv5jxrDyILNzUGolEDV+w/rvMvR3ri3z6OcQ/B8lswgLWz3SZjl1GNUaUW1G
AyAGPBxxTtPUVL8dV8nHcvYq0DCEGrz7Pc7JnhDcI+1vhI88jtiGcTFEvfBf+tl2
w3UJuqZCD/+jfVXdaLMgmd6DZ831WBZW1FdH5rzebwq60slJolO+vuMVqaSz3cyj
Ip4/x8GUCiZzYjQuVh3uRJcsy/kwzW9KOW5XqP+C3YFNEZk9XDkvBFeU6PkCEgP+
r/uLFlNxXWG58QooKlGGfMn5vNO9Egm/l02WY4foSl8geEVrZSAlPJ2T5rqiQBHj
uci/9elxYU769NDtbQ4ER8MFJO+vU7RBkKA/WxwCoWOAZ4rsG8X2GxS5jMOXJVWz
VrsWwOfKybcAibwChcFRJkI5HNJtvy6TLfly16q626x6x0EZR6Mml0CuUdxt7UsC
G3dcidkE1/MLgCvzmLQFH8kMPr+CdsLhv6bhD/g/SQtCV0s3J9yEZi+ymXe3khG1
Oeu3HF0CWDzYNp7kPrEMqZLXZOyBxLQ6GwFJI7pBECKACFbg5mDHThDwwm2FYEon
eXvwXhWtT6YLWjEfnwvRBidF/ZbiiGMVeAwFuTMBlHptonRkvIquCT56cRwQB5Pm
oRErA08HIo32/3NjanWO8jzlcwTp3+siRS7Ehd93Agf3f8unjlI8Bj5bJRotDxOX
AJ21AlXO8uXLqcRr2WMo4kOUhGpvF3vLmRiVrztVa2hO93ySE0qLldXLhM19WCoh
5nyWwOIYT56JRt33eqdNTJwt1GUgg0lcavq/BS8HAFIDqSQ5Ga/kuvkcKQ1iM89L
X0UJU++aqDvllse7IzB7yzkrVVJxE2oPqMgn3lLYFCkXRpNSluH/jBPx8ShaQ4ee
oMfFXDrv4ItV8lhk8MSP+YW1UqL3CfjaLOQtLC258G7ogA0xp8fcuHdfEr/3b4iL
6iNeczgQd6cOvYsnRDoFc8vKnlKgfkp+6LrkZ61KFmgp5VRH7XWQtD68T7yDgDGu
NQwNBr0eE4cpeHZZI2oB6e5bCH+8idmOPW5izuH0JVYtKpMaJORf1yuiZcWKZzp7
4mrYMJs1hnmYvvCvAMETmVS8yV0vL74MAGGSte/ONH8q4KnDe9lqA8Yq9fJufg91
pIh6Fkq0EBvNEIPqCdQpkUacdSLXGLY5d9D/lIjhtAq8IlzWMAOZ7I7ZNwCP4j9E
3fZb9jPwhPUxnUIvz1D48CstWmrMGJ1sjVO8kNpTGH3dkuw2GCPZAxXeMJx0k2ok
fRdXvVnYBZKigLGdCRA0WBvJFxB7Tlt9ecw3dCTfgcXVIYUHYohscqKtqpQbTwMw
VDo4Wg9lHhgigcA8HwgCziIRXVYX/jSxb77rrl8vl7bz5vSjWn09lqSpoS3X7U3P
O/oTyxOi0GMIyQfSQBcWnMG1MMh8qhdHKSmoiK9LmwEEhxUsZrZEPvZPuqz8ZX3c
JiL/HE0ilroExnsEfYGQVFluG6S3ExLqCNK6BdKUYmn2PLe09BGiQczaJ8dCmKfb
Xruc+HHw9y3bnCCuvYM2ZT2H1l4sppoqGHCtnrnHA5DKPIAjxLStkYBFm6RepLQe
T7MZOvzfFwZTdf6TmIoQy7kfz8ll0nAHqwDAKdzntvw/KOm+t41oq4qr0XWJXry+
dxX25al1qVNCwCbiiaxGvs6+F+kt/FcAxJ3Yq6E5egYilAF+RrnNe0WgaFo7D4wB
w8drk6l6P/dcCWnIHcFjQWAMFnOiKT1kuk5/otPscFQRH+7ka73sRBlqQHtjf7zV
FgrrZfCjjK8bRxwVmVDO1JYYiKdemiLATEmSSlD9cA0T+XEVNRfZFV2T2dEi0zdI
6YRm/cBHNCL+iYk/Q22LIyDYzVOQhmsdDUWFLwPgvxXZIJLtgg/Iu0LaMXkksjVj
XLFgmyowHcHWeFs0eOUbN25X7pDC8XWhGiCVW7VZ6MPlNxURaLZCH/4wsF0n9W0Y
mTG8YjWqVf2WSQCu0ti2KC9ovHyKPy7ylsrbDqOcDJR4G3MKBTAMzeho2Xi8ZKOs
R9SvIydJpZFLDnCtm4FiOR2c2Ec1W7UVoDCP4Ozi1zI3mg7A5w2SD1Um1c8OuR4c
iogwUNun48+6zjzWCabqkzVfCJZSRKXSmRwVPjhCI3UyXW4ALyxeFCnI48kpNIta
yXWjDByjcdhU92UJGR6DOtABLpX2Vd09YI7bIafGTWcbc+OkD0NGvKdCWM3nVF6W
2qxvosIJ1X20jwdfCfVlN+yIoY2nIJ+st+yn6CorLW5TDWXMk+EJTIgP3yBHAkcC
jrvhsBvsEItLhwfY9yU4f4xLN5B+0ZEM+nBhuu4rb2SkHeYo6sUkMGlA3ZozPGb3
7wT2DyaO7J8FsoN36b2kcCMNDVm+OF4VyQXRAKcGUdHwha5QRFy6GylE1ntsPEa5
drD9BMZY6Qp5VSGwkuuKH9DwLCmWYU80hkyU9128CoFaBOsBDYFrSzGwcEwChcP1
XL63oNfVApNL1HELYeKI5Y1YPNYS6IyGi97EsaQDFAuo/A+4h36IhkKoGUDME0Vm
/0dG4SiKzoeJGH3X+lSed0ySofMHXXnBkSjWxcT6RM+Rz97GWXta1IfkO+HZg8SG
VQGRDe/XnLPTBwKHSNNs3fYHxdVpfqJXHwvvPfiMn5pGA4H03/TWkvSASo3+gyFZ
iqcNIvezyvvvNA4Sdkk9qmux+w8BaeQlwSnXBNMePfMJ6JIq/MlPh/5ps0po8pEP
7deJY4n1ae7xp/Oul0ttvvUzJT8nhsYgTj7SyX14dOMYnVG6W1CqdSHnZcmLwqP/
4A1k/fVznvwGpl5No6X0BhIfZ3aRPgyrwwrubmM+zue7nerfmACwkp9gZ4hDwCp0
PYTP+VaCilQWGbUl8U79h+bu/tXCDe7/kKYgGPsOw6Pgrzn7S7TiTG/KXqJ4K12o
uqh/vMp+vyf9Uy7HfwOmqesPTEasLJNig6Fys9oWkSR35bLtYOdh2uo2NbFKF0y/
7TTHLVZti+o9FXYFfzQ+CAxNotRGAcCCqNJRM5eGSY0xKtqDRleQQ5FnStrypDg4
/wUPGnml2FIoKtg7sqB6eK4U2Qf+O2YhlLM/KQ9nuwt+/e5bjFmAWN5hGoiTn3wG
xHoqG2Jsc3lx+koTtjEntoiKp570s1swlfp2O7CN61IXUZM7H3H5iv+kjxHKcBT7
OJmqoEbrLpodMJOUAGzUSpOwK6D3zRnhc6ja3QHUV5c/TolxGjy+H0tLiV+f8sr6
b3hu+VSOgGYJuWibmxTOoEfPKICFY7GJzZBSMORdRSV6AZsyWRMrbvLlolz8vVFh
76fCKW+qCTfw27f/IyqhS+wIAZdDehuaov1ifqaBwEBVBVLtlsegwzzPfaICG2Hw
F9TMQ5LDkShBUECaBtsBfAsVdJq4X018dDClHLUijIsYfKD+EjWsnAeOSjb+rZyH
vCgiFgaqeFDhzxHlkm8c6gHmzTaxWMO5tviw6lt2x8Kx5XRjs9B0Z7OCD03/yKM0
cS3tVT4pSW0Q5SCWg7vTfg3YJqNGM549QhtKDZ5vs0XWZ0hCrd5rckmFiqCUDbHz
1+cHF99ERoxS+8i3ULwuKBZhQONyEC6m2JQyDlf4WSJPhYSYMToCA/SUeKx4KIjG
2gLhToFvBzHsAfM5cXI0N99W3UTqUkkoUWsEKyLf+2yFuMkpoJDBNkZDs7s5Yyqf
XTbXSpUH4MPb//mZ7QK6T/n/OGNNLBclXNLs/7gR9DFts9yaMhGS2P+LA4i7Khgi
DIR8AQDMznk/5CMTygH5t0aIxHef8egAr0V3rpDkL6W1fkL+BFyI+fb7XsITzVaB
da+C1qHMi2XtUOgpTir0WN97lNxjeBEkWZt18JA9nz19jWejB5NFgpYqCDIJaqZ8
jofx6BSMRp7PTqNbTDEqkxG9WWiqJAn0rsgh8T+zQifWZceKGUahbu/el2Nq5+PO
7xMpPGL8Q1IJKy08cVxANRJu2zjQrTtNzRbxwxa7EmIwNrmh+6YgVP+PYZVBHtb+
Jmd6qIhnvWA9kpdwEzqCkwggAEK2foHL0zVfxjAbIAMrvsanJnWVEIcyO+LJTo1z
O0GKn+i/D99ZkgWcMBKqXH971g6gQXSNtBEb0kEFT9N9Sr77cnBx57EJkHzoPZpd
DssK49iRD172sJ1XehFg+JSM2/Xa9r7wS9+iBUB4pfZY0WVW55d590UTcKFq0qgY
iu4UEJrpYSqs4IZ8rq8qt9XK9y0VlrwJ6EFvre4yfDu23/RMEY4ah46JmRR5JYm3
28Zs9ucCUPLSLjfngFAdVp5cOQmQ007MmAHQ2DMxmwbXDDoPG88X+RM33NtyqHCM
MpQo7CX0Q7XvNI2zxVlQpm5b2OhLcC4s8+9+ANCJxaScM5Q+hSOL5MGaOX6prw1F
QRhH70uhI3/0AbFMs9pNxNyRt73Ccg0Gio5puaQRnZHXV6sysPHLpUlbE8+0je1p
f4Td1wRlkTAul2HL8kii+gFZ8IbQo87pjqkP7vF7oyieJ1NWt5sZmQHT30oJQK/W
TMafQDww4F4nnf2MnVqYnJ/clCPYetMrjSUNcUjG9mG31XzuQaknqATLifyXFogY
SZQOeuJdE+1Pm4cRsmms9HqCdWUHBIViGRWib9Fi4rIgwpjijNUT+KHvJLL5eWfC
t3IxEwynifC3OZU+4JC7cVTmWFZrSEpncZ5Ekb+2M67cPuCTSNX+WoCFb9zjqz0k
WbdtaZy9TOlitHwQ6jHwe5L3eizefU6Gvis9/5Ke3Wr5/EeDYlgfB6ro+PBf9jHw
JFp2LCbVM/miImC5wG1cRSzAqNqTSJQkxcdc5P31hMGqCe1Nsts/IOYJwAHGh9AP
Y/mjHW5eEsklpniOsmLTKKottZmQ/WVJqAI/CpszFbQrNw4MPZmZrpHcZrInHcgj
Mja9i8UCnIC/77pxyinttZ9dRS+FvvQdSIAfTYJ0s6h+KOaKt/n8dETUJWrCHbh8
LrCh1qNJfMun5l9NcDXXyEGeJnWcHGbJ3UNQd30mmHvp7EIPutYEAmKAS77t0gaz
/jqvutULH6cVklJ472DrQYiN+uaG+UOucyUQw9ibcg8t4Y/vOCYSb52nOjRB0UGx
d+K4QfbB9h9bCqeL7Wk2AtWmwdijp8phH4QledwzNrIBCjY6f/YWsvl5EOw+KMkA
xjolzM9rbHTIh2ybtUlMrlzGjpSQkUaxIaWRYJH4yziSIPF80l03+y3luCc44L3X
1EKlJcwo3IIHmiATIPUoci3oEvuZgcFiW4uGVyNcErt8xR3BkQpX9uR050wCTz93
9r78w9wZuh1ocUwfx38qiF8GBr+4v3qANJH6rCP4UnJ6f5O2+fT0QM8Zj4tttWTk
bce9whHWC958x/cdZ7IS6DLrVMw0SI6dLLcOiymrczl+KLo3tdZAFYtwUCabN/GG
jsXV2mKXSU11oGfK/j+8K49buUpGfNMuAsIEjbjsJBXYvJOJOAswgOAn3+TKfPn0
xdbAT8nE7LLYIvFnkP8vqq6Vvv5SQXYEqLM1clCIRu4W+Dpo+ztIjBttjP1Lirxw
v3nNjzdk4YFAfvQNF9NFG2zdG3JTRfWvzIgAexqRqUH3NMqJzhR5WS9qvIXXa1Fh
gGspIVrmZRXM2MlCWfIGyyBs/AF8QFEm6vNKTZEjuUO4Vx/YnEJuoQejeyA7jIgb
aJkyIgPr+b6kWX6uVb95d+E3EKKZFuriJE0qY2pxRJmOs9mEGunt0vjsnFvgam6O
r/9Fj/D2YSif8gQbuaBSM6UOi2lmYLR8sPim+RROy19oSNNn6F5Rp8OtLT2t2mAj
hrqXaxX3RX0/k8dv++U8Akffrjf/DpQ+redfKsEs/WKa8ZyYr4tI4ziVzaRbgqqA
jQy7y0GFVEdwSu3CpVapp0b+S7thiPeD296hXFiOJQQ9bUjwt+DajP3Pg8CRqCeM
PKzQh7trYVLIN/H0IUk76eAHzNWJThj+SQqpoVRaJlTWQzLYH+XfcUozv30ReYjs
wn5RLtZoEbkUjKSKr94zq9f9aXb9IO5G07F1CaAcR1dhEVu8EZi1qE0J0LMG4CMm
Ypt3PkBl4D01znQFEuZeGYJQou3BMnsANzyN+xDbGKLnvU7bep9QrvuO5AKW/wv/
TH9yiCddNiFk2jxijUuvtPQpp47E6K6t+t55ZfzI/T8a6ckUOd5gjcKR7WT1KYtV
SCeDMhNirf7qg15DpHBpwKei9b6wSSLwYmOqPJwtnmAxtf3l5I3brUftn3Z8xyu1
QhkMukJ7qfWu1dEfWs4CBhVQWXExQHxcH71WkmWJit3H6a3sarZDFmhtpd/drudg
t9dnPyf3R4gROvNXf5abGn5RPErZ673UZcOc7hyZSEEeH+1WzRkcY/ikcxdTEErQ
uDG6r7nOYsT/DdO9fbvl/b1sUHBJRIGnd2XQck31lxEMqcofHZxtOp6c1uwpO9xV
HVfocbcNynbZ23t+1VdmTeFM8FyRfAVXn/jdFS3OI4oBN9LB9bBOBLZydmt1or6X
je3y4dog7YWgLjTlHJbDyk+O+tmAN4e4quQC24qHv8u0pVqvRrlJAkTkblRAWtr/
cJOMzJ5HAHWgVsFRJZSfGs9ObPhVmsWyS1vOVDRZO9V6jYH5DbXgogdjnKws88IS
oHk4iZIzAqCVZbaaZRoniOnIf3dnZGsy8MIfeIoPPqZD2s0dxhgVvy0kuq7vG+99
k9DKHE6e4GyORNjfyb/IxbhA/koHp54HGloKRq751V82QTZiy7KJPaLzJpsai/7X
2HA0UnC0nR9y8P3lrB3GA3rOObhOmwR664amJx4vdkrKuRrO0CtkzwBK4D7fN6oX
XNykDo2Dygy2LgJ6AdIJGpL1ywDEUsJS9JU7d++zP/qItSekrUqkpAS2XuLCz40C
ZZtnep5qih/rudVuZJYInIT3JyA7r/t26UyYSiIA8516OJ9l8a1/dgxRJ5q6aKfx
BcuyCusuj27CbaI74asc8t/X3sFHynJP2FfGFAr2snrQPfvPuGcGQrnB/sdO+hHH
OvKQfD6z8ZOyzV9Tj4XmLuo0XHShswtqjOvSzqQ3GlaEDldbHFMFbuwPUEphOFoz
JxiB6Vl4CXwoZSqURd2D3Yb4DmByD7fMLoEiQlehMj/AI4FYc3XB+XV/vVOtC5n0
/QTRTRQW3h4egGcp/da/+jVWd27YRev63DQjh7iSizG7X82Z0c+ni8tlCb6mgMZy
wGtbZ7rnUj5JBp2hflXye802d2r4oJNrBLUa0m0E1x2TG6Qptxm2Zt3tsjtl2b7R
xfRlIXRxThRT5ZND/dZ96Hout0O5MHbMhTv5oQvM73DPNOcQjkNQ/zfadXljeRWQ
oNm5WSDoJ2vYYfrEOtRX6BFSsD3OnG5UHMH82d42O/iCOQP5tF/VWJvi5pmxbCi9
OdX8Px2vjeYMMDpqo9IDDLv63d47jMC9rG8S78NONc0jVc4hxCKS+uQefxjicDfK
7QcYXnTzMVUk60TAk64xBmiGlvsKhZy3ErEV6YFgKnEivXvwpCGEfssQ1GZ4CcTo
csA16JgR9NJwx8Ck6CREZiq8SorENqeazzDQ5Rvq6d+H7FxLaohO6nQsel5NK//u
EF0ZmFaHeFU8++b3mEsqQjqIXBNmS54mOIc54sE+FaND9LfpofobX7pX1E1er/5U
+9++NrVQolOYsnByeefWlR7jszkRd/zahSbdox2jI++Oi2vgGYkzKkLXUkGXyIar
FhiXFDHqBhyqVuIo/8aRh//4stJGZZPRs18bPzdgVMJ+mPcfwTOBoBw0iYwcfWa2
d2XGxfF0OcMANcWWfnNnEqYmp0/b9sE6LVl+uFTRa0ZWHbSjIluN3OErCz7I4Dcz
5YIbTUyW5CZGeaRiwoSCClysGS0PhJPd8uDI/atp+h91SIWYH+2hw91s/7toMxQi
BzXj1MMfiffYwvrLb5rOeaqY9aruvknzbLIV8fHysOh+tr8sw87XscL8+psHgwjY
KV0eK52XuiCWwIv+PdzwYhA3cIwhKBhapneuxSiylEkJmNXg9Eh+qdYfIgC52my1
qx+FasY5ETydRoCYoG3mPTPjGbNS1UftE4z6tx2APV7y1zG46v0OERPICrplmujU
sFHFnmAtknns7GsQbSmCpXRpVdfXtPjVzM75h44CxhXIXcQUrlakn718qX7g7rbz
WAT442jG2GhYuIPkz5ufK13zO0L3+zndOCY6Jj/czjzQd/A/blInSaluV5ntTfrT
X91cYOmJ5UYB+OrhAY24kN8OVcPLOzshuq1hlDxIEkniMq/CdhcH960HwIBnRf3/
lChlindwcqjLSNSrHaL8k6JwYz0iACS4G7y2GnSTnI1AFh0ucxCx9BzrmwGKzaqA
iCpSqkPviyxJxsdiZvnS09gnMf2UMHd+/e4f/4Z6mwhxX5TzEZBl5UTTjpRxm/GJ
mmjo23D+aRr1e/swlczY2zrTEbRTGciWChiOuPiJuNO0o8kBQQNkrOVMDwBuMr1f
PP5Q2j/OVYsCpztUv8u+PCz92vWhv4cEKRU+J1ZsAR0CLIzvP8cdantutcnKFMCX
N+t3YX0cacaG2YX9tooM5UbfshPFj7wJDWMpBqLeTUsjkApxVfsKpXYo5ZcMHF53
Gk3TjJOXdUBDume3Ou3Q09PYKKe9uvcr3yOsHpxvuExy9zhkdl82/cOAdDoJc3pj
iArAR4VQanPWtSw1VlaM7H27kV0ysH5AZKeoUFdGyt5uohUGcLswU+/QVN+gOHlP
XqzCNgx68p+BJr4bCNYGew62T+kku65moHxa9JRhF0kY0A5DwZ848VQ0gXzoZhfx
1JK3sCwEtdRxtfU8oELWlLbUny4Luq+AYXq9tcWADSMucL1/aXDJ8LM6TQn1YWiT
FFUe5LRJLbNqS28uCqN70JD2C96ezLwe455Gaq1NyvyGzZZ2Pz7uJ0yeSOaT6XEL
hUA6hs937S5oSY9ezdQuXIlyiR1i0meRfaYfh2OXnUxOG3V43jHLSYFfxkuBQWNn
i3Bguk3cOveNCiR2sOwEMuhc+lsgSZd7FQtNeWG35M7VeucgkdAtkAxNAm030zdV
scjtGYzXKcQxt0/Jvk9cGZJ/zthS/wHJWlxKoIjGZDT5jtoIJBadQGcel0cXx65h
D+pRidMFD8pZ9OF5DAKatCV+5ZzLxcIp9Vx+eEljMhn79FTTNNgvNv1GQxIa8i/P
42agbafv8FNPHSYywQngE6HZGArcrM/z+w51hR4dkhTmbyFLpYlhVf+JFAzzehgI
qTtT9QCiALlD4bIItSg0Kktbca3wOa/hgXbdds+IFWhmRvXsxZfNuZ8G3Ie3D66L
V6FnBC1i2MEMetLXuKzPxCWOhLfg37Xp/CeBlcJ9J4TR+RMVqIQjC3AQuN9x1+gJ
oSgXjWpFEkmlxztdSGJkOx0/F+5rj6IeEaHSmgrUWpqYCJ7cEHAHF5tPB1wUqJCX
c1X8EiuSbnm706JI4+9mmL79+cp4hwNamHebgGgQLubC82ZVJNEJq7CM7xF5vbAm
9dzoqXHmiH+zPRd50rq4WJhQSLXUZ0KUAhHfLL+wQbT9hEeW43OC0F6wQ3xV/PkX
lJ7648OKnerPP0gPnA+XV3uzbu0LDVsuETL8npKnI3WFgplijcAB4u6WLvOHA4Pd
C7Pe4Ez9ad0bJW//VVhN3fFWtyHg0B4uF17YCnr4QeuicLprpeIFCZwecOgAjuia
4xnmMXGtLVv8tFbxSTVtC0PL/UDF3jiLr7qEIvl1stp1mK/89eSy1f59tbJqjFg+
4hwuSCZM8uxfUkjwaO9mVkd+CGB+D1ia8g9boExUtQe/7zeXTIEQOzNWQf5TfHsX
Hr0FB4Rno9Lr/JRcv8VK+8T5Ajy2McvGJH7w+IScX8TfeXtwJwdQOzSOp2DI0xE3
mw5gXRxxc3gUFHk6AwhkUkrxbttHmiHIf8/vm7Yo0q29Bpi/qP7TvLsnyvM4FwTN
k4ylutocOPjgueRqkdzb7Ttbk4/kyBuwqmz4ZTKS1/uOhMV8byBvFSpicMXCK44+
Tp4fBjJjER5EXTahy5MAJNhCw9t8H4DwbvF13cpf+T2v6z5zjv3sqCiBUJnt+78o
2G+q/w+SBp41ftNAmmLkAQAnuCi3qfTqaEOiAeLqXbKN/6ZVb2BNGyzAKGYS2JAk
Hcn/To70IBzYuklCHgj5/glUDs3l7+8AcQyax64VE/mX0zbnYR9mVPF7NpPLBCpo
yl+miY68FA28+ezR0jgwCASE8zA5+fR9CajDGD8bLwWG2FyXSkLJSazzIu9Uq8mk
XUEq2obfAG7MXlqCWrGiB3s9ODTw9d28V3jAa7G9WgJJyZfyMvRZRxjHa6XYQPYC
mT/UQkjzRN/3riJYNmhMBNpUqyhTp08LqzbuZ4HDHyriooKbfwVZShR9X5Du2TAT
dugP9Ylsn72yA4wb9Cwr2xxZUNalj36WTAHXtlgXSjR37OVA6oWNTe8p+P2IJz17
41eF/aNWbnp43PzfZz5ERohtEnUEemxM3gQFmU7pdVSqrTCbyzwWzOOKGg7HRE4e
q1hPf4d3g443n11Pk+4LyK8oOIYBLm8uEc5kLF8+b584gz3zz+3An1sV6dWCPZhw
4zIqSSsRNwPwwQeJPl1sTYiAkz9TgDTMMrEEAIICI6QmdV0A9RXrbqifJl4P+pZt
OYAAp/je+U6SM/n7X1FxapnJiCYaa6+6rRicLTE8gAVyYhJA0xhjSEKWLsuh/ko5
KLiC5STA633O9V5g4PLj4CyXbSLOfKz+K9JftZbc44asatCKzxZjx/FWS0q9RhVm
dgj4hmJPdApA82v2xeJYM1EsVM24NGDn1PHkYv/DUz+1JBhN3nfHkyIbAwUH3pqE
hVPsaGuzISnWS6NPTJOtmoytxUIlqFYeiZ+BFk6uFds2IxLWvZ8o8RXoaV6Cdx9N
Cbla6RXHYGz9kxTiCHQlgIXE7RQ/LhyKoJCLsjQEXYgt858Qptvmzvo5uBhh2SNE
Asg6jm1sToXbtq3Nlegk1Qwyn1EkjSL8oyu60xssgdQY5rU3GoCY6y3qvKCFCdcq
KLQcE3U2KLUOsu6F+stZor8GyHiVGCswbIaFR61byjikjExov6Ai9ayzYo25zzkD
VaKTuiDDYRlMrDUjtwkmCLkWBxIwBmMfj0S9yORLPHFkBLWUeSUljLVuMT2cwX+f
8LCwUEnL1XWVLI/4nAvyu7xtmk+Mcc7Wy3LMTnC7Fj1luYt/UwJtM+Y/HMwfHstU
WWK9No2aksQoqO6QdLxmaKDhQpNI+4MEUaKrYYo+41E56oTLYZgikK6ruKbM+lAy
fuwRAUcdMy3p/T986vmNYbMYCFVs56bBf35rfdykFHj1izLrKGyjtKNLiQJTOkJC
GfEfOHa+G4DmPrQlBPDOmowBHvBwzTDpWZc7M88rWbopctnhjfkG8eJ2cEeN7wGn
h/ZLSQboob+zczocvR4BzQf06KdlLRmS/xd8rYvdd0yhbO5uiZ9C25Hvd6Fh/mea
910kbDu4rzSESkel4dIWQz2DeZeiRCAAKczujkZh7S2xZCwXubHvpWDAcrkH0sdl
A9FP2o1CLcdyva/KOoXXER7pLyt+JuZLDM2kQOgBvNnzq07j+p9tkDZwUMRWa/xw
lSOVop6ikjMj4pxefGJsqxzdvRlLbp5NQAuZIR0iqBk5AcCa8s7j+0xT9nwtD8TT
Ezx+MtIMW4ESaCTcI/0lZX64ItZKi6D7B/MdAwX3gjUOkuGgoG2HyHDk/eKsjIMc
yt3Wol4xKZrhNc8Ig84gy/UxMZEGwruzO3GzcGCMUcKHi6uzhPUDrPHnqZDQDArU
G1Bf9ZVAU0xiFEdSVaSrQm3FeOJuTx7Hdn2+3ttmuYDKXhcILvigJGaygCYYyCZG
6M8afqHftiFhqJ8YBdKrvH3JRVYrC1ZT3Iu20TYl3aOVzECk2JDktv1MhDS//cMe
rWPaVCSdgxuGS+SVYwNCAMBgqNMXfFD7KusqkJkEYwBBW451qzpp4BA98dpkaq30
U7eXhYfM3XEIm98OghTA3gQRHPBK0ncS+x72qsy//cWa3BqfO5fXvQd2WU39ySIR
3J78hBtFAeEYNGtSWgBTabNRscy973Je4BsSNsFlogsd24H8D9rXiaQkH/RAbdYY
sjH7CeoUb1Ikl/iFhs1sDXmEqyEzJRsUWjXr3H019hHgchY5hdYUAAuioale9ePf
JX5KDaUYkCvds7l5dcFZY3ApjJp4RFfHa8pChlAtLmSXdIU4Ls4ZWQTu3coS9pE6
vdViunpF9gEpQEL5Iacwv5+YAqbKxUxiqmd/IyZAjhj4B73C+QvvDG0AChJBqsD1
lSBAbL/YteTJCCVilSVLcGQDm2NeoqJYysEeAY9/dZCQzrqVAtQHTAl5BgF3z2Ck
UQWRThmN4oLayfBrTkvXZI9WdZLN6d1HOFiodiEG+1qjYugy7TdbFqzol9vcy1UO
kRrGSKCLYkoF90xZblaoCc0+75sFABWkfjBqT4C3uYGxQXLnu3F7JhVkE/3UU1MP
qcrfTep06dSQ/xf5sntceu8DvBcbssZPIp7fMBlsPAVc3Z/Vs61h656eMC0X8UtF
kRdJ6TeSHOAR0LOU452zF00w84RWZBQBNLDMEQ1G2xC5mAYCYOHctRE9nIqX7ZMu
7fEJUvk4msz8EH9uQzxOx3F4QcT7nYYJR8WvalsQTCdALtUlN/9tCvPHEe/wpTSO
Dy02QnKKH4/Eb53O2w9DR78xI6xHx5Axr/SMCOXFuGGfEz7ncGQOYtI5FDfJNFpy
eZ81wfrANGSaAZ4Wurvh7WPKDob+fYIN3wF69PvvSBocGPuxRcA05Ksd+r/FXJFb
4TXtkCQiJK+XjFUtkhnhyLSvYS/2qNO1YovAK0K15N4WUNCGcZDN17y7rFlrw2fU
jZt+QbM+cmxB7LA3T3BJfMPB/IHxizTzlyWNcApj5aWCHRcH/d6MGphbyEfzEySD
AEIPkYiOJJwVt43r+m9wonX5vVGMZnOb0oDHrfw8hW+vTGXS9bW9lnjEDiPjl/0R
ZWlriXcYSscTI1sBP1DsB/oiruiLADO3d3WIwaScWX1mJYiknmypgCQYRpLJgs+a
KpqMGShQ98EnztLwDCsowADwBzkZsw3bMDPvc+hfm1pn75rjhF2LD+fx3t+Izn+B
pJ92ZUdIdyK6rJUJOOrAKz1c41La6PSHwbSfRKIfV1FUTNoVgVHXQjLKj4se+OlB
rbWV4DhfYw3Hn7RjSnLJkOypiKvPHaBGqQu3I7G8jVEozqbksV6JhId8am7T50sw
tc6bz36Ts4gNTz7eSKBKF2j7OjKj23eZVCGodiH48nkGZmLjqx1q7MgZk0JiJeMj
xMTvHFJrJrpWFj584rMian6oW/f+B6wmt3vy2dj/ZjUhYKCbKC4ymNyFSIdPKZH8
Kqh3rrV+kycjp5BkV3aXOmiYUtxtjdKookLAdMPAqhliMScUVrVSbwQU3htJI9Zj
Ga8qEobJX2k+aly95jCiiFyGfOWK128pHuaI6VOC3Ej3GtpxYKB8FtATozX2DZQr
R6diKI9s+AE3CGf/RyR08evzZoUXH1J2XGnkEjUQ+6W3zusa1nIiLuMrgTpTlbu4
Sdm5i+isinffHP7DP9WTLp/CGSRA+3adBWXhPbw8SXgS5WovgaBpyIRvioa9CGWc
faDq+DL/az13MOixKPxYZBLDX95FWFiQY0So99/cDhhmlZoEHUmMZmPPawQpVvDJ
kqlVi8gdL6gHPL3aSSKukl8gROLW3/1XVqPmQl45PWFOxXQfRe2V1Bbt8r5O9FXO
Wdu9ZUgSgBUbeFVhLPyKQ0hAgg+pjTlD8T1XLH6Ch5UttrBhVRCfXqvADBA99EIq
ExNLiVZ/tcJcvOJLCUhFoJSNNSfKAlSRIAX0jbX6qjXyllj9QtTRbqiBeiTv2jtm
FbuDYUZsYZjhm9jeFFQrzaDVGZZNMzRRDToyK0VDYGFN+HcEDltApAWo1f5nWG+g
x1u74z5RHb6Fdskz3tREOwcFi8smxkBTT8QpFymMXhHLtGX1InSYm6E3ah9cZh9n
3qSO8u7N8AV34vZ4qvg4JG0W67kCVzVxX+bqGSAElI4R/dO9+I/1Ol4pfjhUd5+o
GVHIgIoq53x9MYhOHfbZlf4BCPoCT6SIXLa02u+1IMiYJRosM55h1Dcb5IeZdyov
MduhfPh/0J8bPdQaVc+DkUi7dK7nSHH1FjlUa+vehNEscYAk6hFDeG4HeDhxYcjY
HTAZ2o1CFKOtGT/Wx0PB7axiVDEEwz7v/O0UqajAuqTQ8FBZGXGGpLHT85nednqV
tTEXI2jdppta4Uu3Z8G6fjvmwkdJe2BxVavtTuplPQH02RaAw9jiwHbmlTnTNLxi
3H2NCKDISkh9XnOmK7+ubd3lqmuA+5iA0hck70xkobcxF8m5ZtEWQ5a091tCKVNP
NT+KNnOEZUCaHmZeJIeHsNpDbEDyLuwRUj04+LBAZusERhL4qD4YObjMzRik/MZU
30zAuSFaPo+X9gkOL6xJ6PsMvFD68pfPKHteZWwwz2QGMaxy+fYZFLXnNDWMR+Vt
X8C1F4uqM05I1RGllJeadgoLAyhObfcT9SstURIBG80gMOFdJiAqvA+Rod0N1YDe
UlltQRb0/pl3oNu7HbCcUKC+DCD3WROtSS8IrW8c93gOK7L64r7Aa9b2wZwjqmF0
8oT3vfR2otbxW3724c/6D+1PBBCHS9O7c4LztN2e9v0J2OOUAD4nNa/cgguoO9dt
6wsXzuUEc7umQV7J15i5qDXwo1K2b0lpsPVSQ9M/FntIOO2pybdeb24XT0Jp9bjw
xGoIcCxSQVvLDgZldwaH6pDnf6+GaYzu6pfi62N1JH839ar76ZEacY02aIppcUOk
1Siu9OOBXMpk0j0NBT/68fYFCzEPI2dg7JzA+tFbeBG5JmSOXbsomtSfF4ksXNFH
CfFleX7lmijcn48Si1ljfKkP85qgBBzcWv91CcwY8ybjNrHOhstDVUqXYXLNGExj
HM5Pz04I0Q680W72DkarYgZzswkpbfG5A6r4M3EQCtarBGPV5XzLww6YUvE2ORp0
PYXFeboHEc48x3pucRbnZNj9XBNLeJbFqADUW5FcHGQ5EmNzChHDg30vnH4r84xQ
wKlQOBY/al5yOIf6Oa18OahoopsMNZHdqKHJi3PqlvYBkmTswdLs9fmf0IC1ftpa
uFZFZ+OiYDxZF3URKP/LEsJyiZl7Xyv0QlDYGrYoGvvY1wlm8MIpRxkRN7kWrNa5
5bfBTZyPg4AqAjy9uZvEI/e1X4PrfExdCSJjQP6YFcbj7hg5uU9qyMNbKMG/cyEq
edHu3LeDRRut0rSYxHdXC2yzfmu9DUckCfsUTs+91+Jaet8DY7YxFDOaEfGS4IIC
1K/eQJKW1iNET+Mppzmn0b/UKwzT39SCYHha1APlb/0NfWj85y1r4K8aaiT/vLcW
+jFc3EWLMbDtuWOSdLZrDgLHa4F7qunBoqj/fLC3d8OnYsl+8X9U1GdfdfQ1dWIa
3HI/igA/bKhVdKWsCWdx3S2ZDAd7BiOF+/vDsKeyWsnEwfZXa17BUjeHIpnpc+uR
KyfGH04OpAs9oLQQGfFVtJTgMAL3NEI57iZ3IxS7Fqh78GgYJ5RC46KfjsxkJ1K6
mlOBvoIbreaZZ9FL3JtXWZtvxH4PRrcTmYqNQaw46ZL31b2n7amtCXoBVTby39Bu
WBdaSX0/TY/NTYwzpFquF1Y/h4chpBwb6/jLJp0rR0IWEDLf0aXTzxcPW3jIA6W3
3v/albxOo5RTks+ZHwqnV/dx2FCbYdA99n8UHhAB0qIA46Z7yBgiIO8omB3g/brK
RAanwn9nvVSKkGkmYRLPJ+LNJK52u2/Jlm2dX255jBQ8tvO8lDEDRrbLNJhHPm+A
RMHbgWSIqnylix/wvyfSOdA/8GU/yDNEjMdF+nQcz0yVMFtfhzLl4eFC34nlzQav
wsXVDVuDaovNJbgM2nmMaYejeqPI//XmLfMlX4+qE77UGQDnq7odF58ztiC+ENkx
EB+P6we6glokprLgejFYChiFwsAU4sye8oTFfTlPCsL4kNrZZHCFBl+Z6UVYjG6U
2RPvIRwU8FkQfTfWaI0OFDruWDFr6tKLgEJvwnX6Fvl8KuLCHcH3VQGCJMHDRToC
6luB4k+vefwizEsmeH1ruGyvvU9w4lzaERqpw9kyi4ok5Y7zg2f7QUsH3xXSGWXc
/+ith0PZ5zSzsOBO6aIOBxX+fUKaNaIyluVtSY34HPNY/WEvgrCT9Ve+nGiNmh5X
lpNVZl8YtN55p40Qtdu4wGaMEB303i5TPjY/BdCj5GWvk0p7WXUmqErzb61cwmSL
2z0kMyvd0Sv7BHuSvclRqqYFVFAw4KFrBUWxbxDczkRNUkt/utOFDxngO5kGcLlo
v+/GzOobR41Piq4Jrp9NKR6fxp8bBikxyrNu1R5CJqlfld9ush/vDsBFXhB3TYvD
I8Aw97Snz6ukZ8D4Lj3jFZ1yS6/LfPFf/lnVxYGXD2dpYdM0NAWR6MGuUcG2jWcj
cREWExqzSobanwiHYylxJOq5uaCDPGUULcoFnmSNHu6E+3RpiBuddliWoLPd0iFY
/Do2+8E5j5uNBzWMzeal/XOtILzc+aVLCeoHQ3IuOkKKgc8El/cJ1xXUZerZRELN
YsuGCGhTLjAHmTdL9VKaGim++NfnhSfXW/+gPdVRQmcligpgGpn3YxGZTSqHHcYm
Uq//4IimRKOYSPqitVcrXZ40TWhRpu45HwGImIdfb59+1U7gBayiMlepX/JBaiur
oZERyYBPRwX2hBXsbKAqumntTO9VaIrTTzgGIx1l6J4cjAR8dBhGNKHb3/BaTnTy
Yt5d5s3lmST3kJyE4QbIYgdD1i5CecwZvkZ6vdP+gM0r9eAKU9JvxQo3gz5ckNW7
AMNBjjviGPenwXO84lhUGOFfs+1E/cqKlXkhxxNRtuUAwnAE64Y90orDRa8VT8g9
0c/sSPeef2zLDzqyH3o8+Vg7nt80L0rpHN9d6QmS52LrZFZQLlbejUdUTR7turHS
HcsN5xNcfQIFXnsUNeLMrQp1M0t/DAcndWXR5UQE63mxCO3ef5eAdL7AW+KRRYFG
eFk3HBRjHKigKQVckZyZk6IeUhAyWB0+LcLTPY9lkY55oZiJ8K7JwTIKeWgBFKRS
Nz1Ce7SkUIhDzGcaw1HH0Cvg80bc6KFTqpp3JjH6bZNhQ++8hW6nkWrdN/S07yzi
6uMnpjNQWLVkDBeMdXZxkTLq+X6oC7z1SkdUyVjoA97fo79X/tpY2VZBtAgZKMkf
bTg75QzG7FNPDnyYcYxmL5ROVJbWVwzGWtDpniG0QCW6TKAauhho0Oa6CoLLs+Jr
YUhzDD5YkohjdTnJsjfJWSQcqarySKPCk8nUDfpBfPLtMSq+2xy2bupkhy38mwSs
uTJ0e1bD3xuwvmEdDfNIVNIrpYMV0cNNmW4y2SPW9Ju2Fhz9H5GWZ/BtIcB4bWOr
Avkkqgd1MbPnUQhS64fYSVEBAEtLxXSDUV5180odo390YhpZbAAl+9vDvEmo0eNW
014IAzNnik2fAuC+9vpaeeONlEzGFwoBwNvrGzKKvJlCyD6HR0wLE/iTr+vnsGZW
P9WYAucDpgNkG+ZTq8gv846nrmaG6B6DsKWJeKJlqs+p6WFkh9OswYP+nVH13eVM
o1uF0yx7ha9IV+svU6DENg99hoqTpXzjbmdUgcfGKYzyByKrEpk2/LyYmszgMpN0
Zm08OAWBzqiwYHb0CowP7sMaBS3ixJ6ROz1bzBWjgBPidZZKjPNkz9wK+ow3xv8H
TLTn3t97qFkEsFjuSQqACgVQbq5YBFSQRFd1pXg/KOtUZJr+BGb5tbxIq1P0V8WQ
6XXiEkFZCqDT3XC8mwpb8YD1/re2dHSwNvvP19RHV6ZrDwhnR2DkUNtLnuFcKFFk
qSrMlGorSzEzcseysx2nEuvLz81y/lnWjMyrz6PZ89yhzOL7KsiHSKhYzLDEFwJo
PHQkb6jLshqQoMgGvJnCumUYLybo5LbjD1n74H+DKthZK6ttJvnpaIxRLZbOFI4N
DLaoQEzfk/bsMssccXevu56KLT1qJdBe43AxqLPFMv/UJGGmf/htiPF52+C3zvxe
JR1MMzWXVUvyIbqGJMRgJjQo56N8o4Z0u9lblonqoa3oFn3t1JV+NIVgsBoSu0Lv
DqQ1Up3dQNxhs6AYV0PZlJCerJL3a2IB4bDywL6Zj+twDk93qPJomXZX1A5++76l
qiUd2GSnt9jOWwVoFHq/ZHbr8sTVEnTdoM0mT5Nu6k0K7Ie3fv5jj+ZdREp1lIcK
Hohs+Ughp3QwuaJyryef5NoYTQuDs56b2UDyXBh1zguRJ6Ut2UOMTzQCF3KzfUGT
suuHRF0MarkSAGXUoth2PbmSb/BNHPUEiXYSh5Wgg8DulU9liXH1YEv3StzpBBs/
H47i6A6f5go6dQERY9Je8YwVtTrBUlswJaPNMA5C2IpUQBvzOxiyFkj7bOxihMLq
KnCa0baRmkuojWIUfZHf3TLczOZVc8g+ZoKF7aJmUfTWZDzXT+Ey+S2Jj19xycyL
OBLHl6XwyWPUvJ3WeHtMwz/qOGtua9yNHnhEtwqJcW48dRkGMzxF/IC3O1IaYyVW
C2FtVA4cS+s8ozDZPiT/6s4+SSx6M1OKO3+KK1fso48olRING7adskjqSncWowQj
xlrzgqku+VTKsFU7rlex8XOHToXf8+kSM78Vq6szaad/tgSKPNiDARQFf84YCEEd
DYnuIYWbgJDyfKqiZ3KSs5k468yrU7toewfQOzN+/1DlkiFM1xB01Ij43jGmCBwl
kKlQ8bjAC59LIwJeY+Acl+VKiyjI00x3gGtBP1VZzLwq+jaz9zbQnta/ZNcQFdru
Ji7djiyDyq+iv/wtkyo/m3gJWGkI1gyEjLFxlPoBojwglOOsiwgz66hXJdfXb4ZT
YJ6OJmNyP/8HWd2qLt2BtNRbGvCKpzl4o+lWSJth8hIdQBBURL6wq/VaEVpTNTp8
VAbMutIrtGI4xMlm5mKn0cvQA4Ji8GoRkEmg+08HxZrlFu0J4RKzvkYlOMTaxU+Q
kGbHcq+h2l4x+NktclT5Mr9jt+BWtOoohP0kG4/4RHOC297rxFRb4y/Cf5M1BF8T
/QGm864Fe4uF2konL8wlM8iInHc1LFKp/UeWxOHTPibATLj7oErbnkDQ4Yeg1LXZ
CKRBhrv8F6IUnQBmJ5h2JKgm7zJ+jiCjHVKGarLS+55IIL9X4LCJ1zSFeIm6vcsn
PRVTq6mTsWXom+N3V/hKJniYoBSqxOZAkCxrKBONm1LhyUJe6MM8d7d4XOFbTK/g
8hikQkFWmOwhY+ofY6QKeuplp5Wkg44oVSbbULU105MNcfq0/RjpeDBu3uPJaLdA
Adg9jlheCbbJ3GRfM4iNo+E6j/BOBW77MDisPeIHVziscaPNuQVF45tD9fVzgct7
UBAhOsjFJrY2MjKFghppu9ubIEBLgQKl7H6cKydvO/ZO3uRuNz/UNQ26XiMoR4xU
f/FT3YfaZAV2sBgSW8a3+YjFcq3hhORpjq6oj8JrxVPciCvQdg9y4reB0n56kJV4
66Va6d7bdTTEHzRJ/vrv2Vn8pR6WXvvamcp+D6TIamgSvFLWskE0vmbJc++65FFF
/fv1Fz0ru9Ob7ZqqD1OunbKR90rwoD8vc7tlFATH88rdGqmrdrNj69LRUVQv3eqd
o3l3B1srcfFtoDRpwLQVlK/7rSMzT4+yOw85B96pM/WJHf/mQX4Qz016Fi2eqAAz
lr0NKrZB429mdJcsnPZkInsKBJO/YDuqVGf9z8nZ5PV4ny4og667UCxVowklhOIV
2L6OXuR6OsoVDQmsznha0Cea2DH5fxb/UNf3W60BngY4FufywAfMhnAnU0x6FjaN
LOq5yaE/yuK52HWx2ObAPT5UB6zvvO/GntF47f3H1WvEHHks07SFOHzIypQTiEa1
61TpEi2W+RjbyLW5FECdDBEYnG3dPVFRiuOG97NPZtubSiF2Te7xlfFdfklTS5aZ
f3Ueb796IOff46OUyc7e0xJg6Xii/ZB+vN/cfDiuqdifc8PzzP3bVo01taZ61Guc
Si5HLvInzptGtbyYFn8Kp6Xn5MthIwBze7xsuWJ0nyFbkI3XHrEycA9RJFbr7N+B
xrusuj5iAOEGkv4+2tfJeXh/mn5zBqhQZN4ahMjfAc0MmyOg22SitiP/NeQJQk8i
FyrA0VSI6zAzryazeVLR8RMUXG2CEJeqQhPt36SNIgi5XGsc/XGM8xSVdFHKUOYT
88+O20oAcmDklvJ1j0K+cKGqwIjxj9c3wVGnTeKgc6U83K3bhca46Or0yP/A60S4
b8KxX6oztKOe+E4Xo/N0JsIBKnK/HNWz5Tswsyquf4FV+2zRewGic6Gz0yAhQCWG
NLBaJPpALNGOQX5pN9QtcfxQR1bE7La7cDOEGQ7I/KoJkIcWdNesJ2Gf/z1A2rLS
k681RdQjZRnSQtUoE1Ieb6XdXXhtJuYQLYiuMI+L4r0dhp3Bcf5EW5R//bSo/gWt
BfOYnCAmSY4H+oC05w8xH2sfjhzLGpGntj7EAB1mOk5ij5a16ogzxN3p5TOZk8f1
ovDjkbeRVDrlF5C29HXK2mqx15iEWpFEG5mX+UVsoiWmC8ttNOkTP6+fUC8eQ0xG
Ga33fZX4LV2WX2GNMiv6SaHPZz0SHorm43IL+zpN98fCZrAaNBX5NjmcPJFLIzX+
qXE40UvOIZA1ZclmByiXB9TlJZh47vQw/CnlX5/0STRYkH/+M6XiVFYydTMWUqTa
J30VDMlBHWxizMNLC85avwmsl/js9LgzDzXJpKHGZXn/HC/7eYiXPu25tol61vFw
hQcBcoVmQMO+ZMysDLjQ08wsZvnb1COwCIV2mjvEK7EanIZqxg/sO6ZWGi1OnEuj
7DHpmtdA58dxaPcfYnH/V2dIJA4TbBczJLeajh5VzvwtvlkDAXvv7qDgpbgln/2p
6P3pS8+wnC3VX56v0E9r2CFh8RPSs9fBQPBRI05uUsyLeiDGEivttAqDyaEAWjN1
he6vGGBg25gpp+k/MxwnCBe/44CR7iWKW0olpYYuCw61yCVOpdBqfn8cNPkCOldd
K4IufBxgsOcKlnuxNqjJ1ssxROqpjQqhR2ovjhrQU03LHM8ienVSJEBNgXgXHeyv
oyxiVMa0yHaLX2BO7V8QOy83Bk7S8bUHq9vt9lGaRN9oaNIUDrJrSqgfZH9/EOQk
iXCAOeGejQU0bQun9kOvlkWEirgH5Vf1hh9hKeYF30SG6b87v0eshFVqTnzYtOXs
4viYmFy4+PG+2XenhCu7paIkjwVzxcuGpbYBve+KDz+oirxB7SSRljZMHZzEuHt3
bpLCPy2v7K19drqH+0BiMij7CynV1g/HcmPv29t9y+oTwzSZ+LwkqUPf+SFbKbhR
1mSjQaoOiKotnDNfCP5ilsB+7E6CDPA14bnMya34h9w3SaJW/ucfcfOtL1Hop8Ug
JBSQ7Wmp9wxDTu7JVBJ2kWmoEvQRLbtJ7QXtXFPSreanI4eKdM/30W/i5q8rduxM
O2UVcym23jnk1+7qvh8p+nLkw6mAfV/4BqO1xR9/wa3htFQuRehrgD/T2xgpNHVi
UfCxrtqcq7NcuTuePkR5W5jgIUjeH99KSWGN5IA9xVRLNW/J0kdMYcL+s8a99ZmD
JI/xPF84V3Hk1SSvrUomtTpADNen8qqh1ACrq9MJUpkAehbZOtKozNes27/kC5Wv
zXOvBRzx0Hwt+tQLp6OAfrTHw6amTb0bneIjiR7S81zgcDxJDNQiqdjCy5pJW4qu
nC9k141FDBsMb3ZnD1/LquywWQBVqCsucKgqhvPl8tgBEU8093+wePpqVPLtEwzL
R7cnalsM5d8turQEa3bwz+VRtZ9/QVDZs2YHARnhIGcMY1sPx3mxHhUhmOe9iejS
Iv3jl2oE9qQOiI+lC3JMJMKnniqqn7RPstTp9g1EwNRZhuqd1BmTbMN0Hxg3RZjW
SVTfPEmqcm6ZKoKBvGL+TDpU3UBRil7tk6orbSkQfm/H/wvp3ToRqO2ueInnQFkI
h7xc09Iucaaq6inloC/xC2CzJwFe59FqEK+k2qzOQ58JtERnp8El7fsq9GabxdIq
XURY8YV18HYtkQO9TR1ecSc3spqrAF332cvelSce6vjtWJybEihlq2vwKCmAeK61
UJERExE0DK8Kb0twfuzRaxoOFcu6HVhAIJDuMuscSEFgNsCcN7SY4w0Qtvp4Tln+
3z7nhwOvfA2PC8SH8V+aF5XDP+bGNTu2IjWUhGrs2C0iDnJTngdj5epciYdsGSgZ
/WWVXimf70CVrKv4JvmK5/q6jSYz1Z5D5qgoQDaSljtWB5EPANXQStzPYC09n/rZ
9yBwZeZW1Y2KJgEf5y9IehDndqrVU2w80G9cMOb0RTWqjjv0MbCBMxWvMIFPtqtQ
vDVzaneR/zUNMqJJp4p19iU8yzaOHm9+ox8bzVXviTn/vA4msb6Ac4BvgzdVkWQO
bVTrak7d6AMF8tZGxz7kQOhShOxLQVaFR4pobyV0jeTxzhvZAY4EPqgZaQAY/Yf9
NPEJhLY3ISmxaPvwaGiTVUajXnQjBaqKw0/1lviWx3pzVCAH0ep8OXWVuqnZKE2u
BBtjIGNoMeM2pnuTaqVBKxJANo1A1OudgFajM6yKbkuymuilESiNKqgRV+Ab6cm0
9sr3MQ+r4slnBkNHtMiRUvn7n4Uh0X1fR2B4I88MVZcHkv5xXNJaqFmlyijE6Kmg
uIZZPo18MZoc2UbCKJhrFBQX7/PbUSPOIZPSctAjNNUEX7dldO9EAYcKoUz7+6R3
P90ftKWpFs9dDuFwA1uaF/E8zaSfVq28SFAUdoWbYRYlkyxMQArSwk0JQCq0Rtdr
nw2dH09Y7Oi0fJIXtNihhOhJXcpW7ZIP4lMfcAJiqKuZA4wtNpYBJOBTCcwTY3gv
oZr4PwfSwlKuvdnds5cV2DemWlqsaZNIJNvJMJ2KfKJdnGddXux+cvwryxvh0iL6
YVe7Y28OmUQzRtgs9iQRbJxF3c/te+o6h5If0ImIr/Xio1MMr++7Ys2h1ceMLpsh
eS00ngE3ShYWU8XFExcDX/Nyj1licAVQLHQrVlEC6w0WSLfQEeE45RqlzzXLcnai
1XgMpIpzw+9f6IiTVTQ9BabxjHvTVVAWTnHut68nPkGrmNiktearLkmU8eG/8bOF
cvCxc3svOtpxoHKJx22dsN1hTok0W4pyvPYW/EvIfb8toEY1AMRBHTwziym01WKu
oOtwTpOmvNOCsO12e3etU2zBaC1UG7ZCJfNN6fbChNQ71/mCdiVqpTSpVuFNvMMV
DG9wUqpnirzh/xNbTOI4phYYekZkRrZQVTwsOTCK1zZfVSfGKsWUfHCsul+TXNg1
wpslk0RVOnm+l85MB0GXaufE9nZ1JAZUa/P6JJl97RthOV1P3LpmqkuX7Ph0qBa5
O7rx8mpsDr8hq04B0/KGBJANDD+rZMzx9rIojc28HQVmor0/KUPuNzZXgQIZsmQf
cWzFTwPVfNb4f6TlkrFPELG6QQOM5crj3KMzP56he6QMh3Q7fDIWJKD37tT0K8XU
8R4fidQMDV127mpIL68rjwcD29Ywe8+ykhssuKLh+AR5q7/IwCdzs9DeQRssEygv
dJ7X0I0Ptf0ZrZ+fWmOzb0gdDNLlhiVvMuntUWxT8tHPy9hJJ22BM0Y3s6gt+Vw0
hK+2dMKmMzBUQZ/QcYVCtrc9BsKFbD1rVzlG6dLKSIIa7iK2IuRbjMirUXMWNPKq
ui/a8xgF8mtJzMo8d6/Nra1PWdirp2z1p7RcN4or7FAzDOCzHA9GhThLi3XTOk6V
Laitp7xPXw3sI0ls7C+Vcp39wSZm/fnakRE9OWANNpmu1JpmqM/T/3ScLlL1docC
UaMkeDZtq2Vt27NtqciYPYBvGwBf6O4OdxlVGy7J8A+QO1C0VhH3JJJMQJXKjZbD
XrXRuIGdUMMDsso5nWL5FewoUlUJnwAOgUE9uTYLiG7YUqUZmhJcReYr3uP0r51u
M5L4Zp/o6NQqfUQ/W5rURkiYYneEBrIYILqRhVerjrPW/+//5rIAse0Uio/sSUXv
xZ0fNfP6Mh3fAsUwhaoHxXsmNp/YoptBBNTSXhTETjWhx0HqYF0oEBPToptqFosg
bA7t0Xg+rIyV3p3XfXefT3bLfBIkWnqUEtPQfKQvp/pex9HxiCNhc+VJVeR1grh3
RGBkYaFVK5XUHTGquJR9FGcwS+3c4a5mHkpzYy2dqGdYPEVZudu3zQs4GpmpZKi2
97Tn7X4DeOeVZdrHWfAFW+y3l1C7/fDO7N+tYSEUllLWPKbp5fYRQOvQuwmDLjnj
zphfaN5J4yO/Rswrn3emk5vkJcmima761cECsFZ4ywFA76LHvV1Foc+HajGMJZIE
snWthIAmMOCWR2/mf1+Gi1vawL0kIV3ONQm1Vg71H9+UyND4m0ivAVjOqkKelpiK
+Ce4JkasqJ+ajFBLQnOZVmzd5XbB91aL2HQ4i8c0q4jPr9O1Lr/IDBJO//4Pxutc
0+4+N4Pkgm7Qzd74bK2yiBdsR/sMP4nZSqmfCEW+xgZXvLgDlSA6CBwoo/NDgHDR
2iCAhJucQk0Uw10p1iTkO6vV9cOiwJ25CcKL8Vl/rqtMtD41jUilDRJO6Rm8nzfY
zgBNkhfVRTgGHQQSLiS4/i1MIxXB6MITkUPEbkjtpYNLLgQ0N/z1S9PiuC6ia5zM
TRBM2DwLlQ9L8ZweW0XCP3beT19BNnOt4Lvm1xy4G6OX55BDApdEVc6C6nxyQD3E
4qRRaaEYT7AcJlpb91NAR3Qb4SUXgtVILOUP+3i8vGTRWkZ4aUIjJPccfjyjP7D0
8lv9ItmKTA0EyV5BmU3a7lSoBxdXdYdoMc+/QuZXCAl2ckGTgfIS6iOcxAoKq4Ir
fVsO6Wfx2pmg6dz8KlvMYW+lA4gWxMDIWXWtmjJG+QEemZP6gw8Aa5JFBspwGDl7
5BEMn8PrWmbnsiuP/5blQluzbqmDYjncNqt0b8y0f9jk/02Zh12dYWgJWyPmpQUX
SiM9IoY1Rzl2xJRWsO89EaFH43LcI4zhKeDsBq8xSUxmNdke+aUC6t9oS+Cb9rLu
bYhF4gQgjX/DVkMxNwyYgEWJ3b4SF4tFLFzpvJ326icTUQe6UNNqqpu6imBEvGn9
MtXinp+aTflcOR0X+a8xjxLh7eGidyjVZ3f2hEQPxh3pI1TGcAHd0PhQdO77lZa3
LHO+R/g9qoMytOI262S4ib0CYlGuPALtNmk/Cj8LI2WvjSiDOUA5ykRxUnyhqqQs
1KD5LBGlR1hv2/hnG8wXvvc4ieiZyeYL1b3r47RdegwDyRD1RzMquXHXnal/MlHq
2/cqfVxVTQBNH3lhuPej8EIR1CCoxSWjmBVACCittkgXIIfrZSO5JKr5ZcjeRiIG
qSF3mpgv/N2/UZdyZIsee1lr0E7ypf+bmf7WxpqjIX6wKJ+h1CGl/ncMyslnpkbI
WULWuxmh5bONHGDNRFGFOQFpweS2BenOjDUSORDlDmy+udZxFkn0J1b7BefWS3hb
RDCDG9xPn6ofZY7wbys/Vra/OZIXgzsmjiVcqTqznR8Ey7wp8tD22W9ot6OFAj54
O/oIJeb9Nmrp62tA9Y5PXxOFhue2GCLdIZHIrauKqMu/R0Nhvbckk1RD+QmeemEv
+7zwcDGyr4XnHcdbJEj9j0ol2nMq0UkEf8SmhEGBLU8WfjGpPT8Cna2/m7lrDbNd
NC809uv2g8/FYrrg+MKAl6hwkukPxUq4T7LUihKgKUnkabJ4XoaZRRmUhwwy8D37
ihgRfw7QopWWcpRsI6FhKJDCDvfVeJIfcS/cHKQmDFr20IVIv8d2RZsvNj9G5IPy
g3EHiPxdvEUxNQtSLVsTReYpd7zsh4ydy7wfpQM8kOS7JeFqXHxMQEuy0NzqW3r5
a4+Jn/6+EOtFqOYsT6ZdloJa31MiYgkVk026a3iWOmd395Trqgys6kHs2DILeUd+
hVNVEi74mmbrizXFKuXM8A904N2hEFQ4cL58hEbsT9gMzZI5HzOj3PWzR8hDD6Aq
cg+BBHvIQvcPOPYItHEOIID6o978uSPy45YS7MfPpGW3yesYOUbiNKLq0bPdRbrN
S9L09FMLjsx5ofbongmCna70OKrDNiu0ieQJo5oiq/Zf1DxbqxAqlAwv0USj9p/N
3JlmvReSzggSzhmHPXgObtlEOUVifwOT4U0ggHPyfvzjaM+Gjby1m3/VLsbbEZYj
SoRHx4fZYpcEhCTwMxHeDam/wSSTNklz/ufcfqI5a5gMWZFhiWFkXjdjT8C1mXse
hVMcs1yLyVNOgCHeok6ojg==
`pragma protect end_protected

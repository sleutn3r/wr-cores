-- WRPC LM32 RAM initialization: --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.memory_loader_pkg.all;
use work.genram_pkg.all;

package wrc_bin_pkg is
  constant c_wrc_bin_init : t_ram_fast_load ( 0 to 32767 ) := (
        0 => x"98000000",     1 => x"d0000000",     2 => x"d0200000",
        3 => x"78010000",     4 => x"38210000",     5 => x"d0e10000",
        6 => x"f800003a",     7 => x"34000000",     8 => x"00000000",
        9 => x"00000000",    10 => x"00000000",    11 => x"00000000",
       12 => x"00000000",    13 => x"00000000",    14 => x"00000000",
       15 => x"00000000",    16 => x"00000000",    17 => x"00000000",
       18 => x"00000000",    19 => x"00000000",    20 => x"00000000",
       21 => x"00000000",    22 => x"00000000",    23 => x"00000000",
       24 => x"00000000",    25 => x"00000000",    26 => x"00000000",
       27 => x"00000000",    28 => x"00000000",    29 => x"00000000",
       30 => x"00000000",    31 => x"00000000",    32 => x"57525043",
       33 => x"2d2d2d2d",    34 => x"01234567",    35 => x"89abcdef",
       36 => x"00018f04",    37 => x"00000000",    38 => x"000160a8",
       39 => x"00000000",    40 => x"00000000",    41 => x"00000000",
       42 => x"00000000",    43 => x"00000000",    44 => x"00000000",
       45 => x"00000000",    46 => x"00000000",    47 => x"00000000",
       48 => x"5b9d0000",    49 => x"f800001e",    50 => x"34010002",
       51 => x"f8004619",    52 => x"e000002e",    53 => x"34000000",
       54 => x"34000000",    55 => x"34000000",    56 => x"00000000",
       57 => x"00000000",    58 => x"00000000",    59 => x"00000000",
       60 => x"00000000",    61 => x"00000000",    62 => x"00000000",
       63 => x"00000000",    64 => x"98000000",    65 => x"781c0001",
       66 => x"3b9cfffc",    67 => x"78010001",    68 => x"382174b0",
       69 => x"34020000",    70 => x"78030001",    71 => x"38639280",
       72 => x"c8611800",    73 => x"f8004be6",    74 => x"34010000",
       75 => x"34020000",    76 => x"34030000",    77 => x"f800010e",
       78 => x"e0000000",    79 => x"379cffc4",    80 => x"5b810004",
       81 => x"5b820008",    82 => x"5b83000c",    83 => x"5b840010",
       84 => x"5b850014",    85 => x"5b860018",    86 => x"5b87001c",
       87 => x"5b880020",    88 => x"5b890024",    89 => x"5b8a0028",
       90 => x"5b9e0034",    91 => x"5b9f0038",    92 => x"2b81003c",
       93 => x"5b810030",    94 => x"bb800800",    95 => x"3421003c",
       96 => x"5b81002c",    97 => x"c3a00000",    98 => x"2b810004",
       99 => x"2b820008",   100 => x"2b83000c",   101 => x"2b840010",
      102 => x"2b850014",   103 => x"2b860018",   104 => x"2b87001c",
      105 => x"2b880020",   106 => x"2b890024",   107 => x"2b8a0028",
      108 => x"2b9d0030",   109 => x"2b9e0034",   110 => x"2b9f0038",
      111 => x"2b9c002c",   112 => x"34000000",   113 => x"c3c00000",
      114 => x"90001000",   115 => x"3401fffe",   116 => x"a0410800",
      117 => x"d0010000",   118 => x"90201000",   119 => x"3401fffe",
      120 => x"a0410800",   121 => x"d0210000",   122 => x"c3a00000",
      123 => x"90001000",   124 => x"3401fffe",   125 => x"a0410800",
      126 => x"d0010000",   127 => x"90201000",   128 => x"38420001",
      129 => x"d0220000",   130 => x"38210001",   131 => x"d0010000",
      132 => x"c3a00000",   133 => x"379cfff0",   134 => x"5b8b0008",
      135 => x"5b9d0004",   136 => x"f80037b1",   137 => x"f8004171",
      138 => x"f8004167",   139 => x"78010001",   140 => x"3821368c",
      141 => x"f800312b",   142 => x"34010001",   143 => x"f80036d7",
      144 => x"f8003f18",   145 => x"78010001",   146 => x"38219188",
      147 => x"58200000",   148 => x"f8003e3e",   149 => x"f80038e6",
      150 => x"34010000",   151 => x"f80034b7",   152 => x"34010000",
      153 => x"34020050",   154 => x"f8003b5f",   155 => x"3782000c",
      156 => x"34010000",   157 => x"f8003dcf",   158 => x"3402ffff",
      159 => x"5c220010",   160 => x"78010001",   161 => x"382136a8",
      162 => x"f8003116",   163 => x"34010022",   164 => x"3381000c",
      165 => x"34010033",   166 => x"3381000d",   167 => x"34010044",
      168 => x"3381000e",   169 => x"34010055",   170 => x"3381000f",
      171 => x"34010066",   172 => x"33810010",   173 => x"34010077",
      174 => x"33810011",   175 => x"4384000e",   176 => x"4385000f",
      177 => x"43860010",   178 => x"43870011",   179 => x"4383000d",
      180 => x"4382000c",   181 => x"78010001",   182 => x"382136cc",
      183 => x"f8003101",   184 => x"378b000c",   185 => x"b9600800",
      186 => x"f80032cd",   187 => x"b9600800",   188 => x"f8003913",
      189 => x"34020001",   190 => x"34010001",   191 => x"f800321a",
      192 => x"f800352d",   193 => x"f8003a29",   194 => x"f80002ab",
      195 => x"78020001",   196 => x"384260a0",   197 => x"34010002",
      198 => x"f8003884",   199 => x"f8004643",   200 => x"f8002735",
      201 => x"f800204f",   202 => x"78030001",   203 => x"38635954",
      204 => x"78010001",   205 => x"28620000",   206 => x"382174b0",
      207 => x"58200000",   208 => x"78010001",   209 => x"3821f800",
      210 => x"58220000",   211 => x"34010003",   212 => x"f80002f7",
      213 => x"f80002aa",   214 => x"78020001",   215 => x"34010000",
      216 => x"384274b8",   217 => x"f8003a60",   218 => x"2b9d0004",
      219 => x"2b8b0008",   220 => x"379c0010",   221 => x"c3a00000",
      222 => x"379cfff8",   223 => x"5b8b0008",   224 => x"5b9d0004",
      225 => x"34010000",   226 => x"f8003229",   227 => x"b8205800",
      228 => x"78010001",   229 => x"382160a4",   230 => x"28240000",
      231 => x"7d620000",   232 => x"64830000",   233 => x"a0431800",
      234 => x"4460000d",   235 => x"78010001",   236 => x"38219260",
      237 => x"28210000",   238 => x"34020002",   239 => x"58220004",
      240 => x"f80036e3",   241 => x"f800028e",   242 => x"78010001",
      243 => x"38219258",   244 => x"34020001",   245 => x"58220000",
      246 => x"e0000014",   247 => x"65610000",   248 => x"7c840000",
      249 => x"a0240800",   250 => x"44230012",   251 => x"78010001",
      252 => x"38219260",   253 => x"28210000",   254 => x"34020002",
      255 => x"58220008",   256 => x"78010001",   257 => x"38219258",
      258 => x"58220000",   259 => x"f80002a2",   260 => x"34010002",
      261 => x"34020000",   262 => x"34030001",   263 => x"f800460e",
      264 => x"34010000",   265 => x"f8003a60",   266 => x"34010001",
      267 => x"e0000008",   268 => x"fc411000",   269 => x"78010001",
      270 => x"c8021000",   271 => x"38219258",   272 => x"20420003",
      273 => x"58220000",   274 => x"34010000",   275 => x"78020001",
      276 => x"384260a4",   277 => x"584b0000",   278 => x"2b9d0004",
      279 => x"2b8b0008",   280 => x"379c0008",   281 => x"c3a00000",
      282 => x"379cfffc",   283 => x"5b9d0004",   284 => x"f800365c",
      285 => x"78020001",   286 => x"78030001",   287 => x"386374bc",
      288 => x"384274c0",   289 => x"28640000",   290 => x"28450000",
      291 => x"58610000",   292 => x"340303e8",   293 => x"c8a42000",
      294 => x"b4812000",   295 => x"58440000",   296 => x"34010000",
      297 => x"50640009",   298 => x"78010000",   299 => x"382100a0",
      300 => x"3484fc18",   301 => x"58440000",   302 => x"28220000",
      303 => x"34420001",   304 => x"58220000",   305 => x"34010001",
      306 => x"2b9d0004",   307 => x"379c0004",   308 => x"c3a00000",
      309 => x"379cfffc",   310 => x"5b9d0004",   311 => x"f8003641",
      312 => x"78020001",   313 => x"384274bc",   314 => x"58410000",
      315 => x"2b9d0004",   316 => x"379c0004",   317 => x"c3a00000",
      318 => x"379cfff8",   319 => x"5b8b0008",   320 => x"5b9d0004",
      321 => x"78010001",   322 => x"382174b0",   323 => x"28220000",
      324 => x"34010001",   325 => x"5c41000f",   326 => x"f8001d6b",
      327 => x"b8205800",   328 => x"f80040d8",   329 => x"3402001b",
      330 => x"44220005",   331 => x"78020001",   332 => x"38426098",
      333 => x"28410000",   334 => x"5c200008",   335 => x"f8001fc9",
      336 => x"78020001",   337 => x"384274b0",   338 => x"58400000",
      339 => x"e0000003",   340 => x"f8001fce",   341 => x"b8205800",
      342 => x"b9600800",   343 => x"2b9d0004",   344 => x"2b8b0008",
      345 => x"379c0008",   346 => x"c3a00000",   347 => x"379cffe0",
      348 => x"5b8b001c",   349 => x"5b8c0018",   350 => x"5b8d0014",
      351 => x"5b8e0010",   352 => x"5b8f000c",   353 => x"5b900008",
      354 => x"5b9d0004",   355 => x"780b0001",   356 => x"780c0001",
      357 => x"f800486b",   358 => x"396b735c",   359 => x"398c74ac",
      360 => x"e0000005",   361 => x"29610008",   362 => x"44200002",
      363 => x"d8200000",   364 => x"356b001c",   365 => x"558bfffc",
      366 => x"780b0001",   367 => x"78010001",   368 => x"396b735c",
      369 => x"780f0001",   370 => x"780d0001",   371 => x"38215958",
      372 => x"39ef74ac",   373 => x"39ad74b8",   374 => x"282e0000",
      375 => x"b9608000",   376 => x"e0000025",   377 => x"2961000c",
      378 => x"5c200005",   379 => x"29610010",   380 => x"34210001",
      381 => x"59610010",   382 => x"e000000b",   383 => x"29620004",
      384 => x"44400003",   385 => x"28420000",   386 => x"44400007",
      387 => x"d8200000",   388 => x"29620010",   389 => x"b9606000",
      390 => x"b4411000",   391 => x"59620010",   392 => x"5c200002",
      393 => x"ba006000",   394 => x"34010000",   395 => x"37820020",
      396 => x"f80039ad",   397 => x"2b820020",   398 => x"29a10000",
      399 => x"c8410800",   400 => x"4c200002",   401 => x"b42e0800",
      402 => x"29830018",   403 => x"b4230800",   404 => x"59810018",
      405 => x"51c10006",   406 => x"c82e0800",   407 => x"59810018",
      408 => x"29810014",   409 => x"34210001",   410 => x"59810014",
      411 => x"59a20000",   412 => x"356b001c",   413 => x"55ebffdc",
      414 => x"f8004819",   415 => x"ba005800",   416 => x"e3fffffd",
      417 => x"379cffbc",   418 => x"5b8b0014",   419 => x"5b8c0010",
      420 => x"5b8d000c",   421 => x"5b8e0008",   422 => x"5b9d0004",
      423 => x"5b830030",   424 => x"78030001",   425 => x"386374c4",
      426 => x"5b82002c",   427 => x"5b840034",   428 => x"5b850038",
      429 => x"5b86003c",   430 => x"5b870040",   431 => x"5b880044",
      432 => x"286d0000",   433 => x"b8205800",   434 => x"b8407000",
      435 => x"34030000",   436 => x"44200002",   437 => x"28230018",
      438 => x"b86d1800",   439 => x"0063001c",   440 => x"4460001b",
      441 => x"780c0001",   442 => x"398c74c4",   443 => x"39a10001",
      444 => x"59810000",   445 => x"29610028",   446 => x"37820018",
      447 => x"28230000",   448 => x"b9600800",   449 => x"d8600000",
      450 => x"78030001",   451 => x"3863595c",   452 => x"28620000",
      453 => x"2b81001c",   454 => x"598d0000",   455 => x"296b0334",
      456 => x"f800493b",   457 => x"780c0001",   458 => x"2b830018",
      459 => x"398c3734",   460 => x"b8202000",   461 => x"b9601000",
      462 => x"b9800800",   463 => x"f8002fe9",   464 => x"b9c00800",
      465 => x"37820030",   466 => x"f8002fc4",   467 => x"2b9d0004",
      468 => x"2b8b0014",   469 => x"2b8c0010",   470 => x"2b8d000c",
      471 => x"2b8e0008",   472 => x"379c0044",   473 => x"c3a00000",
      474 => x"379cfffc",   475 => x"5b9d0004",   476 => x"b8402800",
      477 => x"5c600005",   478 => x"78020001",   479 => x"38423750",
      480 => x"b8a01800",   481 => x"e000000c",   482 => x"34020001",
      483 => x"5c620006",   484 => x"78020001",   485 => x"3842376c",
      486 => x"b8a01800",   487 => x"28240008",   488 => x"e0000005",
      489 => x"28240004",   490 => x"78020001",   491 => x"38423784",
      492 => x"b8a01800",   493 => x"fbffffb4",   494 => x"2b9d0004",
      495 => x"379c0004",   496 => x"c3a00000",   497 => x"379cffe8",
      498 => x"5b8b0018",   499 => x"5b8c0014",   500 => x"5b8d0010",
      501 => x"5b8e000c",   502 => x"5b9d0008",   503 => x"b8205800",
      504 => x"b8407000",   505 => x"b8606800",   506 => x"4460001a",
      507 => x"40480000",   508 => x"78020001",   509 => x"384266f4",
      510 => x"2108000f",   511 => x"3d030002",   512 => x"282600e4",
      513 => x"b4431000",   514 => x"28420000",   515 => x"282700e8",
      516 => x"78040001",   517 => x"5b820004",   518 => x"34030001",
      519 => x"34020005",   520 => x"3884379c",   521 => x"b9a02800",
      522 => x"f8000048",   523 => x"34010021",   524 => x"4c2d0006",
      525 => x"b9600800",   526 => x"b9c01000",   527 => x"b9a01800",
      528 => x"f8001613",   529 => x"44200003",   530 => x"340d0000",
      531 => x"340e0000",   532 => x"780c0001",   533 => x"29610000",
      534 => x"398c6584",   535 => x"e000002d",   536 => x"44410003",
      537 => x"358c000c",   538 => x"e000002a",   539 => x"59610004",
      540 => x"2961000c",   541 => x"59600008",   542 => x"44200006",
      543 => x"29820004",   544 => x"b9600800",   545 => x"34030000",
      546 => x"b9a02000",   547 => x"fbffffb7",   548 => x"29840008",
      549 => x"b9a01800",   550 => x"b9600800",   551 => x"b9c01000",
      552 => x"d8800000",   553 => x"b8201800",   554 => x"44200006",
      555 => x"29620334",   556 => x"29840004",   557 => x"78010001",
      558 => x"382137c8",   559 => x"f8002f89",   560 => x"29610004",
      561 => x"29630000",   562 => x"29820004",   563 => x"4461000a",
      564 => x"59610000",   565 => x"34010001",   566 => x"5961000c",
      567 => x"34030002",   568 => x"b9600800",   569 => x"34040000",
      570 => x"fbffffa0",   571 => x"34010000",   572 => x"e000000f",
      573 => x"b9600800",   574 => x"5960000c",   575 => x"34030001",
      576 => x"34040000",   577 => x"fbffff99",   578 => x"29610008",
      579 => x"e0000008",   580 => x"29820000",   581 => x"5c40ffd3",
      582 => x"29620334",   583 => x"78010001",   584 => x"382137e4",
      585 => x"f8002f6f",   586 => x"34012710",   587 => x"2b9d0008",
      588 => x"2b8b0018",   589 => x"2b8c0014",   590 => x"2b8d0010",
      591 => x"2b8e000c",   592 => x"379c0018",   593 => x"c3a00000",
      594 => x"379cffe0",   595 => x"5b8b000c",   596 => x"5b8c0008",
      597 => x"5b9d0004",   598 => x"5b850014",   599 => x"5b840010",
      600 => x"78050001",   601 => x"5b860018",   602 => x"5b87001c",
      603 => x"5b880020",   604 => x"b8604800",   605 => x"b8806000",
      606 => x"38a53804",   607 => x"34030000",   608 => x"44200003",
      609 => x"28250334",   610 => x"28230018",   611 => x"78060001",
      612 => x"38c674c4",   613 => x"28c10000",   614 => x"b8610800",
      615 => x"3c430002",   616 => x"80230800",   617 => x"2021000f",
      618 => x"55210015",   619 => x"78010001",   620 => x"38215a20",
      621 => x"b4231800",   622 => x"78060001",   623 => x"28630000",
      624 => x"780b0001",   625 => x"396b74c8",   626 => x"b8c01000",
      627 => x"3842380c",   628 => x"b9202000",   629 => x"b9600800",
      630 => x"f8002f34",   631 => x"b9600800",   632 => x"f8003f96",
      633 => x"b9600800",   634 => x"b9801000",   635 => x"37830014",
      636 => x"f8002f4b",   637 => x"b9600800",   638 => x"f8003f90",
      639 => x"2b9d0004",   640 => x"2b8b000c",   641 => x"2b8c0008",
      642 => x"379c0020",   643 => x"c3a00000",   644 => x"379cfff8",
      645 => x"5b8b0008",   646 => x"5b9d0004",   647 => x"3402001c",
      648 => x"b8201800",   649 => x"340b0000",   650 => x"3405fffc",
      651 => x"34040003",   652 => x"e0000009",   653 => x"3421ffd0",
      654 => x"202600ff",   655 => x"50860002",   656 => x"e0000008",
      657 => x"bc220800",   658 => x"34630001",   659 => x"b9615800",
      660 => x"3442fffc",   661 => x"40610000",   662 => x"44200007",
      663 => x"5c45fff6",   664 => x"78010001",   665 => x"78020001",
      666 => x"38213818",   667 => x"38425a10",   668 => x"f8002f1c",
      669 => x"b9600800",   670 => x"2b9d0004",   671 => x"2b8b0008",
      672 => x"379c0008",   673 => x"c3a00000",   674 => x"379cfffc",
      675 => x"5b9d0004",   676 => x"34030001",   677 => x"34010003",
      678 => x"34020000",   679 => x"f800446e",   680 => x"34010000",
      681 => x"34020001",   682 => x"f80045ff",   683 => x"34010000",
      684 => x"2b9d0004",   685 => x"379c0004",   686 => x"c3a00000",
      687 => x"379cfff4",   688 => x"5b8b000c",   689 => x"5b8c0008",
      690 => x"5b9d0004",   691 => x"34010000",   692 => x"b8406000",
      693 => x"f800452a",   694 => x"45800005",   695 => x"642c0000",
      696 => x"c80c6000",   697 => x"398c0001",   698 => x"e000000f",
      699 => x"780b0001",   700 => x"396b7548",   701 => x"5c2c0004",
      702 => x"59600000",   703 => x"340cffff",   704 => x"e0000009",
      705 => x"29610000",   706 => x"340c0001",   707 => x"5c200006",
      708 => x"78020001",   709 => x"34010003",   710 => x"384260a0",
      711 => x"f8003683",   712 => x"596c0000",   713 => x"b9800800",
      714 => x"2b9d0004",   715 => x"2b8b000c",   716 => x"2b8c0008",
      717 => x"379c000c",   718 => x"c3a00000",   719 => x"34010000",
      720 => x"c3a00000",   721 => x"379cfffc",   722 => x"5b9d0004",
      723 => x"34010000",   724 => x"34020001",   725 => x"f80045d4",
      726 => x"34010000",   727 => x"2b9d0004",   728 => x"379c0004",
      729 => x"c3a00000",   730 => x"379cfffc",   731 => x"5b9d0004",
      732 => x"282102c8",   733 => x"28210010",   734 => x"2823000c",
      735 => x"44430004",   736 => x"5822000c",   737 => x"b8400800",
      738 => x"f8003887",   739 => x"34010000",   740 => x"2b9d0004",
      741 => x"379c0004",   742 => x"c3a00000",   743 => x"379cfffc",
      744 => x"5b9d0004",   745 => x"f8003879",   746 => x"34020001",
      747 => x"5c200003",   748 => x"f80045ad",   749 => x"7c220000",
      750 => x"b8400800",   751 => x"2b9d0004",   752 => x"379c0004",
      753 => x"c3a00000",   754 => x"379cfff8",   755 => x"5b8b0008",
      756 => x"5b9d0004",   757 => x"b8202800",   758 => x"b8220800",
      759 => x"b8402000",   760 => x"b8605800",   761 => x"44200005",
      762 => x"34010001",   763 => x"b8a01000",   764 => x"b8801800",
      765 => x"f80037fe",   766 => x"45600005",   767 => x"1562001f",
      768 => x"34010002",   769 => x"b9601800",   770 => x"f80037f9",
      771 => x"34010000",   772 => x"2b9d0004",   773 => x"2b8b0008",
      774 => x"379c0008",   775 => x"c3a00000",   776 => x"379cfffc",
      777 => x"5b9d0004",   778 => x"b8201000",   779 => x"3401ffff",
      780 => x"f80044e4",   781 => x"34010000",   782 => x"2b9d0004",
      783 => x"379c0004",   784 => x"c3a00000",   785 => x"379cff24",
      786 => x"5b8b0014",   787 => x"5b8c0010",   788 => x"5b8d000c",
      789 => x"5b8e0008",   790 => x"5b9d0004",   791 => x"b8406000",
      792 => x"28220330",   793 => x"b8807000",   794 => x"37810018",
      795 => x"b8605800",   796 => x"b8a06800",   797 => x"f8001d54",
      798 => x"45c00005",   799 => x"78010001",   800 => x"38216f2c",
      801 => x"28210000",   802 => x"59c10000",   803 => x"45a00003",
      804 => x"2b8100cc",   805 => x"59a10000",   806 => x"2b82006c",
      807 => x"3401fffd",   808 => x"44400013",   809 => x"45800007",
      810 => x"2b820060",   811 => x"2b810058",   812 => x"b4410800",
      813 => x"2b8200a0",   814 => x"b4220800",   815 => x"59810000",
      816 => x"2b820068",   817 => x"3401fffd",   818 => x"44400009",
      819 => x"34010000",   820 => x"45600007",   821 => x"2b830064",
      822 => x"2b82005c",   823 => x"b4621000",   824 => x"2b8300a4",
      825 => x"b4431000",   826 => x"59620000",   827 => x"2b9d0004",
      828 => x"2b8b0014",   829 => x"2b8c0010",   830 => x"2b8d000c",
      831 => x"2b8e0008",   832 => x"379c00dc",   833 => x"c3a00000",
      834 => x"34010000",   835 => x"c3a00000",   836 => x"34010000",
      837 => x"c3a00000",   838 => x"379cffec",   839 => x"5b8b000c",
      840 => x"5b8c0008",   841 => x"5b9d0004",   842 => x"34040000",
      843 => x"b8406000",   844 => x"b8605800",   845 => x"37820010",
      846 => x"37830014",   847 => x"34050000",   848 => x"5b800014",
      849 => x"5b800010",   850 => x"fbffffbf",   851 => x"34010001",
      852 => x"5d810003",   853 => x"2b810010",   854 => x"e0000002",
      855 => x"2b810014",   856 => x"59610000",   857 => x"34010001",
      858 => x"2b9d0004",   859 => x"2b8b000c",   860 => x"2b8c0008",
      861 => x"379c0014",   862 => x"c3a00000",   863 => x"379cfffc",
      864 => x"5b9d0004",   865 => x"f8002feb",   866 => x"34010000",
      867 => x"2b9d0004",   868 => x"379c0004",   869 => x"c3a00000",
      870 => x"379cfffc",   871 => x"5b9d0004",   872 => x"f8002fef",
      873 => x"34010000",   874 => x"2b9d0004",   875 => x"379c0004",
      876 => x"c3a00000",   877 => x"379cfffc",   878 => x"5b9d0004",
      879 => x"f80034ca",   880 => x"f8003e81",   881 => x"f8003e89",
      882 => x"78010001",   883 => x"78020001",   884 => x"384238b8",
      885 => x"38213888",   886 => x"f8002e42",   887 => x"34010000",
      888 => x"2b9d0004",   889 => x"379c0004",   890 => x"c3a00000",
      891 => x"78010001",   892 => x"3821754c",   893 => x"28210000",
      894 => x"c3a00000",   895 => x"379cfff8",   896 => x"5b8b0008",
      897 => x"5b9d0004",   898 => x"78010001",   899 => x"382138d4",
      900 => x"f8002e34",   901 => x"78010001",   902 => x"78020001",
      903 => x"38426754",   904 => x"3821641c",   905 => x"780b0001",
      906 => x"f800199c",   907 => x"396b60a8",   908 => x"34030000",
      909 => x"b9600800",   910 => x"34020000",   911 => x"fbfffe62",
      912 => x"78020001",   913 => x"38426460",   914 => x"58410000",
      915 => x"f80033e5",   916 => x"78020001",   917 => x"38427554",
      918 => x"58410000",   919 => x"296102c8",   920 => x"28210010",
      921 => x"58200068",   922 => x"b9600800",   923 => x"f8000ad5",
      924 => x"78010001",   925 => x"38217550",   926 => x"34020001",
      927 => x"58220000",   928 => x"34010000",   929 => x"2b9d0004",
      930 => x"2b8b0008",   931 => x"379c0008",   932 => x"c3a00000",
      933 => x"379cfff4",   934 => x"5b8b000c",   935 => x"5b8c0008",
      936 => x"5b9d0004",   937 => x"780b0001",   938 => x"396b60a8",
      939 => x"296102c8",   940 => x"282c0010",   941 => x"78010001",
      942 => x"382138e0",   943 => x"f8002e09",   944 => x"29810000",
      945 => x"34020000",   946 => x"28230034",   947 => x"b9600800",
      948 => x"d8600000",   949 => x"78010001",   950 => x"34020000",
      951 => x"340301b8",   952 => x"59800040",   953 => x"31800035",
      954 => x"382161b8",   955 => x"f8004874",   956 => x"78010001",
      957 => x"38217550",   958 => x"58200000",   959 => x"b9600800",
      960 => x"0d60010c",   961 => x"f8000aaf",   962 => x"78010001",
      963 => x"3821641c",   964 => x"f80019ab",   965 => x"34010000",
      966 => x"2b9d0004",   967 => x"2b8b000c",   968 => x"2b8c0008",
      969 => x"379c000c",   970 => x"c3a00000",   971 => x"379cffec",
      972 => x"5b8b0014",   973 => x"5b8c0010",   974 => x"5b8d000c",
      975 => x"5b8e0008",   976 => x"5b9d0004",   977 => x"780b0001",
      978 => x"396b60a8",   979 => x"b8206000",   980 => x"296102c8",
      981 => x"282d0010",   982 => x"78010001",   983 => x"3821754c",
      984 => x"58200000",   985 => x"fbffffcc",   986 => x"34010002",
      987 => x"45810016",   988 => x"34020003",   989 => x"45820026",
      990 => x"34010001",   991 => x"5d81002e",   992 => x"78010001",
      993 => x"31ac0004",   994 => x"38216754",   995 => x"340e0006",
      996 => x"316c001d",   997 => x"302e0000",   998 => x"34020000",
      999 => x"34010001",  1000 => x"34030001",  1001 => x"f800432c",
     1002 => x"29610020",  1003 => x"2821000c",  1004 => x"302e000e",
     1005 => x"b9600800",  1006 => x"f80012ab",  1007 => x"380bea60",
     1008 => x"e000001e",  1009 => x"34010001",  1010 => x"31a10004",
     1011 => x"3161001d",  1012 => x"78010001",  1013 => x"38216754",
     1014 => x"340effbb",  1015 => x"302e0000",  1016 => x"34020000",
     1017 => x"34010002",  1018 => x"34030001",  1019 => x"f800431a",
     1020 => x"29610020",  1021 => x"2821000c",  1022 => x"302e000e",
     1023 => x"b9600800",  1024 => x"f8001299",  1025 => x"340b0fa0",
     1026 => x"e000000c",  1027 => x"31a10004",  1028 => x"3161001d",
     1029 => x"78010001",  1030 => x"38216754",  1031 => x"3402ffff",
     1032 => x"30220000",  1033 => x"34030001",  1034 => x"34010003",
     1035 => x"34020000",  1036 => x"f8004309",  1037 => x"340b0000",
     1038 => x"f800336a",  1039 => x"78020001",  1040 => x"b8207000",
     1041 => x"b8400800",  1042 => x"382138ec",  1043 => x"f8002da5",
     1044 => x"29a20000",  1045 => x"780d0001",  1046 => x"39ad3908",
     1047 => x"28430034",  1048 => x"78020001",  1049 => x"b8400800",
     1050 => x"382160a8",  1051 => x"34020000",  1052 => x"d8600000",
     1053 => x"e000000e",  1054 => x"f80044e4",  1055 => x"340103e8",
     1056 => x"f800335d",  1057 => x"f8003357",  1058 => x"c82e1000",
     1059 => x"51620006",  1060 => x"78010001",  1061 => x"382138f8",
     1062 => x"f8002d92",  1063 => x"340bff8c",  1064 => x"e0000008",
     1065 => x"b9a00800",  1066 => x"f8002d8e",  1067 => x"34010000",
     1068 => x"f80043b3",  1069 => x"5c200002",  1070 => x"5d61fff0",
     1071 => x"340b0000",  1072 => x"78010001",  1073 => x"38214cd8",
     1074 => x"f8002d86",  1075 => x"7d620000",  1076 => x"65810001",
     1077 => x"a0410800",  1078 => x"44200005",  1079 => x"78010001",
     1080 => x"38216754",  1081 => x"34020034",  1082 => x"30220000",
     1083 => x"78010001",  1084 => x"3821754c",  1085 => x"582c0000",
     1086 => x"b9600800",  1087 => x"2b9d0004",  1088 => x"2b8b0014",
     1089 => x"2b8c0010",  1090 => x"2b8d000c",  1091 => x"2b8e0008",
     1092 => x"379c0014",  1093 => x"c3a00000",  1094 => x"379cffec",
     1095 => x"5b8b0014",  1096 => x"5b8c0010",  1097 => x"5b8d000c",
     1098 => x"5b8e0008",  1099 => x"5b9d0004",  1100 => x"78010001",
     1101 => x"38217550",  1102 => x"28210000",  1103 => x"340e0000",
     1104 => x"44200024",  1105 => x"780b0001",  1106 => x"396b60a8",
     1107 => x"29610024",  1108 => x"29620038",  1109 => x"78040001",
     1110 => x"28250008",  1111 => x"3403007c",  1112 => x"b9600800",
     1113 => x"3884618c",  1114 => x"d8a00000",  1115 => x"b8201800",
     1116 => x"4c010005",  1117 => x"29610370",  1118 => x"34210001",
     1119 => x"59610370",  1120 => x"e000000c",  1121 => x"5c20000b",
     1122 => x"780d0001",  1123 => x"f8003315",  1124 => x"39ad7554",
     1125 => x"29a20000",  1126 => x"780c0001",  1127 => x"398c6460",
     1128 => x"c8220800",  1129 => x"29820000",  1130 => x"5441000a",
     1131 => x"e0000011",  1132 => x"78010001",  1133 => x"382160a8",
     1134 => x"28220040",  1135 => x"fbfffd82",  1136 => x"78020001",
     1137 => x"38426460",  1138 => x"58410000",  1139 => x"340e0001",
     1140 => x"b9c00800",  1141 => x"2b9d0004",  1142 => x"2b8b0014",
     1143 => x"2b8c0010",  1144 => x"2b8d000c",  1145 => x"2b8e0008",
     1146 => x"379c0014",  1147 => x"c3a00000",  1148 => x"f80032fc",
     1149 => x"59a10000",  1150 => x"34020000",  1151 => x"b9600800",
     1152 => x"34030000",  1153 => x"fbfffd70",  1154 => x"59810000",
     1155 => x"e3fffff0",  1156 => x"379cffe8",  1157 => x"5b9d0018",
     1158 => x"b8205000",  1159 => x"40610005",  1160 => x"40640000",
     1161 => x"40650001",  1162 => x"40660002",  1163 => x"40670003",
     1164 => x"40680004",  1165 => x"5b810004",  1166 => x"40610006",
     1167 => x"b8404800",  1168 => x"b9401000",  1169 => x"5b810008",
     1170 => x"40610007",  1171 => x"5b81000c",  1172 => x"40610008",
     1173 => x"5b810010",  1174 => x"40610009",  1175 => x"b9201800",
     1176 => x"5b810014",  1177 => x"78010001",  1178 => x"38213910",
     1179 => x"f8002d1d",  1180 => x"2b9d0018",  1181 => x"379c0018",
     1182 => x"c3a00000",  1183 => x"379cffd0",  1184 => x"5b8b0030",
     1185 => x"5b8c002c",  1186 => x"5b8d0028",  1187 => x"5b8e0024",
     1188 => x"5b8f0020",  1189 => x"5b90001c",  1190 => x"5b910018",
     1191 => x"5b920014",  1192 => x"5b930010",  1193 => x"5b94000c",
     1194 => x"5b950008",  1195 => x"5b9d0004",  1196 => x"b8603000",
     1197 => x"b8209800",  1198 => x"b8409000",  1199 => x"78010001",
     1200 => x"b880a800",  1201 => x"38213948",  1202 => x"ba601000",
     1203 => x"ba401800",  1204 => x"b8c02000",  1205 => x"b8a0a000",
     1206 => x"78110001",  1207 => x"f8002d01",  1208 => x"78100001",
     1209 => x"780f0001",  1210 => x"780e0001",  1211 => x"780d0001",
     1212 => x"b8205800",  1213 => x"340c0000",  1214 => x"3a31395c",
     1215 => x"3a103964",  1216 => x"39ef4dfc",  1217 => x"39ce4cd8",
     1218 => x"39ad4b58",  1219 => x"e0000017",  1220 => x"5cc00006",
     1221 => x"ba200800",  1222 => x"ba601000",  1223 => x"ba401800",
     1224 => x"f8002cf0",  1225 => x"b5615800",  1226 => x"b6ac1000",
     1227 => x"40420000",  1228 => x"ba000800",  1229 => x"358c0001",
     1230 => x"f8002cea",  1231 => x"21820003",  1232 => x"b42b5800",
     1233 => x"b9e03000",  1234 => x"5c400005",  1235 => x"2181000f",
     1236 => x"b9c03000",  1237 => x"44220002",  1238 => x"b9a03000",
     1239 => x"b8c00800",  1240 => x"f8002ce0",  1241 => x"b5615800",
     1242 => x"2186000f",  1243 => x"4a8cffe9",  1244 => x"44c00005",
     1245 => x"78010001",  1246 => x"38214cd8",  1247 => x"f8002cd9",
     1248 => x"b42b5800",  1249 => x"b9600800",  1250 => x"2b9d0004",
     1251 => x"2b8b0030",  1252 => x"2b8c002c",  1253 => x"2b8d0028",
     1254 => x"2b8e0024",  1255 => x"2b8f0020",  1256 => x"2b90001c",
     1257 => x"2b910018",  1258 => x"2b920014",  1259 => x"2b930010",
     1260 => x"2b94000c",  1261 => x"2b950008",  1262 => x"379c0030",
     1263 => x"c3a00000",  1264 => x"379cffb8",  1265 => x"5b8b0048",
     1266 => x"5b8c0044",  1267 => x"5b8d0040",  1268 => x"5b8e003c",
     1269 => x"5b8f0038",  1270 => x"5b900034",  1271 => x"5b910030",
     1272 => x"5b92002c",  1273 => x"5b930028",  1274 => x"5b940024",
     1275 => x"5b950020",  1276 => x"5b96001c",  1277 => x"5b970018",
     1278 => x"5b980014",  1279 => x"5b9d0010",  1280 => x"b8608000",
     1281 => x"40430001",  1282 => x"b8206000",  1283 => x"34010002",
     1284 => x"2063000f",  1285 => x"b8406800",  1286 => x"404e0000",
     1287 => x"44610006",  1288 => x"78010001",  1289 => x"b9801000",
     1290 => x"3821396c",  1291 => x"f8002cad",  1292 => x"e000013f",
     1293 => x"40450002",  1294 => x"40460003",  1295 => x"21ce000f",
     1296 => x"3ca50008",  1297 => x"78010001",  1298 => x"b8c52800",
     1299 => x"41a60004",  1300 => x"34030002",  1301 => x"b9c02000",
     1302 => x"344b0022",  1303 => x"3821398c",  1304 => x"b9801000",
     1305 => x"f8002c9f",  1306 => x"41a2000c",  1307 => x"41a1000d",
     1308 => x"41a4000e",  1309 => x"41a30006",  1310 => x"3c420018",
     1311 => x"3c210010",  1312 => x"41a60007",  1313 => x"41a5000f",
     1314 => x"3c840008",  1315 => x"b8220800",  1316 => x"3c630008",
     1317 => x"b8812000",  1318 => x"78010001",  1319 => x"b8c31800",
     1320 => x"b8a42000",  1321 => x"b9801000",  1322 => x"382139b8",
     1323 => x"f8002c8d",  1324 => x"78020001",  1325 => x"b9800800",
     1326 => x"384239dc",  1327 => x"35a30014",  1328 => x"fbffff54",
     1329 => x"41a3001e",  1330 => x"41a4001f",  1331 => x"41a50021",
     1332 => x"3c630008",  1333 => x"78010001",  1334 => x"b8831800",
     1335 => x"41a40020",  1336 => x"382139e4",  1337 => x"b9801000",
     1338 => x"f8002c7e",  1339 => x"3401000c",  1340 => x"55c100d1",
     1341 => x"78010001",  1342 => x"3dce0002",  1343 => x"38215a40",
     1344 => x"b42e0800",  1345 => x"28210000",  1346 => x"c0200000",
     1347 => x"78010001",  1348 => x"b9801000",  1349 => x"38213a10",
     1350 => x"f8002c72",  1351 => x"41620002",  1352 => x"41610003",
     1353 => x"41640004",  1354 => x"3c420018",  1355 => x"3c210010",
     1356 => x"3c840008",  1357 => x"b8220800",  1358 => x"b8812000",
     1359 => x"41620006",  1360 => x"41610007",  1361 => x"41650008",
     1362 => x"3c420018",  1363 => x"3c210010",  1364 => x"3ca50008",
     1365 => x"b8220800",  1366 => x"b8a12800",  1367 => x"78030001",
     1368 => x"78010001",  1369 => x"41670005",  1370 => x"41660009",
     1371 => x"38213a28",  1372 => x"b9801000",  1373 => x"38633a38",
     1374 => x"e000001c",  1375 => x"78010001",  1376 => x"b9801000",
     1377 => x"38213a44",  1378 => x"f8002c56",  1379 => x"41620002",
     1380 => x"41610003",  1381 => x"41640004",  1382 => x"3c420018",
     1383 => x"3c210010",  1384 => x"3c840008",  1385 => x"b8220800",
     1386 => x"b8812000",  1387 => x"41620006",  1388 => x"41610007",
     1389 => x"41650008",  1390 => x"3c420018",  1391 => x"3c210010",
     1392 => x"3ca50008",  1393 => x"b8220800",  1394 => x"41670005",
     1395 => x"41660009",  1396 => x"b8a12800",  1397 => x"78030001",
     1398 => x"78010001",  1399 => x"38213a28",  1400 => x"b9801000",
     1401 => x"38633a60",  1402 => x"b8e42000",  1403 => x"b8c52800",
     1404 => x"f8002c3c",  1405 => x"e000008e",  1406 => x"78010001",
     1407 => x"b9801000",  1408 => x"38213a70",  1409 => x"f8002c37",
     1410 => x"41620002",  1411 => x"41610003",  1412 => x"41640004",
     1413 => x"3c420018",  1414 => x"3c210010",  1415 => x"3c840008",
     1416 => x"b8220800",  1417 => x"b8812000",  1418 => x"41620006",
     1419 => x"41610007",  1420 => x"41650008",  1421 => x"3c420018",
     1422 => x"3c210010",  1423 => x"3ca50008",  1424 => x"b8220800",
     1425 => x"b8a12800",  1426 => x"78030001",  1427 => x"78010001",
     1428 => x"41670005",  1429 => x"41660009",  1430 => x"38213a28",
     1431 => x"b9801000",  1432 => x"38633a8c",  1433 => x"e3ffffe1",
     1434 => x"78010001",  1435 => x"b9801000",  1436 => x"38213a9c",
     1437 => x"f8002c1b",  1438 => x"41620002",  1439 => x"41610003",
     1440 => x"41640004",  1441 => x"3c420018",  1442 => x"3c210010",
     1443 => x"3c840008",  1444 => x"b8220800",  1445 => x"b8812000",
     1446 => x"41620006",  1447 => x"41610007",  1448 => x"41650008",
     1449 => x"3c420018",  1450 => x"3c210010",  1451 => x"41670005",
     1452 => x"41660009",  1453 => x"3ca50008",  1454 => x"b8220800",
     1455 => x"780e0001",  1456 => x"39ce3ab8",  1457 => x"b8a12800",
     1458 => x"78010001",  1459 => x"b9801000",  1460 => x"b9c01800",
     1461 => x"b8e42000",  1462 => x"b8c52800",  1463 => x"38213a28",
     1464 => x"f8002c00",  1465 => x"3563000a",  1466 => x"b9800800",
     1467 => x"b9c01000",  1468 => x"fbfffec8",  1469 => x"340b0036",
     1470 => x"e0000080",  1471 => x"78010001",  1472 => x"b9801000",
     1473 => x"38213acc",  1474 => x"f8002bf6",  1475 => x"41620002",
     1476 => x"41610003",  1477 => x"41640004",  1478 => x"3c420018",
     1479 => x"3c210010",  1480 => x"3c840008",  1481 => x"b8220800",
     1482 => x"b8812000",  1483 => x"41620006",  1484 => x"41610007",
     1485 => x"41650008",  1486 => x"3c420018",  1487 => x"3c210010",
     1488 => x"41670005",  1489 => x"41660009",  1490 => x"3ca50008",
     1491 => x"b8220800",  1492 => x"b8a12800",  1493 => x"78030001",
     1494 => x"78010001",  1495 => x"b8e42000",  1496 => x"b8c52800",
     1497 => x"b9801000",  1498 => x"38633ae8",  1499 => x"38213a28",
     1500 => x"f8002bdc",  1501 => x"41660010",  1502 => x"41670011",
     1503 => x"4165000f",  1504 => x"4164000e",  1505 => x"3cc60008",
     1506 => x"78010001",  1507 => x"78030001",  1508 => x"b8e63000",
     1509 => x"b9801000",  1510 => x"38633b14",  1511 => x"38213b00",
     1512 => x"f8002bd0",  1513 => x"4163000d",  1514 => x"41640012",
     1515 => x"78010001",  1516 => x"b9801000",  1517 => x"38213b38",
     1518 => x"f8002bca",  1519 => x"41610018",  1520 => x"41640013",
     1521 => x"41650014",  1522 => x"41660015",  1523 => x"41670016",
     1524 => x"41680017",  1525 => x"5b810004",  1526 => x"41610019",
     1527 => x"78030001",  1528 => x"b9801000",  1529 => x"5b810008",
     1530 => x"4161001a",  1531 => x"38633b90",  1532 => x"340b0040",
     1533 => x"5b81000c",  1534 => x"78010001",  1535 => x"38213b60",
     1536 => x"f8002bb8",  1537 => x"e000003d",  1538 => x"78010001",
     1539 => x"b9801000",  1540 => x"38213bb0",  1541 => x"f8002bb3",
     1542 => x"78020001",  1543 => x"b9800800",  1544 => x"38423bcc",
     1545 => x"b9601800",  1546 => x"fbfffe7a",  1547 => x"340b002c",
     1548 => x"e0000032",  1549 => x"340b0022",  1550 => x"e0000030",
     1551 => x"55f70009",  1552 => x"78010001",  1553 => x"b9801000",
     1554 => x"ba001800",  1555 => x"b9602000",  1556 => x"b9e02800",
     1557 => x"38213be8",  1558 => x"f8002ba2",  1559 => x"e0000034",
     1560 => x"b5ab7000",  1561 => x"41d60002",  1562 => x"41c10003",
     1563 => x"41c30000",  1564 => x"3ed60008",  1565 => x"41c40001",
     1566 => x"b836b000",  1567 => x"41c10008",  1568 => x"41c50004",
     1569 => x"41c60005",  1570 => x"41c70006",  1571 => x"41c80007",
     1572 => x"5b810004",  1573 => x"41c10009",  1574 => x"3c630008",
     1575 => x"36d10004",  1576 => x"5b810008",  1577 => x"b8831800",
     1578 => x"baa00800",  1579 => x"b9801000",  1580 => x"ba202000",
     1581 => x"f8002b8b",  1582 => x"4df10007",  1583 => x"ba400800",
     1584 => x"b9801000",  1585 => x"ba201800",  1586 => x"b9e02000",
     1587 => x"f8002b85",  1588 => x"e0000008",  1589 => x"b9800800",
     1590 => x"ba801000",  1591 => x"ba601800",  1592 => x"35c4000a",
     1593 => x"36c5fffa",  1594 => x"fbfffe65",  1595 => x"ba207800",
     1596 => x"b56f5800",  1597 => x"e000000b",  1598 => x"78150001",
     1599 => x"78140001",  1600 => x"78130001",  1601 => x"78120001",
     1602 => x"34180002",  1603 => x"34170009",  1604 => x"3ab53c0c",
     1605 => x"3a943c78",  1606 => x"3a733c80",  1607 => x"3a523c4c",
     1608 => x"4d700003",  1609 => x"ca0b7800",  1610 => x"49f8ffc5",
     1611 => x"78020001",  1612 => x"78030001",  1613 => x"b9800800",
     1614 => x"38423c8c",  1615 => x"38633c94",  1616 => x"b9a02000",
     1617 => x"ba002800",  1618 => x"fbfffe4d",  1619 => x"2b9d0010",
     1620 => x"2b8b0048",  1621 => x"2b8c0044",  1622 => x"2b8d0040",
     1623 => x"2b8e003c",  1624 => x"2b8f0038",  1625 => x"2b900034",
     1626 => x"2b910030",  1627 => x"2b92002c",  1628 => x"2b930028",
     1629 => x"2b940024",  1630 => x"2b950020",  1631 => x"2b96001c",
     1632 => x"2b970018",  1633 => x"2b980014",  1634 => x"379c0048",
     1635 => x"c3a00000",  1636 => x"379cfff0",  1637 => x"5b8b0010",
     1638 => x"5b8c000c",  1639 => x"5b8d0008",  1640 => x"5b9d0004",
     1641 => x"b8205800",  1642 => x"b8406800",  1643 => x"b8606000",
     1644 => x"4480000f",  1645 => x"2881000c",  1646 => x"78070001",
     1647 => x"28850000",  1648 => x"28860004",  1649 => x"38e75950",
     1650 => x"5c200003",  1651 => x"78070001",  1652 => x"38e73c9c",
     1653 => x"78010001",  1654 => x"38213ca8",  1655 => x"b9601000",
     1656 => x"b8a01800",  1657 => x"b8a02000",  1658 => x"f8002b3e",
     1659 => x"b9600800",  1660 => x"b9a01000",  1661 => x"b9801800",
     1662 => x"fbfffe72",  1663 => x"34010000",  1664 => x"2b9d0004",
     1665 => x"2b8b0010",  1666 => x"2b8c000c",  1667 => x"2b8d0008",
     1668 => x"379c0010",  1669 => x"c3a00000",  1670 => x"379cffe8",
     1671 => x"5b8b0018",  1672 => x"5b8c0014",  1673 => x"5b8d0010",
     1674 => x"5b8e000c",  1675 => x"5b8f0008",  1676 => x"5b9d0004",
     1677 => x"282d0000",  1678 => x"b8207800",  1679 => x"282e0004",
     1680 => x"b8406000",  1681 => x"340b0000",  1682 => x"34010000",
     1683 => x"34040000",  1684 => x"544d0006",  1685 => x"b9a00800",
     1686 => x"f80044ba",  1687 => x"882c1000",  1688 => x"b9602000",
     1689 => x"c9a26800",  1690 => x"34030000",  1691 => x"34020001",
     1692 => x"e000000b",  1693 => x"3d850001",  1694 => x"3d6b0001",
     1695 => x"f5856000",  1696 => x"3c630001",  1697 => x"b58b5800",
     1698 => x"b8a06000",  1699 => x"3c450001",  1700 => x"f4451000",
     1701 => x"b4431800",  1702 => x"b8a01000",  1703 => x"1565001f",
     1704 => x"c8ac3000",  1705 => x"f4c53000",  1706 => x"c8ab2800",
     1707 => x"c8a62800",  1708 => x"00a5001f",  1709 => x"34060001",
     1710 => x"55ab0004",  1711 => x"5dab0002",  1712 => x"55cc0002",
     1713 => x"34060000",  1714 => x"a0a63000",  1715 => x"5cc0ffea",
     1716 => x"556d000d",  1717 => x"5d6d0002",  1718 => x"558e000b",
     1719 => x"c9cc2800",  1720 => x"f4ae7000",  1721 => x"c9ab6800",
     1722 => x"c9ae6800",  1723 => x"b8a07000",  1724 => x"b4822800",
     1725 => x"f4852000",  1726 => x"b4230800",  1727 => x"b4810800",
     1728 => x"b8a02000",  1729 => x"3c65001f",  1730 => x"00420001",
     1731 => x"00630001",  1732 => x"b8a21000",  1733 => x"b8622800",
     1734 => x"44a00006",  1735 => x"3d65001f",  1736 => x"018c0001",
     1737 => x"016b0001",  1738 => x"b8ac6000",  1739 => x"e3ffffe9",
     1740 => x"59e10000",  1741 => x"b9c00800",  1742 => x"59e40004",
     1743 => x"2b9d0004",  1744 => x"2b8b0018",  1745 => x"2b8c0014",
     1746 => x"2b8d0010",  1747 => x"2b8e000c",  1748 => x"2b8f0008",
     1749 => x"379c0018",  1750 => x"c3a00000",  1751 => x"379cfff8",
     1752 => x"5b8b0008",  1753 => x"5b9d0004",  1754 => x"b8405800",
     1755 => x"f800309d",  1756 => x"b42b0800",  1757 => x"5c200002",
     1758 => x"34010001",  1759 => x"2b9d0004",  1760 => x"2b8b0008",
     1761 => x"379c0008",  1762 => x"c3a00000",  1763 => x"379cfff8",
     1764 => x"5b8b0008",  1765 => x"5b9d0004",  1766 => x"78040001",
     1767 => x"b8405800",  1768 => x"78050001",  1769 => x"34020006",
     1770 => x"34030001",  1771 => x"38843d74",  1772 => x"38a55a74",
     1773 => x"b9603000",  1774 => x"fbfffb64",  1775 => x"45600005",
     1776 => x"1562001f",  1777 => x"34010002",  1778 => x"b9601800",
     1779 => x"f8003408",  1780 => x"34010000",  1781 => x"2b9d0004",
     1782 => x"2b8b0008",  1783 => x"379c0008",  1784 => x"c3a00000",
     1785 => x"379cfff4",  1786 => x"5b8b000c",  1787 => x"5b8c0008",
     1788 => x"5b9d0004",  1789 => x"b8206000",  1790 => x"b8405800",
     1791 => x"b8603000",  1792 => x"44600008",  1793 => x"78040001",
     1794 => x"78050001",  1795 => x"34020006",  1796 => x"34030001",
     1797 => x"38843d80",  1798 => x"38a55a94",  1799 => x"fbfffb4b",
     1800 => x"b9800800",  1801 => x"b9601000",  1802 => x"fbffffd9",
     1803 => x"2b9d0004",  1804 => x"2b8b000c",  1805 => x"2b8c0008",
     1806 => x"379c000c",  1807 => x"c3a00000",  1808 => x"379cfff0",
     1809 => x"5b8b0010",  1810 => x"5b8c000c",  1811 => x"5b8d0008",
     1812 => x"5b9d0004",  1813 => x"b8206800",  1814 => x"44400012",
     1815 => x"284b0000",  1816 => x"284c0004",  1817 => x"34040003",
     1818 => x"1561001f",  1819 => x"b9601000",  1820 => x"b9801800",
     1821 => x"f80033fc",  1822 => x"78040001",  1823 => x"78050001",
     1824 => x"b9a00800",  1825 => x"34020006",  1826 => x"34030001",
     1827 => x"38843dac",  1828 => x"38a55aa8",  1829 => x"b9603000",
     1830 => x"b9803800",  1831 => x"fbfffb2b",  1832 => x"34010000",
     1833 => x"2b9d0004",  1834 => x"2b8b0010",  1835 => x"2b8c000c",
     1836 => x"2b8d0008",  1837 => x"379c0010",  1838 => x"c3a00000",
     1839 => x"379cffe8",  1840 => x"5b8b000c",  1841 => x"5b8c0008",
     1842 => x"5b9d0004",  1843 => x"b8405800",  1844 => x"b8206000",
     1845 => x"37820018",  1846 => x"37810010",  1847 => x"f8003402",
     1848 => x"78020001",  1849 => x"384274c4",  1850 => x"2b860014",
     1851 => x"2b870018",  1852 => x"28410000",  1853 => x"59660000",
     1854 => x"59670004",  1855 => x"20210001",  1856 => x"5c200009",
     1857 => x"78040001",  1858 => x"78050001",  1859 => x"b9800800",
     1860 => x"34020006",  1861 => x"34030002",  1862 => x"38843dac",
     1863 => x"38a55ab8",  1864 => x"fbfffb0a",  1865 => x"34010000",
     1866 => x"2b9d0004",  1867 => x"2b8b000c",  1868 => x"2b8c0008",
     1869 => x"379c0018",  1870 => x"c3a00000",  1871 => x"379cffb0",
     1872 => x"5b8b001c",  1873 => x"5b8c0018",  1874 => x"5b8d0014",
     1875 => x"5b8e0010",  1876 => x"5b8f000c",  1877 => x"5b900008",
     1878 => x"5b9d0004",  1879 => x"28300058",  1880 => x"378c0040",
     1881 => x"b8407800",  1882 => x"b8206800",  1883 => x"78020001",
     1884 => x"340188f7",  1885 => x"b8607000",  1886 => x"0f81004c",
     1887 => x"38425a08",  1888 => x"b9800800",  1889 => x"34030006",
     1890 => x"b8805800",  1891 => x"f800444e",  1892 => x"b9801000",
     1893 => x"ba000800",  1894 => x"b9e01800",  1895 => x"b9c02000",
     1896 => x"37850020",  1897 => x"f80022ac",  1898 => x"b8206000",
     1899 => x"45600011",  1900 => x"2b81003c",  1901 => x"2b870024",
     1902 => x"2b880028",  1903 => x"78040001",  1904 => x"78050001",
     1905 => x"5961000c",  1906 => x"59670000",  1907 => x"59680004",
     1908 => x"59600008",  1909 => x"b9a00800",  1910 => x"34020005",
     1911 => x"34030002",  1912 => x"38843dbc",  1913 => x"38a55ac8",
     1914 => x"b9803000",  1915 => x"fbfffad7",  1916 => x"4c0c0010",
     1917 => x"78010001",  1918 => x"382174c4",  1919 => x"28220000",
     1920 => x"29a10018",  1921 => x"b8410800",  1922 => x"00210014",
     1923 => x"34020001",  1924 => x"2021000f",  1925 => x"50410007",
     1926 => x"78010001",  1927 => x"38213ddc",  1928 => x"b9e01000",
     1929 => x"b9c01800",  1930 => x"b9602000",  1931 => x"fbfffed9",
     1932 => x"b9800800",  1933 => x"2b9d0004",  1934 => x"2b8b001c",
     1935 => x"2b8c0018",  1936 => x"2b8d0014",  1937 => x"2b8e0010",
     1938 => x"2b8f000c",  1939 => x"2b900008",  1940 => x"379c0050",
     1941 => x"c3a00000",  1942 => x"379cffb8",  1943 => x"5b8b0014",
     1944 => x"5b8c0010",  1945 => x"5b8d000c",  1946 => x"5b8e0008",
     1947 => x"5b9d0004",  1948 => x"b8207000",  1949 => x"28210058",
     1950 => x"b8602800",  1951 => x"b8406800",  1952 => x"b8805800",
     1953 => x"37820038",  1954 => x"b8a02000",  1955 => x"b9a01800",
     1956 => x"37850018",  1957 => x"f80021fe",  1958 => x"b8206000",
     1959 => x"4560000b",  1960 => x"2b81001c",  1961 => x"59610000",
     1962 => x"2b810020",  1963 => x"59610004",  1964 => x"2b810024",
     1965 => x"59610008",  1966 => x"2b810034",  1967 => x"5961000c",
     1968 => x"2b810030",  1969 => x"59610010",  1970 => x"4c0c0010",
     1971 => x"78040001",  1972 => x"388474c4",  1973 => x"28820000",
     1974 => x"29c10018",  1975 => x"b8410800",  1976 => x"00210014",
     1977 => x"34020001",  1978 => x"2021000f",  1979 => x"50410007",
     1980 => x"78010001",  1981 => x"38213de4",  1982 => x"b9a01000",
     1983 => x"b9801800",  1984 => x"b9602000",  1985 => x"fbfffea3",
     1986 => x"b9800800",  1987 => x"2b9d0004",  1988 => x"2b8b0014",
     1989 => x"2b8c0010",  1990 => x"2b8d000c",  1991 => x"2b8e0008",
     1992 => x"379c0048",  1993 => x"c3a00000",  1994 => x"379cfffc",
     1995 => x"5b9d0004",  1996 => x"28210058",  1997 => x"f800217c",
     1998 => x"34010000",  1999 => x"2b9d0004",  2000 => x"379c0004",
     2001 => x"c3a00000",  2002 => x"379cffd4",  2003 => x"5b8b0010",
     2004 => x"5b8c000c",  2005 => x"5b8d0008",  2006 => x"5b9d0004",
     2007 => x"b8205800",  2008 => x"28210058",  2009 => x"44200002",
     2010 => x"f800216f",  2011 => x"b9600800",  2012 => x"f8000d2a",
     2013 => x"378c0014",  2014 => x"340188f7",  2015 => x"78020001",
     2016 => x"0f810020",  2017 => x"38425a08",  2018 => x"b9800800",
     2019 => x"34030006",  2020 => x"f80043cd",  2021 => x"78010001",
     2022 => x"b9801000",  2023 => x"38216550",  2024 => x"34030001",
     2025 => x"34040000",  2026 => x"f8002116",  2027 => x"b8206000",
     2028 => x"4420000e",  2029 => x"378d0028",  2030 => x"b9a01000",
     2031 => x"f8002100",  2032 => x"b9a01000",  2033 => x"34030006",
     2034 => x"35610060",  2035 => x"f80043be",  2036 => x"3561004c",
     2037 => x"596c0058",  2038 => x"b9a01000",  2039 => x"34030006",
     2040 => x"f80043b9",  2041 => x"596c0044",  2042 => x"34010000",
     2043 => x"2b9d0004",  2044 => x"2b8b0010",  2045 => x"2b8c000c",
     2046 => x"2b8d0008",  2047 => x"379c002c",  2048 => x"c3a00000",
     2049 => x"379cfff8",  2050 => x"5b8b0008",  2051 => x"5b9d0004",
     2052 => x"78040001",  2053 => x"78050001",  2054 => x"34020002",
     2055 => x"34030002",  2056 => x"38843ed0",  2057 => x"38a55b38",
     2058 => x"b8205800",  2059 => x"fbfffa47",  2060 => x"296302c8",
     2061 => x"28610010",  2062 => x"28220064",  2063 => x"34010000",
     2064 => x"44400010",  2065 => x"34010001",  2066 => x"59610004",
     2067 => x"1061000b",  2068 => x"4062000c",  2069 => x"29640028",
     2070 => x"bc411000",  2071 => x"28830018",  2072 => x"084203e8",
     2073 => x"b9600800",  2074 => x"d8600000",  2075 => x"596102d4",
     2076 => x"296102c8",  2077 => x"28210010",  2078 => x"58200064",
     2079 => x"34010001",  2080 => x"2b9d0004",  2081 => x"2b8b0008",
     2082 => x"379c0008",  2083 => x"c3a00000",  2084 => x"379cfff4",
     2085 => x"5b8b000c",  2086 => x"5b8c0008",  2087 => x"5b9d0004",
     2088 => x"78040001",  2089 => x"78050001",  2090 => x"b8606000",
     2091 => x"34020002",  2092 => x"34030002",  2093 => x"38843ed0",
     2094 => x"38a55a8c",  2095 => x"b8205800",  2096 => x"fbfffa22",
     2097 => x"29820024",  2098 => x"296102c8",  2099 => x"20430003",
     2100 => x"28210010",  2101 => x"7c640000",  2102 => x"58240038",
     2103 => x"20440008",  2104 => x"20420004",  2105 => x"7c840000",
     2106 => x"7c420000",  2107 => x"30230035",  2108 => x"58220044",
     2109 => x"58240040",  2110 => x"29610020",  2111 => x"28220010",
     2112 => x"296102c8",  2113 => x"2c210008",  2114 => x"0c41002c",
     2115 => x"2b9d0004",  2116 => x"2b8b000c",  2117 => x"2b8c0008",
     2118 => x"379c000c",  2119 => x"c3a00000",  2120 => x"379cfff8",
     2121 => x"5b8b0008",  2122 => x"5b9d0004",  2123 => x"282202c8",
     2124 => x"78040001",  2125 => x"78050001",  2126 => x"284b0010",
     2127 => x"34030002",  2128 => x"34020002",  2129 => x"38843ed0",
     2130 => x"38a55b7c",  2131 => x"fbfff9ff",  2132 => x"34010000",
     2133 => x"31600005",  2134 => x"2b9d0004",  2135 => x"2b8b0008",
     2136 => x"379c0008",  2137 => x"c3a00000",  2138 => x"379cfff8",
     2139 => x"5b8b0008",  2140 => x"5b9d0004",  2141 => x"78040001",
     2142 => x"78050001",  2143 => x"b8205800",  2144 => x"34020002",
     2145 => x"34010000",  2146 => x"34030002",  2147 => x"38843ed0",
     2148 => x"38a55b8c",  2149 => x"fbfff9ed",  2150 => x"29610024",
     2151 => x"44200006",  2152 => x"34020000",  2153 => x"34030001",
     2154 => x"34040002",  2155 => x"34060003",  2156 => x"e000001f",
     2157 => x"29610000",  2158 => x"29620040",  2159 => x"58220014",
     2160 => x"e000001d",  2161 => x"29650000",  2162 => x"08410374",
     2163 => x"b4a10800",  2164 => x"29650040",  2165 => x"58250014",
     2166 => x"28250368",  2167 => x"5ca30010",  2168 => x"4025001d",
     2169 => x"44a30004",  2170 => x"282102c8",  2171 => x"5ca40009",
     2172 => x"e0000005",  2173 => x"282102c8",  2174 => x"28210010",
     2175 => x"30230004",  2176 => x"e000000a",  2177 => x"28210010",
     2178 => x"30240004",  2179 => x"e0000007",  2180 => x"28210010",
     2181 => x"30260004",  2182 => x"e0000004",  2183 => x"282102c8",
     2184 => x"28210010",  2185 => x"30200004",  2186 => x"34420001",
     2187 => x"29610024",  2188 => x"4822ffe5",  2189 => x"34010000",
     2190 => x"2b9d0004",  2191 => x"2b8b0008",  2192 => x"379c0008",
     2193 => x"c3a00000",  2194 => x"379cfff4",  2195 => x"5b8b000c",
     2196 => x"5b8c0008",  2197 => x"5b9d0004",  2198 => x"282202c8",
     2199 => x"78040001",  2200 => x"78050001",  2201 => x"284b0010",
     2202 => x"34030002",  2203 => x"34020002",  2204 => x"38843ed0",
     2205 => x"38a55b94",  2206 => x"b8206000",  2207 => x"fbfff9b3",
     2208 => x"41630004",  2209 => x"3401012c",  2210 => x"59610028",
     2211 => x"34020001",  2212 => x"34010bb8",  2213 => x"59610030",
     2214 => x"59600008",  2215 => x"31600035",  2216 => x"59600040",
     2217 => x"59620014",  2218 => x"20630003",  2219 => x"29610000",
     2220 => x"5c620004",  2221 => x"28230034",  2222 => x"b9800800",
     2223 => x"e0000004",  2224 => x"28230034",  2225 => x"34020000",
     2226 => x"b9800800",  2227 => x"d8600000",  2228 => x"34010000",
     2229 => x"2b9d0004",  2230 => x"2b8b000c",  2231 => x"2b8c0008",
     2232 => x"379c000c",  2233 => x"c3a00000",  2234 => x"379cfff0",
     2235 => x"5b8b0010",  2236 => x"5b8c000c",  2237 => x"5b8d0008",
     2238 => x"5b9d0004",  2239 => x"78040001",  2240 => x"78050001",
     2241 => x"2c2d0002",  2242 => x"b8205800",  2243 => x"b8406000",
     2244 => x"34010000",  2245 => x"34020002",  2246 => x"34030002",
     2247 => x"38843ed0",  2248 => x"38a55ad8",  2249 => x"fbfff989",
     2250 => x"34010040",  2251 => x"4c2d0004",  2252 => x"b9600800",
     2253 => x"b9801000",  2254 => x"f8000466",  2255 => x"2b9d0004",
     2256 => x"2b8b0010",  2257 => x"2b8c000c",  2258 => x"2b8d0008",
     2259 => x"379c0010",  2260 => x"c3a00000",  2261 => x"379cfff8",
     2262 => x"5b8b0008",  2263 => x"5b9d0004",  2264 => x"78040001",
     2265 => x"78050001",  2266 => x"34020002",  2267 => x"34030002",
     2268 => x"38843ed0",  2269 => x"38a55afc",  2270 => x"b8205800",
     2271 => x"fbfff973",  2272 => x"296102c8",  2273 => x"34020040",
     2274 => x"28210010",  2275 => x"40210004",  2276 => x"44200006",
     2277 => x"34030002",  2278 => x"44230004",  2279 => x"b9600800",
     2280 => x"f8000409",  2281 => x"3402004e",  2282 => x"b8400800",
     2283 => x"2b9d0004",  2284 => x"2b8b0008",  2285 => x"379c0008",
     2286 => x"c3a00000",  2287 => x"379cfff4",  2288 => x"5b8b000c",
     2289 => x"5b8c0008",  2290 => x"5b9d0004",  2291 => x"78040001",
     2292 => x"78050001",  2293 => x"34030002",  2294 => x"b8406000",
     2295 => x"38843ed0",  2296 => x"34020002",  2297 => x"38a55b10",
     2298 => x"b8205800",  2299 => x"fbfff957",  2300 => x"296102c8",
     2301 => x"34030000",  2302 => x"28210010",  2303 => x"28210008",
     2304 => x"44200007",  2305 => x"35630094",  2306 => x"59800008",
     2307 => x"b9600800",  2308 => x"b9801000",  2309 => x"f80005e9",
     2310 => x"34030001",  2311 => x"b8600800",  2312 => x"2b9d0004",
     2313 => x"2b8b000c",  2314 => x"2b8c0008",  2315 => x"379c000c",
     2316 => x"c3a00000",  2317 => x"379cfff8",  2318 => x"5b8b0008",
     2319 => x"5b9d0004",  2320 => x"78040001",  2321 => x"78050001",
     2322 => x"34020002",  2323 => x"34030002",  2324 => x"38843ed0",
     2325 => x"38a55b24",  2326 => x"b8205800",  2327 => x"fbfff93b",
     2328 => x"296102c8",  2329 => x"28220010",  2330 => x"40410004",
     2331 => x"20210002",  2332 => x"4420000b",  2333 => x"40410035",
     2334 => x"20210001",  2335 => x"44200008",  2336 => x"28410008",
     2337 => x"44200003",  2338 => x"28410040",  2339 => x"5c200004",
     2340 => x"b9600800",  2341 => x"34020009",  2342 => x"f80000a1",
     2343 => x"2b9d0004",  2344 => x"2b8b0008",  2345 => x"379c0008",
     2346 => x"c3a00000",  2347 => x"379cffdc",  2348 => x"5b8b0010",
     2349 => x"5b8c000c",  2350 => x"5b8d0008",  2351 => x"5b9d0004",
     2352 => x"28220020",  2353 => x"78040001",  2354 => x"78050001",
     2355 => x"284d0010",  2356 => x"282202c8",  2357 => x"34030002",
     2358 => x"38843ed0",  2359 => x"284c0010",  2360 => x"38a55b4c",
     2361 => x"34020002",  2362 => x"b8205800",  2363 => x"fbfff917",
     2364 => x"29620318",  2365 => x"2963031c",  2366 => x"37810014",
     2367 => x"f80010df",  2368 => x"29810008",  2369 => x"5c200019",
     2370 => x"296200a0",  2371 => x"44410003",  2372 => x"296100b4",
     2373 => x"5c200008",  2374 => x"78040001",  2375 => x"b9600800",
     2376 => x"34020004",  2377 => x"34030001",  2378 => x"38843edc",
     2379 => x"fbfff907",  2380 => x"e0000013",  2381 => x"b9600800",
     2382 => x"f80011d1",  2383 => x"29a20004",  2384 => x"29810000",
     2385 => x"44400005",  2386 => x"28230034",  2387 => x"34020000",
     2388 => x"b9600800",  2389 => x"e0000004",  2390 => x"28230034",
     2391 => x"34020001",  2392 => x"b9600800",  2393 => x"d8600000",
     2394 => x"29620318",  2395 => x"b9600800",  2396 => x"f80005ac",
     2397 => x"b9600800",  2398 => x"f80005d4",  2399 => x"34010000",
     2400 => x"2b9d0004",  2401 => x"2b8b0010",  2402 => x"2b8c000c",
     2403 => x"2b8d0008",  2404 => x"379c0024",  2405 => x"c3a00000",
     2406 => x"379cfff8",  2407 => x"5b8b0008",  2408 => x"5b9d0004",
     2409 => x"78040001",  2410 => x"78050001",  2411 => x"34020002",
     2412 => x"34030002",  2413 => x"38843ed0",  2414 => x"38a55b5c",
     2415 => x"b8205800",  2416 => x"fbfff8e2",  2417 => x"b9600800",
     2418 => x"f8000523",  2419 => x"34010000",  2420 => x"2b9d0004",
     2421 => x"2b8b0008",  2422 => x"379c0008",  2423 => x"c3a00000",
     2424 => x"379cffd8",  2425 => x"5b8b0010",  2426 => x"5b8c000c",
     2427 => x"5b8d0008",  2428 => x"5b9d0004",  2429 => x"78050001",
     2430 => x"b8806000",  2431 => x"78040001",  2432 => x"b8406800",
     2433 => x"34030002",  2434 => x"34020002",  2435 => x"38843ed0",
     2436 => x"38a55b6c",  2437 => x"b8205800",  2438 => x"fbfff8cc",
     2439 => x"34010001",  2440 => x"45810004",  2441 => x"3401000c",
     2442 => x"5d810036",  2443 => x"e0000022",  2444 => x"296200ec",
     2445 => x"5960031c",  2446 => x"37810024",  2447 => x"4802000c",
     2448 => x"1443001f",  2449 => x"00440010",  2450 => x"3c630010",
     2451 => x"3c420010",  2452 => x"b8641800",  2453 => x"5b820028",
     2454 => x"340203e8",  2455 => x"5b830024",  2456 => x"fbfffcee",
     2457 => x"2b810028",  2458 => x"e000000d",  2459 => x"c8021000",
     2460 => x"1443001f",  2461 => x"00440010",  2462 => x"3c630010",
     2463 => x"3c420010",  2464 => x"b8641800",  2465 => x"5b820028",
     2466 => x"340203e8",  2467 => x"5b830024",  2468 => x"fbfffce2",
     2469 => x"2b810028",  2470 => x"c8010800",  2471 => x"59610318",
     2472 => x"356200e4",  2473 => x"b9600800",  2474 => x"f8001013",
     2475 => x"340c0100",  2476 => x"e0000014",  2477 => x"296102c8",
     2478 => x"b9a01000",  2479 => x"37830014",  2480 => x"28240010",
     2481 => x"b9600800",  2482 => x"340c0100",  2483 => x"3484003c",
     2484 => x"f8000416",  2485 => x"296102c8",  2486 => x"34021000",
     2487 => x"28210010",  2488 => x"2c23003c",  2489 => x"5c620007",
     2490 => x"40210004",  2491 => x"20210001",  2492 => x"44200004",
     2493 => x"b9600800",  2494 => x"34020006",  2495 => x"f8000008",
     2496 => x"b9800800",  2497 => x"2b9d0004",  2498 => x"2b8b0010",
     2499 => x"2b8c000c",  2500 => x"2b8d0008",  2501 => x"379c0028",
     2502 => x"c3a00000",  2503 => x"282302c8",  2504 => x"34040006",
     2505 => x"28630010",  2506 => x"44440004",  2507 => x"34040009",
     2508 => x"5c440008",  2509 => x"e0000004",  2510 => x"34020001",
     2511 => x"30620005",  2512 => x"e0000007",  2513 => x"34020002",
     2514 => x"30620005",  2515 => x"e0000006",  2516 => x"40630005",
     2517 => x"34020001",  2518 => x"5c620003",  2519 => x"34020066",
     2520 => x"e0000002",  2521 => x"34020064",  2522 => x"58220004",
     2523 => x"c3a00000",  2524 => x"379cfff4",  2525 => x"5b8b000c",
     2526 => x"5b8c0008",  2527 => x"5b9d0004",  2528 => x"b8205800",
     2529 => x"282102c8",  2530 => x"78050001",  2531 => x"38a53e2c",
     2532 => x"282c0010",  2533 => x"34010001",  2534 => x"41820005",
     2535 => x"5c410003",  2536 => x"78050001",  2537 => x"38a54314",
     2538 => x"78040001",  2539 => x"b9600800",  2540 => x"34020002",
     2541 => x"34030001",  2542 => x"38843f04",  2543 => x"fbfff863",
     2544 => x"41820005",  2545 => x"34010001",  2546 => x"5c410003",
     2547 => x"34010006",  2548 => x"e0000002",  2549 => x"34010009",
     2550 => x"59610004",  2551 => x"31800005",  2552 => x"2b9d0004",
     2553 => x"2b8b000c",  2554 => x"2b8c0008",  2555 => x"379c000c",
     2556 => x"c3a00000",  2557 => x"379cfffc",  2558 => x"5b9d0004",
     2559 => x"282202c8",  2560 => x"28420010",  2561 => x"4043002c",
     2562 => x"4460000a",  2563 => x"3463ffff",  2564 => x"78040001",
     2565 => x"3043002c",  2566 => x"38843f28",  2567 => x"34020002",
     2568 => x"34030001",  2569 => x"fbfff849",  2570 => x"34010001",
     2571 => x"e0000003",  2572 => x"fbffffd0",  2573 => x"34010000",
     2574 => x"2b9d0004",  2575 => x"379c0004",  2576 => x"c3a00000",
     2577 => x"379cffd8",  2578 => x"5b8b0018",  2579 => x"5b8c0014",
     2580 => x"5b8d0010",  2581 => x"5b8e000c",  2582 => x"5b8f0008",
     2583 => x"5b9d0004",  2584 => x"b8407000",  2585 => x"2824000c",
     2586 => x"282202c8",  2587 => x"b8205800",  2588 => x"b8607800",
     2589 => x"284d0010",  2590 => x"44800004",  2591 => x"34010003",
     2592 => x"31a1002c",  2593 => x"e000000c",  2594 => x"282202e0",
     2595 => x"44440008",  2596 => x"28220028",  2597 => x"28440018",
     2598 => x"34020000",  2599 => x"d8800000",  2600 => x"296202e0",
     2601 => x"c8220800",  2602 => x"4c20003c",  2603 => x"340c0000",
     2604 => x"e0000015",  2605 => x"29610028",  2606 => x"340203e8",
     2607 => x"28240018",  2608 => x"b9600800",  2609 => x"d8800000",
     2610 => x"596102e0",  2611 => x"296102c8",  2612 => x"29620028",
     2613 => x"4025000c",  2614 => x"1021000b",  2615 => x"28440018",
     2616 => x"bca12800",  2617 => x"b9600800",  2618 => x"08a203e8",
     2619 => x"d8800000",  2620 => x"596102d4",  2621 => x"34021000",
     2622 => x"b9600800",  2623 => x"f80003fb",  2624 => x"b8206000",
     2625 => x"45e0000e",  2626 => x"4162030d",  2627 => x"3401000c",
     2628 => x"5c41000b",  2629 => x"b9600800",  2630 => x"b9c01000",
     2631 => x"3783001c",  2632 => x"35a4003c",  2633 => x"f8000381",
     2634 => x"2da2003c",  2635 => x"34011001",  2636 => x"5c410003",
     2637 => x"34010065",  2638 => x"59610004",  2639 => x"5d800004",
     2640 => x"b9600800",  2641 => x"f8000adb",  2642 => x"e0000003",
     2643 => x"34010002",  2644 => x"59610004",  2645 => x"29620004",
     2646 => x"29610000",  2647 => x"44410002",  2648 => x"596002d4",
     2649 => x"296102c8",  2650 => x"28210010",  2651 => x"28210028",
     2652 => x"59610008",  2653 => x"b9800800",  2654 => x"2b9d0004",
     2655 => x"2b8b0018",  2656 => x"2b8c0014",  2657 => x"2b8d0010",
     2658 => x"2b8e000c",  2659 => x"2b8f0008",  2660 => x"379c0028",
     2661 => x"c3a00000",  2662 => x"b9600800",  2663 => x"34020005",
     2664 => x"f800127b",  2665 => x"b9600800",  2666 => x"596002e0",
     2667 => x"fbffff92",  2668 => x"340c0000",  2669 => x"5c20ffc0",
     2670 => x"e3ffffef",  2671 => x"379cffd8",  2672 => x"5b8b0018",
     2673 => x"5b8c0014",  2674 => x"5b8d0010",  2675 => x"5b8e000c",
     2676 => x"5b8f0008",  2677 => x"5b9d0004",  2678 => x"b8407000",
     2679 => x"2824000c",  2680 => x"282202c8",  2681 => x"b8205800",
     2682 => x"b8607800",  2683 => x"284c0010",  2684 => x"44800004",
     2685 => x"34010003",  2686 => x"3181002c",  2687 => x"e000000c",
     2688 => x"282202e0",  2689 => x"44440008",  2690 => x"28220028",
     2691 => x"28440018",  2692 => x"34020000",  2693 => x"d8800000",
     2694 => x"296202e0",  2695 => x"c8220800",  2696 => x"4c200029",
     2697 => x"340d0000",  2698 => x"e000000b",  2699 => x"34021001",
     2700 => x"b9600800",  2701 => x"f80003ad",  2702 => x"b8206800",
     2703 => x"29610028",  2704 => x"34023a98",  2705 => x"28240018",
     2706 => x"b9600800",  2707 => x"d8800000",  2708 => x"596102e0",
     2709 => x"45e0000e",  2710 => x"4162030d",  2711 => x"3401000c",
     2712 => x"5c41000b",  2713 => x"b9600800",  2714 => x"b9c01000",
     2715 => x"3783001c",  2716 => x"3584003c",  2717 => x"f800032d",
     2718 => x"2d82003c",  2719 => x"34011002",  2720 => x"5c410003",
     2721 => x"34010068",  2722 => x"59610004",  2723 => x"45a00003",
     2724 => x"34010002",  2725 => x"59610004",  2726 => x"29810028",
     2727 => x"59610008",  2728 => x"b9a00800",  2729 => x"2b9d0004",
     2730 => x"2b8b0018",  2731 => x"2b8c0014",  2732 => x"2b8d0010",
     2733 => x"2b8e000c",  2734 => x"2b8f0008",  2735 => x"379c0028",
     2736 => x"c3a00000",  2737 => x"b9600800",  2738 => x"34020005",
     2739 => x"f8001230",  2740 => x"b9600800",  2741 => x"596002e0",
     2742 => x"fbffff47",  2743 => x"340d0000",  2744 => x"5c20ffd3",
     2745 => x"e3ffffef",  2746 => x"379cfff4",  2747 => x"5b8b000c",
     2748 => x"5b8c0008",  2749 => x"5b9d0004",  2750 => x"282202c8",
     2751 => x"b8205800",  2752 => x"284c0010",  2753 => x"2822000c",
     2754 => x"44400004",  2755 => x"34010003",  2756 => x"3181002c",
     2757 => x"e000000b",  2758 => x"282302e0",  2759 => x"44620013",
     2760 => x"28220028",  2761 => x"28430018",  2762 => x"34020000",
     2763 => x"d8600000",  2764 => x"296202e0",  2765 => x"c8220800",
     2766 => x"4c200021",  2767 => x"e000000b",  2768 => x"29810000",
     2769 => x"28220000",  2770 => x"b9600800",  2771 => x"d8400000",
     2772 => x"29610028",  2773 => x"34023a98",  2774 => x"28230018",
     2775 => x"b9600800",  2776 => x"d8600000",  2777 => x"596102e0",
     2778 => x"29810000",  2779 => x"34020000",  2780 => x"28230004",
     2781 => x"b9600800",  2782 => x"d8600000",  2783 => x"34020001",
     2784 => x"5c220007",  2785 => x"34010067",  2786 => x"59610004",
     2787 => x"29810000",  2788 => x"28220008",  2789 => x"b9600800",
     2790 => x"d8400000",  2791 => x"29810028",  2792 => x"59610008",
     2793 => x"34010000",  2794 => x"2b9d0004",  2795 => x"2b8b000c",
     2796 => x"2b8c0008",  2797 => x"379c000c",  2798 => x"c3a00000",
     2799 => x"b9600800",  2800 => x"34020005",  2801 => x"f80011f2",
     2802 => x"29810000",  2803 => x"596002e0",  2804 => x"28220008",
     2805 => x"b9600800",  2806 => x"d8400000",  2807 => x"b9600800",
     2808 => x"fbffff05",  2809 => x"5c20ffd7",  2810 => x"e3ffffef",
     2811 => x"379cffd8",  2812 => x"5b8b0018",  2813 => x"5b8c0014",
     2814 => x"5b8d0010",  2815 => x"5b8e000c",  2816 => x"5b8f0008",
     2817 => x"5b9d0004",  2818 => x"b8407000",  2819 => x"2824000c",
     2820 => x"282202c8",  2821 => x"b8205800",  2822 => x"b8607800",
     2823 => x"284c0010",  2824 => x"44800004",  2825 => x"34010003",
     2826 => x"3181002c",  2827 => x"e000000c",  2828 => x"282202e0",
     2829 => x"44440008",  2830 => x"28220028",  2831 => x"28440018",
     2832 => x"34020000",  2833 => x"d8800000",  2834 => x"296202e0",
     2835 => x"c8220800",  2836 => x"4c200029",  2837 => x"340d0000",
     2838 => x"e000000b",  2839 => x"29610028",  2840 => x"29820028",
     2841 => x"28240018",  2842 => x"b9600800",  2843 => x"d8800000",
     2844 => x"596102e0",  2845 => x"34021002",  2846 => x"b9600800",
     2847 => x"f800031b",  2848 => x"b8206800",  2849 => x"45e0000e",
     2850 => x"4162030d",  2851 => x"3401000c",  2852 => x"5c41000b",
     2853 => x"b9600800",  2854 => x"b9c01000",  2855 => x"3783001c",
     2856 => x"3584003c",  2857 => x"f80002a1",  2858 => x"2d82003c",
     2859 => x"34011003",  2860 => x"5c410003",  2861 => x"3401006a",
     2862 => x"59610004",  2863 => x"45a00003",  2864 => x"34010002",
     2865 => x"59610004",  2866 => x"29810028",  2867 => x"59610008",
     2868 => x"b9a00800",  2869 => x"2b9d0004",  2870 => x"2b8b0018",
     2871 => x"2b8c0014",  2872 => x"2b8d0010",  2873 => x"2b8e000c",
     2874 => x"2b8f0008",  2875 => x"379c0028",  2876 => x"c3a00000",
     2877 => x"b9600800",  2878 => x"34020005",  2879 => x"f80011a4",
     2880 => x"b9600800",  2881 => x"596002e0",  2882 => x"fbfffebb",
     2883 => x"340d0000",  2884 => x"5c20ffd3",  2885 => x"e3ffffef",
     2886 => x"379cffec",  2887 => x"5b8b0010",  2888 => x"5b8c000c",
     2889 => x"5b8d0008",  2890 => x"5b9d0004",  2891 => x"282202c8",
     2892 => x"b8206000",  2893 => x"284b0010",  2894 => x"2822000c",
     2895 => x"44400004",  2896 => x"34010003",  2897 => x"3161002c",
     2898 => x"e000000c",  2899 => x"282302e0",  2900 => x"44620008",
     2901 => x"28220028",  2902 => x"28430018",  2903 => x"34020000",
     2904 => x"d8600000",  2905 => x"298202e0",  2906 => x"c8220800",
     2907 => x"4c2000a9",  2908 => x"340d0000",  2909 => x"e0000011",
     2910 => x"29810028",  2911 => x"29620030",  2912 => x"28230018",
     2913 => x"b9800800",  2914 => x"d8600000",  2915 => x"598102e0",
     2916 => x"34021003",  2917 => x"b9800800",  2918 => x"f80002d4",
     2919 => x"b8206800",  2920 => x"3401006c",  2921 => x"31610010",
     2922 => x"29610014",  2923 => x"44200003",  2924 => x"3401006e",
     2925 => x"31610010",  2926 => x"41660010",  2927 => x"78040001",
     2928 => x"78050001",  2929 => x"b9800800",  2930 => x"34020002",
     2931 => x"34030001",  2932 => x"38843f3c",  2933 => x"38a55bc0",
     2934 => x"34c6ff94",  2935 => x"fbfff6db",  2936 => x"41620010",
     2937 => x"34010008",  2938 => x"3442ff94",  2939 => x"204200ff",
     2940 => x"5441007f",  2941 => x"78010001",  2942 => x"3c420002",
     2943 => x"38215b9c",  2944 => x"b4220800",  2945 => x"28210000",
     2946 => x"c0200000",  2947 => x"29610000",  2948 => x"34020000",
     2949 => x"34030000",  2950 => x"2825002c",  2951 => x"34040000",
     2952 => x"b9800800",  2953 => x"d8a00000",  2954 => x"5c200071",
     2955 => x"3401006d",  2956 => x"31610010",  2957 => x"29610000",
     2958 => x"34020001",  2959 => x"28230024",  2960 => x"b9800800",
     2961 => x"d8600000",  2962 => x"5c200069",  2963 => x"3401006e",
     2964 => x"31610010",  2965 => x"29610000",  2966 => x"34020001",
     2967 => x"37830014",  2968 => x"28240028",  2969 => x"b9800800",
     2970 => x"d8800000",  2971 => x"34020001",  2972 => x"5c22005f",
     2973 => x"2b810014",  2974 => x"78040001",  2975 => x"34020002",
     2976 => x"00250010",  2977 => x"3c210010",  2978 => x"5965001c",
     2979 => x"59610018",  2980 => x"34030001",  2981 => x"b9800800",
     2982 => x"38843f50",  2983 => x"fbfff6ab",  2984 => x"29650018",
     2985 => x"78040001",  2986 => x"b9800800",  2987 => x"34020002",
     2988 => x"34030001",  2989 => x"38843f74",  2990 => x"fbfff6a4",
     2991 => x"3401006f",  2992 => x"31610010",  2993 => x"29610000",
     2994 => x"34020001",  2995 => x"28230020",  2996 => x"b9800800",
     2997 => x"d8600000",  2998 => x"5c200045",  2999 => x"34010070",
     3000 => x"31610010",  3001 => x"29610000",  3002 => x"28220030",
     3003 => x"b9800800",  3004 => x"d8400000",  3005 => x"5c20003e",
     3006 => x"34010071",  3007 => x"31610010",  3008 => x"29610000",
     3009 => x"34020002",  3010 => x"28230024",  3011 => x"b9800800",
     3012 => x"d8600000",  3013 => x"5c200036",  3014 => x"34010072",
     3015 => x"31610010",  3016 => x"29610000",  3017 => x"34020002",
     3018 => x"37830014",  3019 => x"28240028",  3020 => x"b9800800",
     3021 => x"d8800000",  3022 => x"34020001",  3023 => x"5c22002c",
     3024 => x"2b850014",  3025 => x"78040001",  3026 => x"b9800800",
     3027 => x"34020002",  3028 => x"34030001",  3029 => x"38843f98",
     3030 => x"fbfff67c",  3031 => x"2b810014",  3032 => x"78040001",
     3033 => x"34020002",  3034 => x"00250010",  3035 => x"3c210010",
     3036 => x"59650024",  3037 => x"59610020",  3038 => x"34030001",
     3039 => x"b9800800",  3040 => x"38843fb0",  3041 => x"fbfff671",
     3042 => x"29650020",  3043 => x"78040001",  3044 => x"b9800800",
     3045 => x"34020002",  3046 => x"34030001",  3047 => x"38843fd4",
     3048 => x"fbfff66a",  3049 => x"34010073",  3050 => x"31610010",
     3051 => x"29610000",  3052 => x"34020002",  3053 => x"28230020",
     3054 => x"b9800800",  3055 => x"d8600000",  3056 => x"5c20000b",
     3057 => x"34010074",  3058 => x"31610010",  3059 => x"b9800800",
     3060 => x"34021004",  3061 => x"f8000245",  3062 => x"b8206800",
     3063 => x"34010069",  3064 => x"59810004",  3065 => x"34010001",
     3066 => x"59610014",  3067 => x"29610028",  3068 => x"59810008",
     3069 => x"b9a00800",  3070 => x"2b9d0004",  3071 => x"2b8b0010",
     3072 => x"2b8c000c",  3073 => x"2b8d0008",  3074 => x"379c0014",
     3075 => x"c3a00000",  3076 => x"b9800800",  3077 => x"34020005",
     3078 => x"f80010dd",  3079 => x"b9800800",  3080 => x"598002e0",
     3081 => x"fbfffdf4",  3082 => x"340d0000",  3083 => x"5c20ff53",
     3084 => x"e3fffff1",  3085 => x"379cffdc",  3086 => x"5b8b0014",
     3087 => x"5b8c0010",  3088 => x"5b8d000c",  3089 => x"5b8e0008",
     3090 => x"5b9d0004",  3091 => x"b8406800",  3092 => x"282202c8",
     3093 => x"b8205800",  3094 => x"b8607000",  3095 => x"284c0010",
     3096 => x"2822000c",  3097 => x"44400006",  3098 => x"28220028",
     3099 => x"28440018",  3100 => x"29820028",  3101 => x"d8800000",
     3102 => x"596102e0",  3103 => x"296102e0",  3104 => x"44200009",
     3105 => x"29610028",  3106 => x"34020000",  3107 => x"28240018",
     3108 => x"b9600800",  3109 => x"d8800000",  3110 => x"296202e0",
     3111 => x"c8220800",  3112 => x"4c200023",  3113 => x"45c00018",
     3114 => x"4162030d",  3115 => x"3401000c",  3116 => x"5c410015",
     3117 => x"b9600800",  3118 => x"b9a01000",  3119 => x"37830018",
     3120 => x"3584003c",  3121 => x"f8000199",  3122 => x"2d81003c",
     3123 => x"34021003",  3124 => x"5c220006",  3125 => x"41820005",
     3126 => x"34010001",  3127 => x"5c41000a",  3128 => x"3401006a",
     3129 => x"e0000007",  3130 => x"34021005",  3131 => x"5c220006",
     3132 => x"41820005",  3133 => x"34010002",  3134 => x"5c410003",
     3135 => x"3401006b",  3136 => x"59610004",  3137 => x"29810028",
     3138 => x"59610008",  3139 => x"34010000",  3140 => x"2b9d0004",
     3141 => x"2b8b0014",  3142 => x"2b8c0010",  3143 => x"2b8d000c",
     3144 => x"2b8e0008",  3145 => x"379c0024",  3146 => x"c3a00000",
     3147 => x"b9600800",  3148 => x"34020005",  3149 => x"f8001096",
     3150 => x"b9600800",  3151 => x"596002e0",  3152 => x"fbfffd8c",
     3153 => x"e3fffff2",  3154 => x"379cffd4",  3155 => x"5b8b001c",
     3156 => x"5b8c0018",  3157 => x"5b8d0014",  3158 => x"5b8e0010",
     3159 => x"5b8f000c",  3160 => x"5b900008",  3161 => x"5b9d0004",
     3162 => x"b8407000",  3163 => x"282202c8",  3164 => x"2824000c",
     3165 => x"b8205800",  3166 => x"284c0010",  3167 => x"b8607800",
     3168 => x"2d8d0048",  3169 => x"7dad0000",  3170 => x"44800004",
     3171 => x"34010003",  3172 => x"3181002c",  3173 => x"e0000012",
     3174 => x"282202e0",  3175 => x"44440022",  3176 => x"28220028",
     3177 => x"28440018",  3178 => x"34020000",  3179 => x"d8800000",
     3180 => x"296202e0",  3181 => x"c8220800",  3182 => x"4c20003f",
     3183 => x"e000001a",  3184 => x"29810000",  3185 => x"28240030",
     3186 => x"b9600800",  3187 => x"d8800000",  3188 => x"b9600800",
     3189 => x"fbfffd88",  3190 => x"4420002d",  3191 => x"45a00008",
     3192 => x"29810000",  3193 => x"34020000",  3194 => x"34030000",
     3195 => x"2825002c",  3196 => x"34040000",  3197 => x"b9600800",
     3198 => x"d8a00000",  3199 => x"2981004c",  3200 => x"29700028",
     3201 => x"340203e8",  3202 => x"f8003ece",  3203 => x"2a050018",
     3204 => x"b8202000",  3205 => x"b8801000",  3206 => x"b9600800",
     3207 => x"d8a00000",  3208 => x"596102e0",  3209 => x"45e00018",
     3210 => x"4162030d",  3211 => x"3401000c",  3212 => x"5c410015",
     3213 => x"b9600800",  3214 => x"b9c01000",  3215 => x"37830020",
     3216 => x"3584003c",  3217 => x"f8000139",  3218 => x"2d82003c",
     3219 => x"34011004",  3220 => x"5c41000d",  3221 => x"45a00005",
     3222 => x"29810000",  3223 => x"28220030",  3224 => x"b9600800",
     3225 => x"d8400000",  3226 => x"41820005",  3227 => x"34010001",
     3228 => x"5c410003",  3229 => x"3401006b",  3230 => x"e0000002",
     3231 => x"34010068",  3232 => x"59610004",  3233 => x"29810028",
     3234 => x"59610008",  3235 => x"34010000",  3236 => x"2b9d0004",
     3237 => x"2b8b001c",  3238 => x"2b8c0018",  3239 => x"2b8d0014",
     3240 => x"2b8e0010",  3241 => x"2b8f000c",  3242 => x"2b900008",
     3243 => x"379c002c",  3244 => x"c3a00000",  3245 => x"b9600800",
     3246 => x"34020005",  3247 => x"f8001034",  3248 => x"596002e0",
     3249 => x"45a0ffc3",  3250 => x"e3ffffbe",  3251 => x"379cfff0",
     3252 => x"5b8b0010",  3253 => x"5b8c000c",  3254 => x"5b8d0008",
     3255 => x"5b9d0004",  3256 => x"282202c8",  3257 => x"340d0001",
     3258 => x"b8206000",  3259 => x"284b0010",  3260 => x"29620000",
     3261 => x"596d0008",  3262 => x"2842000c",  3263 => x"d8400000",
     3264 => x"41610005",  3265 => x"34020000",  3266 => x"5c2d0005",
     3267 => x"34021005",  3268 => x"b9800800",  3269 => x"f8000175",
     3270 => x"b8201000",  3271 => x"34010001",  3272 => x"59610040",
     3273 => x"3401ffff",  3274 => x"5c400009",  3275 => x"41620005",
     3276 => x"34010002",  3277 => x"5c410003",  3278 => x"34010009",
     3279 => x"e0000002",  3280 => x"34010006",  3281 => x"59810004",
     3282 => x"34010000",  3283 => x"2b9d0004",  3284 => x"2b8b0010",
     3285 => x"2b8c000c",  3286 => x"2b8d0008",  3287 => x"379c0010",
     3288 => x"c3a00000",  3289 => x"00430018",  3290 => x"30220003",
     3291 => x"30230000",  3292 => x"00430010",  3293 => x"30230001",
     3294 => x"00430008",  3295 => x"30230002",  3296 => x"c3a00000",
     3297 => x"40220000",  3298 => x"40230003",  3299 => x"3c420018",
     3300 => x"b8621000",  3301 => x"40230001",  3302 => x"40210002",
     3303 => x"3c630010",  3304 => x"3c210008",  3305 => x"b8431000",
     3306 => x"b8410800",  3307 => x"c3a00000",  3308 => x"40220000",
     3309 => x"40210001",  3310 => x"3c420008",  3311 => x"b8410800",
     3312 => x"c3a00000",  3313 => x"379cfff0",  3314 => x"5b8b0010",
     3315 => x"5b8c000c",  3316 => x"5b8d0008",  3317 => x"5b9d0004",
     3318 => x"28230020",  3319 => x"282202c8",  3320 => x"b8205800",
     3321 => x"2863000c",  3322 => x"28420010",  3323 => x"282c003c",
     3324 => x"4064000e",  3325 => x"340300ba",  3326 => x"48830018",
     3327 => x"28420000",  3328 => x"28430004",  3329 => x"34020001",
     3330 => x"d8600000",  3331 => x"ec016800",  3332 => x"b9600800",
     3333 => x"f8000994",  3334 => x"29610020",  3335 => x"c80d6800",
     3336 => x"21ad002e",  3337 => x"2821000c",  3338 => x"35ad0006",
     3339 => x"4021000e",  3340 => x"45a1000a",  3341 => x"78010001",
     3342 => x"b9a01000",  3343 => x"38213ff8",  3344 => x"f80024a8",
     3345 => x"29610020",  3346 => x"21ad00ff",  3347 => x"2821000c",
     3348 => x"302d000e",  3349 => x"318d0030",  3350 => x"3401004e",
     3351 => x"0d810002",  3352 => x"34010003",  3353 => x"0d810040",
     3354 => x"3401000a",  3355 => x"0d810042",  3356 => x"34010800",
     3357 => x"0d810044",  3358 => x"340130de",  3359 => x"0d810046",
     3360 => x"3401ad01",  3361 => x"0d810048",  3362 => x"34012000",
     3363 => x"0d81004a",  3364 => x"296102c8",  3365 => x"28220010",
     3366 => x"28430014",  3367 => x"40410004",  3368 => x"44600002",
     3369 => x"38210004",  3370 => x"28420008",  3371 => x"44400002",
     3372 => x"38210008",  3373 => x"0d81004c",  3374 => x"2b9d0004",
     3375 => x"2b8b0010",  3376 => x"2b8c000c",  3377 => x"2b8d0008",
     3378 => x"379c0010",  3379 => x"c3a00000",  3380 => x"379cfff4",
     3381 => x"5b8b000c",  3382 => x"5b8c0008",  3383 => x"5b9d0004",
     3384 => x"b8205800",  3385 => x"34210040",  3386 => x"b8406000",
     3387 => x"fbffffb1",  3388 => x"2d650044",  3389 => x"2d640046",
     3390 => x"78070001",  3391 => x"3ca50008",  3392 => x"00860008",
     3393 => x"38e75960",  3394 => x"b8a62800",  3395 => x"28e60000",
     3396 => x"64210003",  3397 => x"2d630048",  3398 => x"e4a62800",
     3399 => x"2d62004a",  3400 => x"a0250800",  3401 => x"44200010",
     3402 => x"3c840008",  3403 => x"00610008",  3404 => x"2084ffff",
     3405 => x"b8812000",  3406 => x"206300ff",  3407 => x"3801dead",
     3408 => x"e4812000",  3409 => x"64630001",  3410 => x"a0831800",
     3411 => x"44600006",  3412 => x"34012000",  3413 => x"5c410004",
     3414 => x"3561004c",  3415 => x"fbffff95",  3416 => x"59810024",
     3417 => x"2b9d0004",  3418 => x"2b8b000c",  3419 => x"2b8c0008",
     3420 => x"379c000c",  3421 => x"c3a00000",  3422 => x"379cfff0",
     3423 => x"5b8b0010",  3424 => x"5b8c000c",  3425 => x"5b8d0008",
     3426 => x"5b9d0004",  3427 => x"b8206000",  3428 => x"282102c8",
     3429 => x"204dffff",  3430 => x"28210010",  3431 => x"40250005",
     3432 => x"44a00003",  3433 => x"34012000",  3434 => x"5da1000a",
     3435 => x"78040001",  3436 => x"b9800800",  3437 => x"34020005",
     3438 => x"34030001",  3439 => x"38844010",  3440 => x"b9a03000",
     3441 => x"fbfff4e1",  3442 => x"34010000",  3443 => x"e0000051",
     3444 => x"298b003c",  3445 => x"34030008",  3446 => x"41610000",
     3447 => x"202100f0",  3448 => x"3821000c",  3449 => x"31610000",
     3450 => x"34010005",  3451 => x"31610020",  3452 => x"29820020",
     3453 => x"35610022",  3454 => x"28420014",  3455 => x"f8003e32",
     3456 => x"29810020",  3457 => x"28210014",  3458 => x"2c210008",
     3459 => x"0d6d0036",  3460 => x"00220008",  3461 => x"3161002b",
     3462 => x"34010003",  3463 => x"0d61002c",  3464 => x"34010800",
     3465 => x"0d610030",  3466 => x"340130de",  3467 => x"0d610032",
     3468 => x"3401ad01",  3469 => x"0d610034",  3470 => x"3162002a",
     3471 => x"34011003",  3472 => x"45a10005",  3473 => x"34011004",
     3474 => x"34020008",  3475 => x"5da1002d",  3476 => x"e0000017",
     3477 => x"298102c8",  3478 => x"35620038",  3479 => x"28210010",
     3480 => x"28230014",  3481 => x"44600005",  3482 => x"40210034",
     3483 => x"31610038",  3484 => x"30400001",  3485 => x"e0000007",
     3486 => x"40210034",  3487 => x"3c210008",  3488 => x"38210001",
     3489 => x"00230008",  3490 => x"31630038",  3491 => x"30410001",
     3492 => x"298102c8",  3493 => x"28220010",  3494 => x"3561003a",
     3495 => x"28420030",  3496 => x"fbffff31",  3497 => x"34020014",
     3498 => x"e0000016",  3499 => x"298102c8",  3500 => x"28220010",
     3501 => x"35610038",  3502 => x"2842001c",  3503 => x"fbffff2a",
     3504 => x"298102c8",  3505 => x"28220010",  3506 => x"3561003c",
     3507 => x"28420018",  3508 => x"fbffff25",  3509 => x"298102c8",
     3510 => x"28220010",  3511 => x"35610040",  3512 => x"28420024",
     3513 => x"fbffff20",  3514 => x"298102c8",  3515 => x"28220010",
     3516 => x"35610044",  3517 => x"28420020",  3518 => x"fbffff1b",
     3519 => x"34020018",  3520 => x"34410030",  3521 => x"31600002",
     3522 => x"31610003",  3523 => x"0d62002e",  3524 => x"2b9d0004",
     3525 => x"2b8b0010",  3526 => x"2b8c000c",  3527 => x"2b8d0008",
     3528 => x"379c0010",  3529 => x"c3a00000",  3530 => x"379cffec",
     3531 => x"5b8b0014",  3532 => x"5b8c0010",  3533 => x"5b8d000c",
     3534 => x"5b8e0008",  3535 => x"5b9d0004",  3536 => x"b8405800",
     3537 => x"b8607000",  3538 => x"34420022",  3539 => x"b8206000",
     3540 => x"b8600800",  3541 => x"34030008",  3542 => x"b8806800",
     3543 => x"f8003dda",  3544 => x"3561002a",  3545 => x"fbffff13",
     3546 => x"0dc10008",  3547 => x"3561002c",  3548 => x"fbffff10",
     3549 => x"b8202800",  3550 => x"34040003",  3551 => x"2d630030",
     3552 => x"2d620032",  3553 => x"2d610034",  3554 => x"44a40007",
     3555 => x"78040001",  3556 => x"b9800800",  3557 => x"34020005",
     3558 => x"34030001",  3559 => x"38844044",  3560 => x"e0000022",
     3561 => x"3c650008",  3562 => x"78040001",  3563 => x"00430008",
     3564 => x"38845960",  3565 => x"b8a32800",  3566 => x"28830000",
     3567 => x"44a30007",  3568 => x"78040001",  3569 => x"b9800800",
     3570 => x"34020005",  3571 => x"34030001",  3572 => x"38844094",
     3573 => x"e0000015",  3574 => x"3c450008",  3575 => x"00230008",
     3576 => x"20a5ffff",  3577 => x"b8a32800",  3578 => x"3802dead",
     3579 => x"44a20007",  3580 => x"78040001",  3581 => x"b9800800",
     3582 => x"34020005",  3583 => x"34030001",  3584 => x"388440cc",
     3585 => x"e0000009",  3586 => x"202500ff",  3587 => x"34010001",
     3588 => x"44a10008",  3589 => x"78040001",  3590 => x"b9800800",
     3591 => x"34020005",  3592 => x"34030001",  3593 => x"38844110",
     3594 => x"fbfff448",  3595 => x"e0000028",  3596 => x"2d610036",
     3597 => x"45a00002",  3598 => x"0da10000",  3599 => x"34021003",
     3600 => x"44220004",  3601 => x"34021004",  3602 => x"5c220021",
     3603 => x"e0000012",  3604 => x"298102c8",  3605 => x"356e0038",
     3606 => x"282d0010",  3607 => x"b9c00800",  3608 => x"fbfffed4",
     3609 => x"202100ff",  3610 => x"0da10048",  3611 => x"b9c00800",
     3612 => x"fbfffed0",  3613 => x"00210008",  3614 => x"31a10050",
     3615 => x"3561003a",  3616 => x"fbfffec1",  3617 => x"298202c8",
     3618 => x"28420010",  3619 => x"5841004c",  3620 => x"e000000f",
     3621 => x"298102c8",  3622 => x"282c0010",  3623 => x"35610038",
     3624 => x"fbfffeb9",  3625 => x"59810058",  3626 => x"3561003c",
     3627 => x"fbfffeb6",  3628 => x"59810054",  3629 => x"35610040",
     3630 => x"fbfffeb3",  3631 => x"59810060",  3632 => x"35610044",
     3633 => x"fbfffeb0",  3634 => x"5981005c",  3635 => x"2b9d0004",
     3636 => x"2b8b0014",  3637 => x"2b8c0010",  3638 => x"2b8d000c",
     3639 => x"2b8e0008",  3640 => x"379c0014",  3641 => x"c3a00000",
     3642 => x"379cfff4",  3643 => x"5b8b000c",  3644 => x"5b8c0008",
     3645 => x"5b9d0004",  3646 => x"2042ffff",  3647 => x"b8205800",
     3648 => x"fbffff1e",  3649 => x"b8206000",  3650 => x"29610024",
     3651 => x"29630070",  3652 => x"29620034",  3653 => x"2827000c",
     3654 => x"b5831800",  3655 => x"b9600800",  3656 => x"356400f8",
     3657 => x"34050000",  3658 => x"34060000",  3659 => x"d8e00000",
     3660 => x"78080001",  3661 => x"390866f4",  3662 => x"4c2c000b",
     3663 => x"29050030",  3664 => x"78040001",  3665 => x"b9600800",
     3666 => x"34020005",  3667 => x"34030001",  3668 => x"38844154",
     3669 => x"3406000c",  3670 => x"fbfff3fc",  3671 => x"3401ffff",
     3672 => x"e000000f",  3673 => x"296600f8",  3674 => x"296700fc",
     3675 => x"29080030",  3676 => x"78040001",  3677 => x"b9600800",
     3678 => x"34020005",  3679 => x"34030001",  3680 => x"38844174",
     3681 => x"b9802800",  3682 => x"fbfff3f0",  3683 => x"2961036c",
     3684 => x"34210001",  3685 => x"5961036c",  3686 => x"34010000",
     3687 => x"2b9d0004",  3688 => x"2b8b000c",  3689 => x"2b8c0008",
     3690 => x"379c000c",  3691 => x"c3a00000",  3692 => x"78020001",
     3693 => x"384266f0",  3694 => x"58410000",  3695 => x"c3a00000",
     3696 => x"379cffe8",  3697 => x"5b8b0018",  3698 => x"5b8c0014",
     3699 => x"5b8d0010",  3700 => x"5b8e000c",  3701 => x"5b8f0008",
     3702 => x"5b9d0004",  3703 => x"282b0014",  3704 => x"b8206800",
     3705 => x"45600014",  3706 => x"780c0001",  3707 => x"398c925c",
     3708 => x"29810000",  3709 => x"34020001",  3710 => x"f8001229",
     3711 => x"34020000",  3712 => x"31a0001c",  3713 => x"b9600800",
     3714 => x"34030110",  3715 => x"296f00f0",  3716 => x"296e00f4",
     3717 => x"296d00f8",  3718 => x"f8003da9",  3719 => x"29810000",
     3720 => x"596f00f0",  3721 => x"596e00f4",  3722 => x"596d00f8",
     3723 => x"34020000",  3724 => x"f800121b",  3725 => x"2b9d0004",
     3726 => x"2b8b0018",  3727 => x"2b8c0014",  3728 => x"2b8d0010",
     3729 => x"2b8e000c",  3730 => x"2b8f0008",  3731 => x"379c0018",
     3732 => x"c3a00000",  3733 => x"379cffec",  3734 => x"5b8b0014",
     3735 => x"5b8c0010",  3736 => x"5b8d000c",  3737 => x"5b8e0008",
     3738 => x"5b9d0004",  3739 => x"b8206800",  3740 => x"282102c8",
     3741 => x"780e0001",  3742 => x"39ce925c",  3743 => x"282c0010",
     3744 => x"29c10000",  3745 => x"34020001",  3746 => x"29ab0014",
     3747 => x"f8001204",  3748 => x"29810000",  3749 => x"34020000",
     3750 => x"34030000",  3751 => x"2826001c",  3752 => x"35640028",
     3753 => x"b9a00800",  3754 => x"3565002c",  3755 => x"d8c00000",
     3756 => x"3402ffff",  3757 => x"5c200039",  3758 => x"29810000",
     3759 => x"34020000",  3760 => x"28230034",  3761 => x"b9a00800",
     3762 => x"d8600000",  3763 => x"34030010",  3764 => x"35a20358",
     3765 => x"b9600800",  3766 => x"f8003eab",  3767 => x"29810000",
     3768 => x"596000a8",  3769 => x"28220018",  3770 => x"34010000",
     3771 => x"d8400000",  3772 => x"34010002",  3773 => x"59610014",
     3774 => x"29810058",  3775 => x"2d820054",  3776 => x"59600088",
     3777 => x"3c210010",  3778 => x"b8220800",  3779 => x"59610018",
     3780 => x"29810060",  3781 => x"2d82005c",  3782 => x"3c210010",
     3783 => x"b8220800",  3784 => x"5961001c",  3785 => x"2981001c",
     3786 => x"2d820018",  3787 => x"3c210010",  3788 => x"b8220800",
     3789 => x"59610020",  3790 => x"29810024",  3791 => x"2d820020",
     3792 => x"3c210010",  3793 => x"b8220800",  3794 => x"78020001",
     3795 => x"59610024",  3796 => x"38424198",  3797 => x"356100c0",
     3798 => x"f8003deb",  3799 => x"29610010",  3800 => x"34020000",
     3801 => x"596000b8",  3802 => x"38210001",  3803 => x"59610010",
     3804 => x"78010001",  3805 => x"382166f0",  3806 => x"28210000",
     3807 => x"596100bc",  3808 => x"78010001",  3809 => x"38217a38",
     3810 => x"58200000",  3811 => x"29c10000",  3812 => x"f80011c3",
     3813 => x"34020000",  3814 => x"b8400800",  3815 => x"2b9d0004",
     3816 => x"2b8b0014",  3817 => x"2b8c0010",  3818 => x"2b8d000c",
     3819 => x"2b8e0008",  3820 => x"379c0014",  3821 => x"c3a00000",
     3822 => x"28460000",  3823 => x"28450004",  3824 => x"28440008",
     3825 => x"28210014",  3826 => x"28420010",  3827 => x"58260030",
     3828 => x"58220040",  3829 => x"34020001",  3830 => x"58250034",
     3831 => x"58240038",  3832 => x"5822003c",  3833 => x"28670000",
     3834 => x"28660004",  3835 => x"28650008",  3836 => x"2864000c",
     3837 => x"28630010",  3838 => x"58270044",  3839 => x"58260048",
     3840 => x"5825004c",  3841 => x"58240050",  3842 => x"58230054",
     3843 => x"78010001",  3844 => x"38217a38",  3845 => x"58220000",
     3846 => x"34010000",  3847 => x"c3a00000",  3848 => x"379cfff8",
     3849 => x"5b8b0008",  3850 => x"5b9d0004",  3851 => x"282500b0",
     3852 => x"282400b4",  3853 => x"282300b8",  3854 => x"282b0014",
     3855 => x"282700a8",  3856 => x"282600ac",  3857 => x"59650060",
     3858 => x"59640064",  3859 => x"282500bc",  3860 => x"282400c0",
     3861 => x"59630068",  3862 => x"282300c4",  3863 => x"282100cc",
     3864 => x"59670058",  3865 => x"59640070",  3866 => x"5961007c",
     3867 => x"34010001",  3868 => x"59610078",  3869 => x"1441001f",
     3870 => x"59630074",  3871 => x"5966005c",  3872 => x"5965006c",
     3873 => x"34030000",  3874 => x"340403e8",  3875 => x"f8003bb9",
     3876 => x"1423001f",  3877 => x"2063ffff",  3878 => x"b4621000",
     3879 => x"f4621800",  3880 => x"00420010",  3881 => x"b4610800",
     3882 => x"3c210010",  3883 => x"b8221000",  3884 => x"34010000",
     3885 => x"59620074",  3886 => x"2b9d0004",  3887 => x"2b8b0008",
     3888 => x"379c0008",  3889 => x"c3a00000",  3890 => x"379cffbc",
     3891 => x"5b8b003c",  3892 => x"5b8c0038",  3893 => x"5b8d0034",
     3894 => x"5b8e0030",  3895 => x"5b8f002c",  3896 => x"5b900028",
     3897 => x"5b910024",  3898 => x"5b920020",  3899 => x"5b93001c",
     3900 => x"5b940018",  3901 => x"5b950014",  3902 => x"5b960010",
     3903 => x"5b97000c",  3904 => x"5b980008",  3905 => x"5b9d0004",
     3906 => x"b8206000",  3907 => x"282102c8",  3908 => x"298b0014",
     3909 => x"282e0010",  3910 => x"78010001",  3911 => x"38217a38",
     3912 => x"28210000",  3913 => x"44200283",  3914 => x"2963003c",
     3915 => x"44600007",  3916 => x"29610050",  3917 => x"44200005",
     3918 => x"29610064",  3919 => x"44200003",  3920 => x"29610078",
     3921 => x"5c200011",  3922 => x"78010001",  3923 => x"38217a3c",
     3924 => x"28220000",  3925 => x"34420001",  3926 => x"58220000",
     3927 => x"34010005",  3928 => x"4c220274",  3929 => x"29640050",
     3930 => x"29650064",  3931 => x"29660078",  3932 => x"78010001",
     3933 => x"78020001",  3934 => x"38425aec",  3935 => x"382141b8",
     3936 => x"f8002258",  3937 => x"e000026b",  3938 => x"29c10000",
     3939 => x"28230038",  3940 => x"44600004",  3941 => x"b9600800",
     3942 => x"34020000",  3943 => x"d8600000",  3944 => x"78010001",
     3945 => x"3821925c",  3946 => x"28210000",  3947 => x"34020001",
     3948 => x"f800113b",  3949 => x"78010001",  3950 => x"38217a3c",
     3951 => x"58200000",  3952 => x"296100b8",  3953 => x"356200fc",
     3954 => x"34210001",  3955 => x"596100b8",  3956 => x"29810028",
     3957 => x"28230000",  3958 => x"b9800800",  3959 => x"d8600000",
     3960 => x"78010001",  3961 => x"38217a38",  3962 => x"58200000",
     3963 => x"29660030",  3964 => x"29670034",  3965 => x"29680038",
     3966 => x"2965006c",  3967 => x"29640074",  3968 => x"29610070",
     3969 => x"c8a62800",  3970 => x"c8882000",  3971 => x"c8270800",
     3972 => x"e0000002",  3973 => x"348403e8",  3974 => x"b8201800",
     3975 => x"3421ffff",  3976 => x"4804fffd",  3977 => x"b8a00800",
     3978 => x"78050001",  3979 => x"38a55958",  3980 => x"28a20000",
     3981 => x"e0000002",  3982 => x"b4621800",  3983 => x"b8205000",
     3984 => x"3421ffff",  3985 => x"4803fffd",  3986 => x"29610044",
     3987 => x"29650058",  3988 => x"29620060",  3989 => x"2969005c",
     3990 => x"c8a12800",  3991 => x"2961004c",  3992 => x"c8410800",
     3993 => x"29620048",  3994 => x"c9224800",  3995 => x"e0000002",
     3996 => x"342103e8",  3997 => x"b9201000",  3998 => x"3529ffff",
     3999 => x"4801fffd",  4000 => x"78090001",  4001 => x"39295958",
     4002 => x"292d0000",  4003 => x"e0000002",  4004 => x"b44d1000",
     4005 => x"b8a04800",  4006 => x"34a5ffff",  4007 => x"4802fffd",
     4008 => x"c8810800",  4009 => x"c9495000",  4010 => x"c8622000",
     4011 => x"e0000002",  4012 => x"342103e8",  4013 => x"b8801000",
     4014 => x"3484ffff",  4015 => x"4801fffd",  4016 => x"78040001",
     4017 => x"38845958",  4018 => x"b9401800",  4019 => x"28850000",
     4020 => x"e0000002",  4021 => x"b4451000",  4022 => x"b8602000",
     4023 => x"3463ffff",  4024 => x"4802fffd",  4025 => x"59610094",
     4026 => x"78010001",  4027 => x"382174c4",  4028 => x"59620090",
     4029 => x"28210000",  4030 => x"29820018",  4031 => x"5964008c",
     4032 => x"b8220800",  4033 => x"00210010",  4034 => x"2021000f",
     4035 => x"44200032",  4036 => x"780d0001",  4037 => x"39ad41e8",
     4038 => x"78050001",  4039 => x"b9800800",  4040 => x"34020004",
     4041 => x"34030002",  4042 => x"b9a02000",  4043 => x"38a541f8",
     4044 => x"fbfff286",  4045 => x"29660044",  4046 => x"29670048",
     4047 => x"2968004c",  4048 => x"78050001",  4049 => x"b9800800",
     4050 => x"34020004",  4051 => x"34030002",  4052 => x"b9a02000",
     4053 => x"38a54204",  4054 => x"fbfff27c",  4055 => x"29660058",
     4056 => x"2967005c",  4057 => x"29680060",  4058 => x"78050001",
     4059 => x"b9800800",  4060 => x"34020004",  4061 => x"34030002",
     4062 => x"b9a02000",  4063 => x"38a54210",  4064 => x"fbfff272",
     4065 => x"2966006c",  4066 => x"29670070",  4067 => x"29680074",
     4068 => x"78050001",  4069 => x"b9800800",  4070 => x"34020004",
     4071 => x"34030002",  4072 => x"b9a02000",  4073 => x"38a5421c",
     4074 => x"fbfff268",  4075 => x"2966008c",  4076 => x"29670090",
     4077 => x"29680094",  4078 => x"78050001",  4079 => x"b9800800",
     4080 => x"34020004",  4081 => x"34030002",  4082 => x"b9a02000",
     4083 => x"38a54228",  4084 => x"fbfff25e",  4085 => x"2962008c",
     4086 => x"78050001",  4087 => x"38a55964",  4088 => x"28a40000",
     4089 => x"1441001f",  4090 => x"340300e8",  4091 => x"f8003ae1",
     4092 => x"b8406800",  4093 => x"29620090",  4094 => x"b8207800",
     4095 => x"34030000",  4096 => x"1441001f",  4097 => x"340403e8",
     4098 => x"f8003ada",  4099 => x"29660094",  4100 => x"b5a21800",
     4101 => x"f5a36800",  4102 => x"14c2001f",  4103 => x"b5e10800",
     4104 => x"b4663000",  4105 => x"b5a10800",  4106 => x"f4661800",
     4107 => x"b4220800",  4108 => x"29650018",  4109 => x"29620020",
     4110 => x"2964001c",  4111 => x"b4610800",  4112 => x"29630024",
     4113 => x"b4a21000",  4114 => x"b4441000",  4115 => x"b4431000",
     4116 => x"1444001f",  4117 => x"297600a0",  4118 => x"297400a4",
     4119 => x"596100a0",  4120 => x"596600a4",  4121 => x"48810004",
     4122 => x"5c810005",  4123 => x"54460002",  4124 => x"e0000003",
     4125 => x"596400a0",  4126 => x"596200a4",  4127 => x"296600a4",
     4128 => x"296100a0",  4129 => x"1477001f",  4130 => x"c8c21000",
     4131 => x"f4463000",  4132 => x"c8240800",  4133 => x"c8260800",
     4134 => x"b4652000",  4135 => x"14a6001f",  4136 => x"f4641800",
     4137 => x"b6e6b800",  4138 => x"b477b800",  4139 => x"004d0001",
     4140 => x"3c23001f",  4141 => x"00250001",  4142 => x"b86d6800",
     4143 => x"b48d6800",  4144 => x"f48d2000",  4145 => x"b6e5b800",
     4146 => x"b497b800",  4147 => x"29640028",  4148 => x"1483001f",
     4149 => x"f8003aa7",  4150 => x"14350008",  4151 => x"1421001f",
     4152 => x"b5b5a800",  4153 => x"f5b56800",  4154 => x"b6e10800",
     4155 => x"b5a1b800",  4156 => x"29620030",  4157 => x"29610044",
     4158 => x"29720038",  4159 => x"29630034",  4160 => x"c8411000",
     4161 => x"2961004c",  4162 => x"ca419000",  4163 => x"29610048",
     4164 => x"c8611800",  4165 => x"e0000002",  4166 => x"365203e8",
     4167 => x"b8606800",  4168 => x"3463ffff",  4169 => x"4812fffd",
     4170 => x"78090001",  4171 => x"39295958",  4172 => x"29210000",
     4173 => x"e0000002",  4174 => x"b5a16800",  4175 => x"b8408800",
     4176 => x"3442ffff",  4177 => x"480dfffd",  4178 => x"378f0040",
     4179 => x"340203e8",  4180 => x"b9e00800",  4181 => x"5b970040",
     4182 => x"5b950044",  4183 => x"fbfff62f",  4184 => x"78030001",
     4185 => x"38635958",  4186 => x"28620000",  4187 => x"b8208000",
     4188 => x"b9e00800",  4189 => x"fbfff629",  4190 => x"2b820044",
     4191 => x"b42d6800",  4192 => x"b6509000",  4193 => x"b6221000",
     4194 => x"340103e7",  4195 => x"e0000002",  4196 => x"3652fc18",
     4197 => x"b9a08800",  4198 => x"ba408000",  4199 => x"35ad0001",
     4200 => x"4a41fffc",  4201 => x"78040001",  4202 => x"78050001",
     4203 => x"38845968",  4204 => x"38a5596c",  4205 => x"b8400800",
     4206 => x"28830000",  4207 => x"28a20000",  4208 => x"e0000002",
     4209 => x"b6228800",  4210 => x"b8207800",  4211 => x"ba206800",
     4212 => x"34210001",  4213 => x"4a23fffc",  4214 => x"2961002c",
     4215 => x"340203e8",  4216 => x"b9e0c000",  4217 => x"342103e7",
     4218 => x"f8003a89",  4219 => x"b8209800",  4220 => x"4c110008",
     4221 => x"ba200800",  4222 => x"ba601000",  4223 => x"f8003ab1",
     4224 => x"4420000a",  4225 => x"083003e8",  4226 => x"ca216800",
     4227 => x"b6128000",  4228 => x"4da00006",  4229 => x"78090001",
     4230 => x"39295958",  4231 => x"29210000",  4232 => x"35efffff",
     4233 => x"b5a16800",  4234 => x"3401ffff",  4235 => x"5de10007",
     4236 => x"4c0d0006",  4237 => x"78020001",  4238 => x"3842596c",
     4239 => x"28410000",  4240 => x"340f0000",  4241 => x"b5a16800",
     4242 => x"4da00007",  4243 => x"c8130800",  4244 => x"482d0005",
     4245 => x"5de00004",  4246 => x"b5b36800",  4247 => x"0a73fc18",
     4248 => x"b6138000",  4249 => x"78050001",  4250 => x"38a55964",
     4251 => x"28a40000",  4252 => x"1701001f",  4253 => x"bb001000",
     4254 => x"340300e8",  4255 => x"f8003a3d",  4256 => x"b820c000",
     4257 => x"1621001f",  4258 => x"b8409800",  4259 => x"34030000",
     4260 => x"340403e8",  4261 => x"ba201000",  4262 => x"f8003a36",
     4263 => x"b6621800",  4264 => x"f6639800",  4265 => x"1642001f",
     4266 => x"b7010800",  4267 => x"b4729000",  4268 => x"b6610800",
     4269 => x"b4220800",  4270 => x"f4721800",  4271 => x"78020001",
     4272 => x"384266f0",  4273 => x"b4611800",  4274 => x"28410000",
     4275 => x"596300e8",  4276 => x"34020000",  4277 => x"596100bc",
     4278 => x"29c10000",  4279 => x"597200ec",  4280 => x"597700b0",
     4281 => x"28230004",  4282 => x"597500b4",  4283 => x"b9800800",
     4284 => x"d8600000",  4285 => x"34020001",  4286 => x"4422000c",
     4287 => x"78040001",  4288 => x"b9800800",  4289 => x"34020004",
     4290 => x"34030001",  4291 => x"38844234",  4292 => x"fbfff18e",
     4293 => x"29c10000",  4294 => x"34020000",  4295 => x"28230034",
     4296 => x"b9800800",  4297 => x"d8600000",  4298 => x"29c10000",
     4299 => x"28210010",  4300 => x"d8200000",  4301 => x"5c200007",
     4302 => x"29630010",  4303 => x"3402fffd",  4304 => x"a0621000",
     4305 => x"59620010",  4306 => x"5de10009",  4307 => x"e000000a",
     4308 => x"78040001",  4309 => x"b9800800",  4310 => x"34020004",
     4311 => x"34030001",  4312 => x"38844258",  4313 => x"fbfff179",
     4314 => x"e00000e7",  4315 => x"34010002",  4316 => x"e0000003",
     4317 => x"45af0003",  4318 => x"34010001",  4319 => x"59610014",
     4320 => x"78040001",  4321 => x"b9800800",  4322 => x"34020004",
     4323 => x"b9e02800",  4324 => x"b9a03000",  4325 => x"34030002",
     4326 => x"38844264",  4327 => x"ba003800",  4328 => x"fbfff16a",
     4329 => x"29620014",  4330 => x"78010001",  4331 => x"38215be4",
     4332 => x"3c420002",  4333 => x"78060001",  4334 => x"b4220800",
     4335 => x"28250000",  4336 => x"29610010",  4337 => x"38c65950",
     4338 => x"20210002",  4339 => x"44200003",  4340 => x"78060001",
     4341 => x"38c641a8",  4342 => x"78040001",  4343 => x"b9800800",
     4344 => x"34020004",  4345 => x"34030001",  4346 => x"38844284",
     4347 => x"fbfff157",  4348 => x"29620014",  4349 => x"78010001",
     4350 => x"38215be4",  4351 => x"3c420002",  4352 => x"b4221000",
     4353 => x"28420000",  4354 => x"356100c0",  4355 => x"f8003bbe",
     4356 => x"29620014",  4357 => x"34010004",  4358 => x"3442ffff",
     4359 => x"54410083",  4360 => x"78010001",  4361 => x"3c420002",
     4362 => x"38215bd0",  4363 => x"b4220800",  4364 => x"28210000",
     4365 => x"c0200000",  4366 => x"29c10000",  4367 => x"b9e01000",
     4368 => x"34030000",  4369 => x"28240014",  4370 => x"15e1001f",
     4371 => x"e0000006",  4372 => x"29c10000",  4373 => x"34020000",
     4374 => x"b9a01800",  4375 => x"28240014",  4376 => x"34010000",
     4377 => x"d8800000",  4378 => x"29610010",  4379 => x"38210002",
     4380 => x"59610010",  4381 => x"e0000057",  4382 => x"296500a8",
     4383 => x"78040001",  4384 => x"b9800800",  4385 => x"34020004",
     4386 => x"34030002",  4387 => x"3884429c",  4388 => x"b9a03000",
     4389 => x"ba003800",  4390 => x"fbfff12c",  4391 => x"29c20000",
     4392 => x"296100a8",  4393 => x"28420018",  4394 => x"b6010800",
     4395 => x"596100a8",  4396 => x"d8400000",  4397 => x"29610010",
     4398 => x"38210002",  4399 => x"59610010",  4400 => x"34010005",
     4401 => x"59610014",  4402 => x"e0000058",  4403 => x"78090001",
     4404 => x"39295964",  4405 => x"29240000",  4406 => x"15e1001f",
     4407 => x"b9e01000",  4408 => x"340300e8",  4409 => x"f80039a3",
     4410 => x"b6027800",  4411 => x"1611001f",  4412 => x"f60f8000",
     4413 => x"b6210800",  4414 => x"b6018000",  4415 => x"15a1001f",
     4416 => x"34030000",  4417 => x"b9a01000",  4418 => x"340403e8",
     4419 => x"f8003999",  4420 => x"b5e21800",  4421 => x"f5e37800",
     4422 => x"b6010800",  4423 => x"b5e10800",  4424 => x"c8031000",
     4425 => x"48010002",  4426 => x"b8601000",  4427 => x"3401003b",
     4428 => x"4841000d",  4429 => x"29c10000",  4430 => x"34020001",
     4431 => x"28230034",  4432 => x"b9800800",  4433 => x"d8600000",
     4434 => x"296100b0",  4435 => x"59610080",  4436 => x"296100b4",
     4437 => x"59610084",  4438 => x"34010004",  4439 => x"59610014",
     4440 => x"e0000004",  4441 => x"29610088",  4442 => x"34210001",
     4443 => x"59610088",  4444 => x"29620088",  4445 => x"34010009",
     4446 => x"4c22002c",  4447 => x"59600088",  4448 => x"e0000014",
     4449 => x"296300b4",  4450 => x"29610084",  4451 => x"296400b0",
     4452 => x"29620080",  4453 => x"c8610800",  4454 => x"f4231800",
     4455 => x"596100e4",  4456 => x"78010001",  4457 => x"382166f0",
     4458 => x"c8821000",  4459 => x"28210000",  4460 => x"c8431000",
     4461 => x"596200e0",  4462 => x"4420001c",  4463 => x"1601001f",
     4464 => x"34030078",  4465 => x"98301000",  4466 => x"c8411000",
     4467 => x"4c620003",  4468 => x"34010003",  4469 => x"e3ffffbc",
     4470 => x"0021001e",  4471 => x"29c20000",  4472 => x"b4308000",
     4473 => x"296100a8",  4474 => x"16100002",  4475 => x"28420018",
     4476 => x"b6010800",  4477 => x"596100a8",  4478 => x"d8400000",
     4479 => x"296500a8",  4480 => x"78040001",  4481 => x"b9800800",
     4482 => x"34020006",  4483 => x"34030001",  4484 => x"388442b8",
     4485 => x"fbfff0cd",  4486 => x"296100b0",  4487 => x"59610080",
     4488 => x"296100b4",  4489 => x"59610084",  4490 => x"29620014",
     4491 => x"34010004",  4492 => x"44410004",  4493 => x"296100f0",
     4494 => x"34210001",  4495 => x"596100f0",  4496 => x"296400e8",
     4497 => x"296300ec",  4498 => x"1481001f",  4499 => x"98611800",
     4500 => x"c8611000",  4501 => x"98812000",  4502 => x"f4431800",
     4503 => x"c8810800",  4504 => x"c8230800",  4505 => x"48200005",
     4506 => x"5c200007",  4507 => x"340101f4",  4508 => x"54410002",
     4509 => x"e0000004",  4510 => x"296100f4",  4511 => x"34210001",
     4512 => x"596100f4",  4513 => x"296500a4",  4514 => x"296400a0",
     4515 => x"ca851800",  4516 => x"f4740800",  4517 => x"cac41000",
     4518 => x"c8411000",  4519 => x"48020007",  4520 => x"34010001",
     4521 => x"48400013",  4522 => x"5c400011",  4523 => x"340203e8",
     4524 => x"54620010",  4525 => x"e000000e",  4526 => x"c8140800",
     4527 => x"7c220000",  4528 => x"c8161800",  4529 => x"c8621800",
     4530 => x"c8251000",  4531 => x"f4410800",  4532 => x"c8641800",
     4533 => x"c8611800",  4534 => x"34010001",  4535 => x"48600005",
     4536 => x"5c600003",  4537 => x"340303e8",  4538 => x"54430002",
     4539 => x"34010000",  4540 => x"202100ff",  4541 => x"44200004",
     4542 => x"296100f8",  4543 => x"34210001",  4544 => x"596100f8",
     4545 => x"78010001",  4546 => x"3821925c",  4547 => x"28210000",
     4548 => x"34020000",  4549 => x"f8000ee2",  4550 => x"29c10000",
     4551 => x"28230038",  4552 => x"44600004",  4553 => x"b9600800",
     4554 => x"34020001",  4555 => x"d8600000",  4556 => x"34010000",
     4557 => x"2b9d0004",  4558 => x"2b8b003c",  4559 => x"2b8c0038",
     4560 => x"2b8d0034",  4561 => x"2b8e0030",  4562 => x"2b8f002c",
     4563 => x"2b900028",  4564 => x"2b910024",  4565 => x"2b920020",
     4566 => x"2b93001c",  4567 => x"2b940018",  4568 => x"2b950014",
     4569 => x"2b960010",  4570 => x"2b97000c",  4571 => x"2b980008",
     4572 => x"379c0044",  4573 => x"c3a00000",  4574 => x"379cffe8",
     4575 => x"5b8b0018",  4576 => x"5b8c0014",  4577 => x"5b8d0010",
     4578 => x"5b8e000c",  4579 => x"5b8f0008",  4580 => x"5b9d0004",
     4581 => x"b8407800",  4582 => x"28220020",  4583 => x"b8205800",
     4584 => x"b8607000",  4585 => x"284d0008",  4586 => x"28220024",
     4587 => x"282c02c8",  4588 => x"28440000",  4589 => x"d8800000",
     4590 => x"48010058",  4591 => x"29610020",  4592 => x"34030008",
     4593 => x"2824000c",  4594 => x"4161004c",  4595 => x"30810004",
     4596 => x"4161004d",  4597 => x"30810005",  4598 => x"4161004e",
     4599 => x"30810006",  4600 => x"3401ffff",  4601 => x"30810007",
     4602 => x"3401fffe",  4603 => x"30810008",  4604 => x"4161004f",
     4605 => x"30810009",  4606 => x"41610050",  4607 => x"3081000a",
     4608 => x"41610051",  4609 => x"3081000b",  4610 => x"29610020",
     4611 => x"2824000c",  4612 => x"b9800800",  4613 => x"34820004",
     4614 => x"f80039ab",  4615 => x"29610020",  4616 => x"35620374",
     4617 => x"28210000",  4618 => x"3180000a",  4619 => x"c8410800",
     4620 => x"14210002",  4621 => x"0821d775",  4622 => x"0d810008",
     4623 => x"41a10042",  4624 => x"3181000b",  4625 => x"34010014",
     4626 => x"3181000c",  4627 => x"41a10043",  4628 => x"3181000d",
     4629 => x"34010002",  4630 => x"3181000e",  4631 => x"78010001",
     4632 => x"382166bc",  4633 => x"28240000",  4634 => x"4480000f",
     4635 => x"b9600800",  4636 => x"b9e01000",  4637 => x"b9c01800",
     4638 => x"d8800000",  4639 => x"4420000a",  4640 => x"78040001",
     4641 => x"78050001",  4642 => x"b9600800",  4643 => x"34020002",
     4644 => x"34030001",  4645 => x"38844324",  4646 => x"38a55bfc",
     4647 => x"fbfff02b",  4648 => x"e000001e",  4649 => x"29610020",
     4650 => x"78040001",  4651 => x"34020003",  4652 => x"2825000c",
     4653 => x"34030001",  4654 => x"b9600800",  4655 => x"40a5000e",
     4656 => x"38844340",  4657 => x"fbfff021",  4658 => x"29610020",
     4659 => x"78040001",  4660 => x"34020003",  4661 => x"2825000c",
     4662 => x"34030001",  4663 => x"b9600800",  4664 => x"40a5000f",
     4665 => x"38844354",  4666 => x"fbfff018",  4667 => x"2962003c",
     4668 => x"b9600800",  4669 => x"f8000634",  4670 => x"4162001d",
     4671 => x"34010001",  4672 => x"44410003",  4673 => x"34010004",
     4674 => x"e0000002",  4675 => x"34010006",  4676 => x"59610004",
     4677 => x"e0000003",  4678 => x"340103e8",  4679 => x"59610008",
     4680 => x"34010000",  4681 => x"2b9d0004",  4682 => x"2b8b0018",
     4683 => x"2b8c0014",  4684 => x"2b8d0010",  4685 => x"2b8e000c",
     4686 => x"2b8f0008",  4687 => x"379c0018",  4688 => x"c3a00000",
     4689 => x"379cfff4",  4690 => x"5b8b000c",  4691 => x"5b8c0008",
     4692 => x"5b9d0004",  4693 => x"2822000c",  4694 => x"b8205800",
     4695 => x"44400006",  4696 => x"28220028",  4697 => x"28430018",
     4698 => x"34020fa0",  4699 => x"d8600000",  4700 => x"596102dc",
     4701 => x"296102dc",  4702 => x"44200009",  4703 => x"29610028",
     4704 => x"34020000",  4705 => x"28230018",  4706 => x"b9600800",
     4707 => x"d8600000",  4708 => x"296202dc",  4709 => x"c8220800",
     4710 => x"4c200014",  4711 => x"296c02dc",  4712 => x"34010000",
     4713 => x"4580000a",  4714 => x"29610028",  4715 => x"34020000",
     4716 => x"28230018",  4717 => x"b9600800",  4718 => x"d8600000",
     4719 => x"c9810800",  4720 => x"a4201000",  4721 => x"1442001f",
     4722 => x"a0220800",  4723 => x"59610008",  4724 => x"34010000",
     4725 => x"2b9d0004",  4726 => x"2b8b000c",  4727 => x"2b8c0008",
     4728 => x"379c000c",  4729 => x"c3a00000",  4730 => x"b9600800",
     4731 => x"34020004",  4732 => x"f8000a67",  4733 => x"34010001",
     4734 => x"59610004",  4735 => x"e3fffff5",  4736 => x"340203e8",
     4737 => x"58220008",  4738 => x"34010000",  4739 => x"c3a00000",
     4740 => x"379cfff0",  4741 => x"5b8b0010",  4742 => x"5b8c000c",
     4743 => x"5b8d0008",  4744 => x"5b9d0004",  4745 => x"78040001",
     4746 => x"388466bc",  4747 => x"2884000c",  4748 => x"b8205800",
     4749 => x"b8406800",  4750 => x"b8606000",  4751 => x"44800003",
     4752 => x"d8800000",  4753 => x"5c20001f",  4754 => x"2961000c",
     4755 => x"4420000b",  4756 => x"296102c8",  4757 => x"29630028",
     4758 => x"4022000c",  4759 => x"1021000b",  4760 => x"28630018",
     4761 => x"bc411000",  4762 => x"b9600800",  4763 => x"084203e8",
     4764 => x"d8600000",  4765 => x"596102d4",  4766 => x"4580000f",
     4767 => x"4161030d",  4768 => x"44200008",  4769 => x"3402000b",
     4770 => x"5c22000b",  4771 => x"b9600800",  4772 => x"b9a01000",
     4773 => x"b9801800",  4774 => x"f8000352",  4775 => x"e0000005",
     4776 => x"b9600800",  4777 => x"b9a01000",  4778 => x"b9801800",
     4779 => x"f8000370",  4780 => x"5c200004",  4781 => x"b9600800",
     4782 => x"f800027e",  4783 => x"44200003",  4784 => x"34010002",
     4785 => x"59610004",  4786 => x"29620004",  4787 => x"29610000",
     4788 => x"44410002",  4789 => x"596002d4",  4790 => x"296c02d4",
     4791 => x"34010000",  4792 => x"4580000a",  4793 => x"29610028",
     4794 => x"34020000",  4795 => x"28230018",  4796 => x"b9600800",
     4797 => x"d8600000",  4798 => x"c9810800",  4799 => x"a4201000",
     4800 => x"1442001f",  4801 => x"a0220800",  4802 => x"59610008",
     4803 => x"34010000",  4804 => x"2b9d0004",  4805 => x"2b8b0010",
     4806 => x"2b8c000c",  4807 => x"2b8d0008",  4808 => x"379c0010",
     4809 => x"c3a00000",  4810 => x"34010000",  4811 => x"c3a00000",
     4812 => x"379cffec",  4813 => x"5b8b0014",  4814 => x"5b8c0010",
     4815 => x"5b8d000c",  4816 => x"5b8e0008",  4817 => x"5b9d0004",
     4818 => x"344b00b2",  4819 => x"3d6b0002",  4820 => x"b8407000",
     4821 => x"b42b5800",  4822 => x"29620004",  4823 => x"b8206000",
     4824 => x"340d0000",  4825 => x"44400008",  4826 => x"28220028",
     4827 => x"28430018",  4828 => x"34020000",  4829 => x"d8600000",
     4830 => x"29620004",  4831 => x"c8220800",  4832 => x"4c200009",
     4833 => x"b9a00800",  4834 => x"2b9d0004",  4835 => x"2b8b0014",
     4836 => x"2b8c0010",  4837 => x"2b8d000c",  4838 => x"2b8e0008",
     4839 => x"379c0014",  4840 => x"c3a00000",  4841 => x"b9800800",
     4842 => x"b9c01000",  4843 => x"f80009f8",  4844 => x"340d0001",
     4845 => x"59600004",  4846 => x"e3fffff3",  4847 => x"379cffec",
     4848 => x"5b8b0014",  4849 => x"5b8c0010",  4850 => x"5b8d000c",
     4851 => x"5b8e0008",  4852 => x"5b9d0004",  4853 => x"b8407000",
     4854 => x"2822000c",  4855 => x"b8205800",  4856 => x"b8606800",
     4857 => x"340c0000",  4858 => x"44400014",  4859 => x"282302c8",
     4860 => x"34020001",  4861 => x"1063000d",  4862 => x"f80009f4",
     4863 => x"296302c8",  4864 => x"b9600800",  4865 => x"34020003",
     4866 => x"1063000b",  4867 => x"f80009ef",  4868 => x"29630344",
     4869 => x"34020001",  4870 => x"34010000",  4871 => x"5c620002",
     4872 => x"29610340",  4873 => x"0d61007e",  4874 => x"b9600800",
     4875 => x"f80005d9",  4876 => x"b8206000",  4877 => x"48010047",
     4878 => x"b9600800",  4879 => x"34020001",  4880 => x"fbffffbc",
     4881 => x"44200010",  4882 => x"296302c8",  4883 => x"b9600800",
     4884 => x"34020001",  4885 => x"1063000d",  4886 => x"f80009dc",
     4887 => x"29630344",  4888 => x"34020001",  4889 => x"34010000",
     4890 => x"5c620002",  4891 => x"29610340",  4892 => x"0d61007e",
     4893 => x"b9600800",  4894 => x"f8000613",  4895 => x"48010046",
     4896 => x"340c0000",  4897 => x"b9600800",  4898 => x"34020003",
     4899 => x"fbffffa9",  4900 => x"44200010",  4901 => x"29630344",
     4902 => x"34020001",  4903 => x"34010000",  4904 => x"5c620002",
     4905 => x"29610340",  4906 => x"0d61007e",  4907 => x"b9600800",
     4908 => x"f80005b8",  4909 => x"48010038",  4910 => x"296302c8",
     4911 => x"b9600800",  4912 => x"34020003",  4913 => x"1063000b",
     4914 => x"340c0000",  4915 => x"f80009bf",  4916 => x"45a00020",
     4917 => x"78010001",  4918 => x"382166bc",  4919 => x"28250010",
     4920 => x"4164030d",  4921 => x"44a00007",  4922 => x"b9600800",
     4923 => x"b9c01000",  4924 => x"b9a01800",  4925 => x"d8a00000",
     4926 => x"b8202000",  4927 => x"48010042",  4928 => x"34010001",
     4929 => x"44810010",  4930 => x"3401000b",  4931 => x"44810003",
     4932 => x"5c800010",  4933 => x"e0000006",  4934 => x"b9600800",
     4935 => x"b9c01000",  4936 => x"b9a01800",  4937 => x"f80002af",
     4938 => x"e0000005",  4939 => x"b9600800",  4940 => x"b9c01000",
     4941 => x"b9a01800",  4942 => x"f80002cd",  4943 => x"b8206000",
     4944 => x"e0000004",  4945 => x"b9600800",  4946 => x"356200e4",
     4947 => x"f800066a",  4948 => x"45800006",  4949 => x"34010001",
     4950 => x"4581000f",  4951 => x"3401ffff",  4952 => x"5d81000e",
     4953 => x"e0000029",  4954 => x"29610020",  4955 => x"2821000c",
     4956 => x"4022000e",  4957 => x"340100ff",  4958 => x"44410004",
     4959 => x"4162001d",  4960 => x"34010002",  4961 => x"5c410005",
     4962 => x"34010004",  4963 => x"59610004",  4964 => x"e0000002",
     4965 => x"340c0000",  4966 => x"296e02d8",  4967 => x"340d0000",
     4968 => x"45c0000a",  4969 => x"29610028",  4970 => x"34020000",
     4971 => x"28230018",  4972 => x"b9600800",  4973 => x"d8600000",
     4974 => x"c9c16800",  4975 => x"a5a00800",  4976 => x"1421001f",
     4977 => x"a1a16800",  4978 => x"296e02d0",  4979 => x"34010000",
     4980 => x"45c0000a",  4981 => x"29610028",  4982 => x"34020000",
     4983 => x"28230018",  4984 => x"b9600800",  4985 => x"d8600000",
     4986 => x"c9c10800",  4987 => x"a4201000",  4988 => x"1442001f",
     4989 => x"a0220800",  4990 => x"4da10007",  4991 => x"b9a00800",
     4992 => x"e0000005",  4993 => x"b8206000",  4994 => x"34010002",
     4995 => x"59610004",  4996 => x"340101f4",  4997 => x"59610008",
     4998 => x"b9800800",  4999 => x"2b9d0004",  5000 => x"2b8b0014",
     5001 => x"2b8c0010",  5002 => x"2b8d000c",  5003 => x"2b8e0008",
     5004 => x"379c0014",  5005 => x"c3a00000",  5006 => x"379cfff0",
     5007 => x"5b8b000c",  5008 => x"5b8c0008",  5009 => x"5b9d0004",
     5010 => x"b8406000",  5011 => x"2822000c",  5012 => x"b8205800",
     5013 => x"4440000c",  5014 => x"282202c8",  5015 => x"28250028",
     5016 => x"4044000c",  5017 => x"1042000b",  5018 => x"bc821000",
     5019 => x"28a40018",  5020 => x"084203e8",  5021 => x"5b830010",
     5022 => x"d8800000",  5023 => x"2b830010",  5024 => x"596102d4",
     5025 => x"4460000d",  5026 => x"4161030d",  5027 => x"44200007",
     5028 => x"3402000b",  5029 => x"5c220009",  5030 => x"b9600800",
     5031 => x"b9801000",  5032 => x"f8000250",  5033 => x"e0000004",
     5034 => x"b9600800",  5035 => x"b9801000",  5036 => x"f800026f",
     5037 => x"5c200004",  5038 => x"b9600800",  5039 => x"f800017d",
     5040 => x"44200003",  5041 => x"34010002",  5042 => x"59610004",
     5043 => x"29620004",  5044 => x"29610000",  5045 => x"44410002",
     5046 => x"596002d4",  5047 => x"340103e8",  5048 => x"59610008",
     5049 => x"34010000",  5050 => x"2b9d0004",  5051 => x"2b8b000c",
     5052 => x"2b8c0008",  5053 => x"379c0010",  5054 => x"c3a00000",
     5055 => x"379cfff8",  5056 => x"5b8b0008",  5057 => x"5b9d0004",
     5058 => x"b8205800",  5059 => x"4460000d",  5060 => x"4024030d",
     5061 => x"44800007",  5062 => x"34050008",  5063 => x"44850007",
     5064 => x"3405000b",  5065 => x"5c850007",  5066 => x"f8000198",
     5067 => x"e0000004",  5068 => x"f80001b1",  5069 => x"e0000002",
     5070 => x"f80001e9",  5071 => x"5c200004",  5072 => x"b9600800",
     5073 => x"f800015b",  5074 => x"44200003",  5075 => x"34010002",
     5076 => x"59610004",  5077 => x"340103e8",  5078 => x"59610008",
     5079 => x"34010000",  5080 => x"2b9d0004",  5081 => x"2b8b0008",
     5082 => x"379c0008",  5083 => x"c3a00000",  5084 => x"379cffd4",
     5085 => x"5b8b0014",  5086 => x"5b8c0010",  5087 => x"5b8d000c",
     5088 => x"5b8e0008",  5089 => x"5b9d0004",  5090 => x"b8205800",
     5091 => x"2821000c",  5092 => x"b8407000",  5093 => x"b8606800",
     5094 => x"44200023",  5095 => x"34020000",  5096 => x"34030014",
     5097 => x"35610080",  5098 => x"f8003845",  5099 => x"b9600800",
     5100 => x"f80006da",  5101 => x"78010001",  5102 => x"382166bc",
     5103 => x"28240014",  5104 => x"44800007",  5105 => x"b9600800",
     5106 => x"b9c01000",  5107 => x"b9a01800",  5108 => x"d8800000",
     5109 => x"b8206000",  5110 => x"5c20005f",  5111 => x"4161001c",
     5112 => x"29630028",  5113 => x"202100fd",  5114 => x"3161001c",
     5115 => x"296102c8",  5116 => x"28630018",  5117 => x"4022000c",
     5118 => x"1021000b",  5119 => x"bc411000",  5120 => x"b9600800",
     5121 => x"084203e8",  5122 => x"d8600000",  5123 => x"296302c8",
     5124 => x"596102d4",  5125 => x"34020000",  5126 => x"1063000a",
     5127 => x"b9600800",  5128 => x"f80008ea",  5129 => x"45a00049",
     5130 => x"4161030d",  5131 => x"34020008",  5132 => x"44220012",
     5133 => x"54220003",  5134 => x"5c200044",  5135 => x"e000000a",
     5136 => x"34020009",  5137 => x"44220014",  5138 => x"3402000b",
     5139 => x"5c22003f",  5140 => x"b9600800",  5141 => x"b9c01000",
     5142 => x"b9a01800",  5143 => x"f800014b",  5144 => x"e000000a",
     5145 => x"b9600800",  5146 => x"b9c01000",  5147 => x"b9a01800",
     5148 => x"f8000161",  5149 => x"e0000005",  5150 => x"b9600800",
     5151 => x"b9c01000",  5152 => x"b9a01800",  5153 => x"f8000196",
     5154 => x"b8206000",  5155 => x"5c200032",  5156 => x"e000002e",
     5157 => x"34010035",  5158 => x"340c0001",  5159 => x"4c2d002e",
     5160 => x"378c0018",  5161 => x"b9c00800",  5162 => x"b9801000",
     5163 => x"f80004a2",  5164 => x"296102c8",  5165 => x"37820024",
     5166 => x"34030008",  5167 => x"f8003761",  5168 => x"5c20001c",
     5169 => x"2d6202f2",  5170 => x"2d61032a",  5171 => x"5c410019",
     5172 => x"296102c8",  5173 => x"2c220008",  5174 => x"2f81002c",
     5175 => x"5c410015",  5176 => x"4161001c",  5177 => x"20210001",
     5178 => x"44200012",  5179 => x"b9801000",  5180 => x"356100bc",
     5181 => x"f8000619",  5182 => x"78010001",  5183 => x"382166bc",
     5184 => x"28220018",  5185 => x"44400006",  5186 => x"b9600800",
     5187 => x"d8400000",  5188 => x"b8206000",  5189 => x"5c200010",
     5190 => x"e0000003",  5191 => x"b9600800",  5192 => x"f80006d7",
     5193 => x"4161032d",  5194 => x"316102ee",  5195 => x"e0000007",
     5196 => x"78040001",  5197 => x"b9600800",  5198 => x"34020005",
     5199 => x"34030002",  5200 => x"3884436c",  5201 => x"fbffee01",
     5202 => x"b9600800",  5203 => x"f80000d9",  5204 => x"b8206000",
     5205 => x"296102cc",  5206 => x"44200009",  5207 => x"29610028",
     5208 => x"34020000",  5209 => x"28230018",  5210 => x"b9600800",
     5211 => x"d8600000",  5212 => x"296202cc",  5213 => x"c8220800",
     5214 => x"4c200033",  5215 => x"3401ffff",  5216 => x"45810005",
     5217 => x"7d810001",  5218 => x"c8010800",  5219 => x"a1816000",
     5220 => x"e0000003",  5221 => x"34010002",  5222 => x"59610004",
     5223 => x"29620004",  5224 => x"29610000",  5225 => x"44410005",
     5226 => x"596002d4",  5227 => x"596002cc",  5228 => x"b9600800",
     5229 => x"f8000659",  5230 => x"296e02d4",  5231 => x"340d0000",
     5232 => x"45c0000a",  5233 => x"29610028",  5234 => x"34020000",
     5235 => x"28230018",  5236 => x"b9600800",  5237 => x"d8600000",
     5238 => x"c9c16800",  5239 => x"a5a00800",  5240 => x"1421001f",
     5241 => x"a1a16800",  5242 => x"296e02cc",  5243 => x"b9a00800",
     5244 => x"45c0000a",  5245 => x"29610028",  5246 => x"34020000",
     5247 => x"28230018",  5248 => x"b9600800",  5249 => x"d8600000",
     5250 => x"c9c10800",  5251 => x"a4201000",  5252 => x"1442001f",
     5253 => x"a0220800",  5254 => x"4da10002",  5255 => x"b9a00800",
     5256 => x"59610008",  5257 => x"b9800800",  5258 => x"2b9d0004",
     5259 => x"2b8b0014",  5260 => x"2b8c0010",  5261 => x"2b8d000c",
     5262 => x"2b8e0008",  5263 => x"379c002c",  5264 => x"c3a00000",
     5265 => x"b9600800",  5266 => x"34020000",  5267 => x"f8000850",
     5268 => x"b9600800",  5269 => x"596002cc",  5270 => x"f80004f6",
     5271 => x"29630100",  5272 => x"29620104",  5273 => x"296500f8",
     5274 => x"296400fc",  5275 => x"b8206000",  5276 => x"29610108",
     5277 => x"596300b0",  5278 => x"296302c8",  5279 => x"596200b4",
     5280 => x"596100b8",  5281 => x"596500a8",  5282 => x"596400ac",
     5283 => x"1063000a",  5284 => x"b9600800",  5285 => x"34020000",
     5286 => x"f800084c",  5287 => x"29620020",  5288 => x"356100a8",
     5289 => x"28430008",  5290 => x"b8201000",  5291 => x"34630018",
     5292 => x"f80005bd",  5293 => x"e3ffffb2",  5294 => x"379cfff8",
     5295 => x"5b8b0008",  5296 => x"5b9d0004",  5297 => x"282202c8",
     5298 => x"28240028",  5299 => x"b8205800",  5300 => x"4043000c",
     5301 => x"1042000b",  5302 => x"bc621000",  5303 => x"28830018",
     5304 => x"084203e8",  5305 => x"d8600000",  5306 => x"596102d4",
     5307 => x"2b9d0004",  5308 => x"2b8b0008",  5309 => x"379c0008",
     5310 => x"c3a00000",  5311 => x"379cffe4",  5312 => x"5b8b001c",
     5313 => x"5b8c0018",  5314 => x"5b8d0014",  5315 => x"5b8e0010",
     5316 => x"5b8f000c",  5317 => x"5b900008",  5318 => x"5b9d0004",
     5319 => x"340c0000",  5320 => x"b8205800",  5321 => x"b8407000",
     5322 => x"342f030c",  5323 => x"34300320",  5324 => x"e0000013",
     5325 => x"098d0058",  5326 => x"ba000800",  5327 => x"3403000a",
     5328 => x"35a20110",  5329 => x"b5621000",  5330 => x"f80036be",
     5331 => x"5c20000b",  5332 => x"b56d0800",  5333 => x"b9e01000",
     5334 => x"34030024",  5335 => x"34210144",  5336 => x"f80036d9",
     5337 => x"b56d5800",  5338 => x"b9c00800",  5339 => x"3562011c",
     5340 => x"f80003be",  5341 => x"e0000020",  5342 => x"358c0001",
     5343 => x"2d63010c",  5344 => x"486cffed",  5345 => x"34010004",
     5346 => x"54610003",  5347 => x"34630001",  5348 => x"0d63010c",
     5349 => x"2d6d010c",  5350 => x"35620320",  5351 => x"3403000a",
     5352 => x"35adffff",  5353 => x"09ac0058",  5354 => x"35810110",
     5355 => x"b5610800",  5356 => x"f80036c5",  5357 => x"b56c0800",
     5358 => x"34030024",  5359 => x"b9e01000",  5360 => x"34210144",
     5361 => x"f80036c0",  5362 => x"b56c1000",  5363 => x"b9c00800",
     5364 => x"3442011c",  5365 => x"f80003a5",  5366 => x"78040001",
     5367 => x"b9600800",  5368 => x"34020003",  5369 => x"34030001",
     5370 => x"3884439c",  5371 => x"b9a02800",  5372 => x"fbffed56",
     5373 => x"2b9d0004",  5374 => x"2b8b001c",  5375 => x"2b8c0018",
     5376 => x"2b8d0014",  5377 => x"2b8e0010",  5378 => x"2b8f000c",
     5379 => x"2b900008",  5380 => x"379c001c",  5381 => x"c3a00000",
     5382 => x"4022001e",  5383 => x"34030001",  5384 => x"44430009",
     5385 => x"44400008",  5386 => x"34030002",  5387 => x"5c430008",
     5388 => x"34020012",  5389 => x"58220070",  5390 => x"3402000e",
     5391 => x"58220074",  5392 => x"e0000003",  5393 => x"58200070",
     5394 => x"58200074",  5395 => x"28240070",  5396 => x"2825002c",
     5397 => x"34020000",  5398 => x"b4a42800",  5399 => x"20a30003",
     5400 => x"44600003",  5401 => x"34020004",  5402 => x"c8431000",
     5403 => x"b4a22800",  5404 => x"28260030",  5405 => x"28220074",
     5406 => x"5825003c",  5407 => x"34030000",  5408 => x"b4c23000",
     5409 => x"20c70003",  5410 => x"44e00003",  5411 => x"34030004",
     5412 => x"c8671800",  5413 => x"b4c31800",  5414 => x"c8a42000",
     5415 => x"c8621000",  5416 => x"58230040",  5417 => x"58240034",
     5418 => x"58220038",  5419 => x"c3a00000",  5420 => x"379cfff4",
     5421 => x"5b8b000c",  5422 => x"5b8c0008",  5423 => x"5b9d0004",
     5424 => x"78020001",  5425 => x"384266bc",  5426 => x"28420020",
     5427 => x"b8205800",  5428 => x"44400006",  5429 => x"d8400000",
     5430 => x"b8206000",  5431 => x"34010001",  5432 => x"45810018",
     5433 => x"480c0018",  5434 => x"296102d4",  5435 => x"340c0000",
     5436 => x"44200015",  5437 => x"29610028",  5438 => x"34020000",
     5439 => x"28230018",  5440 => x"b9600800",  5441 => x"d8600000",
     5442 => x"296202d4",  5443 => x"c8220800",  5444 => x"4c200013",
     5445 => x"e000000c",  5446 => x"4162001d",  5447 => x"34010002",
     5448 => x"44410004",  5449 => x"34010006",  5450 => x"59610004",
     5451 => x"e0000006",  5452 => x"34010004",  5453 => x"59610004",
     5454 => x"b9600800",  5455 => x"fbffff5f",  5456 => x"340c0000",
     5457 => x"b9800800",  5458 => x"2b9d0004",  5459 => x"2b8b000c",
     5460 => x"2b8c0008",  5461 => x"379c000c",  5462 => x"c3a00000",
     5463 => x"b9600800",  5464 => x"34020002",  5465 => x"f800078a",
     5466 => x"29610020",  5467 => x"596002d4",  5468 => x"0d60010c",
     5469 => x"2821000c",  5470 => x"4022000e",  5471 => x"340100ff",
     5472 => x"5c41ffe6",  5473 => x"e3ffffeb",  5474 => x"379cfff4",
     5475 => x"5b8b000c",  5476 => x"5b8c0008",  5477 => x"5b9d0004",
     5478 => x"3404003f",  5479 => x"b8205800",  5480 => x"340cffff",
     5481 => x"4c83000e",  5482 => x"fbffff55",  5483 => x"b9600800",
     5484 => x"fbffff42",  5485 => x"b9600800",  5486 => x"f800015a",
     5487 => x"59610004",  5488 => x"78010001",  5489 => x"382166bc",
     5490 => x"28220024",  5491 => x"340c0000",  5492 => x"44400003",
     5493 => x"b9600800",  5494 => x"d8400000",  5495 => x"b9800800",
     5496 => x"2b9d0004",  5497 => x"2b8b000c",  5498 => x"2b8c0008",
     5499 => x"379c000c",  5500 => x"c3a00000",  5501 => x"379cffe0",
     5502 => x"5b8b0014",  5503 => x"5b8c0010",  5504 => x"5b8d000c",
     5505 => x"5b8e0008",  5506 => x"5b9d0004",  5507 => x"b8205800",
     5508 => x"3401002b",  5509 => x"b8407000",  5510 => x"340cffff",
     5511 => x"4c230028",  5512 => x"4161001c",  5513 => x"340c0000",
     5514 => x"20210001",  5515 => x"44200024",  5516 => x"296300ec",
     5517 => x"296200f0",  5518 => x"296100f4",  5519 => x"296500e4",
     5520 => x"296400e8",  5521 => x"5963009c",  5522 => x"596200a0",
     5523 => x"2963031c",  5524 => x"29620318",  5525 => x"596100a4",
     5526 => x"59650094",  5527 => x"356100d0",  5528 => x"59640098",
     5529 => x"f8000485",  5530 => x"41610313",  5531 => x"20210002",
     5532 => x"44200007",  5533 => x"4161001c",  5534 => x"38210002",
     5535 => x"3161001c",  5536 => x"2d61032a",  5537 => x"0d6102ec",
     5538 => x"e000000d",  5539 => x"378d0018",  5540 => x"b9c00800",
     5541 => x"b9a01000",  5542 => x"f80002ed",  5543 => x"4161001c",
     5544 => x"b9a01000",  5545 => x"202100fd",  5546 => x"3161001c",
     5547 => x"35610080",  5548 => x"f80004aa",  5549 => x"b9600800",
     5550 => x"f8000551",  5551 => x"b9800800",  5552 => x"2b9d0004",
     5553 => x"2b8b0014",  5554 => x"2b8c0010",  5555 => x"2b8d000c",
     5556 => x"2b8e0008",  5557 => x"379c0020",  5558 => x"c3a00000",
     5559 => x"379cffe4",  5560 => x"5b8b0010",  5561 => x"5b8c000c",
     5562 => x"5b8d0008",  5563 => x"5b9d0004",  5564 => x"b8205800",
     5565 => x"b8400800",  5566 => x"3402002b",  5567 => x"3404ffff",
     5568 => x"4c430031",  5569 => x"4162001c",  5570 => x"20430001",
     5571 => x"5c600004",  5572 => x"78010001",  5573 => x"382143bc",
     5574 => x"e0000005",  5575 => x"20420002",  5576 => x"5c400007",
     5577 => x"78010001",  5578 => x"382143f8",  5579 => x"78020001",
     5580 => x"38425c0c",  5581 => x"f8001beb",  5582 => x"e0000022",
     5583 => x"2d6402ec",  5584 => x"2d63032a",  5585 => x"44830007",
     5586 => x"78010001",  5587 => x"78020001",  5588 => x"38425c0c",
     5589 => x"38214430",  5590 => x"f8001be2",  5591 => x"e0000019",
     5592 => x"378d0014",  5593 => x"b9a01000",  5594 => x"f80002ec",
     5595 => x"4161001c",  5596 => x"356c0080",  5597 => x"b9a01000",
     5598 => x"202100fd",  5599 => x"3161001c",  5600 => x"b9800800",
     5601 => x"f8000475",  5602 => x"78030001",  5603 => x"386366bc",
     5604 => x"28640028",  5605 => x"44800009",  5606 => x"b9600800",
     5607 => x"b9801000",  5608 => x"356300d0",  5609 => x"d8800000",
     5610 => x"b8202000",  5611 => x"34010001",  5612 => x"44810004",
     5613 => x"48040004",  5614 => x"b9600800",  5615 => x"f8000510",
     5616 => x"34040000",  5617 => x"b8800800",  5618 => x"2b9d0004",
     5619 => x"2b8b0010",  5620 => x"2b8c000c",  5621 => x"2b8d0008",
     5622 => x"379c001c",  5623 => x"c3a00000",  5624 => x"379cfff0",
     5625 => x"5b8b0010",  5626 => x"5b8c000c",  5627 => x"5b8d0008",
     5628 => x"5b9d0004",  5629 => x"b8406800",  5630 => x"3402003f",
     5631 => x"b8205800",  5632 => x"340cffff",  5633 => x"4c430013",
     5634 => x"78040001",  5635 => x"34030002",  5636 => x"38844470",
     5637 => x"34020003",  5638 => x"fbffec4c",  5639 => x"b9a01000",
     5640 => x"b9600800",  5641 => x"fbfffeb6",  5642 => x"b9600800",
     5643 => x"f80000bd",  5644 => x"59610004",  5645 => x"78010001",
     5646 => x"382166bc",  5647 => x"28220024",  5648 => x"340c0000",
     5649 => x"44400003",  5650 => x"b9600800",  5651 => x"d8400000",
     5652 => x"b9800800",  5653 => x"2b9d0004",  5654 => x"2b8b0010",
     5655 => x"2b8c000c",  5656 => x"2b8d0008",  5657 => x"379c0010",
     5658 => x"c3a00000",  5659 => x"34010000",  5660 => x"c3a00000",
     5661 => x"379cfffc",  5662 => x"5b9d0004",  5663 => x"34030008",
     5664 => x"f8003570",  5665 => x"2b9d0004",  5666 => x"379c0004",
     5667 => x"c3a00000",  5668 => x"379cffe0",  5669 => x"5b8b0020",
     5670 => x"5b8c001c",  5671 => x"5b8d0018",  5672 => x"5b8e0014",
     5673 => x"5b8f0010",  5674 => x"5b90000c",  5675 => x"5b910008",
     5676 => x"5b9d0004",  5677 => x"780e0001",  5678 => x"39ce5c2c",
     5679 => x"78040001",  5680 => x"b8406800",  5681 => x"b8606000",
     5682 => x"34020003",  5683 => x"34030002",  5684 => x"38844818",
     5685 => x"b9c02800",  5686 => x"b8207800",  5687 => x"35b10021",
     5688 => x"fbffec1a",  5689 => x"35900021",  5690 => x"ba200800",
     5691 => x"ba001000",  5692 => x"fbffffe1",  5693 => x"5c200033",
     5694 => x"2d81002a",  5695 => x"2dab002a",  5696 => x"c9615800",
     5697 => x"35620001",  5698 => x"34010002",  5699 => x"54410043",
     5700 => x"29e20020",  5701 => x"34030001",  5702 => x"35a10048",
     5703 => x"28420014",  5704 => x"5d63000b",  5705 => x"fbffffd4",
     5706 => x"5c20003c",  5707 => x"78040001",  5708 => x"b9e00800",
     5709 => x"34020003",  5710 => x"34030001",  5711 => x"388444a0",
     5712 => x"b9c02800",  5713 => x"3406008f",  5714 => x"e000000e",
     5715 => x"3403ffff",  5716 => x"358c0048",  5717 => x"5d63000e",
     5718 => x"b9800800",  5719 => x"fbffffc6",  5720 => x"5c20002e",
     5721 => x"78040001",  5722 => x"b9e00800",  5723 => x"34020003",
     5724 => x"34030001",  5725 => x"388444a0",  5726 => x"b9c02800",
     5727 => x"34060098",  5728 => x"fbffebf2",  5729 => x"340b0000",
     5730 => x"e0000024",  5731 => x"b9801000",  5732 => x"fbffffb9",
     5733 => x"b8205800",  5734 => x"5c200020",  5735 => x"78040001",
     5736 => x"b9e00800",  5737 => x"34020003",  5738 => x"34030001",
     5739 => x"388444b0",  5740 => x"b9c02800",  5741 => x"340600a0",
     5742 => x"fbffebe4",  5743 => x"e0000017",  5744 => x"41ab001a",
     5745 => x"4181001a",  5746 => x"5d61000e",  5747 => x"41ab001c",
     5748 => x"4181001c",  5749 => x"5d61000b",  5750 => x"41ab001d",
     5751 => x"4181001d",  5752 => x"5d610008",  5753 => x"2da2001e",
     5754 => x"2d81001e",  5755 => x"340b0000",  5756 => x"5c41000a",
     5757 => x"41ab0020",  5758 => x"41810020",  5759 => x"45610003",
     5760 => x"c9615800",  5761 => x"e0000005",  5762 => x"ba200800",
     5763 => x"ba001000",  5764 => x"fbffff99",  5765 => x"b8205800",
     5766 => x"b9600800",  5767 => x"2b9d0004",  5768 => x"2b8b0020",
     5769 => x"2b8c001c",  5770 => x"2b8d0018",  5771 => x"2b8e0014",
     5772 => x"2b8f0010",  5773 => x"2b90000c",  5774 => x"2b910008",
     5775 => x"379c0020",  5776 => x"c3a00000",  5777 => x"379cfffc",
     5778 => x"5b9d0004",  5779 => x"34020000",  5780 => x"34030014",
     5781 => x"f800359a",  5782 => x"2b9d0004",  5783 => x"379c0004",
     5784 => x"c3a00000",  5785 => x"379cfff0",  5786 => x"5b8b0010",
     5787 => x"5b8c000c",  5788 => x"5b8d0008",  5789 => x"5b9d0004",
     5790 => x"b8206800",  5791 => x"28210020",  5792 => x"282c0014",
     5793 => x"282b000c",  5794 => x"28210010",  5795 => x"0c200000",
     5796 => x"34210004",  5797 => x"fbffffec",  5798 => x"29a10020",
     5799 => x"28210010",  5800 => x"34210018",  5801 => x"fbffffe8",
     5802 => x"b9800800",  5803 => x"34020000",  5804 => x"34030020",
     5805 => x"f8003582",  5806 => x"29610004",  5807 => x"3402ffa0",
     5808 => x"59810000",  5809 => x"29610008",  5810 => x"59810004",
     5811 => x"29610004",  5812 => x"59810010",  5813 => x"29610008",
     5814 => x"59810014",  5815 => x"2d61000e",  5816 => x"0d810018",
     5817 => x"2d610010",  5818 => x"0d81001a",  5819 => x"41610012",
     5820 => x"3181001c",  5821 => x"41610013",  5822 => x"3181001d",
     5823 => x"29a10020",  5824 => x"28210018",  5825 => x"3022001c",
     5826 => x"2b9d0004",  5827 => x"2b8b0010",  5828 => x"2b8c000c",
     5829 => x"2b8d0008",  5830 => x"379c0010",  5831 => x"c3a00000",
     5832 => x"379cff8c",  5833 => x"5b8b0018",  5834 => x"5b8c0014",
     5835 => x"5b8d0010",  5836 => x"5b8e000c",  5837 => x"5b8f0008",
     5838 => x"5b9d0004",  5839 => x"2c22010c",  5840 => x"b8205800",
     5841 => x"340d0000",  5842 => x"340c0001",  5843 => x"5c400014",
     5844 => x"28230000",  5845 => x"b8406800",  5846 => x"34020006",
     5847 => x"5c620010",  5848 => x"fbffffc1",  5849 => x"29610000",
     5850 => x"e0000105",  5851 => x"09820058",  5852 => x"09a30058",
     5853 => x"b9600800",  5854 => x"34420110",  5855 => x"34630110",
     5856 => x"b5621000",  5857 => x"b5631800",  5858 => x"fbffff42",
     5859 => x"48010002",  5860 => x"e0000002",  5861 => x"b9806800",
     5862 => x"358c0001",  5863 => x"2d66010c",  5864 => x"48ccfff3",
     5865 => x"78040001",  5866 => x"b9600800",  5867 => x"34020003",
     5868 => x"34030001",  5869 => x"388444c0",  5870 => x"b9a02800",
     5871 => x"fbffeb63",  5872 => x"1d61010e",  5873 => x"442d0022",
     5874 => x"0d6d010e",  5875 => x"296c0020",  5876 => x"340f0000",
     5877 => x"340e0001",  5878 => x"e0000015",  5879 => x"29820000",
     5880 => x"09c10374",  5881 => x"b4410800",  5882 => x"2c23010c",
     5883 => x"4460000f",  5884 => x"09e40374",  5885 => x"1c23010e",
     5886 => x"b4442000",  5887 => x"1c82010e",  5888 => x"08630058",
     5889 => x"08420058",  5890 => x"34630110",  5891 => x"b4231800",
     5892 => x"34420110",  5893 => x"b4821000",  5894 => x"fbffff1e",
     5895 => x"48010002",  5896 => x"e0000002",  5897 => x"b9c07800",
     5898 => x"35ce0001",  5899 => x"2981000c",  5900 => x"2c21000c",
     5901 => x"482effea",  5902 => x"2981001c",  5903 => x"442f0004",
     5904 => x"34010001",  5905 => x"598f001c",  5906 => x"59810020",
     5907 => x"4162001d",  5908 => x"34010002",  5909 => x"44410063",
     5910 => x"2d61010c",  5911 => x"5c200004",  5912 => x"29620000",
     5913 => x"34010004",  5914 => x"444100c5",  5915 => x"29610020",
     5916 => x"09ac0058",  5917 => x"2821000c",  5918 => x"4023000a",
     5919 => x"4022000b",  5920 => x"40290004",  5921 => x"40280005",
     5922 => x"40270006",  5923 => x"40260007",  5924 => x"40250008",
     5925 => x"40240009",  5926 => x"33830047",  5927 => x"33890041",
     5928 => x"33880042",  5929 => x"33870043",  5930 => x"33860044",
     5931 => x"33850045",  5932 => x"33840046",  5933 => x"33820048",
     5934 => x"2c22000e",  5935 => x"35830110",  5936 => x"b5631800",
     5937 => x"0f82003c",  5938 => x"2c220010",  5939 => x"0f82003e",
     5940 => x"40220012",  5941 => x"3382003a",  5942 => x"40220013",
     5943 => x"0f80004a",  5944 => x"33820040",  5945 => x"28220004",
     5946 => x"5b820068",  5947 => x"28210008",  5948 => x"37820020",
     5949 => x"5b81006c",  5950 => x"b9600800",  5951 => x"fbfffee5",
     5952 => x"4162001d",  5953 => x"34030001",  5954 => x"44430029",
     5955 => x"29620020",  5956 => x"78050001",  5957 => x"38a55c3c",
     5958 => x"2844000c",  5959 => x"1086000e",  5960 => x"48060004",
     5961 => x"48010023",  5962 => x"5c200019",  5963 => x"e0000006",
     5964 => x"48010020",  5965 => x"44200004",  5966 => x"2c81000c",
     5967 => x"5c23000a",  5968 => x"e0000028",  5969 => x"78040001",
     5970 => x"b9600800",  5971 => x"34020003",  5972 => x"34030001",
     5973 => x"388444e0",  5974 => x"fbffeafc",  5975 => x"34010002",
     5976 => x"e0000087",  5977 => x"29630338",  5978 => x"2841001c",
     5979 => x"4461001d",  5980 => x"b56c1000",  5981 => x"37810041",
     5982 => x"34420131",  5983 => x"5b85001c",  5984 => x"fbfffebd",
     5985 => x"2b85001c",  5986 => x"5c20000c",  5987 => x"78040001",
     5988 => x"b9600800",  5989 => x"34020003",  5990 => x"34030001",
     5991 => x"388444ec",  5992 => x"fbffeaea",  5993 => x"34010007",
     5994 => x"e0000075",  5995 => x"4c200003",  5996 => x"b9600800",
     5997 => x"fbffff2c",  5998 => x"78040001",  5999 => x"78050001",
     6000 => x"b9600800",  6001 => x"34020003",  6002 => x"34030001",
     6003 => x"388444fc",  6004 => x"38a55c3c",  6005 => x"fbffeadd",
     6006 => x"34010006",  6007 => x"e0000068",  6008 => x"09a30058",
     6009 => x"29620020",  6010 => x"b5631800",  6011 => x"2c64013a",
     6012 => x"284c0018",  6013 => x"28410014",  6014 => x"28420010",
     6015 => x"34840001",  6016 => x"0c440000",  6017 => x"34620150",
     6018 => x"28450008",  6019 => x"2844000c",  6020 => x"58250000",
     6021 => x"58240004",  6022 => x"2c420010",  6023 => x"0c220008",
     6024 => x"34620128",  6025 => x"404e0009",  6026 => x"4045000f",
     6027 => x"40440010",  6028 => x"404a000a",  6029 => x"4049000b",
     6030 => x"4048000c",  6031 => x"4047000d",  6032 => x"4046000e",
     6033 => x"302e0010",  6034 => x"30250016",  6035 => x"302a0011",
     6036 => x"30290012",  6037 => x"30280013",  6038 => x"30270014",
     6039 => x"30260015",  6040 => x"30240017",  6041 => x"28440004",
     6042 => x"346e0120",  6043 => x"58240018",  6044 => x"41c4000a",
     6045 => x"3024001c",  6046 => x"40420008",  6047 => x"3022001d",
     6048 => x"4061013c",  6049 => x"3181001c",  6050 => x"1dc50008",
     6051 => x"1d810000",  6052 => x"4425000e",  6053 => x"78040001",
     6054 => x"b9600800",  6055 => x"34020003",  6056 => x"34030001",
     6057 => x"38844508",  6058 => x"fbffeaa8",  6059 => x"2dc10008",
     6060 => x"34020000",  6061 => x"0d810000",  6062 => x"29610028",
     6063 => x"28230004",  6064 => x"b9600800",  6065 => x"d8600000",
     6066 => x"09ad0058",  6067 => x"b56d0800",  6068 => x"34210141",
     6069 => x"4022000b",  6070 => x"20420004",  6071 => x"7c420000",
     6072 => x"59820004",  6073 => x"4022000b",  6074 => x"20420002",
     6075 => x"7c420000",  6076 => x"59820008",  6077 => x"4022000b",
     6078 => x"20420001",  6079 => x"5982000c",  6080 => x"4022000b",
     6081 => x"20420010",  6082 => x"7c420000",  6083 => x"59820010",
     6084 => x"4022000b",  6085 => x"20420020",  6086 => x"7c420000",
     6087 => x"59820014",  6088 => x"4021000b",  6089 => x"20210008",
     6090 => x"7c210000",  6091 => x"59810018",  6092 => x"78010001",
     6093 => x"382166bc",  6094 => x"2824001c",  6095 => x"44800007",
     6096 => x"b56d1000",  6097 => x"b8406800",  6098 => x"b9600800",
     6099 => x"34420144",  6100 => x"35a3011c",  6101 => x"d8800000",
     6102 => x"78040001",  6103 => x"78050001",  6104 => x"b9600800",
     6105 => x"34020003",  6106 => x"34030001",  6107 => x"3884451c",
     6108 => x"38a55c3c",  6109 => x"fbffea75",  6110 => x"34010009",
     6111 => x"2b9d0004",  6112 => x"2b8b0018",  6113 => x"2b8c0014",
     6114 => x"2b8d0010",  6115 => x"2b8e000c",  6116 => x"2b8f0008",
     6117 => x"379c0074",  6118 => x"c3a00000",  6119 => x"379cffec",
     6120 => x"5b8b0014",  6121 => x"5b8c0010",  6122 => x"5b8d000c",
     6123 => x"5b8e0008",  6124 => x"5b9d0004",  6125 => x"b8406000",
     6126 => x"28220024",  6127 => x"b8607000",  6128 => x"28230070",
     6129 => x"2847000c",  6130 => x"28220034",  6131 => x"b8806800",
     6132 => x"b5831800",  6133 => x"342400f8",  6134 => x"b9a02800",
     6135 => x"34060000",  6136 => x"b8205800",  6137 => x"d8e00000",
     6138 => x"78070001",  6139 => x"38e766f4",  6140 => x"3dc20002",
     6141 => x"4c2c000c",  6142 => x"b4e23800",  6143 => x"28e50000",
     6144 => x"78040001",  6145 => x"b9600800",  6146 => x"34020005",
     6147 => x"34030001",  6148 => x"38844154",  6149 => x"b9c03000",
     6150 => x"fbffea4c",  6151 => x"3401ffff",  6152 => x"e0000014",
     6153 => x"b4e24000",  6154 => x"296600f8",  6155 => x"296700fc",
     6156 => x"29080000",  6157 => x"78040001",  6158 => x"b9600800",
     6159 => x"34020005",  6160 => x"34030001",  6161 => x"38844174",
     6162 => x"b9802800",  6163 => x"fbffea3f",  6164 => x"34010001",
     6165 => x"5da10003",  6166 => x"29620104",  6167 => x"44400005",
     6168 => x"2961036c",  6169 => x"34210001",  6170 => x"5961036c",
     6171 => x"34010000",  6172 => x"2b9d0004",  6173 => x"2b8b0014",
     6174 => x"2b8c0010",  6175 => x"2b8d000c",  6176 => x"2b8e0008",
     6177 => x"379c0014",  6178 => x"c3a00000",  6179 => x"379cfff0",
     6180 => x"5b8b0010",  6181 => x"5b8c000c",  6182 => x"5b8d0008",
     6183 => x"5b9d0004",  6184 => x"b8205800",  6185 => x"40410000",
     6186 => x"b8406000",  6187 => x"34030002",  6188 => x"00210004",
     6189 => x"356d0320",  6190 => x"3161030c",  6191 => x"40410000",
     6192 => x"2021000f",  6193 => x"3161030d",  6194 => x"40410001",
     6195 => x"2021000f",  6196 => x"3161030e",  6197 => x"2c410002",
     6198 => x"0d610310",  6199 => x"40410004",  6200 => x"34420006",
     6201 => x"31610312",  6202 => x"35610313",  6203 => x"f8003376",
     6204 => x"35820008",  6205 => x"34030004",  6206 => x"3561031c",
     6207 => x"f8003372",  6208 => x"3582000c",  6209 => x"34030004",
     6210 => x"35610318",  6211 => x"f800336e",  6212 => x"35820014",
     6213 => x"34030008",  6214 => x"b9a00800",  6215 => x"f800336a",
     6216 => x"2d81001c",  6217 => x"296202c8",  6218 => x"34030008",
     6219 => x"0d610328",  6220 => x"2d81001e",  6221 => x"0d61032a",
     6222 => x"41810020",  6223 => x"3161032c",  6224 => x"41810021",
     6225 => x"3161032d",  6226 => x"b9a00800",  6227 => x"f800333d",
     6228 => x"3403ffff",  6229 => x"44200015",  6230 => x"29610020",
     6231 => x"28210014",  6232 => x"2c220008",  6233 => x"4440000a",
     6234 => x"b9a01000",  6235 => x"34030008",  6236 => x"f8003334",
     6237 => x"5c200009",  6238 => x"29610020",  6239 => x"28210014",
     6240 => x"2c220008",  6241 => x"2d610328",  6242 => x"5c410004",
     6243 => x"4161001c",  6244 => x"38210001",  6245 => x"e0000003",
     6246 => x"4161001c",  6247 => x"202100fe",  6248 => x"3161001c",
     6249 => x"34030000",  6250 => x"b8600800",  6251 => x"2b9d0004",
     6252 => x"2b8b0010",  6253 => x"2b8c000c",  6254 => x"2b8d0008",
     6255 => x"379c0010",  6256 => x"c3a00000",  6257 => x"379cfff4",
     6258 => x"5b8b000c",  6259 => x"5b8c0008",  6260 => x"5b9d0004",
     6261 => x"30400000",  6262 => x"b8206000",  6263 => x"282102c8",
     6264 => x"b8405800",  6265 => x"34030008",  6266 => x"4021000e",
     6267 => x"30410001",  6268 => x"29810020",  6269 => x"2821000c",
     6270 => x"40210014",  6271 => x"30410004",  6272 => x"34010002",
     6273 => x"30410006",  6274 => x"34410008",  6275 => x"34020000",
     6276 => x"f80033ab",  6277 => x"298202c8",  6278 => x"35610014",
     6279 => x"34030008",  6280 => x"f8003329",  6281 => x"298102c8",
     6282 => x"2c210008",  6283 => x"0d61001c",  6284 => x"3401007f",
     6285 => x"31610021",  6286 => x"2b9d0004",  6287 => x"2b8b000c",
     6288 => x"2b8c0008",  6289 => x"379c000c",  6290 => x"c3a00000",
     6291 => x"2c230022",  6292 => x"0c430004",  6293 => x"28230024",
     6294 => x"58430000",  6295 => x"28210028",  6296 => x"58410008",
     6297 => x"c3a00000",  6298 => x"379cfff4",  6299 => x"5b8b000c",
     6300 => x"5b8c0008",  6301 => x"5b9d0004",  6302 => x"b8205800",
     6303 => x"2c210022",  6304 => x"b8406000",  6305 => x"34030008",
     6306 => x"0c410004",  6307 => x"29610024",  6308 => x"58410000",
     6309 => x"29610028",  6310 => x"58410008",  6311 => x"2d61002c",
     6312 => x"0c41000c",  6313 => x"4161002f",  6314 => x"3041000e",
     6315 => x"41610030",  6316 => x"30410010",  6317 => x"41610031",
     6318 => x"30410011",  6319 => x"2d610032",  6320 => x"0c410012",
     6321 => x"41610034",  6322 => x"30410014",  6323 => x"34410015",
     6324 => x"35620035",  6325 => x"f80032fc",  6326 => x"2d61003d",
     6327 => x"0d81001e",  6328 => x"4161003f",  6329 => x"31810020",
     6330 => x"78010001",  6331 => x"382166bc",  6332 => x"28230030",
     6333 => x"44600004",  6334 => x"b9600800",  6335 => x"b9801000",
     6336 => x"d8600000",  6337 => x"2b9d0004",  6338 => x"2b8b000c",
     6339 => x"2b8c0008",  6340 => x"379c000c",  6341 => x"c3a00000",
     6342 => x"2c230022",  6343 => x"0c430004",  6344 => x"28230024",
     6345 => x"58430000",  6346 => x"28210028",  6347 => x"58410008",
     6348 => x"c3a00000",  6349 => x"379cfff4",  6350 => x"5b8b000c",
     6351 => x"5b8c0008",  6352 => x"5b9d0004",  6353 => x"b8205800",
     6354 => x"2c210022",  6355 => x"b8406000",  6356 => x"34030008",
     6357 => x"0c410004",  6358 => x"29610024",  6359 => x"58410000",
     6360 => x"29610028",  6361 => x"58410008",  6362 => x"3441000c",
     6363 => x"3562002c",  6364 => x"f80032d5",  6365 => x"2d610034",
     6366 => x"0d810014",  6367 => x"2b9d0004",  6368 => x"2b8b000c",
     6369 => x"2b8c0008",  6370 => x"379c000c",  6371 => x"c3a00000",
     6372 => x"379cfff4",  6373 => x"5b8b000c",  6374 => x"5b8c0008",
     6375 => x"5b9d0004",  6376 => x"282b003c",  6377 => x"b8206000",
     6378 => x"34020000",  6379 => x"41610000",  6380 => x"3403000a",
     6381 => x"202100f0",  6382 => x"3821000b",  6383 => x"31610000",
     6384 => x"34010040",  6385 => x"0d610002",  6386 => x"2d810306",
     6387 => x"34210001",  6388 => x"2021ffff",  6389 => x"0d810306",
     6390 => x"0d61001e",  6391 => x"34010005",  6392 => x"31610020",
     6393 => x"298102c8",  6394 => x"4021000b",  6395 => x"31610021",
     6396 => x"35610022",  6397 => x"f8003332",  6398 => x"29810020",
     6399 => x"34030008",  6400 => x"28220018",  6401 => x"28210014",
     6402 => x"2c420000",  6403 => x"0d62002c",  6404 => x"4021001c",
     6405 => x"3161002f",  6406 => x"29810020",  6407 => x"28210014",
     6408 => x"40210018",  6409 => x"31610030",  6410 => x"29810020",
     6411 => x"28210014",  6412 => x"40210019",  6413 => x"31610031",
     6414 => x"29810020",  6415 => x"28210014",  6416 => x"2c22001a",
     6417 => x"0d620032",  6418 => x"4021001d",  6419 => x"31610034",
     6420 => x"29810020",  6421 => x"28220014",  6422 => x"35610035",
     6423 => x"34420010",  6424 => x"f8003299",  6425 => x"29810020",
     6426 => x"28220010",  6427 => x"28210018",  6428 => x"2c420000",
     6429 => x"0d62003d",  6430 => x"4021001c",  6431 => x"34020040",
     6432 => x"3161003f",  6433 => x"78010001",  6434 => x"382166bc",
     6435 => x"2823002c",  6436 => x"44600004",  6437 => x"b9800800",
     6438 => x"d8600000",  6439 => x"b8201000",  6440 => x"b9800800",
     6441 => x"3403000b",  6442 => x"34040000",  6443 => x"fbfffebc",
     6444 => x"2b9d0004",  6445 => x"2b8b000c",  6446 => x"2b8c0008",
     6447 => x"379c000c",  6448 => x"c3a00000",  6449 => x"379cffc8",
     6450 => x"5b8b0018",  6451 => x"5b8c0014",  6452 => x"5b8d0010",
     6453 => x"5b8e000c",  6454 => x"5b8f0008",  6455 => x"5b9d0004",
     6456 => x"28220028",  6457 => x"378c001c",  6458 => x"b8205800",
     6459 => x"28430000",  6460 => x"b9801000",  6461 => x"378f0030",
     6462 => x"d8600000",  6463 => x"b9800800",  6464 => x"b9e01000",
     6465 => x"f8000103",  6466 => x"296c003c",  6467 => x"340efff0",
     6468 => x"340d002c",  6469 => x"41810000",  6470 => x"0d8d0002",
     6471 => x"34020000",  6472 => x"a02e0800",  6473 => x"31810000",
     6474 => x"2d6102f0",  6475 => x"34030008",  6476 => x"34210001",
     6477 => x"2021ffff",  6478 => x"0d6102f0",  6479 => x"31800020",
     6480 => x"0d81001e",  6481 => x"296102c8",  6482 => x"4021000d",
     6483 => x"31810021",  6484 => x"35810008",  6485 => x"f80032da",
     6486 => x"2f810034",  6487 => x"3402002c",  6488 => x"34030000",
     6489 => x"0d810022",  6490 => x"2b810030",  6491 => x"34040001",
     6492 => x"59810024",  6493 => x"2b810038",  6494 => x"59810028",
     6495 => x"b9600800",  6496 => x"fbfffe87",  6497 => x"5c200023",
     6498 => x"29610020",  6499 => x"356c00f8",  6500 => x"b9801000",
     6501 => x"28230008",  6502 => x"b9800800",  6503 => x"34630018",
     6504 => x"f8000101",  6505 => x"b9e01000",  6506 => x"b9800800",
     6507 => x"f80000d9",  6508 => x"2961003c",  6509 => x"34030008",
     6510 => x"34040000",  6511 => x"40220000",  6512 => x"0c2d0002",
     6513 => x"a04e7000",  6514 => x"39ce0008",  6515 => x"302e0000",
     6516 => x"2d6202f0",  6517 => x"0c22001e",  6518 => x"34020002",
     6519 => x"30220020",  6520 => x"296202c8",  6521 => x"4042000d",
     6522 => x"30220021",  6523 => x"2f820034",  6524 => x"0c220022",
     6525 => x"2b820030",  6526 => x"58220024",  6527 => x"2b820038",
     6528 => x"58220028",  6529 => x"b9600800",  6530 => x"3402002c",
     6531 => x"fbfffe64",  6532 => x"2b9d0004",  6533 => x"2b8b0018",
     6534 => x"2b8c0014",  6535 => x"2b8d0010",  6536 => x"2b8e000c",
     6537 => x"2b8f0008",  6538 => x"379c0038",  6539 => x"c3a00000",
     6540 => x"379cffd4",  6541 => x"5b8b000c",  6542 => x"5b8c0008",
     6543 => x"5b9d0004",  6544 => x"28220028",  6545 => x"378b0010",
     6546 => x"b8206000",  6547 => x"28430000",  6548 => x"b9601000",
     6549 => x"d8600000",  6550 => x"37820024",  6551 => x"b9600800",
     6552 => x"f80000ac",  6553 => x"298b003c",  6554 => x"34020000",
     6555 => x"34030008",  6556 => x"41610000",  6557 => x"202100f0",
     6558 => x"38210001",  6559 => x"31610000",  6560 => x"3401002c",
     6561 => x"0d610002",  6562 => x"2d8102f2",  6563 => x"34210001",
     6564 => x"2021ffff",  6565 => x"0d8102f2",  6566 => x"0d61001e",
     6567 => x"34010001",  6568 => x"31610020",  6569 => x"3401007f",
     6570 => x"31610021",  6571 => x"35610008",  6572 => x"f8003283",
     6573 => x"2f810028",  6574 => x"3402002c",  6575 => x"34030001",
     6576 => x"0d610022",  6577 => x"2b810024",  6578 => x"34040001",
     6579 => x"59610024",  6580 => x"2b81002c",  6581 => x"59610028",
     6582 => x"b9800800",  6583 => x"fbfffe30",  6584 => x"2b9d0004",
     6585 => x"2b8b000c",  6586 => x"2b8c0008",  6587 => x"379c002c",
     6588 => x"c3a00000",  6589 => x"379cffe8",  6590 => x"5b8b000c",
     6591 => x"5b8c0008",  6592 => x"5b9d0004",  6593 => x"b8206000",
     6594 => x"b8400800",  6595 => x"37820010",  6596 => x"f8000080",
     6597 => x"298b003c",  6598 => x"34020000",  6599 => x"34030008",
     6600 => x"41610000",  6601 => x"202100f0",  6602 => x"38210009",
     6603 => x"31610000",  6604 => x"34010036",  6605 => x"0d610002",
     6606 => x"41810312",  6607 => x"31610004",  6608 => x"35610008",
     6609 => x"f800325e",  6610 => x"2981031c",  6611 => x"35820320",
     6612 => x"34030008",  6613 => x"59610008",  6614 => x"29810318",
     6615 => x"5961000c",  6616 => x"2d81032a",  6617 => x"0d61001e",
     6618 => x"34010003",  6619 => x"31610020",  6620 => x"298102c8",
     6621 => x"4021000a",  6622 => x"31610021",  6623 => x"2f810014",
     6624 => x"0d610022",  6625 => x"2b810010",  6626 => x"59610024",
     6627 => x"2b810018",  6628 => x"59610028",  6629 => x"3561002c",
     6630 => x"f80031cb",  6631 => x"2d810328",  6632 => x"34020036",
     6633 => x"34030009",  6634 => x"0d610034",  6635 => x"34040000",
     6636 => x"b9800800",  6637 => x"fbfffdfa",  6638 => x"2b9d0004",
     6639 => x"2b8b000c",  6640 => x"2b8c0008",  6641 => x"379c0018",
     6642 => x"c3a00000",  6643 => x"379cfff0",  6644 => x"5b8b0010",
     6645 => x"5b8c000c",  6646 => x"5b8d0008",  6647 => x"5b9d0004",
     6648 => x"78030001",  6649 => x"282d0004",  6650 => x"38635958",
     6651 => x"28620000",  6652 => x"b8205800",  6653 => x"b9a00800",
     6654 => x"f8003105",  6655 => x"78030001",  6656 => x"296c0000",
     6657 => x"38635958",  6658 => x"28620000",  6659 => x"b42c6000",
     6660 => x"596c0000",  6661 => x"b9a00800",  6662 => x"f800312a",
     6663 => x"59610004",  6664 => x"4c0c0007",  6665 => x"4c20000f",
     6666 => x"358cffff",  6667 => x"78030001",  6668 => x"596c0000",
     6669 => x"38635958",  6670 => x"e0000007",  6671 => x"45800009",
     6672 => x"4c010008",  6673 => x"358c0001",  6674 => x"78030001",
     6675 => x"596c0000",  6676 => x"3863596c",  6677 => x"28620000",
     6678 => x"b4220800",  6679 => x"59610004",  6680 => x"2b9d0004",
     6681 => x"2b8b0010",  6682 => x"2b8c000c",  6683 => x"2b8d0008",
     6684 => x"379c0010",  6685 => x"c3a00000",  6686 => x"379cffe8",
     6687 => x"5b8b0008",  6688 => x"5b9d0004",  6689 => x"5b82000c",
     6690 => x"5b830010",  6691 => x"5b830014",  6692 => x"5b820018",
     6693 => x"b8205800",  6694 => x"4c600006",  6695 => x"78010001",
     6696 => x"78020001",  6697 => x"3821459c",  6698 => x"38425c50",
     6699 => x"f800178d",  6700 => x"2b810018",  6701 => x"38028000",
     6702 => x"2b830014",  6703 => x"b4221000",  6704 => x"f4220800",
     6705 => x"00420010",  6706 => x"b4230800",  6707 => x"3c230010",
     6708 => x"00210010",  6709 => x"b8431000",  6710 => x"78030001",
     6711 => x"38635958",  6712 => x"5b820018",  6713 => x"28620000",
     6714 => x"5b810014",  6715 => x"37810014",  6716 => x"fbffec4a",
     6717 => x"59610004",  6718 => x"2b810018",  6719 => x"59610000",
     6720 => x"2b9d0004",  6721 => x"2b8b0008",  6722 => x"379c0018",
     6723 => x"c3a00000",  6724 => x"379cfffc",  6725 => x"5b9d0004",
     6726 => x"28230000",  6727 => x"48030003",  6728 => x"28210004",
     6729 => x"4c200006",  6730 => x"78010001",  6731 => x"382145c8",
     6732 => x"f800176c",  6733 => x"3401ffff",  6734 => x"e0000005",
     6735 => x"58410008",  6736 => x"58430000",  6737 => x"0c400004",
     6738 => x"34010000",  6739 => x"2b9d0004",  6740 => x"379c0004",
     6741 => x"c3a00000",  6742 => x"379cfffc",  6743 => x"5b9d0004",
     6744 => x"78050001",  6745 => x"38a55970",  6746 => x"28430000",
     6747 => x"28a40000",  6748 => x"54640006",  6749 => x"28420008",
     6750 => x"58230000",  6751 => x"58220004",  6752 => x"34010000",
     6753 => x"e0000005",  6754 => x"78010001",  6755 => x"38214604",
     6756 => x"f8001754",  6757 => x"3401ffff",  6758 => x"2b9d0004",
     6759 => x"379c0004",  6760 => x"c3a00000",  6761 => x"379cfffc",
     6762 => x"5b9d0004",  6763 => x"28660000",  6764 => x"28450000",
     6765 => x"28630004",  6766 => x"28420004",  6767 => x"b4c52800",
     6768 => x"58250000",  6769 => x"b4621000",  6770 => x"58220004",
     6771 => x"fbffff80",  6772 => x"2b9d0004",  6773 => x"379c0004",
     6774 => x"c3a00000",  6775 => x"379cfffc",  6776 => x"5b9d0004",
     6777 => x"28460000",  6778 => x"28650000",  6779 => x"c8c52800",
     6780 => x"58250000",  6781 => x"28450004",  6782 => x"28620004",
     6783 => x"c8a21000",  6784 => x"58220004",  6785 => x"fbffff72",
     6786 => x"2b9d0004",  6787 => x"379c0004",  6788 => x"c3a00000",
     6789 => x"379cfffc",  6790 => x"5b9d0004",  6791 => x"78040001",
     6792 => x"38845974",  6793 => x"28230000",  6794 => x"28820000",
     6795 => x"a0621000",  6796 => x"4c400005",  6797 => x"3442ffff",
     6798 => x"3404fffe",  6799 => x"b8441000",  6800 => x"34420001",
     6801 => x"78050001",  6802 => x"38a55958",  6803 => x"28a40000",
     6804 => x"88441000",  6805 => x"28240004",  6806 => x"b4441000",
     6807 => x"0064001f",  6808 => x"b4831800",  6809 => x"14630001",
     6810 => x"58230000",  6811 => x"0043001f",  6812 => x"b4621000",
     6813 => x"14420001",  6814 => x"58220004",  6815 => x"fbffff54",
     6816 => x"2b9d0004",  6817 => x"379c0004",  6818 => x"c3a00000",
     6819 => x"379cfff8",  6820 => x"5b8b0008",  6821 => x"5b9d0004",
     6822 => x"28250000",  6823 => x"78030001",  6824 => x"b8201000",
     6825 => x"38634654",  6826 => x"4805000a",  6827 => x"78030001",
     6828 => x"38634dfc",  6829 => x"5ca00007",  6830 => x"28210004",
     6831 => x"78030001",  6832 => x"38634654",  6833 => x"48a10003",
     6834 => x"78030001",  6835 => x"38634dfc",  6836 => x"28410004",
     6837 => x"14a4001f",  6838 => x"780b0001",  6839 => x"1426001f",
     6840 => x"98853800",  6841 => x"396b7a40",  6842 => x"98c12800",
     6843 => x"78020001",  6844 => x"b9600800",  6845 => x"38424658",
     6846 => x"c8e42000",  6847 => x"c8a62800",  6848 => x"f80016ea",
     6849 => x"b9600800",  6850 => x"2b9d0004",  6851 => x"2b8b0008",
     6852 => x"379c0008",  6853 => x"c3a00000",  6854 => x"379cfff8",
     6855 => x"5b8b0008",  6856 => x"5b9d0004",  6857 => x"28220020",
     6858 => x"28240028",  6859 => x"b8205800",  6860 => x"28430004",
     6861 => x"58600038",  6862 => x"28430014",  6863 => x"0c20010c",
     6864 => x"0c600008",  6865 => x"28830014",  6866 => x"44600013",
     6867 => x"d8600000",  6868 => x"3402ffff",  6869 => x"5c220008",
     6870 => x"78040001",  6871 => x"b9600800",  6872 => x"34020004",
     6873 => x"34030001",  6874 => x"38844664",  6875 => x"fbffe777",
     6876 => x"34010000",  6877 => x"29620020",  6878 => x"c8010800",
     6879 => x"3c21000a",  6880 => x"28420004",  6881 => x"1423001f",
     6882 => x"5841002c",  6883 => x"58430028",  6884 => x"e000000d",
     6885 => x"28420008",  6886 => x"28420038",  6887 => x"20420001",
     6888 => x"5c430005",  6889 => x"28840008",  6890 => x"34020000",
     6891 => x"34030000",  6892 => x"d8800000",  6893 => x"29610020",
     6894 => x"28210004",  6895 => x"58200028",  6896 => x"5820002c",
     6897 => x"29610020",  6898 => x"78040001",  6899 => x"34020004",
     6900 => x"28260004",  6901 => x"34030001",  6902 => x"b9600800",
     6903 => x"28c50028",  6904 => x"28c6002c",  6905 => x"38844680",
     6906 => x"fbffe758",  6907 => x"2b9d0004",  6908 => x"2b8b0008",
     6909 => x"379c0008",  6910 => x"c3a00000",  6911 => x"379cfff0",
     6912 => x"5b8b0010",  6913 => x"5b8c000c",  6914 => x"5b8d0008",
     6915 => x"5b9d0004",  6916 => x"b8205800",  6917 => x"28210020",
     6918 => x"35620094",  6919 => x"35630080",  6920 => x"282d0004",
     6921 => x"356c00d0",  6922 => x"b9a00800",  6923 => x"fbffff6c",
     6924 => x"b9a01000",  6925 => x"b9801800",  6926 => x"b9a00800",
     6927 => x"fbffff68",  6928 => x"b9800800",  6929 => x"fbffff92",
     6930 => x"78040001",  6931 => x"b8202800",  6932 => x"34020004",
     6933 => x"b9600800",  6934 => x"34030003",  6935 => x"388446a0",
     6936 => x"fbffe73a",  6937 => x"2b9d0004",  6938 => x"2b8b0010",
     6939 => x"2b8c000c",  6940 => x"2b8d0008",  6941 => x"379c0010",
     6942 => x"c3a00000",  6943 => x"379cffb8",  6944 => x"5b8b0024",
     6945 => x"5b8c0020",  6946 => x"5b8d001c",  6947 => x"5b8e0018",
     6948 => x"5b8f0014",  6949 => x"5b900010",  6950 => x"5b91000c",
     6951 => x"5b920008",  6952 => x"5b9d0004",  6953 => x"28220020",
     6954 => x"b8205800",  6955 => x"284d0004",  6956 => x"284c0010",
     6957 => x"28220080",  6958 => x"5c400008",  6959 => x"28230084",
     6960 => x"5c620006",  6961 => x"78040001",  6962 => x"34020004",
     6963 => x"34030002",  6964 => x"388446b8",  6965 => x"e000006e",
     6966 => x"35af0014",  6967 => x"357000bc",  6968 => x"357100a8",
     6969 => x"b9e00800",  6970 => x"ba001000",  6971 => x"ba201800",
     6972 => x"fbffff3b",  6973 => x"357200d0",  6974 => x"b9e01000",
     6975 => x"ba401800",  6976 => x"b9e00800",  6977 => x"fbffff36",
     6978 => x"ba400800",  6979 => x"fbffff60",  6980 => x"78040001",
     6981 => x"b8202800",  6982 => x"34020004",  6983 => x"34030003",
     6984 => x"388446d8",  6985 => x"b9600800",  6986 => x"fbffe708",
     6987 => x"35610080",  6988 => x"fbffff57",  6989 => x"78040001",
     6990 => x"b8202800",  6991 => x"34020004",  6992 => x"34030002",
     6993 => x"388446f0",  6994 => x"b9600800",  6995 => x"fbffe6ff",
     6996 => x"35610094",  6997 => x"fbffff4e",  6998 => x"78040001",
     6999 => x"b8202800",  7000 => x"34020004",  7001 => x"34030002",
     7002 => x"388446f8",  7003 => x"b9600800",  7004 => x"fbffe6f6",
     7005 => x"ba200800",  7006 => x"fbffff45",  7007 => x"78040001",
     7008 => x"b8202800",  7009 => x"34020004",  7010 => x"34030002",
     7011 => x"38844700",  7012 => x"b9600800",  7013 => x"fbffe6ed",
     7014 => x"ba000800",  7015 => x"fbffff3c",  7016 => x"78040001",
     7017 => x"b8202800",  7018 => x"34020004",  7019 => x"34030002",
     7020 => x"38844708",  7021 => x"b9600800",  7022 => x"fbffe6e4",
     7023 => x"b9a00800",  7024 => x"fbffff33",  7025 => x"78040001",
     7026 => x"b8202800",  7027 => x"34020004",  7028 => x"34030001",
     7029 => x"38844710",  7030 => x"b9600800",  7031 => x"fbffe6db",
     7032 => x"b9e00800",  7033 => x"fbffff2a",  7034 => x"78040001",
     7035 => x"b8202800",  7036 => x"38844728",  7037 => x"b9600800",
     7038 => x"34020004",  7039 => x"34030001",  7040 => x"fbffe6d2",
     7041 => x"29610020",  7042 => x"358e0018",  7043 => x"28220004",
     7044 => x"b9c00800",  7045 => x"34430014",  7046 => x"fbfffee3",
     7047 => x"b9c00800",  7048 => x"fbfffefd",  7049 => x"b9c00800",
     7050 => x"fbffff19",  7051 => x"78040001",  7052 => x"b8202800",
     7053 => x"34020004",  7054 => x"b9600800",  7055 => x"34030001",
     7056 => x"38844740",  7057 => x"fbffe6c1",  7058 => x"29610020",
     7059 => x"28220010",  7060 => x"28260004",  7061 => x"28420018",
     7062 => x"5c400142",  7063 => x"28210008",  7064 => x"28270030",
     7065 => x"44e2013c",  7066 => x"28c20000",  7067 => x"5c400003",
     7068 => x"28c30014",  7069 => x"44620008",  7070 => x"78040001",
     7071 => x"b9600800",  7072 => x"34020004",  7073 => x"34030001",
     7074 => x"38844754",  7075 => x"fbffe6af",  7076 => x"e0000134",
     7077 => x"28c50004",  7078 => x"48a70003",  7079 => x"28c20018",
     7080 => x"4ce2012d",  7081 => x"28c60018",  7082 => x"78040001",
     7083 => x"b9600800",  7084 => x"34020004",  7085 => x"34030001",
     7086 => x"38844780",  7087 => x"fbffe6a3",  7088 => x"e0000128",
     7089 => x"2982001c",  7090 => x"59a20034",  7091 => x"1c220040",
     7092 => x"29a10034",  7093 => x"3444ffff",  7094 => x"1423001f",
     7095 => x"98612800",  7096 => x"c8a32800",  7097 => x"3403001f",
     7098 => x"c8621800",  7099 => x"94a33800",  7100 => x"34820001",
     7101 => x"34630001",  7102 => x"3484ffff",  7103 => x"5ce0fffc",
     7104 => x"34030001",  7105 => x"bc621000",  7106 => x"4c460002",
     7107 => x"59a20038",  7108 => x"29a30038",  7109 => x"4c620003",
     7110 => x"34630001",  7111 => x"59a30038",  7112 => x"2982001c",
     7113 => x"4c400002",  7114 => x"5981001c",  7115 => x"2982001c",
     7116 => x"4c400002",  7117 => x"5980001c",  7118 => x"2985001c",
     7119 => x"08210003",  7120 => x"4c25000d",  7121 => x"78040001",
     7122 => x"b9600800",  7123 => x"34020004",  7124 => x"34030001",
     7125 => x"388447c4",  7126 => x"fbffe67c",  7127 => x"29a10034",
     7128 => x"29a20038",  7129 => x"3c210001",  7130 => x"34420001",
     7131 => x"b4410800",  7132 => x"5981001c",  7133 => x"29af0038",
     7134 => x"29a20034",  7135 => x"35900004",  7136 => x"35e1ffff",
     7137 => x"88220800",  7138 => x"2982001c",  7139 => x"b4220800",
     7140 => x"b9e01000",  7141 => x"f8002f1e",  7142 => x"59a10034",
     7143 => x"78040001",  7144 => x"b8203000",  7145 => x"b9e02800",
     7146 => x"388447dc",  7147 => x"5981001c",  7148 => x"34020004",
     7149 => x"b9600800",  7150 => x"34030001",  7151 => x"fbffe663",
     7152 => x"b9a01000",  7153 => x"b9c01800",  7154 => x"ba000800",
     7155 => x"fbfffe84",  7156 => x"ba000800",  7157 => x"fbfffeae",
     7158 => x"78040001",  7159 => x"b8202800",  7160 => x"34020004",
     7161 => x"b9600800",  7162 => x"34030001",  7163 => x"38844800",
     7164 => x"fbffe656",  7165 => x"296f0020",  7166 => x"29e10008",
     7167 => x"2825002c",  7168 => x"44a00011",  7169 => x"29820004",
     7170 => x"44400007",  7171 => x"78040001",  7172 => x"b9600800",
     7173 => x"34020004",  7174 => x"34030001",  7175 => x"3884481c",
     7176 => x"e3ffff9b",  7177 => x"29820008",  7178 => x"4ca20007",
     7179 => x"78040001",  7180 => x"b9600800",  7181 => x"34020004",
     7182 => x"34030001",  7183 => x"3884484c",  7184 => x"e00000c3",
     7185 => x"29820004",  7186 => x"44400031",  7187 => x"28220038",
     7188 => x"20410001",  7189 => x"5c2000c3",  7190 => x"20420002",
     7191 => x"5c410019",  7192 => x"296300c4",  7193 => x"296200c8",
     7194 => x"296100cc",  7195 => x"5b830030",  7196 => x"29e30010",
     7197 => x"296500bc",  7198 => x"296400c0",  7199 => x"378c0028",
     7200 => x"5b820034",  7201 => x"5b810038",  7202 => x"b9801000",
     7203 => x"b9800800",  7204 => x"34630018",  7205 => x"5b850028",
     7206 => x"5b84002c",  7207 => x"fbfffe42",  7208 => x"29610028",
     7209 => x"b9801000",  7210 => x"28230004",  7211 => x"b9600800",
     7212 => x"d8600000",  7213 => x"b9600800",  7214 => x"fbfffe98",
     7215 => x"e00000a9",  7216 => x"29820008",  7217 => x"78030001",
     7218 => x"38635978",  7219 => x"28610000",  7220 => x"ec021000",
     7221 => x"78050001",  7222 => x"c8021000",  7223 => x"38a5597c",
     7224 => x"a0411000",  7225 => x"28a10000",  7226 => x"b4411000",
     7227 => x"29610028",  7228 => x"c8021000",  7229 => x"28230010",
     7230 => x"5c600002",  7231 => x"2823000c",  7232 => x"b9600800",
     7233 => x"d8600000",  7234 => x"e0000096",  7235 => x"29830008",
     7236 => x"29ed0004",  7237 => x"78050001",  7238 => x"1462001f",
     7239 => x"29b0002c",  7240 => x"00640016",  7241 => x"3c63000a",
     7242 => x"29ae0028",  7243 => x"3c42000a",  7244 => x"b4708000",
     7245 => x"b8821000",  7246 => x"f4701800",  7247 => x"b44e1000",
     7248 => x"b4627000",  7249 => x"1c22003e",  7250 => x"38a5597c",
     7251 => x"28a40000",  7252 => x"1441001f",  7253 => x"34030000",
     7254 => x"59ae0028",  7255 => x"59b0002c",  7256 => x"f8002e84",
     7257 => x"00430016",  7258 => x"3c21000a",  7259 => x"3c42000a",
     7260 => x"b8610800",  7261 => x"49c1000b",  7262 => x"5dc10002",
     7263 => x"56020009",  7264 => x"c8021000",  7265 => x"7c430000",
     7266 => x"c8010800",  7267 => x"c8230800",  7268 => x"482e0004",
     7269 => x"5c2e0005",  7270 => x"54500002",  7271 => x"e0000003",
     7272 => x"59a10028",  7273 => x"59a2002c",  7274 => x"29a10028",
     7275 => x"29a2002c",  7276 => x"48200003",  7277 => x"5c200004",
     7278 => x"44410003",  7279 => x"340d0000",  7280 => x"e0000002",
     7281 => x"340dffff",  7282 => x"5b810044",  7283 => x"5b820048",
     7284 => x"45a00007",  7285 => x"c8021000",  7286 => x"7c430000",
     7287 => x"c8010800",  7288 => x"c8230800",  7289 => x"5b810044",
     7290 => x"5b820048",  7291 => x"29e20008",  7292 => x"37810044",
     7293 => x"1c42003e",  7294 => x"fbffea08",  7295 => x"45a00009",
     7296 => x"2b810048",  7297 => x"2b820044",  7298 => x"c8010800",
     7299 => x"7c230000",  7300 => x"c8021000",  7301 => x"c8431000",
     7302 => x"5b820044",  7303 => x"5b810048",  7304 => x"29820008",
     7305 => x"1441001f",  7306 => x"00430016",  7307 => x"3c21000a",
     7308 => x"ec026000",  7309 => x"3c42000a",  7310 => x"b8610800",
     7311 => x"c80c6000",  7312 => x"5b81003c",  7313 => x"5b820040",
     7314 => x"45800007",  7315 => x"c8021000",  7316 => x"7c430000",
     7317 => x"c8010800",  7318 => x"c8230800",  7319 => x"5b81003c",
     7320 => x"5b820040",  7321 => x"29610020",  7322 => x"28220008",
     7323 => x"3781003c",  7324 => x"1c42003c",  7325 => x"fbffe9e9",
     7326 => x"45800009",  7327 => x"2b810040",  7328 => x"2b82003c",
     7329 => x"c8010800",  7330 => x"7c230000",  7331 => x"c8021000",
     7332 => x"c8431000",  7333 => x"5b82003c",  7334 => x"5b810040",
     7335 => x"2b830048",  7336 => x"2b820040",  7337 => x"2b81003c",
     7338 => x"2b840044",  7339 => x"b4621000",  7340 => x"f4621800",
     7341 => x"b4810800",  7342 => x"b4610800",  7343 => x"48200003",
     7344 => x"5c200006",  7345 => x"44410005",  7346 => x"3c210016",
     7347 => x"0042000a",  7348 => x"b8221000",  7349 => x"e0000009",
     7350 => x"c8021000",  7351 => x"7c430000",  7352 => x"c8010800",
     7353 => x"c8230800",  7354 => x"3c210016",  7355 => x"0042000a",
     7356 => x"b8221000",  7357 => x"c8021000",  7358 => x"29610020",
     7359 => x"28210008",  7360 => x"28250038",  7361 => x"20a50001",
     7362 => x"5ca00008",  7363 => x"29640028",  7364 => x"c8021000",
     7365 => x"28830010",  7366 => x"5c650002",  7367 => x"2883000c",
     7368 => x"b9600800",  7369 => x"d8600000",  7370 => x"29610020",
     7371 => x"78040001",  7372 => x"34020004",  7373 => x"28210004",
     7374 => x"34030002",  7375 => x"38844888",  7376 => x"2825002c",
     7377 => x"b9600800",  7378 => x"14a5000a",  7379 => x"fbffe57f",
     7380 => x"e0000004",  7381 => x"29a60038",  7382 => x"4c06fedb",
     7383 => x"e3fffedc",  7384 => x"2b9d0004",  7385 => x"2b8b0024",
     7386 => x"2b8c0020",  7387 => x"2b8d001c",  7388 => x"2b8e0018",
     7389 => x"2b8f0014",  7390 => x"2b900010",  7391 => x"2b91000c",
     7392 => x"2b920008",  7393 => x"379c0048",  7394 => x"c3a00000",
     7395 => x"379cfffc",  7396 => x"5b9d0004",  7397 => x"78030001",
     7398 => x"3c420002",  7399 => x"38636734",  7400 => x"b4622800",
     7401 => x"28a50000",  7402 => x"78040001",  7403 => x"34020006",
     7404 => x"34030001",  7405 => x"388448a0",  7406 => x"fbffe564",
     7407 => x"2b9d0004",  7408 => x"379c0004",  7409 => x"c3a00000",
     7410 => x"379cfff0",  7411 => x"5b8b0010",  7412 => x"5b8c000c",
     7413 => x"5b8d0008",  7414 => x"5b9d0004",  7415 => x"b8205800",
     7416 => x"78010001",  7417 => x"38217a58",  7418 => x"b8406800",
     7419 => x"28220000",  7420 => x"5c400005",  7421 => x"29620020",
     7422 => x"2844000c",  7423 => x"28820008",  7424 => x"58220000",
     7425 => x"78040001",  7426 => x"78010001",  7427 => x"38847a58",
     7428 => x"38215980",  7429 => x"28260000",  7430 => x"28850000",
     7431 => x"340c0190",  7432 => x"bd836000",  7433 => x"88a62800",
     7434 => x"b9801000",  7435 => x"34a53039",  7436 => x"00a10010",
     7437 => x"88a62800",  7438 => x"202107ff",  7439 => x"34a53039",
     7440 => x"58850000",  7441 => x"00a50010",  7442 => x"3c24000a",
     7443 => x"20a103ff",  7444 => x"b8240800",  7445 => x"f8002e4b",
     7446 => x"3d820001",  7447 => x"b4221000",  7448 => x"29610028",
     7449 => x"28230018",  7450 => x"b9600800",  7451 => x"d8600000",
     7452 => x"35a200b2",  7453 => x"3c420002",  7454 => x"b5625800",
     7455 => x"59610004",  7456 => x"2b9d0004",  7457 => x"2b8b0010",
     7458 => x"2b8c000c",  7459 => x"2b8d0008",  7460 => x"379c0010",
     7461 => x"c3a00000",  7462 => x"379cfff0",  7463 => x"5b8b0010",
     7464 => x"5b8c000c",  7465 => x"5b8d0008",  7466 => x"5b9d0004",
     7467 => x"282b000c",  7468 => x"b8206000",  7469 => x"34010001",
     7470 => x"59610000",  7471 => x"29810024",  7472 => x"48200002",
     7473 => x"34010001",  7474 => x"0d61000c",  7475 => x"29810008",
     7476 => x"5c200002",  7477 => x"59820008",  7478 => x"298d0008",
     7479 => x"3561000e",  7480 => x"34030004",  7481 => x"b9a01000",
     7482 => x"f8002e77",  7483 => x"2d62000c",  7484 => x"34010001",
     7485 => x"5c410004",  7486 => x"29810000",  7487 => x"4021001d",
     7488 => x"64210002",  7489 => x"59610018",  7490 => x"41a10044",
     7491 => x"2d67000c",  7492 => x"34060002",  7493 => x"31610012",
     7494 => x"41a10045",  7495 => x"34050001",  7496 => x"3404ffff",
     7497 => x"31610013",  7498 => x"41a10046",  7499 => x"31610014",
     7500 => x"34010000",  7501 => x"e000000c",  7502 => x"08220374",
     7503 => x"29880000",  7504 => x"b5021000",  7505 => x"44600004",
     7506 => x"4043001d",  7507 => x"44660002",  7508 => x"59600018",
     7509 => x"58410338",  7510 => x"58450000",  7511 => x"0c44010e",
     7512 => x"34210001",  7513 => x"29630018",  7514 => x"48e1fff4",
     7515 => x"44600006",  7516 => x"78010001",  7517 => x"38214930",
     7518 => x"f800145a",  7519 => x"3401ffff",  7520 => x"3161000e",
     7521 => x"78010001",  7522 => x"382166bc",  7523 => x"28230004",
     7524 => x"34010000",  7525 => x"44600004",  7526 => x"b9800800",
     7527 => x"b9a01000",  7528 => x"d8600000",  7529 => x"2b9d0004",
     7530 => x"2b8b0010",  7531 => x"2b8c000c",  7532 => x"2b8d0008",
     7533 => x"379c0010",  7534 => x"c3a00000",  7535 => x"379cfffc",
     7536 => x"5b9d0004",  7537 => x"78020001",  7538 => x"384266bc",
     7539 => x"28430008",  7540 => x"34020000",  7541 => x"44600003",
     7542 => x"d8600000",  7543 => x"b8201000",  7544 => x"b8400800",
     7545 => x"2b9d0004",  7546 => x"379c0004",  7547 => x"c3a00000",
     7548 => x"78010001",  7549 => x"382167a0",  7550 => x"28220000",
     7551 => x"78010001",  7552 => x"38216584",  7553 => x"e0000004",
     7554 => x"28440000",  7555 => x"44640004",  7556 => x"3421000c",
     7557 => x"28230000",  7558 => x"5c60fffc",  7559 => x"28210004",
     7560 => x"c3a00000",  7561 => x"379cfff4",  7562 => x"5b9d0004",
     7563 => x"5b810008",  7564 => x"5b82000c",  7565 => x"b8401800",
     7566 => x"5c20000b",  7567 => x"78020001",  7568 => x"38425968",
     7569 => x"28410000",  7570 => x"54610007",  7571 => x"78010001",
     7572 => x"78020001",  7573 => x"38424954",  7574 => x"38217a60",
     7575 => x"f8001413",  7576 => x"e000000d",  7577 => x"78030001",
     7578 => x"38635958",  7579 => x"28620000",  7580 => x"37810008",
     7581 => x"fbffe8e9",  7582 => x"2b83000c",  7583 => x"b8202000",
     7584 => x"78020001",  7585 => x"78010001",  7586 => x"38217a60",
     7587 => x"38424958",  7588 => x"f8001406",  7589 => x"78010001",
     7590 => x"38217a60",  7591 => x"2b9d0004",  7592 => x"379c000c",
     7593 => x"c3a00000",  7594 => x"379cff18",  7595 => x"5b8b000c",
     7596 => x"5b8c0008",  7597 => x"5b9d0004",  7598 => x"78010001",
     7599 => x"382167a0",  7600 => x"28210000",  7601 => x"282b0014",
     7602 => x"78010001",  7603 => x"38219248",  7604 => x"28220000",
     7605 => x"34010000",  7606 => x"444000ce",  7607 => x"780c0001",
     7608 => x"398c7a5c",  7609 => x"29810000",  7610 => x"5c200008",
     7611 => x"f80019bd",  7612 => x"78020001",  7613 => x"38426098",
     7614 => x"28420000",  7615 => x"a4401000",  7616 => x"b4410800",
     7617 => x"59810000",  7618 => x"78010001",  7619 => x"38218ee4",
     7620 => x"28210000",  7621 => x"296200b8",  7622 => x"5c220007",
     7623 => x"78010001",  7624 => x"3821754c",  7625 => x"28230000",
     7626 => x"34020003",  7627 => x"34010000",  7628 => x"446200b8",
     7629 => x"f80019ab",  7630 => x"78030001",  7631 => x"78020001",
     7632 => x"38636098",  7633 => x"38427a5c",  7634 => x"28630000",
     7635 => x"28420000",  7636 => x"b4621000",  7637 => x"c8220800",
     7638 => x"4c200007",  7639 => x"78010001",  7640 => x"3821754c",
     7641 => x"28230000",  7642 => x"34020003",  7643 => x"34010000",
     7644 => x"5c6200a8",  7645 => x"f800199b",  7646 => x"78020001",
     7647 => x"38427a5c",  7648 => x"58410000",  7649 => x"296200b8",
     7650 => x"78010001",  7651 => x"38218ee4",  7652 => x"58220000",
     7653 => x"378100d8",  7654 => x"378200e0",  7655 => x"f8001d52",
     7656 => x"34020000",  7657 => x"37810010",  7658 => x"f8000287",
     7659 => x"378100e8",  7660 => x"378200e4",  7661 => x"f8001972",
     7662 => x"2b8300e4",  7663 => x"2b8400e8",  7664 => x"2b82003c",
     7665 => x"78010001",  7666 => x"38214960",  7667 => x"f80013c5",
     7668 => x"2b820044",  7669 => x"78010001",  7670 => x"38214974",
     7671 => x"7c420000",  7672 => x"f80013c0",  7673 => x"fbffff83",
     7674 => x"b8201000",  7675 => x"78010001",  7676 => x"38214980",
     7677 => x"f80013bb",  7678 => x"78010001",  7679 => x"3821754c",
     7680 => x"28220000",  7681 => x"34010003",  7682 => x"5c41000a",
     7683 => x"29620010",  7684 => x"78010001",  7685 => x"38214988",
     7686 => x"20420001",  7687 => x"f80013b1",  7688 => x"78010001",
     7689 => x"38214990",  7690 => x"356200c0",  7691 => x"f80013ad",
     7692 => x"34010000",  7693 => x"f8002ac2",  7694 => x"b8201000",
     7695 => x"78010001",  7696 => x"3821499c",  7697 => x"f80013a7",
     7698 => x"2b8200dc",  7699 => x"2b8300e0",  7700 => x"78010001",
     7701 => x"382149a4",  7702 => x"f80013a2",  7703 => x"78010001",
     7704 => x"3821754c",  7705 => x"28220000",  7706 => x"34010003",
     7707 => x"5c41004b",  7708 => x"296200a4",  7709 => x"296100a0",
     7710 => x"fbffff6b",  7711 => x"b8201000",  7712 => x"78010001",
     7713 => x"382149b4",  7714 => x"f8001396",  7715 => x"296200b4",
     7716 => x"296100b0",  7717 => x"fbffff64",  7718 => x"b8201000",
     7719 => x"78010001",  7720 => x"382149bc",  7721 => x"f800138f",
     7722 => x"29620018",  7723 => x"2963001c",  7724 => x"78010001",
     7725 => x"382149c4",  7726 => x"f800138a",  7727 => x"29620020",
     7728 => x"29630024",  7729 => x"78010001",  7730 => x"382149d8",
     7731 => x"f8001385",  7732 => x"296200b4",  7733 => x"296300a4",
     7734 => x"78010001",  7735 => x"3c420001",  7736 => x"382149ec",
     7737 => x"c8621000",  7738 => x"f800137e",  7739 => x"29620018",
     7740 => x"296100a4",  7741 => x"296300a0",  7742 => x"1444001f",
     7743 => x"c8221000",  7744 => x"f4410800",  7745 => x"c8641800",
     7746 => x"c8611800",  7747 => x"2961001c",  7748 => x"1424001f",
     7749 => x"c8410800",  7750 => x"f4221000",  7751 => x"c8641800",
     7752 => x"c8621000",  7753 => x"29630020",  7754 => x"1464001f",
     7755 => x"c8231800",  7756 => x"f4610800",  7757 => x"c8441000",
     7758 => x"c8410800",  7759 => x"29620024",  7760 => x"1444001f",
     7761 => x"c8621000",  7762 => x"f4431800",  7763 => x"c8240800",
     7764 => x"c8230800",  7765 => x"fbffff34",  7766 => x"b8201000",
     7767 => x"78010001",  7768 => x"382149f8",  7769 => x"f800135f",
     7770 => x"296200ec",  7771 => x"78010001",  7772 => x"38214a04",
     7773 => x"f800135b",  7774 => x"296200a8",  7775 => x"78010001",
     7776 => x"38214a0c",  7777 => x"f8001357",  7778 => x"296200b8",
     7779 => x"78010001",  7780 => x"38214a18",  7781 => x"f8001353",
     7782 => x"3401ffff",  7783 => x"f8002a73",  7784 => x"b8206000",
     7785 => x"34010000",  7786 => x"f8002a70",  7787 => x"b8205800",
     7788 => x"34010001",  7789 => x"f8002a6d",  7790 => x"78050001",
     7791 => x"b8202000",  7792 => x"b8a00800",  7793 => x"b9801000",
     7794 => x"b9601800",  7795 => x"38214a24",  7796 => x"f8001344",
     7797 => x"78010001",  7798 => x"38214a38",  7799 => x"f8001bbd",
     7800 => x"2023ffff",  7801 => x"08632710",  7802 => x"b8201000",
     7803 => x"14420010",  7804 => x"14630010",  7805 => x"78010001",
     7806 => x"38214a3c",  7807 => x"f8001339",  7808 => x"78010001",
     7809 => x"38214cd8",  7810 => x"f8001336",  7811 => x"34010001",
     7812 => x"2b9d0004",  7813 => x"2b8b000c",  7814 => x"2b8c0008",
     7815 => x"379c00e8",  7816 => x"c3a00000",  7817 => x"379cfff4",
     7818 => x"5b8b000c",  7819 => x"5b8c0008",  7820 => x"5b9d0004",
     7821 => x"780b0001",  7822 => x"396b67a0",  7823 => x"29610000",
     7824 => x"78020001",  7825 => x"38424a4c",  7826 => x"282c0014",
     7827 => x"34010004",  7828 => x"f80008f5",  7829 => x"fbfffee7",
     7830 => x"78020001",  7831 => x"b8201800",  7832 => x"38424a5c",
     7833 => x"34010007",  7834 => x"f80008ef",  7835 => x"29810010",
     7836 => x"44200005",  7837 => x"29610000",  7838 => x"28220000",
     7839 => x"34010009",  7840 => x"44410007",  7841 => x"78020001",
     7842 => x"34010001",  7843 => x"38424a60",  7844 => x"f80008e5",
     7845 => x"34010000",  7846 => x"e0000006",  7847 => x"78020001",
     7848 => x"34010004",  7849 => x"38424a78",  7850 => x"f80008df",
     7851 => x"34010001",  7852 => x"2b9d0004",  7853 => x"2b8b000c",
     7854 => x"2b8c0008",  7855 => x"379c000c",  7856 => x"c3a00000",
     7857 => x"379cfef0",  7858 => x"5b8b0018",  7859 => x"5b8c0014",
     7860 => x"5b8d0010",  7861 => x"5b8e000c",  7862 => x"5b8f0008",
     7863 => x"5b9d0004",  7864 => x"78010001",  7865 => x"382167a0",
     7866 => x"28210000",  7867 => x"780c0001",  7868 => x"398c7a7c",
     7869 => x"282b0014",  7870 => x"29810000",  7871 => x"5c200008",
     7872 => x"f80018b8",  7873 => x"78020001",  7874 => x"38426098",
     7875 => x"28420000",  7876 => x"a4401000",  7877 => x"b4410800",
     7878 => x"59810000",  7879 => x"f80018b1",  7880 => x"78030001",
     7881 => x"78020001",  7882 => x"38636098",  7883 => x"38427a7c",
     7884 => x"28630000",  7885 => x"28420000",  7886 => x"b4621000",
     7887 => x"c8220800",  7888 => x"4c200007",  7889 => x"78010001",
     7890 => x"38217a78",  7891 => x"28210000",  7892 => x"296200b8",
     7893 => x"340d0000",  7894 => x"44220192",  7895 => x"f80018a1",
     7896 => x"78020001",  7897 => x"38427a7c",  7898 => x"58410000",
     7899 => x"296200b8",  7900 => x"78010001",  7901 => x"38217a78",
     7902 => x"58220000",  7903 => x"f80008f0",  7904 => x"78040001",
     7905 => x"34010001",  7906 => x"34020001",  7907 => x"34030004",
     7908 => x"38844a94",  7909 => x"f80008c3",  7910 => x"78040001",
     7911 => x"38844ab4",  7912 => x"34030087",  7913 => x"34010002",
     7914 => x"34020001",  7915 => x"f80008bd",  7916 => x"378100fc",
     7917 => x"37820108",  7918 => x"f8001c4b",  7919 => x"78020001",
     7920 => x"34010004",  7921 => x"38424ac0",  7922 => x"f8000897",
     7923 => x"2b820100",  7924 => x"2b8100fc",  7925 => x"34030000",
     7926 => x"f80007e2",  7927 => x"78020001",  7928 => x"b8201800",
     7929 => x"38424a5c",  7930 => x"34010007",  7931 => x"f800088e",
     7932 => x"34020000",  7933 => x"37810020",  7934 => x"f8000173",
     7935 => x"78040001",  7936 => x"34010004",  7937 => x"34020001",
     7938 => x"34030004",  7939 => x"38844ae0",  7940 => x"f80008a4",
     7941 => x"78040001",  7942 => x"78050001",  7943 => x"34010006",
     7944 => x"34020001",  7945 => x"34030007",  7946 => x"38844af0",
     7947 => x"38a54af8",  7948 => x"f800089c",  7949 => x"2b81004c",
     7950 => x"44200005",  7951 => x"78020001",  7952 => x"34010002",
     7953 => x"38424b00",  7954 => x"e0000004",  7955 => x"78020001",
     7956 => x"34010001",  7957 => x"38424b0c",  7958 => x"f8000873",
     7959 => x"2b81004c",  7960 => x"4420014c",  7961 => x"37810110",
     7962 => x"3782010c",  7963 => x"f8001844",  7964 => x"2b83010c",
     7965 => x"2b840110",  7966 => x"78020001",  7967 => x"34010087",
     7968 => x"38424b18",  7969 => x"780c0001",  7970 => x"f8000867",
     7971 => x"398c67a0",  7972 => x"29810000",  7973 => x"282102c8",
     7974 => x"28210010",  7975 => x"282e0008",  7976 => x"5dc00039",
     7977 => x"78020001",  7978 => x"34010001",  7979 => x"38424b34",
     7980 => x"f800085d",  7981 => x"fbffff5c",  7982 => x"340d0001",
     7983 => x"442e0139",  7984 => x"78020001",  7985 => x"34010087",
     7986 => x"38424b3c",  7987 => x"f8000856",  7988 => x"29810000",
     7989 => x"28210020",  7990 => x"28240010",  7991 => x"28830004",
     7992 => x"4460000b",  7993 => x"78020001",  7994 => x"38424b5c",
     7995 => x"28840008",  7996 => x"4c030003",  7997 => x"34010007",
     7998 => x"e0000003",  7999 => x"34010007",  8000 => x"c8042000",
     8001 => x"f8000848",  8002 => x"e0000126",  8003 => x"28830008",
     8004 => x"780b0001",  8005 => x"396b4b68",  8006 => x"b9601000",
     8007 => x"34010007",  8008 => x"f8000841",  8009 => x"78020001",
     8010 => x"34010087",  8011 => x"38424b70",  8012 => x"f800083d",
     8013 => x"29810000",  8014 => x"b9601000",  8015 => x"28210020",
     8016 => x"28230010",  8017 => x"34010007",  8018 => x"2863001c",
     8019 => x"f8000836",  8020 => x"78020001",  8021 => x"34010087",
     8022 => x"38424b90",  8023 => x"f8000832",  8024 => x"29810000",
     8025 => x"b9601000",  8026 => x"28210020",  8027 => x"28240004",
     8028 => x"34010007",  8029 => x"28830028",  8030 => x"2884002c",
     8031 => x"f800082a",  8032 => x"e0000108",  8033 => x"78010001",
     8034 => x"3821754c",  8035 => x"28210000",  8036 => x"34020001",
     8037 => x"4841000e",  8038 => x"34020002",  8039 => x"4c410004",
     8040 => x"34020003",  8041 => x"5c22000a",  8042 => x"e0000005",
     8043 => x"78020001",  8044 => x"34010007",  8045 => x"38424bb0",
     8046 => x"e0000008",  8047 => x"78020001",  8048 => x"34010007",
     8049 => x"38424bbc",  8050 => x"e0000004",  8051 => x"78020001",
     8052 => x"34010001",  8053 => x"38424bc8",  8054 => x"f8000813",
     8055 => x"2b810054",  8056 => x"44200005",  8057 => x"78020001",
     8058 => x"34010002",  8059 => x"38424bd8",  8060 => x"e0000004",
     8061 => x"78020001",  8062 => x"34010001",  8063 => x"38424be4",
     8064 => x"f8000809",  8065 => x"2b810070",  8066 => x"44200007",
     8067 => x"2b810074",  8068 => x"44200005",  8069 => x"78020001",
     8070 => x"34010002",  8071 => x"38424bf0",  8072 => x"e0000004",
     8073 => x"78020001",  8074 => x"34010001",  8075 => x"38424c00",
     8076 => x"f80007fd",  8077 => x"78020001",  8078 => x"38424c10",
     8079 => x"34010007",  8080 => x"f80007f9",  8081 => x"378c0104",
     8082 => x"b9800800",  8083 => x"f8000b85",  8084 => x"378300e8",
     8085 => x"b8600800",  8086 => x"b9801000",  8087 => x"5b83001c",
     8088 => x"f80006a9",  8089 => x"78010001",  8090 => x"38217d48",
     8091 => x"28210000",  8092 => x"34020001",  8093 => x"2b83001c",
     8094 => x"4422000a",  8095 => x"44200004",  8096 => x"34020002",
     8097 => x"5c22000f",  8098 => x"e000000a",  8099 => x"78020001",
     8100 => x"34010001",  8101 => x"38424c18",  8102 => x"f80007e3",
     8103 => x"e0000009",  8104 => x"78020001",  8105 => x"34010002",
     8106 => x"38424c28",  8107 => x"e0000004",  8108 => x"78020001",
     8109 => x"34010002",  8110 => x"38424c38",  8111 => x"f80007da",
     8112 => x"fbfffed9",  8113 => x"340d0001",  8114 => x"442000b6",
     8115 => x"78020001",  8116 => x"34010087",  8117 => x"38424c50",
     8118 => x"f80007d3",  8119 => x"78020001",  8120 => x"34010007",
     8121 => x"38424818",  8122 => x"356300c0",  8123 => x"f80007ce",
     8124 => x"78020001",  8125 => x"34010087",  8126 => x"38424c6c",
     8127 => x"f80007ca",  8128 => x"296100bc",  8129 => x"44200005",
     8130 => x"78020001",  8131 => x"34010002",  8132 => x"38424c88",
     8133 => x"e0000004",  8134 => x"78020001",  8135 => x"34010001",
     8136 => x"38424c8c",  8137 => x"f80007c0",  8138 => x"78020001",
     8139 => x"34010087",  8140 => x"38424c94",  8141 => x"f80007bc",
     8142 => x"34010000",  8143 => x"f8002900",  8144 => x"b8206000",
     8145 => x"20210001",  8146 => x"44200005",  8147 => x"78020001",
     8148 => x"34010002",  8149 => x"38424cb0",  8150 => x"f80007b3",
     8151 => x"218c0002",  8152 => x"45800005",  8153 => x"78020001",
     8154 => x"34010002",  8155 => x"38424cb8",  8156 => x"f80007ad",
     8157 => x"78010001",  8158 => x"38214cd8",  8159 => x"f80011d9",
     8160 => x"78020001",  8161 => x"34010004",  8162 => x"38424cc4",
     8163 => x"f80007a6",  8164 => x"78020001",  8165 => x"34010087",
     8166 => x"38424cdc",  8167 => x"f80007a2",  8168 => x"296200a4",
     8169 => x"296100a0",  8170 => x"780d0001",  8171 => x"39ad4cf8",
     8172 => x"fbfffd9d",  8173 => x"b8201800",  8174 => x"b9a01000",
     8175 => x"34010007",  8176 => x"f8000799",  8177 => x"78020001",
     8178 => x"34010087",  8179 => x"38424d00",  8180 => x"f8000795",
     8181 => x"296200b4",  8182 => x"296100b0",  8183 => x"780c0001",
     8184 => x"398c4d38",  8185 => x"fbfffd90",  8186 => x"b8201800",
     8187 => x"b9a01000",  8188 => x"34010007",  8189 => x"f800078c",
     8190 => x"78020001",  8191 => x"34010087",  8192 => x"38424d1c",
     8193 => x"f8000788",  8194 => x"29630018",  8195 => x"2964001c",
     8196 => x"b9801000",  8197 => x"34010007",  8198 => x"f8000783",
     8199 => x"78020001",  8200 => x"34010087",  8201 => x"38424d50",
     8202 => x"f800077f",  8203 => x"29640024",  8204 => x"29630020",
     8205 => x"b9801000",  8206 => x"34010007",  8207 => x"f800077a",
     8208 => x"296e00b4",  8209 => x"296100a4",  8210 => x"78020001",
     8211 => x"3dce0001",  8212 => x"38424d6c",  8213 => x"c82e7000",
     8214 => x"780c0001",  8215 => x"34010087",  8216 => x"f8000771",
     8217 => x"398c4d88",  8218 => x"b9c01800",  8219 => x"34010007",
     8220 => x"b9801000",  8221 => x"f800076c",  8222 => x"29610018",
     8223 => x"296200a4",  8224 => x"296f00a0",  8225 => x"1423001f",
     8226 => x"c8410800",  8227 => x"f4221000",  8228 => x"c9e37800",
     8229 => x"c9e27800",  8230 => x"2962001c",  8231 => x"296e0024",
     8232 => x"1443001f",  8233 => x"c8221000",  8234 => x"f4410800",
     8235 => x"c9e37800",  8236 => x"c9e17800",  8237 => x"29610020",
     8238 => x"1423001f",  8239 => x"c8410800",  8240 => x"f4221000",
     8241 => x"c9e37800",  8242 => x"15c3001f",  8243 => x"c82e7000",
     8244 => x"c9e27800",  8245 => x"f5c10800",  8246 => x"c9e37800",
     8247 => x"78020001",  8248 => x"c9e17800",  8249 => x"38424d90",
     8250 => x"34010087",  8251 => x"f800074e",  8252 => x"b9c01000",
     8253 => x"b9e00800",  8254 => x"fbfffd4b",  8255 => x"b8201800",
     8256 => x"b9a01000",  8257 => x"34010007",  8258 => x"f8000747",
     8259 => x"78020001",  8260 => x"34010087",  8261 => x"38424dac",
     8262 => x"f8000743",  8263 => x"296300ec",  8264 => x"34010007",
     8265 => x"b9801000",  8266 => x"f800073f",  8267 => x"78020001",
     8268 => x"34010087",  8269 => x"38424dc8",  8270 => x"f800073b",
     8271 => x"296300a8",  8272 => x"34010007",  8273 => x"b9801000",
     8274 => x"f8000737",  8275 => x"78020001",  8276 => x"34010087",
     8277 => x"38424de4",  8278 => x"f8000733",  8279 => x"296300e4",
     8280 => x"34010007",  8281 => x"b9801000",  8282 => x"f800072f",
     8283 => x"78020001",  8284 => x"34010087",  8285 => x"38424e00",
     8286 => x"f800072b",  8287 => x"296300b8",  8288 => x"78020001",
     8289 => x"34010007",  8290 => x"38424e1c",  8291 => x"f8000726",
     8292 => x"78010001",  8293 => x"38214e24",  8294 => x"f8001152",
     8295 => x"340d0001",  8296 => x"b9a00800",  8297 => x"2b9d0004",
     8298 => x"2b8b0018",  8299 => x"2b8c0014",  8300 => x"2b8d0010",
     8301 => x"2b8e000c",  8302 => x"2b8f0008",  8303 => x"379c0110",
     8304 => x"c3a00000",  8305 => x"379cfff4",  8306 => x"5b8b0008",
     8307 => x"5b9d0004",  8308 => x"b8205800",  8309 => x"fbffe306",
     8310 => x"34020003",  8311 => x"5c220003",  8312 => x"34010002",
     8313 => x"e0000002",  8314 => x"34010001",  8315 => x"59610028",
     8316 => x"3562004c",  8317 => x"35610048",  8318 => x"f80012b5",
     8319 => x"34010000",  8320 => x"59600040",  8321 => x"59600044",
     8322 => x"59600088",  8323 => x"5960008c",  8324 => x"3782000c",
     8325 => x"34030000",  8326 => x"f80027be",  8327 => x"44200006",
     8328 => x"2b81000c",  8329 => x"596100a0",  8330 => x"34010001",
     8331 => x"596100a4",  8332 => x"e0000003",  8333 => x"596000a0",
     8334 => x"596000a4",  8335 => x"34010000",  8336 => x"f800127b",
     8337 => x"5961002c",  8338 => x"34010001",  8339 => x"59610054",
     8340 => x"59610050",  8341 => x"34010000",  8342 => x"f8002749",
     8343 => x"59610034",  8344 => x"34011f40",  8345 => x"596100b4",
     8346 => x"78010001",  8347 => x"382160a0",  8348 => x"28210000",
     8349 => x"596100b8",  8350 => x"596100bc",  8351 => x"35610014",
     8352 => x"f8001220",  8353 => x"34010000",  8354 => x"5960001c",
     8355 => x"2b9d0004",  8356 => x"2b8b0008",  8357 => x"379c000c",
     8358 => x"c3a00000",  8359 => x"c3a00000",  8360 => x"379cfffc",
     8361 => x"5b9d0004",  8362 => x"b8201000",  8363 => x"78010001",
     8364 => x"38214e38",  8365 => x"f800110b",  8366 => x"2b9d0004",
     8367 => x"379c0004",  8368 => x"c3a00000",  8369 => x"379cffcc",
     8370 => x"5b8b0010",  8371 => x"5b8c000c",  8372 => x"5b8d0008",
     8373 => x"5b9d0004",  8374 => x"378b0014",  8375 => x"34020000",
     8376 => x"34030024",  8377 => x"b9600800",  8378 => x"f8002b75",
     8379 => x"78030001",  8380 => x"b9600800",  8381 => x"34040000",
     8382 => x"34020000",  8383 => x"38637a80",  8384 => x"34080020",
     8385 => x"34070008",  8386 => x"e0000004",  8387 => x"34840001",
     8388 => x"34210004",  8389 => x"44870017",  8390 => x"b4432800",
     8391 => x"e0000004",  8392 => x"30a00000",  8393 => x"34420001",
     8394 => x"34a50001",  8395 => x"40a60000",  8396 => x"44c8fffc",
     8397 => x"44c0000d",  8398 => x"b4432800",  8399 => x"58250000",
     8400 => x"e0000002",  8401 => x"34420001",  8402 => x"b4432800",
     8403 => x"40a50000",  8404 => x"7ca90000",  8405 => x"7ca60020",
     8406 => x"a1263000",  8407 => x"5cc0fffa",  8408 => x"5ca6ffeb",
     8409 => x"e0000003",  8410 => x"340c0000",  8411 => x"448c0021",
     8412 => x"2b810014",  8413 => x"340c0000",  8414 => x"40220000",
     8415 => x"34010023",  8416 => x"4441001c",  8417 => x"780b0001",
     8418 => x"780c0001",  8419 => x"396b7298",  8420 => x"398c7350",
     8421 => x"e0000011",  8422 => x"29610000",  8423 => x"f8002b89",
     8424 => x"b8206800",  8425 => x"5c20000c",  8426 => x"29620004",
     8427 => x"37810018",  8428 => x"d8400000",  8429 => x"b8206000",
     8430 => x"4c2d000e",  8431 => x"29620000",  8432 => x"78010001",
     8433 => x"b9801800",  8434 => x"38214e40",  8435 => x"f80010c5",
     8436 => x"e0000008",  8437 => x"356b0008",  8438 => x"2b820014",
     8439 => x"558bffef",  8440 => x"78010001",  8441 => x"38214e58",
     8442 => x"f80010be",  8443 => x"340cffea",  8444 => x"b9800800",
     8445 => x"2b9d0004",  8446 => x"2b8b0010",  8447 => x"2b8c000c",
     8448 => x"2b8d0008",  8449 => x"379c0034",  8450 => x"c3a00000",
     8451 => x"379cfff8",  8452 => x"5b8b0008",  8453 => x"5b9d0004",
     8454 => x"780b0001",  8455 => x"396b7ad4",  8456 => x"29650000",
     8457 => x"78020001",  8458 => x"34240001",  8459 => x"b8201800",
     8460 => x"38427a80",  8461 => x"b4220800",  8462 => x"c8a31800",
     8463 => x"b4821000",  8464 => x"f8002ada",  8465 => x"29610000",
     8466 => x"3421ffff",  8467 => x"59610000",  8468 => x"2b9d0004",
     8469 => x"2b8b0008",  8470 => x"379c0008",  8471 => x"c3a00000",
     8472 => x"78010001",  8473 => x"38217adc",  8474 => x"58200000",
     8475 => x"78010001",  8476 => x"38217ad4",  8477 => x"58200000",
     8478 => x"78010001",  8479 => x"38217ad8",  8480 => x"58200000",
     8481 => x"c3a00000",  8482 => x"379cfff4",  8483 => x"5b8b000c",
     8484 => x"5b8c0008",  8485 => x"5b9d0004",  8486 => x"780b0001",
     8487 => x"396b7ad8",  8488 => x"29610000",  8489 => x"340c0001",
     8490 => x"442c0010",  8491 => x"34020002",  8492 => x"4422009d",
     8493 => x"34020000",  8494 => x"5c2000a5",  8495 => x"78010001",
     8496 => x"38214e74",  8497 => x"f8001087",  8498 => x"78010001",
     8499 => x"38217adc",  8500 => x"58200000",  8501 => x"78010001",
     8502 => x"38217ad4",  8503 => x"58200000",  8504 => x"596c0000",
     8505 => x"e000008e",  8506 => x"f80020e6",  8507 => x"34020000",
     8508 => x"48010097",  8509 => x"3402001b",  8510 => x"44220008",
     8511 => x"78020001",  8512 => x"38427ae0",  8513 => x"28430000",
     8514 => x"6424005b",  8515 => x"00650010",  8516 => x"a0a42000",
     8517 => x"44800006",  8518 => x"78010001",  8519 => x"38217ae0",
     8520 => x"78020001",  8521 => x"58220000",  8522 => x"e0000003",
     8523 => x"b8230800",  8524 => x"58410000",  8525 => x"78010001",
     8526 => x"38217ae0",  8527 => x"282b0000",  8528 => x"34020001",
     8529 => x"216100ff",  8530 => x"44200081",  8531 => x"3401007e",
     8532 => x"4561002e",  8533 => x"49610006",  8534 => x"34010009",
     8535 => x"4561006d",  8536 => x"3401000d",  8537 => x"5d610042",
     8538 => x"e0000020",  8539 => x"78020001",  8540 => x"38425984",
     8541 => x"28410000",  8542 => x"45610010",  8543 => x"78020001",
     8544 => x"38425988",  8545 => x"28410000",  8546 => x"45610004",
     8547 => x"3401007f",  8548 => x"5d610037",  8549 => x"e0000027",
     8550 => x"78010001",  8551 => x"38217adc",  8552 => x"28220000",
     8553 => x"4c02005b",  8554 => x"3442ffff",  8555 => x"58220000",
     8556 => x"34010044",  8557 => x"e000000b",  8558 => x"78010001",
     8559 => x"78020001",  8560 => x"38217adc",  8561 => x"38427ad4",
     8562 => x"28230000",  8563 => x"28420000",  8564 => x"4c620050",
     8565 => x"34630001",  8566 => x"58230000",  8567 => x"34010043",
     8568 => x"fbffff30",  8569 => x"e000004b",  8570 => x"78010001",
     8571 => x"38214cd8",  8572 => x"f800103c",  8573 => x"78010001",
     8574 => x"38217ad8",  8575 => x"34020002",  8576 => x"58220000",
     8577 => x"e0000043",  8578 => x"78010001",  8579 => x"78020001",
     8580 => x"38217adc",  8581 => x"38427ad4",  8582 => x"28210000",
     8583 => x"28420000",  8584 => x"4422003c",  8585 => x"fbffff7a",
     8586 => x"34010050",  8587 => x"e3ffffed",  8588 => x"780b0001",
     8589 => x"396b7adc",  8590 => x"29610000",  8591 => x"4c010035",
     8592 => x"34010044",  8593 => x"fbffff17",  8594 => x"34010050",
     8595 => x"fbffff15",  8596 => x"29610000",  8597 => x"3421ffff",
     8598 => x"fbffff6d",  8599 => x"29610000",  8600 => x"3421ffff",
     8601 => x"59610000",  8602 => x"e000002a",  8603 => x"78010001",
     8604 => x"a1610800",  8605 => x"5c200027",  8606 => x"78010001",
     8607 => x"38217ad4",  8608 => x"28240000",  8609 => x"3401004f",
     8610 => x"48810022",  8611 => x"78010001",  8612 => x"38217adc",
     8613 => x"28230000",  8614 => x"44640008",  8615 => x"78020001",
     8616 => x"34610001",  8617 => x"38427a80",  8618 => x"b4220800",
     8619 => x"b4621000",  8620 => x"c8831800",  8621 => x"f8002a3d",
     8622 => x"78010001",  8623 => x"38217adc",  8624 => x"28230000",
     8625 => x"78020001",  8626 => x"38427a80",  8627 => x"b4431000",
     8628 => x"304b0000",  8629 => x"34620001",  8630 => x"58220000",
     8631 => x"78010001",  8632 => x"38217ad4",  8633 => x"28220000",
     8634 => x"34420001",  8635 => x"58220000",  8636 => x"34010040",
     8637 => x"fbfffeeb",  8638 => x"78020001",  8639 => x"38427ae0",
     8640 => x"28420000",  8641 => x"78010001",  8642 => x"38214e7c",
     8643 => x"f8000ff5",  8644 => x"78010001",  8645 => x"38217ae0",
     8646 => x"58200000",  8647 => x"34020001",  8648 => x"e000000b",
     8649 => x"78020001",  8650 => x"38427ad4",  8651 => x"28420000",
     8652 => x"78010001",  8653 => x"38217a80",  8654 => x"b4220800",
     8655 => x"30200000",  8656 => x"fbfffee1",  8657 => x"59600000",
     8658 => x"e3fffff5",  8659 => x"b8400800",  8660 => x"2b9d0004",
     8661 => x"2b8b000c",  8662 => x"2b8c0008",  8663 => x"379c000c",
     8664 => x"c3a00000",  8665 => x"34030000",  8666 => x"34070009",
     8667 => x"34050005",  8668 => x"e0000014",  8669 => x"3486ffd0",
     8670 => x"20c800ff",  8671 => x"55070004",  8672 => x"3c630004",
     8673 => x"b4c31800",  8674 => x"e000000d",  8675 => x"3486ffbf",
     8676 => x"20c600ff",  8677 => x"54c50004",  8678 => x"3c630004",
     8679 => x"3484ffc9",  8680 => x"e0000006",  8681 => x"3486ff9f",
     8682 => x"20c600ff",  8683 => x"54c50007",  8684 => x"3c630004",
     8685 => x"3484ffa9",  8686 => x"b4831800",  8687 => x"34210001",
     8688 => x"40240000",  8689 => x"5c80ffec",  8690 => x"58430000",
     8691 => x"c3a00000",  8692 => x"34030000",  8693 => x"34050009",
     8694 => x"e0000007",  8695 => x"3484ffd0",  8696 => x"208600ff",
     8697 => x"54c50006",  8698 => x"0863000a",  8699 => x"34210001",
     8700 => x"b4831800",  8701 => x"40240000",  8702 => x"5c80fff9",
     8703 => x"58430000",  8704 => x"c3a00000",  8705 => x"379cffec",
     8706 => x"5b8b0014",  8707 => x"5b8c0010",  8708 => x"5b8d000c",
     8709 => x"5b8e0008",  8710 => x"5b9d0004",  8711 => x"78010001",
     8712 => x"38218eb4",  8713 => x"40210000",  8714 => x"4420001b",
     8715 => x"780b0001",  8716 => x"780e0001",  8717 => x"780d0001",
     8718 => x"340c0000",  8719 => x"396b7a80",  8720 => x"39ce7ad4",
     8721 => x"39ad4e98",  8722 => x"b9600800",  8723 => x"34020050",
     8724 => x"b9801800",  8725 => x"f8001bfc",  8726 => x"59c10000",
     8727 => x"48200006",  8728 => x"5d80000d",  8729 => x"78010001",
     8730 => x"38214e80",  8731 => x"f8000f9d",  8732 => x"e0000009",
     8733 => x"b5610800",  8734 => x"3020ffff",  8735 => x"b9601000",
     8736 => x"b9a00800",  8737 => x"f8000f97",  8738 => x"fbfffe8f",
     8739 => x"340c0001",  8740 => x"e3ffffee",  8741 => x"2b9d0004",
     8742 => x"2b8b0014",  8743 => x"2b8c0010",  8744 => x"2b8d000c",
     8745 => x"2b8e0008",  8746 => x"379c0014",  8747 => x"c3a00000",
     8748 => x"379cfff8",  8749 => x"5b8b0008",  8750 => x"5b9d0004",
     8751 => x"78010001",  8752 => x"38219260",  8753 => x"28210000",
     8754 => x"78030001",  8755 => x"38636088",  8756 => x"28620000",
     8757 => x"282b000c",  8758 => x"78030001",  8759 => x"78010001",
     8760 => x"38634ec0",  8761 => x"38214ea8",  8762 => x"f8000f7e",
     8763 => x"78050001",  8764 => x"78030001",  8765 => x"78040001",
     8766 => x"38a5608c",  8767 => x"38636090",  8768 => x"38846094",
     8769 => x"28a20000",  8770 => x"28630000",  8771 => x"28840000",
     8772 => x"78010001",  8773 => x"38214ee0",  8774 => x"f8000f72",
     8775 => x"216b000f",  8776 => x"356b0001",  8777 => x"78010001",
     8778 => x"34020080",  8779 => x"3d6b0004",  8780 => x"38214ef4",
     8781 => x"34030800",  8782 => x"f8000f6a",  8783 => x"3561ff80",
     8784 => x"3402000f",  8785 => x"50410006",  8786 => x"78010001",
     8787 => x"38214f1c",  8788 => x"b9601000",  8789 => x"35630010",
     8790 => x"f8000f62",  8791 => x"34010000",  8792 => x"2b9d0004",
     8793 => x"2b8b0008",  8794 => x"379c0008",  8795 => x"c3a00000",
     8796 => x"379cfff8",  8797 => x"5b8b0008",  8798 => x"5b9d0004",
     8799 => x"b8205800",  8800 => x"28210000",  8801 => x"78020001",
     8802 => x"38424f4c",  8803 => x"f8002a0d",  8804 => x"5c200003",
     8805 => x"fbffe11a",  8806 => x"e0000008",  8807 => x"29610000",
     8808 => x"78020001",  8809 => x"38424f54",  8810 => x"f8002a06",
     8811 => x"3402ffea",  8812 => x"5c200003",  8813 => x"fbffe138",
     8814 => x"b8201000",  8815 => x"b8400800",  8816 => x"2b9d0004",
     8817 => x"2b8b0008",  8818 => x"379c0008",  8819 => x"c3a00000",
     8820 => x"379cfff8",  8821 => x"5b8b0008",  8822 => x"5b9d0004",
     8823 => x"b8205800",  8824 => x"28210000",  8825 => x"78020001",
     8826 => x"38424f5c",  8827 => x"f80029f5",  8828 => x"34020001",
     8829 => x"44200018",  8830 => x"29610000",  8831 => x"78020001",
     8832 => x"38424314",  8833 => x"f80029ef",  8834 => x"34020002",
     8835 => x"44200012",  8836 => x"29610000",  8837 => x"78020001",
     8838 => x"38423e2c",  8839 => x"f80029e9",  8840 => x"34020003",
     8841 => x"4420000c",  8842 => x"fbffe0f1",  8843 => x"3c210002",
     8844 => x"78020001",  8845 => x"38425c68",  8846 => x"b4411000",
     8847 => x"28420000",  8848 => x"78010001",  8849 => x"38214818",
     8850 => x"f8000f26",  8851 => x"34010000",  8852 => x"e0000003",
     8853 => x"b8400800",  8854 => x"fbffe135",  8855 => x"2b9d0004",
     8856 => x"2b8b0008",  8857 => x"379c0008",  8858 => x"c3a00000",
     8859 => x"379cfff0",  8860 => x"5b8b0010",  8861 => x"5b8c000c",
     8862 => x"5b8d0008",  8863 => x"5b9d0004",  8864 => x"78010001",
     8865 => x"38214f74",  8866 => x"780b0001",  8867 => x"780d0001",
     8868 => x"780c0001",  8869 => x"f8000f13",  8870 => x"396b7298",
     8871 => x"39ad7350",  8872 => x"398c4f8c",  8873 => x"e0000005",
     8874 => x"29620000",  8875 => x"b9800800",  8876 => x"356b0008",
     8877 => x"f8000f0b",  8878 => x"55abfffc",  8879 => x"34010000",
     8880 => x"2b9d0004",  8881 => x"2b8b0010",  8882 => x"2b8c000c",
     8883 => x"2b8d0008",  8884 => x"379c0010",  8885 => x"c3a00000",
     8886 => x"379cffec",  8887 => x"5b8b0010",  8888 => x"5b8c000c",
     8889 => x"5b8d0008",  8890 => x"5b9d0004",  8891 => x"340b0000",
     8892 => x"b8406800",  8893 => x"340c0006",  8894 => x"37820014",
     8895 => x"fbffff1a",  8896 => x"2b830014",  8897 => x"b5ab1000",
     8898 => x"356b0001",  8899 => x"30430000",  8900 => x"40220000",
     8901 => x"6442003a",  8902 => x"b4220800",  8903 => x"5d6cfff7",
     8904 => x"2b9d0004",  8905 => x"2b8b0010",  8906 => x"2b8c000c",
     8907 => x"2b8d0008",  8908 => x"379c0014",  8909 => x"c3a00000",
     8910 => x"379cfff8",  8911 => x"5b8b0008",  8912 => x"5b9d0004",
     8913 => x"b8404000",  8914 => x"41030000",  8915 => x"41040001",
     8916 => x"41050002",  8917 => x"41060003",  8918 => x"41070004",
     8919 => x"41080005",  8920 => x"78020001",  8921 => x"38424f9c",
     8922 => x"b8205800",  8923 => x"f8000ecf",  8924 => x"b9600800",
     8925 => x"2b9d0004",  8926 => x"2b8b0008",  8927 => x"379c0008",
     8928 => x"c3a00000",  8929 => x"379cffd0",  8930 => x"5b8b0008",
     8931 => x"5b9d0004",  8932 => x"b8205800",  8933 => x"28210000",
     8934 => x"44200005",  8935 => x"78020001",  8936 => x"38424fbc",
     8937 => x"f8002987",  8938 => x"5c200004",  8939 => x"3781002c",
     8940 => x"f8000fd4",  8941 => x"e000002b",  8942 => x"29610000",
     8943 => x"78020001",  8944 => x"38424fc0",  8945 => x"f800297f",
     8946 => x"5c200008",  8947 => x"378b002c",  8948 => x"b9600800",
     8949 => x"f8000fcb",  8950 => x"b9601000",  8951 => x"34010000",
     8952 => x"f8001b74",  8953 => x"e000001f",  8954 => x"29610000",
     8955 => x"78020001",  8956 => x"38424fc8",  8957 => x"f8002973",
     8958 => x"5c20000b",  8959 => x"29630004",  8960 => x"44610009",
     8961 => x"378b002c",  8962 => x"b8600800",  8963 => x"b9601000",
     8964 => x"fbffffb2",  8965 => x"b9600800",  8966 => x"f8000fa6",
     8967 => x"f80010a1",  8968 => x"e0000010",  8969 => x"29610000",
     8970 => x"78020001",  8971 => x"38424fcc",  8972 => x"f8002964",
     8973 => x"b8201800",  8974 => x"3402ffea",  8975 => x"5c200011",
     8976 => x"29610004",  8977 => x"4423000f",  8978 => x"378b002c",
     8979 => x"b9601000",  8980 => x"fbffffa2",  8981 => x"34010000",
     8982 => x"b9601000",  8983 => x"f8001b4c",  8984 => x"3782002c",
     8985 => x"3781000c",  8986 => x"fbffffb4",  8987 => x"b8201000",
     8988 => x"78010001",  8989 => x"38214fd4",  8990 => x"f8000e9a",
     8991 => x"34020000",  8992 => x"b8400800",  8993 => x"2b9d0004",
     8994 => x"2b8b0008",  8995 => x"379c0030",  8996 => x"c3a00000",
     8997 => x"379cffe8",  8998 => x"5b8b0018",  8999 => x"5b8c0014",
     9000 => x"5b8d0010",  9001 => x"5b8e000c",  9002 => x"5b8f0008",
     9003 => x"5b9d0004",  9004 => x"28210000",  9005 => x"44200010",
     9006 => x"78020001",  9007 => x"38424fec",  9008 => x"f8002940",
     9009 => x"5c20000c",  9010 => x"78010001",  9011 => x"78020001",
     9012 => x"3821735c",  9013 => x"384274ac",  9014 => x"e0000005",
     9015 => x"58200018",  9016 => x"58200014",  9017 => x"58200010",
     9018 => x"3421001c",  9019 => x"5441fffc",  9020 => x"e0000018",
     9021 => x"78010001",  9022 => x"38214ff4",  9023 => x"780b0001",
     9024 => x"780d0001",  9025 => x"780c0001",  9026 => x"f8000e76",
     9027 => x"396b735c",  9028 => x"39ad74ac",  9029 => x"398c501c",
     9030 => x"e000000d",  9031 => x"29610018",  9032 => x"340203e8",
     9033 => x"296f0010",  9034 => x"f8002806",  9035 => x"296e0014",
     9036 => x"29650000",  9037 => x"b8202000",  9038 => x"b9e01000",
     9039 => x"b9800800",  9040 => x"b9c01800",  9041 => x"f8000e67",
     9042 => x"356b001c",  9043 => x"55abfff4",  9044 => x"34010000",
     9045 => x"2b9d0004",  9046 => x"2b8b0018",  9047 => x"2b8c0014",
     9048 => x"2b8d0010",  9049 => x"2b8e000c",  9050 => x"2b8f0008",
     9051 => x"379c0018",  9052 => x"c3a00000",  9053 => x"379cfff8",
     9054 => x"5b9d0004",  9055 => x"b8201000",  9056 => x"28210000",
     9057 => x"4420000d",  9058 => x"28420004",  9059 => x"5c40000b",
     9060 => x"37820008",  9061 => x"fbfffe8f",  9062 => x"2b820008",
     9063 => x"78010001",  9064 => x"38216098",  9065 => x"084203e8",
     9066 => x"58220000",  9067 => x"78010001",  9068 => x"38214cd8",
     9069 => x"e0000003",  9070 => x"78010001",  9071 => x"3821503c",
     9072 => x"f8000e48",  9073 => x"34010000",  9074 => x"2b9d0004",
     9075 => x"379c0008",  9076 => x"c3a00000",  9077 => x"379cfff8",
     9078 => x"5b8b0008",  9079 => x"5b9d0004",  9080 => x"b8205800",
     9081 => x"28210000",  9082 => x"5c200011",  9083 => x"78010001",
     9084 => x"38219248",  9085 => x"28220000",  9086 => x"340b0000",
     9087 => x"64420000",  9088 => x"58220000",  9089 => x"78010001",
     9090 => x"38218ee4",  9091 => x"28230000",  9092 => x"3463ffff",
     9093 => x"58230000",  9094 => x"5c4b002b",  9095 => x"78010001",
     9096 => x"38215060",  9097 => x"f8000e2f",  9098 => x"e0000027",
     9099 => x"78020001",  9100 => x"38425074",  9101 => x"f80028e3",
     9102 => x"5c200007",  9103 => x"f8000f9a",  9104 => x"b8201000",
     9105 => x"78010001",  9106 => x"382156bc",  9107 => x"f8000e25",
     9108 => x"e000001c",  9109 => x"29610000",  9110 => x"78020001",
     9111 => x"38423ecc",  9112 => x"f80028d8",  9113 => x"5c20000b",
     9114 => x"78010001",  9115 => x"38219248",  9116 => x"34020001",
     9117 => x"58220000",  9118 => x"78010001",  9119 => x"38218ee4",
     9120 => x"28220000",  9121 => x"3442ffff",  9122 => x"58220000",
     9123 => x"e000000d",  9124 => x"29610000",  9125 => x"78020001",
     9126 => x"38425078",  9127 => x"f80028c9",  9128 => x"340bffea",
     9129 => x"5c200008",  9130 => x"78010001",  9131 => x"38219248",
     9132 => x"58200000",  9133 => x"78010001",  9134 => x"38215060",
     9135 => x"f8000e09",  9136 => x"340b0000",  9137 => x"b9600800",
     9138 => x"2b9d0004",  9139 => x"2b8b0008",  9140 => x"379c0008",
     9141 => x"c3a00000",  9142 => x"379cffb8",  9143 => x"5b8b0028",
     9144 => x"5b8c0024",  9145 => x"5b8d0020",  9146 => x"5b8e001c",
     9147 => x"5b8f0018",  9148 => x"5b900014",  9149 => x"5b910010",
     9150 => x"5b92000c",  9151 => x"5b930008",  9152 => x"5b9d0004",
     9153 => x"b8205800",  9154 => x"28210000",  9155 => x"442000c8",
     9156 => x"78020001",  9157 => x"38425098",  9158 => x"f80028aa",
     9159 => x"5c200008",  9160 => x"f8001852",  9161 => x"3403ffff",
     9162 => x"34020000",  9163 => x"5c2300c4",  9164 => x"78010001",
     9165 => x"382150a0",  9166 => x"e000003c",  9167 => x"29610010",
     9168 => x"44200045",  9169 => x"29610000",  9170 => x"78020001",
     9171 => x"384250b4",  9172 => x"f800289c",  9173 => x"5c200040",
     9174 => x"29610004",  9175 => x"34020010",  9176 => x"356c0004",
     9177 => x"f80029bb",  9178 => x"3c210018",  9179 => x"34030000",
     9180 => x"14210018",  9181 => x"3784002c",  9182 => x"e0000007",
     9183 => x"29820000",  9184 => x"b4832800",  9185 => x"b4431000",
     9186 => x"40420000",  9187 => x"34630001",  9188 => x"30a20000",
     9189 => x"b0601000",  9190 => x"4822fff9",  9191 => x"b4820800",
     9192 => x"34030020",  9193 => x"3404000f",  9194 => x"e0000005",
     9195 => x"34420001",  9196 => x"30230000",  9197 => x"b0401000",
     9198 => x"34210001",  9199 => x"4c82fffc",  9200 => x"29610008",
     9201 => x"f80003e6",  9202 => x"5b810040",  9203 => x"2961000c",
     9204 => x"f80003e3",  9205 => x"5b810044",  9206 => x"29610010",
     9207 => x"f80003e0",  9208 => x"5b81003c",  9209 => x"34020001",
     9210 => x"3781002c",  9211 => x"34030000",  9212 => x"f8001837",
     9213 => x"3c220018",  9214 => x"3401fffe",  9215 => x"14420018",
     9216 => x"5c410006",  9217 => x"78010001",  9218 => x"382150b8",
     9219 => x"f8000db5",  9220 => x"3402ffe4",  9221 => x"e000008a",
     9222 => x"3401ffff",  9223 => x"5c410006",  9224 => x"78010001",
     9225 => x"382150c8",  9226 => x"f8000dae",  9227 => x"3402fffb",
     9228 => x"e0000083",  9229 => x"4c400004",  9230 => x"78010001",
     9231 => x"382150d4",  9232 => x"e0000023",  9233 => x"78010001",
     9234 => x"382150f0",  9235 => x"f8000da5",  9236 => x"e0000075",
     9237 => x"29610000",  9238 => x"78020001",  9239 => x"38425100",
     9240 => x"f8002858",  9241 => x"5c200030",  9242 => x"78100001",
     9243 => x"780f0001",  9244 => x"780e0001",  9245 => x"340c0000",
     9246 => x"34110000",  9247 => x"3792002c",  9248 => x"3a10511c",
     9249 => x"3793003c",  9250 => x"39ef4e7c",  9251 => x"39ce5124",
     9252 => x"ba400800",  9253 => x"34020000",  9254 => x"b9801800",
     9255 => x"f800180c",  9256 => x"3c2b0018",  9257 => x"156b0018",
     9258 => x"5d600005",  9259 => x"78010001",  9260 => x"38215108",
     9261 => x"f8000d8b",  9262 => x"e000005b",  9263 => x"4d600007",
     9264 => x"78010001",  9265 => x"382150d4",  9266 => x"b9601000",
     9267 => x"f8000d85",  9268 => x"3402fff2",  9269 => x"e000005a",
     9270 => x"358c0001",  9271 => x"ba000800",  9272 => x"b9801000",
     9273 => x"f8000d7f",  9274 => x"ba406800",  9275 => x"41a20000",
     9276 => x"b9e00800",  9277 => x"35ad0001",  9278 => x"f8000d7a",
     9279 => x"5db3fffc",  9280 => x"2b820040",  9281 => x"2b830044",
     9282 => x"2b84003c",  9283 => x"36310001",  9284 => x"b9c00800",
     9285 => x"b2208800",  9286 => x"f8000d72",  9287 => x"4971ffdd",
     9288 => x"e0000041",  9289 => x"29610000",  9290 => x"78020001",
     9291 => x"38425144",  9292 => x"f8002824",  9293 => x"5c200032",
     9294 => x"f8001385",  9295 => x"3c2c0018",  9296 => x"3401ffed",
     9297 => x"158c0018",  9298 => x"5d810006",  9299 => x"78010001",
     9300 => x"3821514c",  9301 => x"f8000d63",  9302 => x"3402ffed",
     9303 => x"e0000038",  9304 => x"780b0001",  9305 => x"396b8eec",
     9306 => x"780d0001",  9307 => x"3401fffb",  9308 => x"356e0010",
     9309 => x"39ad4e7c",  9310 => x"5d810004",  9311 => x"78010001",
     9312 => x"38215158",  9313 => x"e3ffffa9",  9314 => x"41620000",
     9315 => x"b9a00800",  9316 => x"356b0001",  9317 => x"f8000d53",
     9318 => x"5d6efffc",  9319 => x"78010001",  9320 => x"38214cd8",
     9321 => x"f8000d4f",  9322 => x"3401fffa",  9323 => x"5d810006",
     9324 => x"78010001",  9325 => x"38215168",  9326 => x"f8000d4a",
     9327 => x"3402fffa",  9328 => x"e000001f",  9329 => x"78020001",
     9330 => x"78030001",  9331 => x"78040001",  9332 => x"38428e80",
     9333 => x"38638e84",  9334 => x"38846f2c",  9335 => x"28420000",
     9336 => x"28630000",  9337 => x"28840000",  9338 => x"78010001",
     9339 => x"38215180",  9340 => x"f8000d3c",  9341 => x"b9801000",
     9342 => x"e0000011",  9343 => x"29610004",  9344 => x"4420000b",
     9345 => x"29610000",  9346 => x"78020001",  9347 => x"384251a8",
     9348 => x"f80027ec",  9349 => x"5c200006",  9350 => x"29610004",
     9351 => x"f8000350",  9352 => x"f8000eee",  9353 => x"34020000",
     9354 => x"e0000005",  9355 => x"78010001",  9356 => x"38215084",
     9357 => x"f8000d2b",  9358 => x"3402ffea",  9359 => x"b8400800",
     9360 => x"2b9d0004",  9361 => x"2b8b0028",  9362 => x"2b8c0024",
     9363 => x"2b8d0020",  9364 => x"2b8e001c",  9365 => x"2b8f0018",
     9366 => x"2b900014",  9367 => x"2b910010",  9368 => x"2b92000c",
     9369 => x"2b930008",  9370 => x"379c0048",  9371 => x"c3a00000",
     9372 => x"379cffe8",  9373 => x"5b8b0010",  9374 => x"5b8c000c",
     9375 => x"5b8d0008",  9376 => x"5b9d0004",  9377 => x"b8205800",
     9378 => x"28210000",  9379 => x"78020001",  9380 => x"384251b0",
     9381 => x"f80027cb",  9382 => x"5c200011",  9383 => x"2963000c",
     9384 => x"3402ffea",  9385 => x"44610086",  9386 => x"29610004",
     9387 => x"f800032c",  9388 => x"b8206800",  9389 => x"29610008",
     9390 => x"f8000329",  9391 => x"b8206000",  9392 => x"2961000c",
     9393 => x"f8000326",  9394 => x"b8201800",  9395 => x"b9801000",
     9396 => x"b9a00800",  9397 => x"f8002260",  9398 => x"e0000078",
     9399 => x"29610000",  9400 => x"78020001",  9401 => x"384251b8",
     9402 => x"f80027b6",  9403 => x"b8201800",  9404 => x"5c200007",
     9405 => x"29610004",  9406 => x"3402ffea",  9407 => x"44230070",
     9408 => x"f8000317",  9409 => x"f800231e",  9410 => x"e0000060",
     9411 => x"29610000",  9412 => x"78020001",  9413 => x"3842507c",
     9414 => x"f80027aa",  9415 => x"5c200003",  9416 => x"f80023b1",
     9417 => x"e0000065",  9418 => x"29610000",  9419 => x"78020001",
     9420 => x"384251bc",  9421 => x"f80027a3",  9422 => x"5c20000d",
     9423 => x"29630008",  9424 => x"3402ffea",  9425 => x"4461005e",
     9426 => x"29610004",  9427 => x"f8000304",  9428 => x"b8206000",
     9429 => x"29610008",  9430 => x"f8000301",  9431 => x"b8201000",
     9432 => x"b9800800",  9433 => x"f8002317",  9434 => x"e0000054",
     9435 => x"29610000",  9436 => x"78020001",  9437 => x"384251c0",
     9438 => x"f8002792",  9439 => x"b8201800",  9440 => x"5c20000e",
     9441 => x"29610004",  9442 => x"3402ffea",  9443 => x"4423004c",
     9444 => x"f80002f3",  9445 => x"37820018",  9446 => x"37830014",
     9447 => x"f8002331",  9448 => x"2b820018",  9449 => x"2b830014",
     9450 => x"78010001",  9451 => x"382151c4",  9452 => x"f8000ccc",
     9453 => x"e0000041",  9454 => x"29610000",  9455 => x"78020001",
     9456 => x"38424f4c",  9457 => x"f800277f",  9458 => x"b8201800",
     9459 => x"5c200007",  9460 => x"29610004",  9461 => x"3402ffea",
     9462 => x"44230039",  9463 => x"f80002e0",  9464 => x"f80022c9",
     9465 => x"e0000035",  9466 => x"29610000",  9467 => x"78020001",
     9468 => x"38424f54",  9469 => x"f8002773",  9470 => x"b8201800",
     9471 => x"5c200007",  9472 => x"29610004",  9473 => x"3402ffea",
     9474 => x"4423002d",  9475 => x"f80002d4",  9476 => x"f80022ce",
     9477 => x"e0000029",  9478 => x"29610000",  9479 => x"78020001",
     9480 => x"384251cc",  9481 => x"f8002767",  9482 => x"5c20000d",
     9483 => x"29630008",  9484 => x"3402ffea",  9485 => x"44610022",
     9486 => x"29610004",  9487 => x"f80002c8",  9488 => x"b8206000",
     9489 => x"29610008",  9490 => x"f80002c5",  9491 => x"b8201000",
     9492 => x"b9800800",  9493 => x"f80023d4",  9494 => x"e0000018",
     9495 => x"29610000",  9496 => x"78020001",  9497 => x"384251d4",
     9498 => x"f8002756",  9499 => x"b8201800",  9500 => x"5c20000b",
     9501 => x"29610004",  9502 => x"3402ffea",  9503 => x"44230010",
     9504 => x"f80002b7",  9505 => x"f80023b9",  9506 => x"b8201000",
     9507 => x"78010001",  9508 => x"38214e54",  9509 => x"f8000c93",
     9510 => x"e0000008",  9511 => x"29610000",  9512 => x"78020001",
     9513 => x"384251dc",  9514 => x"f8002746",  9515 => x"3402ffea",
     9516 => x"5c200003",  9517 => x"f800246b",  9518 => x"34020000",
     9519 => x"b8400800",  9520 => x"2b9d0004",  9521 => x"2b8b0010",
     9522 => x"2b8c000c",  9523 => x"2b8d0008",  9524 => x"379c0018",
     9525 => x"c3a00000",  9526 => x"379cfff0",  9527 => x"5b8b000c",
     9528 => x"5b8c0008",  9529 => x"5b9d0004",  9530 => x"b8205800",
     9531 => x"28210000",  9532 => x"4420000b",  9533 => x"78020001",
     9534 => x"384251ec",  9535 => x"f8002731",  9536 => x"b8206000",
     9537 => x"5c200006",  9538 => x"37810010",  9539 => x"f80013db",
     9540 => x"340bffff",  9541 => x"49810021",  9542 => x"e000001c",
     9543 => x"29610000",  9544 => x"340b0000",  9545 => x"5c20001d",
     9546 => x"37810010",  9547 => x"34020000",  9548 => x"f80017c0",
     9549 => x"4d61000a",  9550 => x"2b820010",  9551 => x"78010001",
     9552 => x"382151f4",  9553 => x"f8000c67",  9554 => x"2b820010",
     9555 => x"78010001",  9556 => x"382160a0",  9557 => x"58220000",
     9558 => x"e0000010",  9559 => x"78010001",  9560 => x"3821521c",
     9561 => x"f8000c5f",  9562 => x"37810010",  9563 => x"f80013c3",
     9564 => x"340bffff",  9565 => x"48010009",  9566 => x"2b820010",
     9567 => x"78010001",  9568 => x"382160a0",  9569 => x"58220000",
     9570 => x"37810010",  9571 => x"34020001",  9572 => x"f80017a8",
     9573 => x"b8205800",  9574 => x"b9600800",  9575 => x"2b9d0004",
     9576 => x"2b8b000c",  9577 => x"2b8c0008",  9578 => x"379c0010",
     9579 => x"c3a00000",  9580 => x"379cffe8",  9581 => x"5b8b000c",
     9582 => x"5b8c0008",  9583 => x"5b9d0004",  9584 => x"b8205800",
     9585 => x"37820018",  9586 => x"37810010",  9587 => x"f80015c6",
     9588 => x"29610008",  9589 => x"44200014",  9590 => x"29610000",
     9591 => x"78020001",  9592 => x"38424fc8",  9593 => x"f80026f7",
     9594 => x"5c20000f",  9595 => x"fbffde00",  9596 => x"34030003",
     9597 => x"3402fff0",  9598 => x"44230040",  9599 => x"29610004",
     9600 => x"f8000257",  9601 => x"b8206000",  9602 => x"29610008",
     9603 => x"f8000254",  9604 => x"b8201800",  9605 => x"b9801000",
     9606 => x"1581001f",  9607 => x"34040003",  9608 => x"e0000020",
     9609 => x"29610000",  9610 => x"4420000f",  9611 => x"78020001",
     9612 => x"38425250",  9613 => x"f80026e3",  9614 => x"5c20000b",
     9615 => x"fbffddec",  9616 => x"34020003",  9617 => x"44220023",
     9618 => x"29610004",  9619 => x"f8000244",  9620 => x"b8201000",
     9621 => x"34030000",  9622 => x"1421001f",  9623 => x"34040001",
     9624 => x"e0000010",  9625 => x"29610000",  9626 => x"44200010",
     9627 => x"78020001",  9628 => x"38425258",  9629 => x"f80026d3",
     9630 => x"5c20000c",  9631 => x"fbffdddc",  9632 => x"34020003",
     9633 => x"44220013",  9634 => x"29610004",  9635 => x"f8000234",
     9636 => x"b8201800",  9637 => x"34020000",  9638 => x"34010000",
     9639 => x"34040002",  9640 => x"f8001571",  9641 => x"e0000014",
     9642 => x"29610000",  9643 => x"44200009",  9644 => x"78020001",
     9645 => x"38425260",  9646 => x"f80026c2",  9647 => x"5c200005",
     9648 => x"78010001",  9649 => x"382151c4",  9650 => x"2b820014",
     9651 => x"e0000008",  9652 => x"2b820014",  9653 => x"2b810010",
     9654 => x"34030000",  9655 => x"f8000121",  9656 => x"b8201000",
     9657 => x"78010001",  9658 => x"38215264",  9659 => x"2b830018",
     9660 => x"f8000bfc",  9661 => x"34020000",  9662 => x"b8400800",
     9663 => x"2b9d0004",  9664 => x"2b8b000c",  9665 => x"2b8c0008",
     9666 => x"379c0018",  9667 => x"c3a00000",  9668 => x"78010001",
     9669 => x"382174b0",  9670 => x"34020001",  9671 => x"58220000",
     9672 => x"34010000",  9673 => x"c3a00000",  9674 => x"379cfffc",
     9675 => x"5b9d0004",  9676 => x"f800123b",  9677 => x"34010000",
     9678 => x"2b9d0004",  9679 => x"379c0004",  9680 => x"c3a00000",
     9681 => x"379cfff8",  9682 => x"5b8b0008",  9683 => x"5b9d0004",
     9684 => x"b8205800",  9685 => x"28210000",  9686 => x"4420000c",
     9687 => x"78020001",  9688 => x"38425294",  9689 => x"f8002697",
     9690 => x"5c200008",  9691 => x"34010001",  9692 => x"fbffe890",
     9693 => x"78010001",  9694 => x"3821609c",  9695 => x"34020001",
     9696 => x"58220000",  9697 => x"e000000b",  9698 => x"29610000",
     9699 => x"44200009",  9700 => x"78020001",  9701 => x"3842529c",
     9702 => x"f800268a",  9703 => x"5c200005",  9704 => x"fbffe884",
     9705 => x"78010001",  9706 => x"3821609c",  9707 => x"58200000",
     9708 => x"78010001",  9709 => x"3821609c",  9710 => x"28210000",
     9711 => x"78020001",  9712 => x"38425290",  9713 => x"44200003",
     9714 => x"78020001",  9715 => x"3842528c",  9716 => x"78010001",
     9717 => x"382152a4",  9718 => x"f8000bc2",  9719 => x"34010000",
     9720 => x"2b9d0004",  9721 => x"2b8b0008",  9722 => x"379c0008",
     9723 => x"c3a00000",  9724 => x"379cfff8",  9725 => x"5b8b0008",
     9726 => x"5b9d0004",  9727 => x"b8205800",  9728 => x"28210000",
     9729 => x"78020001",  9730 => x"384251b0",  9731 => x"f800266d",
     9732 => x"5c200003",  9733 => x"f8001384",  9734 => x"e000001d",
     9735 => x"29610000",  9736 => x"78020001",  9737 => x"384252c0",
     9738 => x"f8002666",  9739 => x"5c200003",  9740 => x"f8001388",
     9741 => x"e0000016",  9742 => x"29610000",  9743 => x"78020001",
     9744 => x"384252c8",  9745 => x"f800265f",  9746 => x"5c200003",
     9747 => x"f8001387",  9748 => x"e000000f",  9749 => x"29610000",
     9750 => x"78020001",  9751 => x"384252cc",  9752 => x"f8002658",
     9753 => x"5c200003",  9754 => x"f8001386",  9755 => x"e0000008",
     9756 => x"29610000",  9757 => x"78020001",  9758 => x"38424f4c",
     9759 => x"f8002651",  9760 => x"3402ffea",  9761 => x"5c200003",
     9762 => x"f8001384",  9763 => x"34020000",  9764 => x"b8400800",
     9765 => x"2b9d0004",  9766 => x"2b8b0008",  9767 => x"379c0008",
     9768 => x"c3a00000",  9769 => x"379cffec",  9770 => x"5b8b0010",
     9771 => x"5b8c000c",  9772 => x"5b8d0008",  9773 => x"5b9d0004",
     9774 => x"340b0000",  9775 => x"b8406800",  9776 => x"340c0004",
     9777 => x"37820014",  9778 => x"fbfffbc2",  9779 => x"2b830014",
     9780 => x"b5ab1000",  9781 => x"356b0001",  9782 => x"30430000",
     9783 => x"40220000",  9784 => x"6442002e",  9785 => x"b4220800",
     9786 => x"5d6cfff7",  9787 => x"2b9d0004",  9788 => x"2b8b0010",
     9789 => x"2b8c000c",  9790 => x"2b8d0008",  9791 => x"379c0014",
     9792 => x"c3a00000",  9793 => x"379cfff8",  9794 => x"5b8b0008",
     9795 => x"5b9d0004",  9796 => x"b8403000",  9797 => x"40c30000",
     9798 => x"40c40001",  9799 => x"40c50002",  9800 => x"40c60003",
     9801 => x"78020001",  9802 => x"384252d4",  9803 => x"b8205800",
     9804 => x"f8000b5e",  9805 => x"b9600800",  9806 => x"2b9d0004",
     9807 => x"2b8b0008",  9808 => x"379c0008",  9809 => x"c3a00000",
     9810 => x"379cffe0",  9811 => x"5b8b0008",  9812 => x"5b9d0004",
     9813 => x"b8205800",  9814 => x"28210000",  9815 => x"44200005",
     9816 => x"78020001",  9817 => x"38424fbc",  9818 => x"f8002616",
     9819 => x"5c200004",  9820 => x"37810020",  9821 => x"f80004bb",
     9822 => x"e0000012",  9823 => x"29610000",  9824 => x"78020001",
     9825 => x"38424fc8",  9826 => x"f800260e",  9827 => x"b8201800",
     9828 => x"3402ffea",  9829 => x"5c200024",  9830 => x"29610004",
     9831 => x"44230022",  9832 => x"78020001",  9833 => x"38427d48",
     9834 => x"34030002",  9835 => x"58430000",  9836 => x"37820020",
     9837 => x"fbffffbc",  9838 => x"37810020",  9839 => x"f80004b2",
     9840 => x"378b000c",  9841 => x"37820020",  9842 => x"b9600800",
     9843 => x"fbffffce",  9844 => x"78010001",  9845 => x"38217d48",
     9846 => x"28210000",  9847 => x"34020001",  9848 => x"44220009",
     9849 => x"44200004",  9850 => x"34020002",  9851 => x"5c22000d",
     9852 => x"e0000008",  9853 => x"78010001",  9854 => x"382152e0",
     9855 => x"f8000b39",  9856 => x"e0000008",  9857 => x"78010001",
     9858 => x"382152fc",  9859 => x"e0000003",  9860 => x"78010001",
     9861 => x"3821531c",  9862 => x"b9601000",  9863 => x"f8000b31",
     9864 => x"34020000",  9865 => x"b8400800",  9866 => x"2b9d0004",
     9867 => x"2b8b0008",  9868 => x"379c0020",  9869 => x"c3a00000",
     9870 => x"379cfffc",  9871 => x"5b9d0004",  9872 => x"28210000",
     9873 => x"44200005",  9874 => x"fbffdbf2",  9875 => x"78020001",
     9876 => x"384274c4",  9877 => x"58410000",  9878 => x"78020001",
     9879 => x"384274c4",  9880 => x"28420000",  9881 => x"78010001",
     9882 => x"38215344",  9883 => x"f8000b1d",  9884 => x"34010000",
     9885 => x"2b9d0004",  9886 => x"379c0004",  9887 => x"c3a00000",
     9888 => x"379cfff4",  9889 => x"5b8b000c",  9890 => x"5b8c0008",
     9891 => x"5b9d0004",  9892 => x"b8205800",  9893 => x"28210000",
     9894 => x"4420000b",  9895 => x"78020001",  9896 => x"38425098",
     9897 => x"f80025c7",  9898 => x"b8206000",  9899 => x"5c200006",
     9900 => x"f8001695",  9901 => x"4c2c0025",  9902 => x"78010001",
     9903 => x"38215364",  9904 => x"e000000e",  9905 => x"29610004",
     9906 => x"44200011",  9907 => x"29610000",  9908 => x"78020001",
     9909 => x"384250b4",  9910 => x"f80025ba",  9911 => x"b8206000",
     9912 => x"5c20000b",  9913 => x"b9600800",  9914 => x"f800169c",
     9915 => x"4c2c0005",  9916 => x"78010001",  9917 => x"38215384",
     9918 => x"f8000afa",  9919 => x"e0000013",  9920 => x"78010001",
     9921 => x"382153a0",  9922 => x"e3fffffc",  9923 => x"29610000",
     9924 => x"44200007",  9925 => x"78020001",  9926 => x"38425100",
     9927 => x"f80025a9",  9928 => x"5c200003",  9929 => x"f8001707",
     9930 => x"e0000008",  9931 => x"29610000",  9932 => x"44200006",
     9933 => x"78020001",  9934 => x"384253a8",  9935 => x"f80025a1",
     9936 => x"5c200002",  9937 => x"fbfffb30",  9938 => x"34010000",
     9939 => x"2b9d0004",  9940 => x"2b8b000c",  9941 => x"2b8c0008",
     9942 => x"379c000c",  9943 => x"c3a00000",  9944 => x"379cffd0",
     9945 => x"5b8b0030",  9946 => x"5b8c002c",  9947 => x"5b8d0028",
     9948 => x"5b8e0024",  9949 => x"5b8f0020",  9950 => x"5b90001c",
     9951 => x"5b910018",  9952 => x"5b920014",  9953 => x"5b930010",
     9954 => x"5b94000c",  9955 => x"5b9d0008",  9956 => x"b8609000",
     9957 => x"78030001",  9958 => x"3863598c",  9959 => x"b8406000",
     9960 => x"b8400800",  9961 => x"28620000",  9962 => x"f8002476",
     9963 => x"78030001",  9964 => x"3863598c",  9965 => x"28620000",
     9966 => x"b8205800",  9967 => x"b9800800",  9968 => x"f8002460",
     9969 => x"b820a000",  9970 => x"3402003c",  9971 => x"b9600800",
     9972 => x"f800246c",  9973 => x"34020e10",  9974 => x"b8207800",
     9975 => x"b9600800",  9976 => x"f8002468",  9977 => x"3402003c",
     9978 => x"f8002456",  9979 => x"b8208000",  9980 => x"34020e10",
     9981 => x"b9600800",  9982 => x"f8002452",  9983 => x"b8208800",
     9984 => x"ba807000",  9985 => x"340b07b2",  9986 => x"e000000f",
     9987 => x"3402016d",  9988 => x"5d80000b",  9989 => x"34020064",
     9990 => x"b9600800",  9991 => x"f8002429",  9992 => x"3402016e",
     9993 => x"5c2c0006",  9994 => x"34020190",  9995 => x"b9600800",
     9996 => x"f8002424",  9997 => x"64220000",  9998 => x"3442016d",
     9999 => x"c9c27000", 10000 => x"356b0001", 10001 => x"216c0003",
    10002 => x"3402016d", 10003 => x"5d80000b", 10004 => x"34020064",
    10005 => x"b9600800", 10006 => x"f800241a", 10007 => x"3402016e",
    10008 => x"5c2c0006", 10009 => x"34020190", 10010 => x"b9600800",
    10011 => x"f8002415", 10012 => x"64220000", 10013 => x"3442016d",
    10014 => x"51c2ffe5", 10015 => x"34020064", 10016 => x"b9600800",
    10017 => x"f800240f", 10018 => x"34020190", 10019 => x"b8209800",
    10020 => x"b9600800", 10021 => x"f800240b", 10022 => x"78020001",
    10023 => x"340d0000", 10024 => x"64250000", 10025 => x"38425c78",
    10026 => x"e000000d", 10027 => x"34040000", 10028 => x"5d800004",
    10029 => x"34040001", 10030 => x"5e6c0002", 10031 => x"b8a02000",
    10032 => x"0884000c", 10033 => x"b48d2000", 10034 => x"3c840002",
    10035 => x"35ad0001", 10036 => x"b4442000", 10037 => x"28810000",
    10038 => x"c9c17000", 10039 => x"34040000", 10040 => x"5d800004",
    10041 => x"34040001", 10042 => x"5e6c0002", 10043 => x"b8a02000",
    10044 => x"0884000c", 10045 => x"b48d2000", 10046 => x"3c840002",
    10047 => x"b4442000", 10048 => x"28810000", 10049 => x"51c1ffea",
    10050 => x"34010001", 10051 => x"35ce0001", 10052 => x"4641001d",
    10053 => x"780c0001", 10054 => x"34010002", 10055 => x"398c7ae4",
    10056 => x"46410028", 10057 => x"36810004", 10058 => x"34020007",
    10059 => x"f8002415", 10060 => x"3c210002", 10061 => x"78130001",
    10062 => x"78020001", 10063 => x"3dad0002", 10064 => x"38425cf4",
    10065 => x"3a735cd8", 10066 => x"b6619800", 10067 => x"b44d6800",
    10068 => x"78120001", 10069 => x"2a630000", 10070 => x"29a40000",
    10071 => x"3a5253b0", 10072 => x"b9800800", 10073 => x"ba401000",
    10074 => x"b9c02800", 10075 => x"b9603000", 10076 => x"ba203800",
    10077 => x"ba004000", 10078 => x"5b8f0004", 10079 => x"f8000a4b",
    10080 => x"e000001a", 10081 => x"78010001", 10082 => x"3dad0002",
    10083 => x"38215cf4", 10084 => x"b42d6800", 10085 => x"29a30000",
    10086 => x"78010001", 10087 => x"78020001", 10088 => x"384253d0",
    10089 => x"b9c02000", 10090 => x"ba202800", 10091 => x"ba003000",
    10092 => x"b9e03800", 10093 => x"38217ae4", 10094 => x"f8000a3c",
    10095 => x"e000000b", 10096 => x"78020001", 10097 => x"b9800800",
    10098 => x"384253e8", 10099 => x"b9601800", 10100 => x"35a40001",
    10101 => x"b9c02800", 10102 => x"ba203000", 10103 => x"ba003800",
    10104 => x"b9e04000", 10105 => x"f8000a31", 10106 => x"78010001",
    10107 => x"38217ae4", 10108 => x"2b9d0008", 10109 => x"2b8b0030",
    10110 => x"2b8c002c", 10111 => x"2b8d0028", 10112 => x"2b8e0024",
    10113 => x"2b8f0020", 10114 => x"2b90001c", 10115 => x"2b910018",
    10116 => x"2b920014", 10117 => x"2b930010", 10118 => x"2b94000c",
    10119 => x"379c0030", 10120 => x"c3a00000", 10121 => x"379cffdc",
    10122 => x"5b8b0008", 10123 => x"5b9d0004", 10124 => x"5b840014",
    10125 => x"20240080", 10126 => x"64840000", 10127 => x"5b830010",
    10128 => x"78030001", 10129 => x"b8204800", 10130 => x"b8600800",
    10131 => x"34030002", 10132 => x"5b82000c", 10133 => x"b8405800",
    10134 => x"38215408", 10135 => x"c8641000", 10136 => x"2123007f",
    10137 => x"5b850018", 10138 => x"5b86001c", 10139 => x"5b870020",
    10140 => x"5b880024", 10141 => x"f8000a1b", 10142 => x"37820010",
    10143 => x"b9600800", 10144 => x"f80009f6", 10145 => x"78010001",
    10146 => x"38215414", 10147 => x"f8000a15", 10148 => x"2b9d0004",
    10149 => x"2b8b0008", 10150 => x"379c0024", 10151 => x"c3a00000",
    10152 => x"379cffe0", 10153 => x"5b8b000c", 10154 => x"5b8c0008",
    10155 => x"5b9d0004", 10156 => x"b8404800", 10157 => x"78020001",
    10158 => x"b8205000", 10159 => x"b8400800", 10160 => x"b8605800",
    10161 => x"b9401000", 10162 => x"b9201800", 10163 => x"38215418",
    10164 => x"b8806000", 10165 => x"5b840010", 10166 => x"5b850014",
    10167 => x"5b860018", 10168 => x"5b87001c", 10169 => x"5b880020",
    10170 => x"f80009fe", 10171 => x"21620080", 10172 => x"78030001",
    10173 => x"64420000", 10174 => x"b8600800", 10175 => x"34030002",
    10176 => x"c8621000", 10177 => x"38215408", 10178 => x"2163007f",
    10179 => x"f80009f5", 10180 => x"37820014", 10181 => x"b9800800",
    10182 => x"f80009d0", 10183 => x"78010001", 10184 => x"38215414",
    10185 => x"f80009ef", 10186 => x"2b9d0004", 10187 => x"2b8b000c",
    10188 => x"2b8c0008", 10189 => x"379c0020", 10190 => x"c3a00000",
    10191 => x"379cfffc", 10192 => x"5b9d0004", 10193 => x"78010001",
    10194 => x"38215424", 10195 => x"f80009e5", 10196 => x"2b9d0004",
    10197 => x"379c0004", 10198 => x"c3a00000", 10199 => x"40240000",
    10200 => x"3402002d", 10201 => x"34030001", 10202 => x"5c820003",
    10203 => x"34210001", 10204 => x"3403ffff", 10205 => x"34020000",
    10206 => x"34050009", 10207 => x"e0000004", 10208 => x"0842000a",
    10209 => x"34210001", 10210 => x"b4821000", 10211 => x"40240000",
    10212 => x"3484ffd0", 10213 => x"208600ff", 10214 => x"50a6fffa",
    10215 => x"88430800", 10216 => x"c3a00000", 10217 => x"379cfff4",
    10218 => x"5b8b000c", 10219 => x"5b8c0008", 10220 => x"5b9d0004",
    10221 => x"b8206000", 10222 => x"f8000f8a", 10223 => x"342b0001",
    10224 => x"f8000f88", 10225 => x"5c2bffff", 10226 => x"b9800800",
    10227 => x"e0000002", 10228 => x"3421ffff", 10229 => x"4820ffff",
    10230 => x"f8000f82", 10231 => x"c82b0800", 10232 => x"2b9d0004",
    10233 => x"2b8b000c", 10234 => x"2b8c0008", 10235 => x"379c000c",
    10236 => x"c3a00000", 10237 => x"379cfff0", 10238 => x"5b8b0010",
    10239 => x"5b8c000c", 10240 => x"5b8d0008", 10241 => x"5b9d0004",
    10242 => x"340b0400", 10243 => x"340c0400", 10244 => x"e0000003",
    10245 => x"b58b6000", 10246 => x"3d6b0001", 10247 => x"b9800800",
    10248 => x"fbffffe1", 10249 => x"4420fffc", 10250 => x"158c0001",
    10251 => x"156b0002", 10252 => x"e0000009", 10253 => x"b56c6800",
    10254 => x"b9a00800", 10255 => x"fbffffda", 10256 => x"5c200002",
    10257 => x"b9a06000", 10258 => x"0161001f", 10259 => x"b42b5800",
    10260 => x"156b0001", 10261 => x"5d60fff8", 10262 => x"78010001",
    10263 => x"38217b24", 10264 => x"582c0000", 10265 => x"78010001",
    10266 => x"b9801000", 10267 => x"3821547c", 10268 => x"f800099c",
    10269 => x"2b9d0004", 10270 => x"2b8b0010", 10271 => x"2b8c000c",
    10272 => x"2b8d0008", 10273 => x"379c0010", 10274 => x"c3a00000",
    10275 => x"379cfffc", 10276 => x"5b9d0004", 10277 => x"78020001",
    10278 => x"38427b24", 10279 => x"28430000", 10280 => x"34042710",
    10281 => x"0865000a", 10282 => x"e0000004", 10283 => x"3442ffff",
    10284 => x"4840ffff", 10285 => x"3421d8f0", 10286 => x"50810003",
    10287 => x"b8a01000", 10288 => x"e3fffffc", 10289 => x"88230800",
    10290 => x"340203e8", 10291 => x"f800231d", 10292 => x"e0000002",
    10293 => x"3421ffff", 10294 => x"4820ffff", 10295 => x"34010000",
    10296 => x"2b9d0004", 10297 => x"379c0004", 10298 => x"c3a00000",
    10299 => x"b8202800", 10300 => x"5c800002", 10301 => x"b8602000",
    10302 => x"b8803000", 10303 => x"50640002", 10304 => x"b8603000",
    10305 => x"b4260800", 10306 => x"e000000e", 10307 => x"2c460002",
    10308 => x"2847000c", 10309 => x"b4e63800", 10310 => x"40e60000",
    10311 => x"30a60000", 10312 => x"2c470002", 10313 => x"2c460006",
    10314 => x"34a50001", 10315 => x"34e70001", 10316 => x"20e7ffff",
    10317 => x"0c470002", 10318 => x"5cc70002", 10319 => x"0c400002",
    10320 => x"5ca1fff3", 10321 => x"5083000b", 10322 => x"2c410002",
    10323 => x"b4610800", 10324 => x"c8242000", 10325 => x"0c440002",
    10326 => x"2c410006", 10327 => x"e0000003", 10328 => x"c8812000",
    10329 => x"0c440002", 10330 => x"2c440002", 10331 => x"5481fffd",
    10332 => x"b8600800", 10333 => x"c3a00000", 10334 => x"b4432800",
    10335 => x"e000000d", 10336 => x"2c240000", 10337 => x"2826000c",
    10338 => x"40470000", 10339 => x"34420001", 10340 => x"b4c43000",
    10341 => x"30c70000", 10342 => x"34840001", 10343 => x"2c260006",
    10344 => x"2084ffff", 10345 => x"0c240000", 10346 => x"5cc40002",
    10347 => x"0c200000", 10348 => x"5c45fff4", 10349 => x"b8600800",
    10350 => x"c3a00000", 10351 => x"379cffc8", 10352 => x"5b8b001c",
    10353 => x"5b8c0018", 10354 => x"5b8d0014", 10355 => x"5b8e0010",
    10356 => x"5b8f000c", 10357 => x"5b900008", 10358 => x"5b9d0004",
    10359 => x"780b0001", 10360 => x"780c0001", 10361 => x"396b7d38",
    10362 => x"398c7b58", 10363 => x"b9600800", 10364 => x"b9801000",
    10365 => x"340301e0", 10366 => x"37840020", 10367 => x"f8000d94",
    10368 => x"b8206800", 10369 => x"340f0000", 10370 => x"4c010061",
    10371 => x"2d62000c", 10372 => x"0f800038", 10373 => x"38018100",
    10374 => x"5c41000e", 10375 => x"b9801000", 10376 => x"34030002",
    10377 => x"37810038", 10378 => x"f8002327", 10379 => x"78010001",
    10380 => x"78020001", 10381 => x"38217d44", 10382 => x"38427b5a",
    10383 => x"34030002", 10384 => x"780c0001", 10385 => x"f8002320",
    10386 => x"35adfffc", 10387 => x"398c7b5c", 10388 => x"78010001",
    10389 => x"2f820038", 10390 => x"382174b4", 10391 => x"28210000",
    10392 => x"20420fff", 10393 => x"340f0000", 10394 => x"5c410049",
    10395 => x"41820000", 10396 => x"34010045", 10397 => x"34030000",
    10398 => x"5c410008", 10399 => x"41820009", 10400 => x"34010011",
    10401 => x"5c410005", 10402 => x"41830016", 10403 => x"41810017",
    10404 => x"3c630008", 10405 => x"b8611800", 10406 => x"78010001",
    10407 => x"78020001", 10408 => x"38217d38", 10409 => x"38427b28",
    10410 => x"2c27000c", 10411 => x"34460030", 10412 => x"34040000",
    10413 => x"340b0000", 10414 => x"e000000c", 10415 => x"28410000",
    10416 => x"44200009", 10417 => x"2c25000c", 10418 => x"5ca70007",
    10419 => x"2c25000e", 10420 => x"5c600003", 10421 => x"44a30038",
    10422 => x"e0000003", 10423 => x"5ca30002", 10424 => x"b8202000",
    10425 => x"34420004", 10426 => x"5c46fff5", 10427 => x"44800002",
    10428 => x"b8805800", 10429 => x"340f0001", 10430 => x"45600025",
    10431 => x"2d700028", 10432 => x"35a10028", 10433 => x"48300022",
    10434 => x"356e0024", 10435 => x"3782003a", 10436 => x"34030002",
    10437 => x"b9c00800", 10438 => x"0f8d003a", 10439 => x"fbffff97",
    10440 => x"ca016800", 10441 => x"21adffff", 10442 => x"0d6d0028",
    10443 => x"37820020", 10444 => x"34030018", 10445 => x"b9c00800",
    10446 => x"fbffff90", 10447 => x"c9a16800", 10448 => x"21adffff",
    10449 => x"78020001", 10450 => x"0d6d0028", 10451 => x"38427d38",
    10452 => x"3403000e", 10453 => x"b9c00800", 10454 => x"fbffff88",
    10455 => x"c9a16800", 10456 => x"2f83003a", 10457 => x"21adffff",
    10458 => x"0d6d0028", 10459 => x"b9c00800", 10460 => x"b9801000",
    10461 => x"fbffff81", 10462 => x"c9a10800", 10463 => x"0d610028",
    10464 => x"2d61002c", 10465 => x"34210001", 10466 => x"0d61002c",
    10467 => x"b9e00800", 10468 => x"2b9d0004", 10469 => x"2b8b001c",
    10470 => x"2b8c0018", 10471 => x"2b8d0014", 10472 => x"2b8e0010",
    10473 => x"2b8f000c", 10474 => x"2b900008", 10475 => x"379c0038",
    10476 => x"c3a00000", 10477 => x"b8205800", 10478 => x"e3ffffcb",
    10479 => x"379cfffc", 10480 => x"5b9d0004", 10481 => x"b8400800",
    10482 => x"f80009ce", 10483 => x"34010000", 10484 => x"2b9d0004",
    10485 => x"379c0004", 10486 => x"c3a00000", 10487 => x"78020001",
    10488 => x"38427b28", 10489 => x"34430030", 10490 => x"e0000004",
    10491 => x"28440000", 10492 => x"34420004", 10493 => x"5881001c",
    10494 => x"5c43fffd", 10495 => x"c3a00000", 10496 => x"379cff24",
    10497 => x"5b8b0014", 10498 => x"5b8c0010", 10499 => x"5b8d000c",
    10500 => x"5b8e0008", 10501 => x"5b9d0004", 10502 => x"78050001",
    10503 => x"b8205800", 10504 => x"b8406000", 10505 => x"b8607000",
    10506 => x"b8806800", 10507 => x"38a57b28", 10508 => x"34010000",
    10509 => x"3402000c", 10510 => x"28a30000", 10511 => x"34a50004",
    10512 => x"5c600009", 10513 => x"3c220002", 10514 => x"78050001",
    10515 => x"38a57b28", 10516 => x"b4a22800", 10517 => x"58ab0000",
    10518 => x"3402000c", 10519 => x"5c22000a", 10520 => x"e0000003",
    10521 => x"34210001", 10522 => x"5c22fff4", 10523 => x"78010001",
    10524 => x"78020001", 10525 => x"38425d24", 10526 => x"38215494",
    10527 => x"f8000899", 10528 => x"e0000020", 10529 => x"78020001",
    10530 => x"37810018", 10531 => x"384254b0", 10532 => x"fbfff74d",
    10533 => x"4801001b", 10534 => x"b9600800", 10535 => x"34020000",
    10536 => x"34030012", 10537 => x"f8002306", 10538 => x"45800005",
    10539 => x"b9600800", 10540 => x"b9801000", 10541 => x"34030012",
    10542 => x"f8002283", 10543 => x"0d60000e", 10544 => x"5dc00004",
    10545 => x"34010800", 10546 => x"0d61000c", 10547 => x"0d6d000e",
    10548 => x"35610012", 10549 => x"f800098b", 10550 => x"2b8100d0",
    10551 => x"0d600026", 10552 => x"0d600024", 10553 => x"5961001c",
    10554 => x"2b8100b8", 10555 => x"0d60002c", 10556 => x"59610020",
    10557 => x"2d61002a", 10558 => x"0d610028", 10559 => x"e0000002",
    10560 => x"340b0000", 10561 => x"b9600800", 10562 => x"2b9d0004",
    10563 => x"2b8b0014", 10564 => x"2b8c0010", 10565 => x"2b8d000c",
    10566 => x"2b8e0008", 10567 => x"379c00dc", 10568 => x"c3a00000",
    10569 => x"78020001", 10570 => x"38427b28", 10571 => x"34430030",
    10572 => x"e0000005", 10573 => x"28440000", 10574 => x"5c810002",
    10575 => x"58400000", 10576 => x"34420004", 10577 => x"5c43fffc",
    10578 => x"34010000", 10579 => x"c3a00000", 10580 => x"379cffe8",
    10581 => x"5b8b0018", 10582 => x"5b8c0014", 10583 => x"5b8d0010",
    10584 => x"5b8e000c", 10585 => x"5b8f0008", 10586 => x"5b9d0004",
    10587 => x"b8205800", 10588 => x"59620010", 10589 => x"b8407000",
    10590 => x"b8807800", 10591 => x"b8a06000", 10592 => x"282d0008",
    10593 => x"44600005", 10594 => x"b8a00800", 10595 => x"3402fc18",
    10596 => x"f800219f", 10597 => x"b42d6800", 10598 => x"c9cf2000",
    10599 => x"b8801800", 10600 => x"4c800002", 10601 => x"b48c1800",
    10602 => x"0181001f", 10603 => x"b42c0800", 10604 => x"14210001",
    10605 => x"b4242000", 10606 => x"4c800002", 10607 => x"b48c2000",
    10608 => x"49840002", 10609 => x"c88c2000", 10610 => x"09820003",
    10611 => x"1445001f", 10612 => x"00a5001e", 10613 => x"b4a21000",
    10614 => x"14420002", 10615 => x"48620006", 10616 => x"1582001f",
    10617 => x"0042001e", 10618 => x"b44c1000", 10619 => x"14420002",
    10620 => x"4c62000d", 10621 => x"b4812000", 10622 => x"596d0008",
    10623 => x"5964000c", 10624 => x"4984000a", 10625 => x"c88c2000",
    10626 => x"5964000c", 10627 => x"b9800800", 10628 => x"340203e8",
    10629 => x"f800217e", 10630 => x"b5a10800", 10631 => x"59610008",
    10632 => x"e0000002", 10633 => x"5963000c", 10634 => x"78030001",
    10635 => x"38635968", 10636 => x"29610008", 10637 => x"28620000",
    10638 => x"4c41000d", 10639 => x"78030001", 10640 => x"3863596c",
    10641 => x"28620000", 10642 => x"29630000", 10643 => x"b4220800",
    10644 => x"29620004", 10645 => x"59610008", 10646 => x"34410001",
    10647 => x"f4411000", 10648 => x"59610004", 10649 => x"b4431000",
    10650 => x"59620000", 10651 => x"2b9d0004", 10652 => x"2b8b0018",
    10653 => x"2b8c0014", 10654 => x"2b8d0010", 10655 => x"2b8e000c",
    10656 => x"2b8f0008", 10657 => x"379c0018", 10658 => x"c3a00000",
    10659 => x"379cffb4", 10660 => x"5b8b0024", 10661 => x"5b8c0020",
    10662 => x"5b8d001c", 10663 => x"5b8e0018", 10664 => x"5b8f0014",
    10665 => x"5b900010", 10666 => x"5b91000c", 10667 => x"5b920008",
    10668 => x"5b9d0004", 10669 => x"b8406800", 10670 => x"2c22002c",
    10671 => x"b8a05800", 10672 => x"b8206000", 10673 => x"b8609000",
    10674 => x"b8807800", 10675 => x"34050000", 10676 => x"44400055",
    10677 => x"342e0024", 10678 => x"2c310028", 10679 => x"3442ffff",
    10680 => x"0c22002c", 10681 => x"34030002", 10682 => x"b9c01000",
    10683 => x"34040000", 10684 => x"3781004e", 10685 => x"fbfffe7e",
    10686 => x"b6218800", 10687 => x"2231ffff", 10688 => x"0d910028",
    10689 => x"b9c01000", 10690 => x"34030018", 10691 => x"34040000",
    10692 => x"37810028", 10693 => x"fbfffe76", 10694 => x"b6218800",
    10695 => x"2231ffff", 10696 => x"37900040", 10697 => x"0d910028",
    10698 => x"b9c01000", 10699 => x"3403000e", 10700 => x"34040000",
    10701 => x"ba000800", 10702 => x"fbfffe6d", 10703 => x"b6218800",
    10704 => x"2f83004e", 10705 => x"2231ffff", 10706 => x"b9c01000",
    10707 => x"b9e02000", 10708 => x"0d910028", 10709 => x"ba400800",
    10710 => x"fbfffe65", 10711 => x"b6210800", 10712 => x"0d810028",
    10713 => x"2f81004c", 10714 => x"78030001", 10715 => x"386374b4",
    10716 => x"0da1000c", 10717 => x"28610000", 10718 => x"37820046",
    10719 => x"34030006", 10720 => x"0da10010", 10721 => x"b9a00800",
    10722 => x"f80021cf", 10723 => x"35a10006", 10724 => x"ba001000",
    10725 => x"34030006", 10726 => x"f80021cb", 10727 => x"4560001e",
    10728 => x"2b810038", 10729 => x"59610014", 10730 => x"2b81002c",
    10731 => x"59610018", 10732 => x"34010000", 10733 => x"f8001eac",
    10734 => x"b8206800", 10735 => x"35620010", 10736 => x"34030000",
    10737 => x"34010000", 10738 => x"f8001e52", 10739 => x"2b810030",
    10740 => x"43820028", 10741 => x"2b83002c", 10742 => x"59610000",
    10743 => x"2b810034", 10744 => x"2984001c", 10745 => x"5960000c",
    10746 => x"59610004", 10747 => x"2b810038", 10748 => x"34051f40",
    10749 => x"59610008", 10750 => x"21a100ff", 10751 => x"64210000",
    10752 => x"a0220800", 10753 => x"29620010", 10754 => x"5961001c",
    10755 => x"b9600800", 10756 => x"fbffff50", 10757 => x"2f81004e",
    10758 => x"b9e02800", 10759 => x"502f0002", 10760 => x"b8202800",
    10761 => x"b8a00800", 10762 => x"2b9d0004", 10763 => x"2b8b0024",
    10764 => x"2b8c0020", 10765 => x"2b8d001c", 10766 => x"2b8e0018",
    10767 => x"2b8f0014", 10768 => x"2b900010", 10769 => x"2b91000c",
    10770 => x"2b920008", 10771 => x"379c004c", 10772 => x"c3a00000",
    10773 => x"379cffc0", 10774 => x"5b8b0014", 10775 => x"5b8c0010",
    10776 => x"5b8d000c", 10777 => x"5b8e0008", 10778 => x"5b9d0004",
    10779 => x"b8206000", 10780 => x"b8607000", 10781 => x"37810030",
    10782 => x"34030006", 10783 => x"b8a05800", 10784 => x"b8806800",
    10785 => x"f8002190", 10786 => x"37810036", 10787 => x"35820012",
    10788 => x"34030006", 10789 => x"f800218c", 10790 => x"78010001",
    10791 => x"382174b4", 10792 => x"28250000", 10793 => x"2d81000c",
    10794 => x"44a00009", 10795 => x"34028100", 10796 => x"0f82003c",
    10797 => x"2d820018", 10798 => x"0f810040", 10799 => x"3c42000d",
    10800 => x"b8452800", 10801 => x"0f85003e", 10802 => x"e0000002",
    10803 => x"0f81003c", 10804 => x"37810030", 10805 => x"b9c01000",
    10806 => x"b9a01800", 10807 => x"37840018", 10808 => x"f8000c86",
    10809 => x"4560000a", 10810 => x"2b820020", 10811 => x"5960000c",
    10812 => x"59620000", 10813 => x"2b820024", 10814 => x"59620004",
    10815 => x"2b820028", 10816 => x"59620008", 10817 => x"43820018",
    10818 => x"5962001c", 10819 => x"2b9d0004", 10820 => x"2b8b0014",
    10821 => x"2b8c0010", 10822 => x"2b8d000c", 10823 => x"2b8e0008",
    10824 => x"379c0040", 10825 => x"c3a00000", 10826 => x"c3a00000",
    10827 => x"379cffe4", 10828 => x"5b8b0008", 10829 => x"5b9d0004",
    10830 => x"78010001", 10831 => x"34020000", 10832 => x"34030000",
    10833 => x"34040044", 10834 => x"382167a4", 10835 => x"fbfffead",
    10836 => x"78020001", 10837 => x"38427d4c", 10838 => x"58410000",
    10839 => x"78010001", 10840 => x"34040025", 10841 => x"34020000",
    10842 => x"34030000", 10843 => x"382167d8", 10844 => x"fbfffea4",
    10845 => x"78020001", 10846 => x"378b000c", 10847 => x"38427d5c",
    10848 => x"58410000", 10849 => x"34030012", 10850 => x"b9600800",
    10851 => x"34020000", 10852 => x"f80021cb", 10853 => x"34010800",
    10854 => x"0f810018", 10855 => x"78010001", 10856 => x"b9601000",
    10857 => x"34030001", 10858 => x"34040000", 10859 => x"3821680c",
    10860 => x"fbfffe94", 10861 => x"78020001", 10862 => x"38427d58",
    10863 => x"58410000", 10864 => x"fbffffda", 10865 => x"2b9d0004",
    10866 => x"2b8b0008", 10867 => x"379c001c", 10868 => x"c3a00000",
    10869 => x"34010000", 10870 => x"c3a00000", 10871 => x"379cfe34",
    10872 => x"5b8b001c", 10873 => x"5b8c0018", 10874 => x"5b8d0014",
    10875 => x"5b8e0010", 10876 => x"5b8f000c", 10877 => x"5b900008",
    10878 => x"5b9d0004", 10879 => x"78010001", 10880 => x"38219258",
    10881 => x"28220000", 10882 => x"34010001", 10883 => x"5c410006",
    10884 => x"78010001", 10885 => x"38217d48", 10886 => x"28230000",
    10887 => x"5c620002", 10888 => x"58200000", 10889 => x"78020001",
    10890 => x"38427d4c", 10891 => x"28410000", 10892 => x"378b0020",
    10893 => x"378201b0", 10894 => x"34040190", 10895 => x"b9601800",
    10896 => x"34050000", 10897 => x"fbffff12", 10898 => x"78040001",
    10899 => x"38847d48", 10900 => x"b8201000", 10901 => x"28810000",
    10902 => x"340c0000", 10903 => x"5c200023", 10904 => x"4c220003",
    10905 => x"b9600800", 10906 => x"f800027a", 10907 => x"f8000cdd",
    10908 => x"78020001", 10909 => x"38427d50", 10910 => x"28430000",
    10911 => x"5c600003", 10912 => x"58410000", 10913 => x"e0000006",
    10914 => x"346303e8", 10915 => x"c8230800", 10916 => x"340c0000",
    10917 => x"48010015", 10918 => x"58430000", 10919 => x"78010001",
    10920 => x"38217d54", 10921 => x"28230000", 10922 => x"378c01b0",
    10923 => x"378b0020", 10924 => x"34630001", 10925 => x"58230000",
    10926 => x"b9601000", 10927 => x"b9800800", 10928 => x"f8000200",
    10929 => x"78050001", 10930 => x"38a57d4c", 10931 => x"b8202000",
    10932 => x"28a10000", 10933 => x"b9801000", 10934 => x"b9601800",
    10935 => x"34050000", 10936 => x"fbffff5d", 10937 => x"340c0001",
    10938 => x"780b0001", 10939 => x"396b7d58", 10940 => x"29610000",
    10941 => x"378e01b0", 10942 => x"378d0020", 10943 => x"34040080",
    10944 => x"b9c01000", 10945 => x"b9a01800", 10946 => x"34050000",
    10947 => x"fbfffee0", 10948 => x"b8202000", 10949 => x"340f0000",
    10950 => x"4c010010", 10951 => x"78030001", 10952 => x"38637d48",
    10953 => x"28610000", 10954 => x"4420000c", 10955 => x"b8801000",
    10956 => x"b9a00800", 10957 => x"f8000108", 10958 => x"b8202000",
    10959 => x"340f0001", 10960 => x"4c010006", 10961 => x"29610000",
    10962 => x"b9c01000", 10963 => x"b9a01800", 10964 => x"34050000",
    10965 => x"fbffff40", 10966 => x"780b0001", 10967 => x"396b7d5c",
    10968 => x"29610000", 10969 => x"379001b0", 10970 => x"378d0020",
    10971 => x"ba001000", 10972 => x"b9a01800", 10973 => x"34040020",
    10974 => x"34050000", 10975 => x"fbfffec4", 10976 => x"340e0000",
    10977 => x"4c010019", 10978 => x"378101c4", 10979 => x"34020000",
    10980 => x"f8001055", 10981 => x"78020001", 10982 => x"38425990",
    10983 => x"28410000", 10984 => x"2b8201c8", 10985 => x"34030004",
    10986 => x"340e0001", 10987 => x"b4410800", 10988 => x"5b8101cc",
    10989 => x"378201cc", 10990 => x"3781003c", 10991 => x"f80020c2",
    10992 => x"b9a00800", 10993 => x"34020020", 10994 => x"34030000",
    10995 => x"f8000143", 10996 => x"29610000", 10997 => x"ba001000",
    10998 => x"b9a01800", 10999 => x"34040020", 11000 => x"34050000",
    11001 => x"fbffff1c", 11002 => x"fbffff7b", 11003 => x"b5ec6000",
    11004 => x"b5810800", 11005 => x"b42e7000", 11006 => x"7dc10000",
    11007 => x"2b9d0004", 11008 => x"2b8b001c", 11009 => x"2b8c0018",
    11010 => x"2b8d0014", 11011 => x"2b8e0010", 11012 => x"2b8f000c",
    11013 => x"2b900008", 11014 => x"379c01cc", 11015 => x"c3a00000",
    11016 => x"34030000", 11017 => x"34040000", 11018 => x"e0000005",
    11019 => x"2c250000", 11020 => x"34840001", 11021 => x"34210002",
    11022 => x"b4651800", 11023 => x"4844fffc", 11024 => x"00610010",
    11025 => x"2063ffff", 11026 => x"b4611800", 11027 => x"00610010",
    11028 => x"b4231800", 11029 => x"a4600800", 11030 => x"2021ffff",
    11031 => x"c3a00000", 11032 => x"379cfffc", 11033 => x"5b9d0004",
    11034 => x"78020001", 11035 => x"38427d60", 11036 => x"34030004",
    11037 => x"f8002094", 11038 => x"2b9d0004", 11039 => x"379c0004",
    11040 => x"c3a00000", 11041 => x"379cfff0", 11042 => x"5b8b0010",
    11043 => x"5b8c000c", 11044 => x"5b8d0008", 11045 => x"5b9d0004",
    11046 => x"78030001", 11047 => x"780b0001", 11048 => x"396b7d60",
    11049 => x"b8206000", 11050 => x"38639270", 11051 => x"286d0000",
    11052 => x"b9600800", 11053 => x"b9801000", 11054 => x"34030004",
    11055 => x"f8002082", 11056 => x"41620000", 11057 => x"41610001",
    11058 => x"3c420018", 11059 => x"3c210010", 11060 => x"b8411000",
    11061 => x"41610003", 11062 => x"b8411000", 11063 => x"41610002",
    11064 => x"3c210008", 11065 => x"b8415800", 11066 => x"29a10018",
    11067 => x"b9800800", 11068 => x"f8000ea7", 11069 => x"5d600004",
    11070 => x"78010001", 11071 => x"38217d48", 11072 => x"58200000",
    11073 => x"78010001", 11074 => x"38217d54", 11075 => x"58200000",
    11076 => x"2b9d0004", 11077 => x"2b8b0010", 11078 => x"2b8c000c",
    11079 => x"2b8d0008", 11080 => x"379c0010", 11081 => x"c3a00000",
    11082 => x"379cfffc", 11083 => x"5b9d0004", 11084 => x"b8201000",
    11085 => x"3401ffff", 11086 => x"44400006", 11087 => x"34410010",
    11088 => x"78020001", 11089 => x"38427d60", 11090 => x"34030004",
    11091 => x"f800203d", 11092 => x"2b9d0004", 11093 => x"379c0004",
    11094 => x"c3a00000", 11095 => x"379cff34", 11096 => x"5b8b0028",
    11097 => x"5b8c0024", 11098 => x"5b8d0020", 11099 => x"5b8e001c",
    11100 => x"5b8f0018", 11101 => x"5b900014", 11102 => x"5b910010",
    11103 => x"5b92000c", 11104 => x"5b930008", 11105 => x"5b9d0004",
    11106 => x"78010001", 11107 => x"38217d48", 11108 => x"28210000",
    11109 => x"340b0000", 11110 => x"44200047", 11111 => x"780c0001",
    11112 => x"398c8044", 11113 => x"29810000", 11114 => x"378f00ac",
    11115 => x"378e002c", 11116 => x"b9e01000", 11117 => x"b9c01800",
    11118 => x"34040080", 11119 => x"34050000", 11120 => x"fbfffe33",
    11121 => x"4c01003c", 11122 => x"3402001b", 11123 => x"340b0001",
    11124 => x"4c410039", 11125 => x"378d00c8", 11126 => x"b9a00800",
    11127 => x"fbffffa1", 11128 => x"43810032", 11129 => x"5c200034",
    11130 => x"43810033", 11131 => x"5c2b0032", 11132 => x"37900044",
    11133 => x"ba000800", 11134 => x"b9a01000", 11135 => x"34030004",
    11136 => x"f8002010", 11137 => x"5c20002c", 11138 => x"379100c0",
    11139 => x"37930034", 11140 => x"ba601000", 11141 => x"34030006",
    11142 => x"ba200800", 11143 => x"f800202a", 11144 => x"3792003a",
    11145 => x"ba401000", 11146 => x"34030004", 11147 => x"378100cc",
    11148 => x"f8002025", 11149 => x"34010008", 11150 => x"3381002e",
    11151 => x"34010006", 11152 => x"33810030", 11153 => x"34010004",
    11154 => x"33810031", 11155 => x"34010002", 11156 => x"33810033",
    11157 => x"ba600800", 11158 => x"3380002c", 11159 => x"338b002d",
    11160 => x"3380002f", 11161 => x"33800032", 11162 => x"f8000726",
    11163 => x"b9a01000", 11164 => x"34030004", 11165 => x"ba400800",
    11166 => x"f8002013", 11167 => x"ba201000", 11168 => x"34030006",
    11169 => x"3781003e", 11170 => x"f800200f", 11171 => x"378200cc",
    11172 => x"34030004", 11173 => x"ba000800", 11174 => x"f800200b",
    11175 => x"29810000", 11176 => x"b9e01000", 11177 => x"b9c01800",
    11178 => x"3404001c", 11179 => x"34050000", 11180 => x"fbfffe69",
    11181 => x"b9600800", 11182 => x"2b9d0004", 11183 => x"2b8b0028",
    11184 => x"2b8c0024", 11185 => x"2b8d0020", 11186 => x"2b8e001c",
    11187 => x"2b8f0018", 11188 => x"2b900014", 11189 => x"2b910010",
    11190 => x"2b92000c", 11191 => x"2b930008", 11192 => x"379c00cc",
    11193 => x"c3a00000", 11194 => x"379cffe4", 11195 => x"5b8b0008",
    11196 => x"5b9d0004", 11197 => x"378b000c", 11198 => x"b9600800",
    11199 => x"34020000", 11200 => x"34030012", 11201 => x"f800206e",
    11202 => x"b9600800", 11203 => x"340200ff", 11204 => x"34030006",
    11205 => x"f800206a", 11206 => x"34010806", 11207 => x"0f810018",
    11208 => x"78010001", 11209 => x"b9601000", 11210 => x"34030001",
    11211 => x"34040000", 11212 => x"38216840", 11213 => x"fbfffd33",
    11214 => x"78020001", 11215 => x"38428044", 11216 => x"58410000",
    11217 => x"2b9d0004", 11218 => x"2b8b0008", 11219 => x"379c001c",
    11220 => x"c3a00000", 11221 => x"379cffe0", 11222 => x"5b8b0018",
    11223 => x"5b8c0014", 11224 => x"5b8d0010", 11225 => x"5b8e000c",
    11226 => x"5b8f0008", 11227 => x"5b9d0004", 11228 => x"378d001c",
    11229 => x"b8205800", 11230 => x"b9a00800", 11231 => x"fbffff39",
    11232 => x"41620000", 11233 => x"34010045", 11234 => x"340c0000",
    11235 => x"5c41004a", 11236 => x"356e0010", 11237 => x"b9a01000",
    11238 => x"b9c00800", 11239 => x"34030004", 11240 => x"f8001fa8",
    11241 => x"b8201000", 11242 => x"5c200043", 11243 => x"41640009",
    11244 => x"34030001", 11245 => x"416d0002", 11246 => x"41610003",
    11247 => x"b8406000", 11248 => x"5c83003d", 11249 => x"41630014",
    11250 => x"34020008", 11251 => x"5c62003a", 11252 => x"3dad0008",
    11253 => x"b9a16800", 11254 => x"35adffe8", 11255 => x"34010040",
    11256 => x"4c2d0002", 11257 => x"340d0040", 11258 => x"356f000c",
    11259 => x"b9e01000", 11260 => x"34030004", 11261 => x"37810020",
    11262 => x"f8001fb3", 11263 => x"35ac0018", 11264 => x"34010045",
    11265 => x"31610000", 11266 => x"15810008", 11267 => x"3782001c",
    11268 => x"31610002", 11269 => x"3401003f", 11270 => x"31610008",
    11271 => x"34010001", 11272 => x"31610009", 11273 => x"34030004",
    11274 => x"31600001", 11275 => x"316c0003", 11276 => x"31600004",
    11277 => x"31600005", 11278 => x"31600006", 11279 => x"31600007",
    11280 => x"3160000a", 11281 => x"3160000b", 11282 => x"b9e00800",
    11283 => x"f8001f9e", 11284 => x"34030004", 11285 => x"37820020",
    11286 => x"b9c00800", 11287 => x"f8001f9a", 11288 => x"35ad0005",
    11289 => x"01a1001f", 11290 => x"31600014", 11291 => x"b42d6800",
    11292 => x"15a20001", 11293 => x"31600015", 11294 => x"31600016",
    11295 => x"31600017", 11296 => x"35610014", 11297 => x"fbfffee7",
    11298 => x"2021ffff", 11299 => x"00220008", 11300 => x"31610017",
    11301 => x"31620016", 11302 => x"b9600800", 11303 => x"3402000a",
    11304 => x"fbfffee0", 11305 => x"2021ffff", 11306 => x"00220008",
    11307 => x"3161000b", 11308 => x"3162000a", 11309 => x"b9800800",
    11310 => x"2b9d0004", 11311 => x"2b8b0018", 11312 => x"2b8c0014",
    11313 => x"2b8d0010", 11314 => x"2b8e000c", 11315 => x"2b8f0008",
    11316 => x"379c0020", 11317 => x"c3a00000", 11318 => x"379cffcc",
    11319 => x"5b8b0028", 11320 => x"5b8c0024", 11321 => x"5b8d0020",
    11322 => x"5b8e001c", 11323 => x"5b8f0018", 11324 => x"5b900014",
    11325 => x"5b910010", 11326 => x"5b92000c", 11327 => x"5b930008",
    11328 => x"5b9d0004", 11329 => x"b8205800", 11330 => x"b8406800",
    11331 => x"b8606000", 11332 => x"5c600012", 11333 => x"3562000c",
    11334 => x"34030004", 11335 => x"37810030", 11336 => x"f8001f69",
    11337 => x"378c002c", 11338 => x"35620010", 11339 => x"34030004",
    11340 => x"b9800800", 11341 => x"f8001f64", 11342 => x"35620014",
    11343 => x"34030002", 11344 => x"37810036", 11345 => x"f8001f60",
    11346 => x"37810034", 11347 => x"35620016", 11348 => x"34030002",
    11349 => x"f8001f5c", 11350 => x"35700008", 11351 => x"b9801000",
    11352 => x"34030004", 11353 => x"ba000800", 11354 => x"f8001f57",
    11355 => x"35b1ffec", 11356 => x"356f000c", 11357 => x"358e0004",
    11358 => x"b9c01000", 11359 => x"34030004", 11360 => x"16320008",
    11361 => x"b9e00800", 11362 => x"f8001f4f", 11363 => x"34010011",
    11364 => x"225200ff", 11365 => x"223100ff", 11366 => x"31610011",
    11367 => x"35820008", 11368 => x"34030002", 11369 => x"31600010",
    11370 => x"31720012", 11371 => x"31710013", 11372 => x"35610014",
    11373 => x"f8001f44", 11374 => x"34030002", 11375 => x"3582000a",
    11376 => x"35610016", 11377 => x"f8001f40", 11378 => x"b56d0800",
    11379 => x"31720018", 11380 => x"31710019", 11381 => x"3160001a",
    11382 => x"3160001b", 11383 => x"35a2fff9", 11384 => x"30200000",
    11385 => x"0041001f", 11386 => x"35730010", 11387 => x"b4221000",
    11388 => x"14420001", 11389 => x"ba000800", 11390 => x"fbfffe8a",
    11391 => x"2023ffff", 11392 => x"5c600002", 11393 => x"3803ffff",
    11394 => x"00610008", 11395 => x"3163001b", 11396 => x"3161001a",
    11397 => x"34010045", 11398 => x"31610000", 11399 => x"15a10008",
    11400 => x"b9801000", 11401 => x"31610002", 11402 => x"3401003f",
    11403 => x"31610008", 11404 => x"34010011", 11405 => x"31610009",
    11406 => x"31600001", 11407 => x"316d0003", 11408 => x"31600004",
    11409 => x"31600005", 11410 => x"31600006", 11411 => x"31600007",
    11412 => x"3160000a", 11413 => x"3160000b", 11414 => x"b9e00800",
    11415 => x"34030004", 11416 => x"f8001f19", 11417 => x"b9c01000",
    11418 => x"34030004", 11419 => x"ba600800", 11420 => x"f8001f15",
    11421 => x"b9600800", 11422 => x"3402000a", 11423 => x"fbfffe69",
    11424 => x"2021ffff", 11425 => x"00220008", 11426 => x"3161000b",
    11427 => x"3162000a", 11428 => x"2b9d0004", 11429 => x"2b8b0028",
    11430 => x"2b8c0024", 11431 => x"2b8d0020", 11432 => x"2b8e001c",
    11433 => x"2b8f0018", 11434 => x"2b900014", 11435 => x"2b910010",
    11436 => x"2b92000c", 11437 => x"2b930008", 11438 => x"379c0034",
    11439 => x"c3a00000", 11440 => x"379cffe4", 11441 => x"5b8b0010",
    11442 => x"5b8c000c", 11443 => x"5b8d0008", 11444 => x"5b9d0004",
    11445 => x"b8405800", 11446 => x"b8206800", 11447 => x"34020001",
    11448 => x"34010006", 11449 => x"3162001c", 11450 => x"3162001d",
    11451 => x"3161001e", 11452 => x"3160001f", 11453 => x"35610020",
    11454 => x"b8606000", 11455 => x"f8000601", 11456 => x"41620024",
    11457 => x"41610020", 11458 => x"34030002", 11459 => x"98410800",
    11460 => x"31610020", 11461 => x"41620025", 11462 => x"41610021",
    11463 => x"316c0025", 11464 => x"98410800", 11465 => x"31610021",
    11466 => x"41610022", 11467 => x"15820008", 11468 => x"98410800",
    11469 => x"31610022", 11470 => x"41610023", 11471 => x"31620024",
    11472 => x"34020000", 11473 => x"982c0800", 11474 => x"31610023",
    11475 => x"35610026", 11476 => x"f8001f5b", 11477 => x"35610028",
    11478 => x"34020000", 11479 => x"34030004", 11480 => x"f8001f57",
    11481 => x"3561002c", 11482 => x"34020000", 11483 => x"34030004",
    11484 => x"f8001f53", 11485 => x"35610030", 11486 => x"34020000",
    11487 => x"34030004", 11488 => x"f8001f4f", 11489 => x"35610034",
    11490 => x"34020000", 11491 => x"34030004", 11492 => x"f8001f4b",
    11493 => x"356c0038", 11494 => x"34020000", 11495 => x"34030010",
    11496 => x"b9800800", 11497 => x"f8001f46", 11498 => x"b9800800",
    11499 => x"f80005d5", 11500 => x"35610048", 11501 => x"34020000",
    11502 => x"34030040", 11503 => x"f8001f40", 11504 => x"35610088",
    11505 => x"34020000", 11506 => x"34030080", 11507 => x"f8001f3c",
    11508 => x"35610108", 11509 => x"34020000", 11510 => x"34030040",
    11511 => x"f8001f38", 11512 => x"378c0014", 11513 => x"b9800800",
    11514 => x"34020000", 11515 => x"34030004", 11516 => x"f8001f33",
    11517 => x"37810018", 11518 => x"340200ff", 11519 => x"34030004",
    11520 => x"f8001f2f", 11521 => x"34010044", 11522 => x"0f81001c",
    11523 => x"34010043", 11524 => x"0f81001e", 11525 => x"b9801800",
    11526 => x"b9600800", 11527 => x"34020148", 11528 => x"fbffff2e",
    11529 => x"b9a00800", 11530 => x"340200ff", 11531 => x"34030006",
    11532 => x"f8001f23", 11533 => x"34010148", 11534 => x"2b9d0004",
    11535 => x"2b8b0010", 11536 => x"2b8c000c", 11537 => x"2b8d0008",
    11538 => x"379c001c", 11539 => x"c3a00000", 11540 => x"379cffe0",
    11541 => x"5b8b0014", 11542 => x"5b8c0010", 11543 => x"5b8d000c",
    11544 => x"5b8e0008", 11545 => x"5b9d0004", 11546 => x"378d0018",
    11547 => x"b8205800", 11548 => x"b9a00800", 11549 => x"b8407000",
    11550 => x"f80005a2", 11551 => x"34010148", 11552 => x"340c0000",
    11553 => x"5dc1001b", 11554 => x"41610014", 11555 => x"5c200019",
    11556 => x"41620015", 11557 => x"34010043", 11558 => x"5c410016",
    11559 => x"35610038", 11560 => x"b9a01000", 11561 => x"34030006",
    11562 => x"f8001e66", 11563 => x"5c200011", 11564 => x"78010001",
    11565 => x"34020001", 11566 => x"38217d48", 11567 => x"58220000",
    11568 => x"3561002c", 11569 => x"fbfffdf0", 11570 => x"37810020",
    11571 => x"fbfffde5", 11572 => x"43820020", 11573 => x"43830021",
    11574 => x"43840022", 11575 => x"43850023", 11576 => x"78010001",
    11577 => x"382154c8", 11578 => x"f800047e", 11579 => x"340c0001",
    11580 => x"b9800800", 11581 => x"2b9d0004", 11582 => x"2b8b0014",
    11583 => x"2b8c0010", 11584 => x"2b8d000c", 11585 => x"2b8e0008",
    11586 => x"379c0020", 11587 => x"c3a00000", 11588 => x"379cfffc",
    11589 => x"5b8b0004", 11590 => x"78040001", 11591 => x"38845d5c",
    11592 => x"3442ffff", 11593 => x"348a001c", 11594 => x"34030000",
    11595 => x"340900fd", 11596 => x"340800f9", 11597 => x"340700ff",
    11598 => x"3406ffa2", 11599 => x"e0000011", 11600 => x"40850000",
    11601 => x"5ca90004", 11602 => x"b4232800", 11603 => x"30a60000",
    11604 => x"e000000a", 11605 => x"5ca80005", 11606 => x"b4232800",
    11607 => x"40a50000", 11608 => x"b4651800", 11609 => x"e0000005",
    11610 => x"5ca70004", 11611 => x"b4232800", 11612 => x"c8435800",
    11613 => x"30ab0000", 11614 => x"34630001", 11615 => x"34840001",
    11616 => x"5c8afff0", 11617 => x"2b8b0004", 11618 => x"379c0004",
    11619 => x"c3a00000", 11620 => x"379cfff8", 11621 => x"5b8b0008",
    11622 => x"5b9d0004", 11623 => x"40230006", 11624 => x"34040020",
    11625 => x"4c830002", 11626 => x"34030020", 11627 => x"206b00ff",
    11628 => x"b42b1800", 11629 => x"3404ffa2", 11630 => x"30640007",
    11631 => x"4063000a", 11632 => x"34040004", 11633 => x"4c830002",
    11634 => x"34030004", 11635 => x"b5635800", 11636 => x"216b00ff",
    11637 => x"b42b1800", 11638 => x"3062000d", 11639 => x"34020001",
    11640 => x"30620010", 11641 => x"40620016", 11642 => x"34030028",
    11643 => x"4c620002", 11644 => x"34020028", 11645 => x"b5621000",
    11646 => x"204200ff", 11647 => x"b4221800", 11648 => x"34420019",
    11649 => x"34040005", 11650 => x"204b00ff", 11651 => x"30640017",
    11652 => x"30600018", 11653 => x"b9601000", 11654 => x"fbffffbe",
    11655 => x"b9600800", 11656 => x"2b9d0004", 11657 => x"2b8b0008",
    11658 => x"379c0008", 11659 => x"c3a00000", 11660 => x"379cfefc",
    11661 => x"5b8b0028", 11662 => x"5b8c0024", 11663 => x"5b8d0020",
    11664 => x"5b8e001c", 11665 => x"5b8f0018", 11666 => x"5b900014",
    11667 => x"5b910010", 11668 => x"5b92000c", 11669 => x"5b930008",
    11670 => x"5b9d0004", 11671 => x"78010001", 11672 => x"382180c8",
    11673 => x"28210000", 11674 => x"378b002c", 11675 => x"378200f4",
    11676 => x"b9601800", 11677 => x"340400c8", 11678 => x"34050000",
    11679 => x"fbfffc04", 11680 => x"34020038", 11681 => x"340c0000",
    11682 => x"504100a6", 11683 => x"b9600800", 11684 => x"fbfffda6",
    11685 => x"5c2000a3", 11686 => x"78010001", 11687 => x"78020001",
    11688 => x"38219250", 11689 => x"38425d5c", 11690 => x"78030001",
    11691 => x"40250000", 11692 => x"344e001c", 11693 => x"b9600800",
    11694 => x"34040000", 11695 => x"340d0006", 11696 => x"38635d40",
    11697 => x"340b00a0", 11698 => x"340a00a1", 11699 => x"340900a3",
    11700 => x"34080001", 11701 => x"e0000028", 11702 => x"40460000",
    11703 => x"34c70007", 11704 => x"20e700ff", 11705 => x"54ed0014",
    11706 => x"3ce70002", 11707 => x"b4673800", 11708 => x"28e60000",
    11709 => x"c0c00000", 11710 => x"b4813000", 11711 => x"40c6001c",
    11712 => x"b4862000", 11713 => x"e000001a", 11714 => x"b4812800",
    11715 => x"40a5001c", 11716 => x"51050017", 11717 => x"e000000b",
    11718 => x"b4813000", 11719 => x"40c6001c", 11720 => x"44cb000e",
    11721 => x"44ca000f", 11722 => x"44c90010", 11723 => x"5d800010",
    11724 => x"e0000004", 11725 => x"b4813800", 11726 => x"40e7001c",
    11727 => x"44e6000c", 11728 => x"78010001", 11729 => x"38219250",
    11730 => x"30250000", 11731 => x"34020005", 11732 => x"37810048",
    11733 => x"e000005b", 11734 => x"340c0002", 11735 => x"e0000004",
    11736 => x"340c0004", 11737 => x"e0000002", 11738 => x"340c0001",
    11739 => x"34840001", 11740 => x"34420001", 11741 => x"5c4effd9",
    11742 => x"78010001", 11743 => x"38219250", 11744 => x"30250000",
    11745 => x"37810048", 11746 => x"b4246800", 11747 => x"780b0001",
    11748 => x"34840001", 11749 => x"b4247800", 11750 => x"396b6894",
    11751 => x"21930003", 11752 => x"21900004", 11753 => x"39920008",
    11754 => x"e000003f", 11755 => x"41b10000", 11756 => x"46600002",
    11757 => x"5431003b", 11758 => x"222200ff", 11759 => x"50220002",
    11760 => x"b8208800", 11761 => x"29610000", 11762 => x"223100ff",
    11763 => x"b9e01000", 11764 => x"ba201800", 11765 => x"f8001d9b",
    11766 => x"3c250018", 11767 => x"b9807000", 11768 => x"14a50018",
    11769 => x"4600000a", 11770 => x"48a00007", 11771 => x"4163000c",
    11772 => x"41a10000", 11773 => x"64a20000", 11774 => x"f0610800",
    11775 => x"a0410800", 11776 => x"44200003", 11777 => x"4171000c",
    11778 => x"ba407000", 11779 => x"4163000c", 11780 => x"64a10000",
    11781 => x"e4711000", 11782 => x"a0411000", 11783 => x"5c400003",
    11784 => x"21c10008", 11785 => x"4422001e", 11786 => x"5e000003",
    11787 => x"21c10008", 11788 => x"44300004", 11789 => x"29620000",
    11790 => x"b9e00800", 11791 => x"f8001da2", 11792 => x"29650004",
    11793 => x"29630008", 11794 => x"b9a00800", 11795 => x"ba201000",
    11796 => x"b9c02000", 11797 => x"d8a00000", 11798 => x"4c01000c",
    11799 => x"5e000003", 11800 => x"21ce0008", 11801 => x"45d00005",
    11802 => x"41a30000", 11803 => x"4162000c", 11804 => x"b4621000",
    11805 => x"31a20000", 11806 => x"4164000c", 11807 => x"b5e47800",
    11808 => x"b5e17800", 11809 => x"e000000a", 11810 => x"44200006",
    11811 => x"c8011000", 11812 => x"204200ff", 11813 => x"37810048",
    11814 => x"e000000a", 11815 => x"48a10007", 11816 => x"356b0010",
    11817 => x"4161000c", 11818 => x"5c20ffc1", 11819 => x"45600003",
    11820 => x"4161000c", 11821 => x"5c200006", 11822 => x"37810048",
    11823 => x"34020002", 11824 => x"fbffff34", 11825 => x"b8205800",
    11826 => x"e0000007", 11827 => x"37810048", 11828 => x"c9e15800",
    11829 => x"b9601000", 11830 => x"fbffff0e", 11831 => x"340c0000",
    11832 => x"480b0010", 11833 => x"378c002c", 11834 => x"356b001c",
    11835 => x"b9800800", 11836 => x"b9601000", 11837 => x"34030000",
    11838 => x"fbfffdf8", 11839 => x"78050001", 11840 => x"38a580c8",
    11841 => x"28a10000", 11842 => x"b9801800", 11843 => x"378200f4",
    11844 => x"b9602000", 11845 => x"34050000", 11846 => x"fbfffbcf",
    11847 => x"340c0001", 11848 => x"b9800800", 11849 => x"2b9d0004",
    11850 => x"2b8b0028", 11851 => x"2b8c0024", 11852 => x"2b8d0020",
    11853 => x"2b8e001c", 11854 => x"2b8f0018", 11855 => x"2b900014",
    11856 => x"2b910010", 11857 => x"2b92000c", 11858 => x"2b930008",
    11859 => x"379c0104", 11860 => x"c3a00000", 11861 => x"379cffec",
    11862 => x"5b8b0010", 11863 => x"5b8c000c", 11864 => x"5b8d0008",
    11865 => x"5b9d0004", 11866 => x"b8403000", 11867 => x"40c50011",
    11868 => x"40220000", 11869 => x"b8606000", 11870 => x"402b0001",
    11871 => x"3404fffd", 11872 => x"5ca2001e", 11873 => x"34220002",
    11874 => x"34010004", 11875 => x"44a10013", 11876 => x"34010042",
    11877 => x"44a10004", 11878 => x"34010002", 11879 => x"34040000",
    11880 => x"5ca10016", 11881 => x"340d0004", 11882 => x"3404fffd",
    11883 => x"556d0013", 11884 => x"37810014", 11885 => x"b9601800",
    11886 => x"5b800014", 11887 => x"f8001d42", 11888 => x"2b810014",
    11889 => x"c9ab6800", 11890 => x"3dad0003", 11891 => x"802d6800",
    11892 => x"598d0000", 11893 => x"e0000008", 11894 => x"40c10013",
    11895 => x"55610007", 11896 => x"b8600800", 11897 => x"b58b6000",
    11898 => x"b9601800", 11899 => x"f8001d36", 11900 => x"31800000",
    11901 => x"35640002", 11902 => x"b8800800", 11903 => x"2b9d0004",
    11904 => x"2b8b0010", 11905 => x"2b8c000c", 11906 => x"2b8d0008",
    11907 => x"379c0014", 11908 => x"c3a00000", 11909 => x"379cfffc",
    11910 => x"5b9d0004", 11911 => x"40430012", 11912 => x"2844000c",
    11913 => x"b4831800", 11914 => x"fbffffcb", 11915 => x"2b9d0004",
    11916 => x"379c0004", 11917 => x"c3a00000", 11918 => x"379cffcc",
    11919 => x"5b8b0020", 11920 => x"5b8c001c", 11921 => x"5b8d0018",
    11922 => x"5b8e0014", 11923 => x"5b8f0010", 11924 => x"5b90000c",
    11925 => x"5b910008", 11926 => x"5b9d0004", 11927 => x"402e0000",
    11928 => x"204200ff", 11929 => x"208400ff", 11930 => x"344c0001",
    11931 => x"c9c27000", 11932 => x"20820001", 11933 => x"b8207800",
    11934 => x"b42c6000", 11935 => x"3401fffc", 11936 => x"5c400068",
    11937 => x"208d0004", 11938 => x"7dad0000", 11939 => x"20900008",
    11940 => x"7e100000", 11941 => x"b8605800", 11942 => x"21b100ff",
    11943 => x"e0000023", 11944 => x"b9c01800", 11945 => x"4c2e0002",
    11946 => x"b8201800", 11947 => x"29610000", 11948 => x"b9801000",
    11949 => x"206300ff", 11950 => x"f8001ce2", 11951 => x"5e00000a",
    11952 => x"b0200800", 11953 => x"64220000", 11954 => x"a0511800",
    11955 => x"44700003", 11956 => x"41630010", 11957 => x"4c6e0004",
    11958 => x"68210000", 11959 => x"a2210800", 11960 => x"4420000b",
    11961 => x"29620000", 11962 => x"41630010", 11963 => x"b9800800",
    11964 => x"340e0000", 11965 => x"f8001cf4", 11966 => x"41610010",
    11967 => x"34020001", 11968 => x"b5810800", 11969 => x"30220000",
    11970 => x"e000000d", 11971 => x"44410006", 11972 => x"41610010",
    11973 => x"34210001", 11974 => x"45c10006", 11975 => x"45a00002",
    11976 => x"49c10006", 11977 => x"356b0014", 11978 => x"41610010",
    11979 => x"5c20ffdd", 11980 => x"b9a07000", 11981 => x"e0000002",
    11982 => x"340e0001", 11983 => x"41620010", 11984 => x"34010000",
    11985 => x"44400037", 11986 => x"41610011", 11987 => x"33820034",
    11988 => x"5b8c0024", 11989 => x"33810035", 11990 => x"2961000c",
    11991 => x"5b810030", 11992 => x"45c00004", 11993 => x"41810001",
    11994 => x"34210001", 11995 => x"31810001", 11996 => x"41610010",
    11997 => x"29630004", 11998 => x"37910024", 11999 => x"34210001",
    12000 => x"b5810800", 12001 => x"ba201000", 12002 => x"d8600000",
    12003 => x"64230000", 12004 => x"a06e7000", 12005 => x"45c00019",
    12006 => x"356b0014", 12007 => x"41630010", 12008 => x"34010000",
    12009 => x"4460001f", 12010 => x"29620000", 12011 => x"b9800800",
    12012 => x"f8001cc5", 12013 => x"41610010", 12014 => x"34020001",
    12015 => x"b5810800", 12016 => x"30220000", 12017 => x"41620011",
    12018 => x"41610010", 12019 => x"29630004", 12020 => x"33820035",
    12021 => x"2962000c", 12022 => x"33810034", 12023 => x"34210001",
    12024 => x"5b820030", 12025 => x"b5810800", 12026 => x"ba201000",
    12027 => x"d8600000", 12028 => x"5c200003", 12029 => x"e000000b",
    12030 => x"5c6e0009", 12031 => x"48010009", 12032 => x"41620010",
    12033 => x"ba0d6800", 12034 => x"34420001", 12035 => x"b4220800",
    12036 => x"45a00004", 12037 => x"31e20000", 12038 => x"e0000002",
    12039 => x"34010000", 12040 => x"2b9d0004", 12041 => x"2b8b0020",
    12042 => x"2b8c001c", 12043 => x"2b8d0018", 12044 => x"2b8e0014",
    12045 => x"2b8f0010", 12046 => x"2b90000c", 12047 => x"2b910008",
    12048 => x"379c0034", 12049 => x"c3a00000", 12050 => x"379cffd0",
    12051 => x"5b8b0030", 12052 => x"5b8c002c", 12053 => x"5b8d0028",
    12054 => x"5b8e0024", 12055 => x"5b8f0020", 12056 => x"5b90001c",
    12057 => x"5b910018", 12058 => x"5b920014", 12059 => x"5b930010",
    12060 => x"5b94000c", 12061 => x"5b950008", 12062 => x"5b9d0004",
    12063 => x"208400ff", 12064 => x"40310000", 12065 => x"204200ff",
    12066 => x"008d0003", 12067 => x"344e0001", 12068 => x"208f0004",
    12069 => x"b8208000", 12070 => x"ca228800", 12071 => x"b42e7000",
    12072 => x"21ad0001", 12073 => x"b8605800", 12074 => x"340c0000",
    12075 => x"20950003", 12076 => x"20940001", 12077 => x"7df30000",
    12078 => x"e0000034", 12079 => x"b8a09000", 12080 => x"5da00005",
    12081 => x"ba209000", 12082 => x"4cb10002", 12083 => x"b8a09000",
    12084 => x"225200ff", 12085 => x"46a00002", 12086 => x"5e25002b",
    12087 => x"5da0000c", 12088 => x"29610000", 12089 => x"b9c01000",
    12090 => x"ba401800", 12091 => x"f8001c55", 12092 => x"3c2c0018",
    12093 => x"158c0018", 12094 => x"5d8d0006", 12095 => x"45ec0009",
    12096 => x"41610010", 12097 => x"5c320007", 12098 => x"e000001f",
    12099 => x"45800005", 12100 => x"69810000", 12101 => x"a0331000",
    12102 => x"5c400002", 12103 => x"45a20019", 12104 => x"45e00007",
    12105 => x"29620000", 12106 => x"41630010", 12107 => x"b9c00800",
    12108 => x"f8001c65", 12109 => x"41610010", 12110 => x"32010000",
    12111 => x"46800008", 12112 => x"29630008", 12113 => x"44600014",
    12114 => x"41610010", 12115 => x"b9601000", 12116 => x"b5c10800",
    12117 => x"d8600000", 12118 => x"48010012", 12119 => x"41610010",
    12120 => x"29630004", 12121 => x"b9601000", 12122 => x"b5c10800",
    12123 => x"d8600000", 12124 => x"44200005", 12125 => x"41620010",
    12126 => x"b4220800", 12127 => x"e0000009", 12128 => x"5c2d0007",
    12129 => x"356b0014", 12130 => x"41650010", 12131 => x"5ca0ffcc",
    12132 => x"e0000003", 12133 => x"3401fffc", 12134 => x"e0000002",
    12135 => x"34010000", 12136 => x"2b9d0004", 12137 => x"2b8b0030",
    12138 => x"2b8c002c", 12139 => x"2b8d0028", 12140 => x"2b8e0024",
    12141 => x"2b8f0020", 12142 => x"2b90001c", 12143 => x"2b910018",
    12144 => x"2b920014", 12145 => x"2b930010", 12146 => x"2b94000c",
    12147 => x"2b950008", 12148 => x"379c0030", 12149 => x"c3a00000",
    12150 => x"379cffe4", 12151 => x"5b8b0010", 12152 => x"5b8c000c",
    12153 => x"5b8d0008", 12154 => x"5b9d0004", 12155 => x"b8206000",
    12156 => x"342d0002", 12157 => x"30220000", 12158 => x"34010043",
    12159 => x"b8605800", 12160 => x"54410008", 12161 => x"34010041",
    12162 => x"50410009", 12163 => x"34010002", 12164 => x"44410007",
    12165 => x"34010004", 12166 => x"5c410029", 12167 => x"e000001c",
    12168 => x"34010046", 12169 => x"5c410026", 12170 => x"e0000009",
    12171 => x"29610000", 12172 => x"3782001c", 12173 => x"34030004",
    12174 => x"5b81001c", 12175 => x"b9a00800", 12176 => x"f8001c21",
    12177 => x"34010004", 12178 => x"e000000f", 12179 => x"78010001",
    12180 => x"38219250", 12181 => x"40210000", 12182 => x"34020000",
    12183 => x"44200019", 12184 => x"28610000", 12185 => x"37820014",
    12186 => x"5b810014", 12187 => x"28610004", 12188 => x"34030008",
    12189 => x"5b810018", 12190 => x"b9a00800", 12191 => x"f8001c12",
    12192 => x"34010008", 12193 => x"31810001", 12194 => x"e000000a",
    12195 => x"b8600800", 12196 => x"3402001f", 12197 => x"f8001def",
    12198 => x"202300ff", 12199 => x"31830001", 12200 => x"b9a00800",
    12201 => x"b9601000", 12202 => x"34630001", 12203 => x"f8001c06",
    12204 => x"41820001", 12205 => x"34420002", 12206 => x"e0000002",
    12207 => x"34020000", 12208 => x"b8400800", 12209 => x"2b9d0004",
    12210 => x"2b8b0010", 12211 => x"2b8c000c", 12212 => x"2b8d0008",
    12213 => x"379c001c", 12214 => x"c3a00000", 12215 => x"379cff98",
    12216 => x"5b8b0034", 12217 => x"5b8c0030", 12218 => x"5b8d002c",
    12219 => x"5b8e0028", 12220 => x"5b8f0024", 12221 => x"5b900020",
    12222 => x"5b91001c", 12223 => x"5b920018", 12224 => x"5b930014",
    12225 => x"5b940010", 12226 => x"5b95000c", 12227 => x"5b960008",
    12228 => x"5b9d0004", 12229 => x"b8208000", 12230 => x"28410000",
    12231 => x"b8407000", 12232 => x"340d0000", 12233 => x"40360001",
    12234 => x"402c0000", 12235 => x"340b0001", 12236 => x"378f0038",
    12237 => x"3415ffff", 12238 => x"34140002", 12239 => x"34130003",
    12240 => x"34120004", 12241 => x"34110005", 12242 => x"21a300ff",
    12243 => x"b9e00800", 12244 => x"34020000", 12245 => x"f8000c5e",
    12246 => x"b8201800", 12247 => x"4420001c", 12248 => x"4435001b",
    12249 => x"5ecb000d", 12250 => x"5d940009", 12251 => x"378b0058",
    12252 => x"34030010", 12253 => x"b9600800", 12254 => x"b9e01000",
    12255 => x"f8001bd2", 12256 => x"b9601800", 12257 => x"33800068",
    12258 => x"e000000d", 12259 => x"45930007", 12260 => x"45920008",
    12261 => x"45910009", 12262 => x"356b0001", 12263 => x"35ad0001",
    12264 => x"4c6bffea", 12265 => x"e000000a", 12266 => x"3783004c",
    12267 => x"e0000004", 12268 => x"37830050", 12269 => x"e0000002",
    12270 => x"37830048", 12271 => x"41c20011", 12272 => x"ba000800",
    12273 => x"fbffff85", 12274 => x"e0000002", 12275 => x"34010000",
    12276 => x"2b9d0004", 12277 => x"2b8b0034", 12278 => x"2b8c0030",
    12279 => x"2b8d002c", 12280 => x"2b8e0028", 12281 => x"2b8f0024",
    12282 => x"2b900020", 12283 => x"2b91001c", 12284 => x"2b920018",
    12285 => x"2b930014", 12286 => x"2b940010", 12287 => x"2b95000c",
    12288 => x"2b960008", 12289 => x"379c0068", 12290 => x"c3a00000",
    12291 => x"379cffe8", 12292 => x"5b8b0010", 12293 => x"5b8c000c",
    12294 => x"5b8d0008", 12295 => x"5b9d0004", 12296 => x"b8405800",
    12297 => x"2842000c", 12298 => x"34030001", 12299 => x"b8206800",
    12300 => x"44430019", 12301 => x"34030002", 12302 => x"5c43002e",
    12303 => x"78020001", 12304 => x"384280cc", 12305 => x"28430000",
    12306 => x"286400b4", 12307 => x"286500b0", 12308 => x"c8042000",
    12309 => x"7c820000", 12310 => x"c8052800", 12311 => x"c8a22800",
    12312 => x"3c820001", 12313 => x"3ca50001", 12314 => x"f4822000",
    12315 => x"b4852000", 12316 => x"286500a0", 12317 => x"286300a4",
    12318 => x"b4852000", 12319 => x"b4431800", 12320 => x"f4431000",
    12321 => x"5b830018", 12322 => x"b4441000", 12323 => x"5b820014",
    12324 => x"e0000014", 12325 => x"78020001", 12326 => x"384280cc",
    12327 => x"284c0000", 12328 => x"78050001", 12329 => x"38a55958",
    12330 => x"298200fc", 12331 => x"28a40000", 12332 => x"34030000",
    12333 => x"1441001f", 12334 => x"f8001aae", 12335 => x"29830100",
    12336 => x"1464001f", 12337 => x"b4431800", 12338 => x"f4431000",
    12339 => x"b4242000", 12340 => x"b4442000", 12341 => x"5b840014",
    12342 => x"5b830018", 12343 => x"b9a00800", 12344 => x"41620011",
    12345 => x"37830014", 12346 => x"fbffff3c", 12347 => x"e0000002",
    12348 => x"3401ffff", 12349 => x"2b9d0004", 12350 => x"2b8b0010",
    12351 => x"2b8c000c", 12352 => x"2b8d0008", 12353 => x"379c0018",
    12354 => x"c3a00000", 12355 => x"379cfff8", 12356 => x"5b9d0004",
    12357 => x"2843000c", 12358 => x"40450011", 12359 => x"40420012",
    12360 => x"28630000", 12361 => x"b4621000", 12362 => x"28440000",
    12363 => x"28430004", 12364 => x"4880000e", 12365 => x"5c800005",
    12366 => x"78060001", 12367 => x"38c65970", 12368 => x"28c20000",
    12369 => x"54620009", 12370 => x"3402ffff", 12371 => x"4844000b",
    12372 => x"5c82000b", 12373 => x"78040001", 12374 => x"38845974",
    12375 => x"28820000", 12376 => x"54430006", 12377 => x"e0000006",
    12378 => x"78060001", 12379 => x"38c65994", 12380 => x"28c30000",
    12381 => x"e0000002", 12382 => x"78038000", 12383 => x"5b830008",
    12384 => x"b8a01000", 12385 => x"37830008", 12386 => x"fbffff14",
    12387 => x"2b9d0004", 12388 => x"379c0008", 12389 => x"c3a00000",
    12390 => x"379cfffc", 12391 => x"5b9d0004", 12392 => x"2844000c",
    12393 => x"40430012", 12394 => x"40420011", 12395 => x"28840000",
    12396 => x"b4831800", 12397 => x"fbffff09", 12398 => x"2b9d0004",
    12399 => x"379c0004", 12400 => x"c3a00000", 12401 => x"379cfffc",
    12402 => x"5b9d0004", 12403 => x"2844000c", 12404 => x"40430012",
    12405 => x"40420011", 12406 => x"b4831800", 12407 => x"fbfffeff",
    12408 => x"2b9d0004", 12409 => x"379c0004", 12410 => x"c3a00000",
    12411 => x"379cfff0", 12412 => x"5b8b000c", 12413 => x"5b8c0008",
    12414 => x"5b9d0004", 12415 => x"b8405800", 12416 => x"2842000c",
    12417 => x"b8206000", 12418 => x"34010001", 12419 => x"5c41000a",
    12420 => x"34010000", 12421 => x"f8000286", 12422 => x"34220001",
    12423 => x"5b820010", 12424 => x"41620011", 12425 => x"b9800800",
    12426 => x"37830010", 12427 => x"fbfffeeb", 12428 => x"e0000002",
    12429 => x"3401ffff", 12430 => x"2b9d0004", 12431 => x"2b8b000c",
    12432 => x"2b8c0008", 12433 => x"379c0010", 12434 => x"c3a00000",
    12435 => x"379cfff4", 12436 => x"5b8b000c", 12437 => x"5b8c0008",
    12438 => x"5b9d0004", 12439 => x"284b000c", 12440 => x"b9601800",
    12441 => x"fbfffdbc", 12442 => x"b8206000", 12443 => x"4c01000a",
    12444 => x"29620000", 12445 => x"34010001", 12446 => x"5c410005",
    12447 => x"fbffd306", 12448 => x"fbffd2df", 12449 => x"34010064",
    12450 => x"e0000002", 12451 => x"340100c8", 12452 => x"59610000",
    12453 => x"b9800800", 12454 => x"2b9d0004", 12455 => x"2b8b000c",
    12456 => x"2b8c0008", 12457 => x"379c000c", 12458 => x"c3a00000",
    12459 => x"379cfff0", 12460 => x"5b8b0010", 12461 => x"5b8c000c",
    12462 => x"5b8d0008", 12463 => x"5b9d0004", 12464 => x"284b000c",
    12465 => x"b9601800", 12466 => x"fbfffda3", 12467 => x"b8206800",
    12468 => x"4c010050", 12469 => x"29620000", 12470 => x"34010002",
    12471 => x"4441001e", 12472 => x"48410004", 12473 => x"34010001",
    12474 => x"5c410048", 12475 => x"e0000020", 12476 => x"34010003",
    12477 => x"44410004", 12478 => x"34010032", 12479 => x"5c410043",
    12480 => x"e000003d", 12481 => x"78020001", 12482 => x"384280d0",
    12483 => x"28410014", 12484 => x"78030001", 12485 => x"38638e80",
    12486 => x"58610000", 12487 => x"28410018", 12488 => x"78030001",
    12489 => x"38638e84", 12490 => x"58610000", 12491 => x"28410010",
    12492 => x"78030001", 12493 => x"38636f2c", 12494 => x"58610000",
    12495 => x"78010001", 12496 => x"382154f0", 12497 => x"f80000e7",
    12498 => x"fbffd2d3", 12499 => x"fbffd2ac", 12500 => x"e000002c",
    12501 => x"78010001", 12502 => x"78020001", 12503 => x"382180d0",
    12504 => x"38428eec", 12505 => x"34030010", 12506 => x"f8001ad7",
    12507 => x"780c0001", 12508 => x"398c80d0", 12509 => x"41810000",
    12510 => x"5c200003", 12511 => x"340100cb", 12512 => x"e0000023",
    12513 => x"34020010", 12514 => x"b9800800", 12515 => x"f8001cb1",
    12516 => x"b8201000", 12517 => x"3403000f", 12518 => x"34010020",
    12519 => x"e0000004", 12520 => x"b44c2000", 12521 => x"30810000",
    12522 => x"34420001", 12523 => x"4c62fffd", 12524 => x"34020001",
    12525 => x"b9800800", 12526 => x"34030000", 12527 => x"f8000b44",
    12528 => x"b8201000", 12529 => x"3401fffe", 12530 => x"5c410003",
    12531 => x"340100ca", 12532 => x"e000000f", 12533 => x"3401ffff",
    12534 => x"5c410003", 12535 => x"340100c9", 12536 => x"e000000b",
    12537 => x"f80006da", 12538 => x"44200006", 12539 => x"34010065",
    12540 => x"e0000007", 12541 => x"f8000b1d", 12542 => x"3402ffff",
    12543 => x"44220003", 12544 => x"34010064", 12545 => x"e0000002",
    12546 => x"340100c8", 12547 => x"59610000", 12548 => x"b9a00800",
    12549 => x"2b9d0004", 12550 => x"2b8b0010", 12551 => x"2b8c000c",
    12552 => x"2b8d0008", 12553 => x"379c0010", 12554 => x"c3a00000",
    12555 => x"379cffc8", 12556 => x"5b8b0024", 12557 => x"5b8c0020",
    12558 => x"5b8d001c", 12559 => x"5b8e0018", 12560 => x"5b8f0014",
    12561 => x"5b900010", 12562 => x"5b91000c", 12563 => x"5b920008",
    12564 => x"5b9d0004", 12565 => x"b8207800", 12566 => x"28410000",
    12567 => x"b8406800", 12568 => x"340c0001", 12569 => x"40320001",
    12570 => x"402e0000", 12571 => x"34010000", 12572 => x"f8000938",
    12573 => x"b8202000", 12574 => x"34110002", 12575 => x"34100003",
    12576 => x"e0000025", 12577 => x"5e4c0020", 12578 => x"288b0004",
    12579 => x"5dd10007", 12580 => x"28830000", 12581 => x"78020001",
    12582 => x"37810028", 12583 => x"38424a5c", 12584 => x"f8000082",
    12585 => x"e000001f", 12586 => x"5dd00017", 12587 => x"78018000",
    12588 => x"5d610006", 12589 => x"78020001", 12590 => x"37810028",
    12591 => x"3842551c", 12592 => x"f800007a", 12593 => x"e0000017",
    12594 => x"4d600006", 12595 => x"78020001", 12596 => x"37810028",
    12597 => x"38424654", 12598 => x"c80b5800", 12599 => x"f8000073",
    12600 => x"2164ffff", 12601 => x"08842710", 12602 => x"78020001",
    12603 => x"15630010", 12604 => x"00840010", 12605 => x"37810028",
    12606 => x"38425524", 12607 => x"f800006b", 12608 => x"e0000008",
    12609 => x"b8800800", 12610 => x"f8000912", 12611 => x"b8202000",
    12612 => x"358c0001", 12613 => x"5c80ffdc", 12614 => x"34010000",
    12615 => x"e0000005", 12616 => x"41a20011", 12617 => x"b9e00800",
    12618 => x"37830028", 12619 => x"fbfffe2b", 12620 => x"2b9d0004",
    12621 => x"2b8b0024", 12622 => x"2b8c0020", 12623 => x"2b8d001c",
    12624 => x"2b8e0018", 12625 => x"2b8f0014", 12626 => x"2b900010",
    12627 => x"2b91000c", 12628 => x"2b920008", 12629 => x"379c0038",
    12630 => x"c3a00000", 12631 => x"379cffe4", 12632 => x"5b8b0010",
    12633 => x"5b8c000c", 12634 => x"5b8d0008", 12635 => x"5b9d0004",
    12636 => x"284d000c", 12637 => x"b8206000", 12638 => x"b8405800",
    12639 => x"21a10002", 12640 => x"44200009", 12641 => x"f8000617",
    12642 => x"3402000a", 12643 => x"f80019ed", 12644 => x"5b81001c",
    12645 => x"41620011", 12646 => x"b9800800", 12647 => x"3783001c",
    12648 => x"e0000013", 12649 => x"21a20004", 12650 => x"44410004",
    12651 => x"37810014", 12652 => x"34020000", 12653 => x"f80009cc",
    12654 => x"21ad0001", 12655 => x"45a00009", 12656 => x"2b820018",
    12657 => x"2b810014", 12658 => x"34030002", 12659 => x"fbfff565",
    12660 => x"b8201800", 12661 => x"41620011", 12662 => x"b9800800",
    12663 => x"e0000004", 12664 => x"41620011", 12665 => x"b9800800",
    12666 => x"37830014", 12667 => x"fbfffdfb", 12668 => x"2b9d0004",
    12669 => x"2b8b0010", 12670 => x"2b8c000c", 12671 => x"2b8d0008",
    12672 => x"379c001c", 12673 => x"c3a00000", 12674 => x"379cfffc",
    12675 => x"5b9d0004", 12676 => x"78010001", 12677 => x"34020000",
    12678 => x"34030000", 12679 => x"340400a1", 12680 => x"38216924",
    12681 => x"fbfff777", 12682 => x"78020001", 12683 => x"384280c8",
    12684 => x"58410000", 12685 => x"78010001", 12686 => x"382160a8",
    12687 => x"28210014", 12688 => x"78020001", 12689 => x"384280cc",
    12690 => x"58410000", 12691 => x"2b9d0004", 12692 => x"379c0004",
    12693 => x"c3a00000", 12694 => x"379cfff4", 12695 => x"5b8b000c",
    12696 => x"5b8c0008", 12697 => x"5b9d0004", 12698 => x"780b0001",
    12699 => x"b8202000", 12700 => x"396b81f8", 12701 => x"b8401800",
    12702 => x"b9600800", 12703 => x"b8801000", 12704 => x"f8000027",
    12705 => x"b8206000", 12706 => x"b9600800", 12707 => x"f800106b",
    12708 => x"b9800800", 12709 => x"2b9d0004", 12710 => x"2b8b000c",
    12711 => x"2b8c0008", 12712 => x"379c000c", 12713 => x"c3a00000",
    12714 => x"379cffe0", 12715 => x"5b9d0004", 12716 => x"5b83000c",
    12717 => x"3783000c", 12718 => x"5b820008", 12719 => x"5b840010",
    12720 => x"5b850014", 12721 => x"5b860018", 12722 => x"5b87001c",
    12723 => x"5b880020", 12724 => x"f8000013", 12725 => x"2b9d0004",
    12726 => x"379c0020", 12727 => x"c3a00000", 12728 => x"379cffdc",
    12729 => x"5b9d0004", 12730 => x"5b82000c", 12731 => x"3782000c",
    12732 => x"5b810008", 12733 => x"5b830010", 12734 => x"5b840014",
    12735 => x"5b850018", 12736 => x"5b86001c", 12737 => x"5b870020",
    12738 => x"5b880024", 12739 => x"fbffffd3", 12740 => x"2b9d0004",
    12741 => x"379c0024", 12742 => x"c3a00000", 12743 => x"379cff94",
    12744 => x"5b8b0044", 12745 => x"5b8c0040", 12746 => x"5b8d003c",
    12747 => x"5b8e0038", 12748 => x"5b8f0034", 12749 => x"5b900030",
    12750 => x"5b91002c", 12751 => x"5b920028", 12752 => x"5b930024",
    12753 => x"5b940020", 12754 => x"5b95001c", 12755 => x"5b960018",
    12756 => x"5b970014", 12757 => x"5b980010", 12758 => x"5b99000c",
    12759 => x"5b9b0008", 12760 => x"5b9d0004", 12761 => x"78160001",
    12762 => x"b820c800", 12763 => x"b840a000", 12764 => x"b8209800",
    12765 => x"34180025", 12766 => x"34090069", 12767 => x"34080070",
    12768 => x"34070058", 12769 => x"34060063", 12770 => x"34050064",
    12771 => x"341b002a", 12772 => x"340a0030", 12773 => x"34170010",
    12774 => x"37950060", 12775 => x"3ad6554c", 12776 => x"e0000093",
    12777 => x"34110001", 12778 => x"34100020", 12779 => x"340e000a",
    12780 => x"44380004", 12781 => x"32610000", 12782 => x"e0000038",
    12783 => x"34100030", 12784 => x"36940001", 12785 => x"42810000",
    12786 => x"4429003c", 12787 => x"5429000d", 12788 => x"44270037",
    12789 => x"54270008", 12790 => x"443b0018", 12791 => x"543b0004",
    12792 => x"44200085", 12793 => x"5c380017", 12794 => x"e000002b",
    12795 => x"5c2a0015", 12796 => x"e3fffff3", 12797 => x"44260019",
    12798 => x"5c250012", 12799 => x"e000002f", 12800 => x"4428002b",
    12801 => x"54280006", 12802 => x"3402006e", 12803 => x"44220077",
    12804 => x"3404006f", 12805 => x"5c24000b", 12806 => x"e0000022",
    12807 => x"34020075", 12808 => x"44220026", 12809 => x"34040078",
    12810 => x"44240021", 12811 => x"34020073", 12812 => x"5c220004",
    12813 => x"e000000e", 12814 => x"286e0000", 12815 => x"34630004",
    12816 => x"3422ffcf", 12817 => x"204200ff", 12818 => x"34040008",
    12819 => x"5444ffdd", 12820 => x"3431ffd0", 12821 => x"e3ffffdb",
    12822 => x"28610000", 12823 => x"34630004", 12824 => x"32610000",
    12825 => x"36730001", 12826 => x"e0000060", 12827 => x"b8600800",
    12828 => x"28210000", 12829 => x"34630004", 12830 => x"e0000004",
    12831 => x"32620000", 12832 => x"34210001", 12833 => x"36730001",
    12834 => x"40220000", 12835 => x"5c40fffc", 12836 => x"e0000056",
    12837 => x"32780000", 12838 => x"36730001", 12839 => x"e0000053",
    12840 => x"3401000a", 12841 => x"45c10004", 12842 => x"e0000004",
    12843 => x"340e0010", 12844 => x"e0000002", 12845 => x"340e0008",
    12846 => x"286d0000", 12847 => x"34720004", 12848 => x"65c3000a",
    12849 => x"01a4001f", 12850 => x"340f0000", 12851 => x"a0831800",
    12852 => x"44600003", 12853 => x"c80d6800", 12854 => x"340f0001",
    12855 => x"340c0010", 12856 => x"e0000019", 12857 => x"b9a00800",
    12858 => x"b9c01000", 12859 => x"5b85004c", 12860 => x"5b860050",
    12861 => x"5b870054", 12862 => x"5b880058", 12863 => x"5b89005c",
    12864 => x"5b8a0048", 12865 => x"f800191f", 12866 => x"b6c11800",
    12867 => x"40630000", 12868 => x"358cffff", 12869 => x"b6ac5800",
    12870 => x"b9a00800", 12871 => x"31630000", 12872 => x"b9c01000",
    12873 => x"f8001907", 12874 => x"2b8a0048", 12875 => x"2b89005c",
    12876 => x"2b880058", 12877 => x"2b870054", 12878 => x"2b860050",
    12879 => x"2b85004c", 12880 => x"b8206800", 12881 => x"7d840000",
    12882 => x"7da30000", 12883 => x"a0831800", 12884 => x"5c60ffe5",
    12885 => x"5d970004", 12886 => x"34020030", 12887 => x"3382006f",
    12888 => x"340c000f", 12889 => x"66020020", 12890 => x"a1e21000",
    12891 => x"4440000b", 12892 => x"358cffff", 12893 => x"b6ac1000",
    12894 => x"3403002d", 12895 => x"30430000", 12896 => x"340f0000",
    12897 => x"e0000005", 12898 => x"358cffff", 12899 => x"b6ac1000",
    12900 => x"30500000", 12901 => x"e0000003", 12902 => x"caf10800",
    12903 => x"b42f0800", 12904 => x"4981fffa", 12905 => x"45e00005",
    12906 => x"358cffff", 12907 => x"b6ac0800", 12908 => x"3402002d",
    12909 => x"30220000", 12910 => x"caec1800", 12911 => x"ba600800",
    12912 => x"3404000f", 12913 => x"e0000006", 12914 => x"b6ac1000",
    12915 => x"40420000", 12916 => x"358c0001", 12917 => x"30220000",
    12918 => x"34210001", 12919 => x"4c8cfffb", 12920 => x"b6639800",
    12921 => x"ba401800", 12922 => x"36940001", 12923 => x"42810000",
    12924 => x"5c20ff6d", 12925 => x"ca790800", 12926 => x"32600000",
    12927 => x"2b9d0004", 12928 => x"2b8b0044", 12929 => x"2b8c0040",
    12930 => x"2b8d003c", 12931 => x"2b8e0038", 12932 => x"2b8f0034",
    12933 => x"2b900030", 12934 => x"2b91002c", 12935 => x"2b920028",
    12936 => x"2b930024", 12937 => x"2b940020", 12938 => x"2b95001c",
    12939 => x"2b960018", 12940 => x"2b970014", 12941 => x"2b980010",
    12942 => x"2b99000c", 12943 => x"2b9b0008", 12944 => x"379c006c",
    12945 => x"c3a00000", 12946 => x"78020001", 12947 => x"14210002",
    12948 => x"38429264", 12949 => x"28420000", 12950 => x"202100ff",
    12951 => x"3c210010", 12952 => x"5841002c", 12953 => x"28410030",
    12954 => x"4c20ffff", 12955 => x"28410030", 12956 => x"2021ffff",
    12957 => x"c3a00000", 12958 => x"14210002", 12959 => x"78030001",
    12960 => x"38639264", 12961 => x"202100ff", 12962 => x"28630000",
    12963 => x"2042ffff", 12964 => x"78048000", 12965 => x"3c210010",
    12966 => x"b8441000", 12967 => x"b8411000", 12968 => x"5862002c",
    12969 => x"28610030", 12970 => x"4c20ffff", 12971 => x"c3a00000",
    12972 => x"40240002", 12973 => x"40230003", 12974 => x"78020001",
    12975 => x"3c840018", 12976 => x"3c630010", 12977 => x"38429264",
    12978 => x"b8831800", 12979 => x"40240005", 12980 => x"28420000",
    12981 => x"b8641800", 12982 => x"40240004", 12983 => x"3c840008",
    12984 => x"b8641800", 12985 => x"58430028", 12986 => x"40230001",
    12987 => x"40210000", 12988 => x"3c210008", 12989 => x"b8610800",
    12990 => x"58410024", 12991 => x"c3a00000", 12992 => x"78020001",
    12993 => x"38429264", 12994 => x"28430000", 12995 => x"28630028",
    12996 => x"30230005", 12997 => x"28430000", 12998 => x"28630028",
    12999 => x"00630008", 13000 => x"30230004", 13001 => x"28430000",
    13002 => x"28630028", 13003 => x"00630010", 13004 => x"30230003",
    13005 => x"28430000", 13006 => x"28630028", 13007 => x"00630018",
    13008 => x"30230002", 13009 => x"28430000", 13010 => x"28630024",
    13011 => x"30230001", 13012 => x"28420000", 13013 => x"28420024",
    13014 => x"00420008", 13015 => x"30220000", 13016 => x"c3a00000",
    13017 => x"379cfff4", 13018 => x"5b8b000c", 13019 => x"5b8c0008",
    13020 => x"5b9d0004", 13021 => x"780b0001", 13022 => x"b8406000",
    13023 => x"396b9264", 13024 => x"5c200004", 13025 => x"29610000",
    13026 => x"58200000", 13027 => x"e0000022", 13028 => x"29610000",
    13029 => x"58200000", 13030 => x"28220034", 13031 => x"78010001",
    13032 => x"38215560", 13033 => x"fbfffecf", 13034 => x"f80000be",
    13035 => x"29610000", 13036 => x"340200e0", 13037 => x"58220000",
    13038 => x"78010001", 13039 => x"38218278", 13040 => x"34020800",
    13041 => x"582c0000", 13042 => x"34010000", 13043 => x"fbffffab",
    13044 => x"340100c8", 13045 => x"f8000488", 13046 => x"34010000",
    13047 => x"38028000", 13048 => x"fbffffa6", 13049 => x"34010000",
    13050 => x"34020000", 13051 => x"fbffffa3", 13052 => x"34010010",
    13053 => x"34020000", 13054 => x"fbffffa0", 13055 => x"7d820000",
    13056 => x"34010000", 13057 => x"c8021000", 13058 => x"20421200",
    13059 => x"34420140", 13060 => x"fbffff9a", 13061 => x"34010000",
    13062 => x"2b9d0004", 13063 => x"2b8b000c", 13064 => x"2b8c0008",
    13065 => x"379c000c", 13066 => x"c3a00000", 13067 => x"379cfff0",
    13068 => x"5b8b000c", 13069 => x"5b8c0008", 13070 => x"5b9d0004",
    13071 => x"78020001", 13072 => x"38428278", 13073 => x"284b0000",
    13074 => x"b8206000", 13075 => x"34010004", 13076 => x"fbffff7e",
    13077 => x"7d6b0000", 13078 => x"0f810012", 13079 => x"34010004",
    13080 => x"c80b5800", 13081 => x"fbffff79", 13082 => x"216b0020",
    13083 => x"0f810012", 13084 => x"356b0004", 13085 => x"45800004",
    13086 => x"34010014", 13087 => x"fbffff73", 13088 => x"0d810000",
    13089 => x"2f810012", 13090 => x"a1610800", 13091 => x"e42b0800",
    13092 => x"2b9d0004", 13093 => x"2b8b000c", 13094 => x"2b8c0008",
    13095 => x"379c0010", 13096 => x"c3a00000", 13097 => x"379cfffc",
    13098 => x"5b9d0004", 13099 => x"34010040", 13100 => x"fbffff66",
    13101 => x"00210004", 13102 => x"2021001f", 13103 => x"08210320",
    13104 => x"2b9d0004", 13105 => x"379c0004", 13106 => x"c3a00000",
    13107 => x"379cfff4", 13108 => x"5b8b000c", 13109 => x"5b8c0008",
    13110 => x"5b9d0004", 13111 => x"78030001", 13112 => x"38638e80",
    13113 => x"b8405800", 13114 => x"28620000", 13115 => x"58220000",
    13116 => x"78010001", 13117 => x"38218e84", 13118 => x"282c0000",
    13119 => x"34010040", 13120 => x"fbffff52", 13121 => x"00210004",
    13122 => x"2021001f", 13123 => x"08210320", 13124 => x"b42c0800",
    13125 => x"59610000", 13126 => x"34010000", 13127 => x"2b9d0004",
    13128 => x"2b8b000c", 13129 => x"2b8c0008", 13130 => x"379c000c",
    13131 => x"c3a00000", 13132 => x"379cfffc", 13133 => x"5b9d0004",
    13134 => x"34010040", 13135 => x"fbffff43", 13136 => x"38220001",
    13137 => x"34010040", 13138 => x"fbffff4c", 13139 => x"34010000",
    13140 => x"2b9d0004", 13141 => x"379c0004", 13142 => x"c3a00000",
    13143 => x"379cfffc", 13144 => x"5b9d0004", 13145 => x"34010040",
    13146 => x"fbffff38", 13147 => x"3402fffe", 13148 => x"a0221000",
    13149 => x"34010040", 13150 => x"fbffff40", 13151 => x"34010000",
    13152 => x"2b9d0004", 13153 => x"379c0004", 13154 => x"c3a00000",
    13155 => x"379cfff8", 13156 => x"5b8b0008", 13157 => x"5b9d0004",
    13158 => x"780b0001", 13159 => x"396b9264", 13160 => x"29610000",
    13161 => x"28220004", 13162 => x"38420010", 13163 => x"58220004",
    13164 => x"34010001", 13165 => x"f8000410", 13166 => x"29610000",
    13167 => x"28210004", 13168 => x"20210020", 13169 => x"7c210000",
    13170 => x"2b9d0004", 13171 => x"2b8b0008", 13172 => x"379c0008",
    13173 => x"c3a00000", 13174 => x"379cfff8", 13175 => x"5b8b0008",
    13176 => x"5b9d0004", 13177 => x"b8205800", 13178 => x"34010044",
    13179 => x"fbffff17", 13180 => x"38220020", 13181 => x"45600003",
    13182 => x"3402ffdf", 13183 => x"a0221000", 13184 => x"34010044",
    13185 => x"fbffff1d", 13186 => x"34010000", 13187 => x"2b9d0004",
    13188 => x"2b8b0008", 13189 => x"379c0008", 13190 => x"c3a00000",
    13191 => x"379cfff8", 13192 => x"5b8b0008", 13193 => x"5b9d0004",
    13194 => x"78020001", 13195 => x"38428ee0", 13196 => x"28420000",
    13197 => x"780b0001", 13198 => x"396b9264", 13199 => x"59620000",
    13200 => x"fbffff1c", 13201 => x"34010001", 13202 => x"fbffffe4",
    13203 => x"78020001", 13204 => x"38425998", 13205 => x"28410000",
    13206 => x"78040001", 13207 => x"3884599c", 13208 => x"58200000",
    13209 => x"29610000", 13210 => x"28830000", 13211 => x"34020003",
    13212 => x"58200000", 13213 => x"5822000c", 13214 => x"58230008",
    13215 => x"78030001", 13216 => x"386359a0", 13217 => x"58220004",
    13218 => x"28620000", 13219 => x"5822003c", 13220 => x"2b9d0004",
    13221 => x"2b8b0008", 13222 => x"379c0008", 13223 => x"c3a00000",
    13224 => x"379cffec", 13225 => x"5b8b000c", 13226 => x"5b8c0008",
    13227 => x"5b9d0004", 13228 => x"78010001", 13229 => x"382174b4",
    13230 => x"28220000", 13231 => x"78010001", 13232 => x"38216f0c",
    13233 => x"44400003", 13234 => x"78010001", 13235 => x"38216f14",
    13236 => x"282b0000", 13237 => x"5d600004", 13238 => x"78010001",
    13239 => x"38215568", 13240 => x"e0000036", 13241 => x"78030001",
    13242 => x"386359a4", 13243 => x"282c0004", 13244 => x"29620000",
    13245 => x"28610000", 13246 => x"44410011", 13247 => x"b9600800",
    13248 => x"780400ff", 13249 => x"e000000d", 13250 => x"28230000",
    13251 => x"3c660018", 13252 => x"00650018", 13253 => x"b8c52800",
    13254 => x"a0643000", 13255 => x"00c60008", 13256 => x"2063ff00",
    13257 => x"3c630008", 13258 => x"b8a62800", 13259 => x"b8a31800",
    13260 => x"58230000", 13261 => x"34210004", 13262 => x"5581fff4",
    13263 => x"78040001", 13264 => x"388459a4", 13265 => x"29630000",
    13266 => x"28810000", 13267 => x"44610005", 13268 => x"78010001",
    13269 => x"38215580", 13270 => x"fbfffde2", 13271 => x"e000008c",
    13272 => x"78010001", 13273 => x"3821827c", 13274 => x"28220000",
    13275 => x"356b0004", 13276 => x"5c400016", 13277 => x"29630008",
    13278 => x"34021234", 13279 => x"0063000d", 13280 => x"2063ffff",
    13281 => x"5c62000b", 13282 => x"29630010", 13283 => x"34025678",
    13284 => x"0063000d", 13285 => x"2063ffff", 13286 => x"5c620006",
    13287 => x"29630018", 13288 => x"34424444", 13289 => x"0063000d",
    13290 => x"2063ffff", 13291 => x"44620005", 13292 => x"78010001",
    13293 => x"382155a8", 13294 => x"fbfffdca", 13295 => x"e0000074",
    13296 => x"34020001", 13297 => x"58220000", 13298 => x"37810010",
    13299 => x"fbfffecd", 13300 => x"78050001", 13301 => x"38a559a8",
    13302 => x"28a20000", 13303 => x"29640008", 13304 => x"29630010",
    13305 => x"29610018", 13306 => x"a0822000", 13307 => x"a0621800",
    13308 => x"a0220800", 13309 => x"59640008", 13310 => x"59630010",
    13311 => x"59610018", 13312 => x"43850010", 13313 => x"43860011",
    13314 => x"3ca50008", 13315 => x"b8a62800", 13316 => x"3ca5000d",
    13317 => x"3806cafe", 13318 => x"b8852000", 13319 => x"59640008",
    13320 => x"43840012", 13321 => x"43850013", 13322 => x"3c840008",
    13323 => x"b8852000", 13324 => x"3c84000d", 13325 => x"34050001",
    13326 => x"b8641800", 13327 => x"59630010", 13328 => x"43830014",
    13329 => x"43840015", 13330 => x"3c630008", 13331 => x"b8641800",
    13332 => x"3c63000d", 13333 => x"b8230800", 13334 => x"78030001",
    13335 => x"386359ac", 13336 => x"59610018", 13337 => x"28640000",
    13338 => x"b9600800", 13339 => x"e000000b", 13340 => x"28230000",
    13341 => x"0067000d", 13342 => x"20e7ffff", 13343 => x"5ce60006",
    13344 => x"20670007", 13345 => x"5ce50004", 13346 => x"a0621800",
    13347 => x"b8641800", 13348 => x"58230000", 13349 => x"34210008",
    13350 => x"5581fff6", 13351 => x"78040001", 13352 => x"388459a8",
    13353 => x"78030001", 13354 => x"b9600800", 13355 => x"34020000",
    13356 => x"34070aaa", 13357 => x"34060007", 13358 => x"28850000",
    13359 => x"386374b4", 13360 => x"e0000010", 13361 => x"28240000",
    13362 => x"0088000d", 13363 => x"2108ffff", 13364 => x"5d07000b",
    13365 => x"00880007", 13366 => x"2108001f", 13367 => x"5d060008",
    13368 => x"a0852000", 13369 => x"58240000", 13370 => x"28620000",
    13371 => x"3c42000d", 13372 => x"b8442000", 13373 => x"58240000",
    13374 => x"b8201000", 13375 => x"34210008", 13376 => x"5581fff1",
    13377 => x"78010001", 13378 => x"38219264", 13379 => x"28210000",
    13380 => x"34030000", 13381 => x"58200014", 13382 => x"e000000f",
    13383 => x"29640000", 13384 => x"29660004", 13385 => x"356b0008",
    13386 => x"20850fff", 13387 => x"3cc60014", 13388 => x"0084000c",
    13389 => x"58250018", 13390 => x"b8c42000", 13391 => x"3c840008",
    13392 => x"2066003f", 13393 => x"38840040", 13394 => x"b8862000",
    13395 => x"58240014", 13396 => x"34630001", 13397 => x"558bfff2",
    13398 => x"4440000b", 13399 => x"78050001", 13400 => x"38a559a8",
    13401 => x"28440000", 13402 => x"28a30000", 13403 => x"78050001",
    13404 => x"38a559b0", 13405 => x"a0831800", 13406 => x"28a40000",
    13407 => x"b8641800", 13408 => x"58430000", 13409 => x"34020080",
    13410 => x"58220014", 13411 => x"2b9d0004", 13412 => x"2b8b000c",
    13413 => x"2b8c0008", 13414 => x"379c0014", 13415 => x"c3a00000",
    13416 => x"78030001", 13417 => x"38639260", 13418 => x"44400004",
    13419 => x"28620000", 13420 => x"58410004", 13421 => x"c3a00000",
    13422 => x"28620000", 13423 => x"58410008", 13424 => x"c3a00000",
    13425 => x"78030001", 13426 => x"38639260", 13427 => x"44400004",
    13428 => x"28620000", 13429 => x"58410004", 13430 => x"c3a00000",
    13431 => x"28620000", 13432 => x"58410008", 13433 => x"c3a00000",
    13434 => x"3401012c", 13435 => x"34000000", 13436 => x"3421ffff",
    13437 => x"5c20fffe", 13438 => x"c3a00000", 13439 => x"379cfff8",
    13440 => x"5b8b0008", 13441 => x"5b9d0004", 13442 => x"202100ff",
    13443 => x"3c2b0003", 13444 => x"78020001", 13445 => x"38426f1c",
    13446 => x"b44b5800", 13447 => x"29610004", 13448 => x"34020000",
    13449 => x"fbffffdf", 13450 => x"fbfffff0", 13451 => x"29610000",
    13452 => x"34020000", 13453 => x"fbffffdb", 13454 => x"fbffffec",
    13455 => x"2b9d0004", 13456 => x"2b8b0008", 13457 => x"379c0008",
    13458 => x"c3a00000", 13459 => x"379cfff8", 13460 => x"5b8b0008",
    13461 => x"5b9d0004", 13462 => x"202100ff", 13463 => x"3c2b0003",
    13464 => x"78020001", 13465 => x"38426f1c", 13466 => x"b44b5800",
    13467 => x"29610004", 13468 => x"34020001", 13469 => x"fbffffcb",
    13470 => x"fbffffdc", 13471 => x"29610000", 13472 => x"34020001",
    13473 => x"fbffffc7", 13474 => x"fbffffd8", 13475 => x"29610004",
    13476 => x"34020000", 13477 => x"fbffffc3", 13478 => x"fbffffd4",
    13479 => x"29610000", 13480 => x"34020000", 13481 => x"fbffffbf",
    13482 => x"fbffffd0", 13483 => x"2b9d0004", 13484 => x"2b8b0008",
    13485 => x"379c0008", 13486 => x"c3a00000", 13487 => x"379cfff8",
    13488 => x"5b8b0008", 13489 => x"5b9d0004", 13490 => x"202100ff",
    13491 => x"3c2b0003", 13492 => x"78020001", 13493 => x"38426f1c",
    13494 => x"b44b5800", 13495 => x"29610004", 13496 => x"34020000",
    13497 => x"fbffffaf", 13498 => x"fbffffc0", 13499 => x"29610000",
    13500 => x"34020001", 13501 => x"fbffffab", 13502 => x"fbffffbc",
    13503 => x"29610004", 13504 => x"34020001", 13505 => x"fbffffa7",
    13506 => x"fbffffb8", 13507 => x"2b9d0004", 13508 => x"2b8b0008",
    13509 => x"379c0008", 13510 => x"c3a00000", 13511 => x"379cffec",
    13512 => x"5b8b0014", 13513 => x"5b8c0010", 13514 => x"5b8d000c",
    13515 => x"5b8e0008", 13516 => x"5b9d0004", 13517 => x"202100ff",
    13518 => x"78030001", 13519 => x"3c2b0003", 13520 => x"38636f1c",
    13521 => x"204e00ff", 13522 => x"340d0008", 13523 => x"b46b5800",
    13524 => x"29610004", 13525 => x"21c20080", 13526 => x"35adffff",
    13527 => x"fbffff91", 13528 => x"fbffffa2", 13529 => x"29610000",
    13530 => x"34020001", 13531 => x"3dce0001", 13532 => x"fbffff8c",
    13533 => x"fbffff9d", 13534 => x"29610000", 13535 => x"34020000",
    13536 => x"21ad00ff", 13537 => x"fbffff87", 13538 => x"356c0004",
    13539 => x"fbffff97", 13540 => x"21ce00ff", 13541 => x"5da0ffef",
    13542 => x"29810000", 13543 => x"34020001", 13544 => x"fbffff80",
    13545 => x"fbffff91", 13546 => x"29610000", 13547 => x"34020001",
    13548 => x"fbffff7c", 13549 => x"fbffff8d", 13550 => x"78010001",
    13551 => x"38219260", 13552 => x"28210000", 13553 => x"298d0000",
    13554 => x"34020000", 13555 => x"28210004", 13556 => x"a02d6800",
    13557 => x"29610000", 13558 => x"fbffff72", 13559 => x"fbffff83",
    13560 => x"29810000", 13561 => x"34020000", 13562 => x"fbffff6e",
    13563 => x"fbffff7f", 13564 => x"7da10000", 13565 => x"2b9d0004",
    13566 => x"2b8b0014", 13567 => x"2b8c0010", 13568 => x"2b8d000c",
    13569 => x"2b8e0008", 13570 => x"379c0014", 13571 => x"c3a00000",
    13572 => x"379cffe0", 13573 => x"5b8b0020", 13574 => x"5b8c001c",
    13575 => x"5b8d0018", 13576 => x"5b8e0014", 13577 => x"5b8f0010",
    13578 => x"5b90000c", 13579 => x"5b910008", 13580 => x"5b9d0004",
    13581 => x"202100ff", 13582 => x"3c2b0003", 13583 => x"78040001",
    13584 => x"38846f1c", 13585 => x"b48b5800", 13586 => x"29610004",
    13587 => x"b8407800", 13588 => x"34020001", 13589 => x"207000ff",
    13590 => x"fbffff52", 13591 => x"fbffff63", 13592 => x"29610000",
    13593 => x"34020000", 13594 => x"780d0001", 13595 => x"fbffff4d",
    13596 => x"340c0000", 13597 => x"fbffff5d", 13598 => x"340e0000",
    13599 => x"39ad9260", 13600 => x"34110008", 13601 => x"29610000",
    13602 => x"34020001", 13603 => x"3d8c0001", 13604 => x"fbffff44",
    13605 => x"fbffff55", 13606 => x"29a10000", 13607 => x"29620004",
    13608 => x"218c00ff", 13609 => x"28210004", 13610 => x"a0220800",
    13611 => x"44200002", 13612 => x"398c0001", 13613 => x"29610000",
    13614 => x"34020000", 13615 => x"35ce0001", 13616 => x"fbffff38",
    13617 => x"fbffff49", 13618 => x"5dd1ffef", 13619 => x"46000004",
    13620 => x"29610004", 13621 => x"34020001", 13622 => x"e0000003",
    13623 => x"29610004", 13624 => x"34020000", 13625 => x"fbffff2f",
    13626 => x"fbffff40", 13627 => x"29610000", 13628 => x"34020001",
    13629 => x"fbffff2b", 13630 => x"fbffff3c", 13631 => x"29610000",
    13632 => x"34020000", 13633 => x"fbffff27", 13634 => x"fbffff38",
    13635 => x"31ec0000", 13636 => x"2b9d0004", 13637 => x"2b8b0020",
    13638 => x"2b8c001c", 13639 => x"2b8d0018", 13640 => x"2b8e0014",
    13641 => x"2b8f0010", 13642 => x"2b90000c", 13643 => x"2b910008",
    13644 => x"379c0020", 13645 => x"c3a00000", 13646 => x"379cfff8",
    13647 => x"5b8b0008", 13648 => x"5b9d0004", 13649 => x"202100ff",
    13650 => x"3c2b0003", 13651 => x"78020001", 13652 => x"38426f1c",
    13653 => x"b44b5800", 13654 => x"29610000", 13655 => x"34020001",
    13656 => x"fbffff10", 13657 => x"fbffff21", 13658 => x"29610004",
    13659 => x"34020001", 13660 => x"fbffff0c", 13661 => x"fbffff1d",
    13662 => x"2b9d0004", 13663 => x"2b8b0008", 13664 => x"379c0008",
    13665 => x"c3a00000", 13666 => x"379cfff4", 13667 => x"5b8b000c",
    13668 => x"5b8c0008", 13669 => x"5b9d0004", 13670 => x"202b00ff",
    13671 => x"b9600800", 13672 => x"204c00ff", 13673 => x"fbffff16",
    13674 => x"3d820001", 13675 => x"b9600800", 13676 => x"204200fe",
    13677 => x"fbffff5a", 13678 => x"b8206000", 13679 => x"b9600800",
    13680 => x"fbffff3f", 13681 => x"65810000", 13682 => x"2b9d0004",
    13683 => x"2b8b000c", 13684 => x"2b8c0008", 13685 => x"379c000c",
    13686 => x"c3a00000", 13687 => x"379cffe8", 13688 => x"5b8b0018",
    13689 => x"5b8c0014", 13690 => x"5b8d0010", 13691 => x"5b8e000c",
    13692 => x"5b8f0008", 13693 => x"5b9d0004", 13694 => x"780b0001",
    13695 => x"396b9214", 13696 => x"296d000c", 13697 => x"296f0004",
    13698 => x"b8206000", 13699 => x"3dad0002", 13700 => x"c84f0800",
    13701 => x"b9a01000", 13702 => x"b8607000", 13703 => x"f80015d9",
    13704 => x"b42f1000", 13705 => x"b5af6800", 13706 => x"b44e0800",
    13707 => x"542d0006", 13708 => x"b9800800", 13709 => x"b9c01800",
    13710 => x"f8001623", 13711 => x"b8206000", 13712 => x"e0000009",
    13713 => x"c9a26800", 13714 => x"b9a01800", 13715 => x"b9800800",
    13716 => x"f800161d", 13717 => x"29620004", 13718 => x"b58d0800",
    13719 => x"c9cd1800", 13720 => x"f8001619", 13721 => x"b9800800",
    13722 => x"2b9d0004", 13723 => x"2b8b0018", 13724 => x"2b8c0014",
    13725 => x"2b8d0010", 13726 => x"2b8e000c", 13727 => x"2b8f0008",
    13728 => x"379c0018", 13729 => x"c3a00000", 13730 => x"379cffe8",
    13731 => x"5b8b0018", 13732 => x"5b8c0014", 13733 => x"5b8d0010",
    13734 => x"5b8e000c", 13735 => x"5b8f0008", 13736 => x"5b9d0004",
    13737 => x"780b0001", 13738 => x"396b9214", 13739 => x"296f000c",
    13740 => x"296e0004", 13741 => x"b8406800", 13742 => x"3def0002",
    13743 => x"c82e0800", 13744 => x"b9e01000", 13745 => x"f80015af",
    13746 => x"b42e6000", 13747 => x"b58d0800", 13748 => x"b5ee7000",
    13749 => x"542e0006", 13750 => x"b9800800", 13751 => x"34020000",
    13752 => x"b9a01800", 13753 => x"f8001676", 13754 => x"e000000b",
    13755 => x"c9cc7000", 13756 => x"34020000", 13757 => x"b9c01800",
    13758 => x"b9800800", 13759 => x"f8001670", 13760 => x"29610004",
    13761 => x"34020000", 13762 => x"c9ae1800", 13763 => x"f800166c",
    13764 => x"b9800800", 13765 => x"2b9d0004", 13766 => x"2b8b0018",
    13767 => x"2b8c0014", 13768 => x"2b8d0010", 13769 => x"2b8e000c",
    13770 => x"2b8f0008", 13771 => x"379c0018", 13772 => x"c3a00000",
    13773 => x"379cfff4", 13774 => x"5b8b000c", 13775 => x"5b8c0008",
    13776 => x"5b9d0004", 13777 => x"780c0001", 13778 => x"398c9274",
    13779 => x"29810000", 13780 => x"780b0001", 13781 => x"396b9214",
    13782 => x"58200000", 13783 => x"34020200", 13784 => x"78010001",
    13785 => x"38218680", 13786 => x"5962000c", 13787 => x"34020800",
    13788 => x"59610004", 13789 => x"59610000", 13790 => x"fbffffc4",
    13791 => x"29620004", 13792 => x"29810000", 13793 => x"58220008",
    13794 => x"2962000c", 13795 => x"5822000c", 13796 => x"34020002",
    13797 => x"5822004c", 13798 => x"34020400", 13799 => x"58220000",
    13800 => x"2b9d0004", 13801 => x"2b8b000c", 13802 => x"2b8c0008",
    13803 => x"379c000c", 13804 => x"c3a00000", 13805 => x"379cfff4",
    13806 => x"5b8b000c", 13807 => x"5b8c0008", 13808 => x"5b9d0004",
    13809 => x"780b0001", 13810 => x"396b9274", 13811 => x"29630000",
    13812 => x"340c0002", 13813 => x"78010001", 13814 => x"586c0040",
    13815 => x"78020001", 13816 => x"586c004c", 13817 => x"38219214",
    13818 => x"38428680", 13819 => x"58220004", 13820 => x"00420002",
    13821 => x"34040800", 13822 => x"5824000c", 13823 => x"344401ff",
    13824 => x"3c840010", 13825 => x"2042ffff", 13826 => x"b8821000",
    13827 => x"58620020", 13828 => x"78020001", 13829 => x"38428280",
    13830 => x"58220014", 13831 => x"34020100", 13832 => x"5822001c",
    13833 => x"58200020", 13834 => x"58200024", 13835 => x"fbffffc2",
    13836 => x"29610000", 13837 => x"582c0044", 13838 => x"2b9d0004",
    13839 => x"2b8b000c", 13840 => x"2b8c0008", 13841 => x"379c000c",
    13842 => x"c3a00000", 13843 => x"379cffc8", 13844 => x"5b8b0024",
    13845 => x"5b8c0020", 13846 => x"5b8d001c", 13847 => x"5b8e0018",
    13848 => x"5b8f0014", 13849 => x"5b900010", 13850 => x"5b91000c",
    13851 => x"5b920008", 13852 => x"5b9d0004", 13853 => x"b8805800",
    13854 => x"78040001", 13855 => x"38849274", 13856 => x"b8608000",
    13857 => x"28830000", 13858 => x"b8209000", 13859 => x"b8408800",
    13860 => x"2861004c", 13861 => x"340d0000", 13862 => x"20210002",
    13863 => x"4420008b", 13864 => x"780e0001", 13865 => x"39ce9214",
    13866 => x"29c20000", 13867 => x"28440000", 13868 => x"4804000a",
    13869 => x"28610000", 13870 => x"20210200", 13871 => x"5c200005",
    13872 => x"78010001", 13873 => x"382155d0", 13874 => x"b8801800",
    13875 => x"fbfffb85", 13876 => x"fbffff99", 13877 => x"e000007d",
    13878 => x"20810001", 13879 => x"208c0ffe", 13880 => x"c9816000",
    13881 => x"358f0003", 13882 => x"01ef0002", 13883 => x"78034000",
    13884 => x"a0831800", 13885 => x"35ef0001", 13886 => x"340dffff",
    13887 => x"5c600054", 13888 => x"7d610000", 13889 => x"0084001d",
    13890 => x"a0812000", 13891 => x"4483003e", 13892 => x"b44c1000",
    13893 => x"34030004", 13894 => x"37810034", 13895 => x"fbffff30",
    13896 => x"29c30000", 13897 => x"358dfffa", 13898 => x"358cfffe",
    13899 => x"b46c1000", 13900 => x"3781003a", 13901 => x"34030002",
    13902 => x"fbffff29", 13903 => x"78010001", 13904 => x"382159b4",
    13905 => x"282c0000", 13906 => x"37820030", 13907 => x"37810028",
    13908 => x"2b8e0034", 13909 => x"f80004e4", 13910 => x"78020001",
    13911 => x"384259b8", 13912 => x"28410000", 13913 => x"a1cc6000",
    13914 => x"01ce001c", 13915 => x"502c000e", 13916 => x"78030001",
    13917 => x"386359bc", 13918 => x"2b820030", 13919 => x"28610000",
    13920 => x"54410009", 13921 => x"2b82002c", 13922 => x"2b810028",
    13923 => x"3444ffff", 13924 => x"f4441000", 13925 => x"3421ffff",
    13926 => x"b4410800", 13927 => x"5b810028", 13928 => x"5b84002c",
    13929 => x"78020001", 13930 => x"38425994", 13931 => x"28410000",
    13932 => x"2b82002c", 13933 => x"2183000f", 13934 => x"c86e1800",
    13935 => x"a0410800", 13936 => x"5961000c", 13937 => x"6461fff1",
    13938 => x"64630001", 13939 => x"59600008", 13940 => x"b8231800",
    13941 => x"44600004", 13942 => x"34010001", 13943 => x"59610004",
    13944 => x"e0000002", 13945 => x"59600004", 13946 => x"2f81003a",
    13947 => x"3d8c0003", 13948 => x"20210800", 13949 => x"64210000",
    13950 => x"596c0010", 13951 => x"31610000", 13952 => x"b9a06000",
    13953 => x"358dfff2", 13954 => x"520d0002", 13955 => x"ba006800",
    13956 => x"780b0001", 13957 => x"396b9214", 13958 => x"29610024",
    13959 => x"29620000", 13960 => x"3403000e", 13961 => x"34210001",
    13962 => x"59610024", 13963 => x"34420004", 13964 => x"ba400800",
    13965 => x"fbfffeea", 13966 => x"29630000", 13967 => x"ba200800",
    13968 => x"34620012", 13969 => x"b9a01800", 13970 => x"fbfffee5",
    13971 => x"780b0001", 13972 => x"396b9214", 13973 => x"3dee0002",
    13974 => x"29610000", 13975 => x"b9c01000", 13976 => x"fbffff0a",
    13977 => x"78030001", 13978 => x"38639274", 13979 => x"286c0000",
    13980 => x"29610000", 13981 => x"598f0010", 13982 => x"2962000c",
    13983 => x"296f0004", 13984 => x"3c420002", 13985 => x"c82f0800",
    13986 => x"b42e0800", 13987 => x"f80014bd", 13988 => x"b42f0800",
    13989 => x"59610000", 13990 => x"29820010", 13991 => x"28210000",
    13992 => x"4801000a", 13993 => x"29810000", 13994 => x"20210200",
    13995 => x"44200002", 13996 => x"fbffff21", 13997 => x"78010001",
    13998 => x"38219274", 13999 => x"28210000", 14000 => x"34020002",
    14001 => x"5822004c", 14002 => x"b9a00800", 14003 => x"2b9d0004",
    14004 => x"2b8b0024", 14005 => x"2b8c0020", 14006 => x"2b8d001c",
    14007 => x"2b8e0018", 14008 => x"2b8f0014", 14009 => x"2b900010",
    14010 => x"2b91000c", 14011 => x"2b920008", 14012 => x"379c0038",
    14013 => x"c3a00000", 14014 => x"379cffd4", 14015 => x"5b8b0020",
    14016 => x"5b8c001c", 14017 => x"5b8d0018", 14018 => x"5b8e0014",
    14019 => x"5b8f0010", 14020 => x"5b90000c", 14021 => x"5b910008",
    14022 => x"5b9d0004", 14023 => x"780b0001", 14024 => x"78050001",
    14025 => x"396b9214", 14026 => x"38a59274", 14027 => x"b8208000",
    14028 => x"34010100", 14029 => x"5961001c", 14030 => x"59610018",
    14031 => x"b8806000", 14032 => x"28a10000", 14033 => x"78040001",
    14034 => x"38848280", 14035 => x"2e0e000c", 14036 => x"59640014",
    14037 => x"59640010", 14038 => x"58240004", 14039 => x"38018100",
    14040 => x"fdc17000", 14041 => x"3401fffc", 14042 => x"c80e7000",
    14043 => x"a1c17000", 14044 => x"35ce0012", 14045 => x"b5c36800",
    14046 => x"b8800800", 14047 => x"b8408800", 14048 => x"b8607800",
    14049 => x"34020000", 14050 => x"35a30004", 14051 => x"f800154c",
    14052 => x"29610010", 14053 => x"b9c01800", 14054 => x"ba001000",
    14055 => x"34210004", 14056 => x"f80014c9", 14057 => x"29610010",
    14058 => x"35ce0004", 14059 => x"ba201000", 14060 => x"b42e0800",
    14061 => x"b9e01800", 14062 => x"f80014c3", 14063 => x"3401003b",
    14064 => x"502d0002", 14065 => x"e0000002", 14066 => x"340d003c",
    14067 => x"35a30001", 14068 => x"7d810000", 14069 => x"00630001",
    14070 => x"3c21001e", 14071 => x"78048000", 14072 => x"b8642000",
    14073 => x"b8812000", 14074 => x"78010001", 14075 => x"38219214",
    14076 => x"28220010", 14077 => x"3c630002", 14078 => x"78010001",
    14079 => x"58440000", 14080 => x"38219274", 14081 => x"b4431000",
    14082 => x"58400000", 14083 => x"28220000", 14084 => x"340b0000",
    14085 => x"b8207800", 14086 => x"28430000", 14087 => x"341003e8",
    14088 => x"38630001", 14089 => x"58430000", 14090 => x"29e10000",
    14091 => x"282e0000", 14092 => x"21c10002", 14093 => x"5c200009",
    14094 => x"34010001", 14095 => x"356b0001", 14096 => x"f800006d",
    14097 => x"5d70fff9", 14098 => x"78010001", 14099 => x"382155f0",
    14100 => x"b9c01000", 14101 => x"fbfffaa3", 14102 => x"4580003e",
    14103 => x"780b0001", 14104 => x"340e0000", 14105 => x"396b9274",
    14106 => x"340f0064", 14107 => x"29610000", 14108 => x"28220000",
    14109 => x"20420800", 14110 => x"5c40000a", 14111 => x"34010001",
    14112 => x"35ce0001", 14113 => x"f800005c", 14114 => x"5dcffff9",
    14115 => x"78010001", 14116 => x"38215620", 14117 => x"fbfffa93",
    14118 => x"340e0000", 14119 => x"e0000003", 14120 => x"282e0014",
    14121 => x"21ce0001", 14122 => x"78010001", 14123 => x"38219274",
    14124 => x"28210000", 14125 => x"78020001", 14126 => x"384259b4",
    14127 => x"282b0018", 14128 => x"28210014", 14129 => x"28410000",
    14130 => x"3782002c", 14131 => x"a1615800", 14132 => x"37810024",
    14133 => x"f8000404", 14134 => x"78030001", 14135 => x"386359b8",
    14136 => x"28610000", 14137 => x"502b000e", 14138 => x"78030001",
    14139 => x"386359bc", 14140 => x"2b82002c", 14141 => x"28610000",
    14142 => x"54410009", 14143 => x"2b830028", 14144 => x"2b820024",
    14145 => x"3461ffff", 14146 => x"f4611800", 14147 => x"3442ffff",
    14148 => x"b4621000", 14149 => x"5b820024", 14150 => x"5b810028",
    14151 => x"2b810024", 14152 => x"318e0000", 14153 => x"3d6b0003",
    14154 => x"59810008", 14155 => x"2b810028", 14156 => x"59800004",
    14157 => x"598b0010", 14158 => x"5981000c", 14159 => x"78010001",
    14160 => x"38219214", 14161 => x"28220020", 14162 => x"34420001",
    14163 => x"58220020", 14164 => x"b9a00800", 14165 => x"2b9d0004",
    14166 => x"2b8b0020", 14167 => x"2b8c001c", 14168 => x"2b8d0018",
    14169 => x"2b8e0014", 14170 => x"2b8f0010", 14171 => x"2b90000c",
    14172 => x"2b910008", 14173 => x"379c002c", 14174 => x"c3a00000",
    14175 => x"78030001", 14176 => x"38639214", 14177 => x"28640020",
    14178 => x"58240000", 14179 => x"28610024", 14180 => x"58410000",
    14181 => x"c3a00000", 14182 => x"78020001", 14183 => x"38429278",
    14184 => x"28420000", 14185 => x"78030001", 14186 => x"38639260",
    14187 => x"58620000", 14188 => x"44200005", 14189 => x"28430010",
    14190 => x"78018000", 14191 => x"b8610800", 14192 => x"e0000006",
    14193 => x"78040001", 14194 => x"38845994", 14195 => x"28430010",
    14196 => x"28810000", 14197 => x"a0610800", 14198 => x"58410010",
    14199 => x"c3a00000", 14200 => x"78010001", 14201 => x"38219260",
    14202 => x"28210000", 14203 => x"28210014", 14204 => x"c3a00000",
    14205 => x"78020001", 14206 => x"38429260", 14207 => x"28420000",
    14208 => x"28430014", 14209 => x"b4230800", 14210 => x"28430014",
    14211 => x"c8611800", 14212 => x"4803fffe", 14213 => x"c3a00000",
    14214 => x"78010001", 14215 => x"38219260", 14216 => x"28210000",
    14217 => x"28210004", 14218 => x"20210080", 14219 => x"64210000",
    14220 => x"c3a00000", 14221 => x"379cffe0", 14222 => x"5b8b001c",
    14223 => x"5b8c0018", 14224 => x"5b8d0014", 14225 => x"5b8e0010",
    14226 => x"5b8f000c", 14227 => x"5b900008", 14228 => x"5b9d0004",
    14229 => x"b8208000", 14230 => x"34010001", 14231 => x"fbfffdb7",
    14232 => x"34010001", 14233 => x"fbfffce6", 14234 => x"340200a0",
    14235 => x"34010001", 14236 => x"fbfffd2b", 14237 => x"34020000",
    14238 => x"34010001", 14239 => x"fbfffd28", 14240 => x"34010001",
    14241 => x"fbfffcf2", 14242 => x"340200a1", 14243 => x"34010001",
    14244 => x"fbfffd23", 14245 => x"378d0023", 14246 => x"b9a01000",
    14247 => x"34030001", 14248 => x"34010001", 14249 => x"fbfffd5b",
    14250 => x"34010001", 14251 => x"fbfffd04", 14252 => x"34010001",
    14253 => x"438c0023", 14254 => x"fbfffcd1", 14255 => x"34010001",
    14256 => x"340200a1", 14257 => x"fbfffd16", 14258 => x"340bffd9",
    14259 => x"340f000f", 14260 => x"340e0017", 14261 => x"34030000",
    14262 => x"34010001", 14263 => x"b9a01000", 14264 => x"fbfffd4c",
    14265 => x"43830023", 14266 => x"b5836000", 14267 => x"218c00ff",
    14268 => x"556f0003", 14269 => x"b60b0800", 14270 => x"30230000",
    14271 => x"356b0001", 14272 => x"5d6efff5", 14273 => x"37820023",
    14274 => x"34030001", 14275 => x"34010001", 14276 => x"fbfffd40",
    14277 => x"34010001", 14278 => x"fbfffce9", 14279 => x"43810023",
    14280 => x"fc2c6000", 14281 => x"c80c0800", 14282 => x"2b9d0004",
    14283 => x"2b8b001c", 14284 => x"2b8c0018", 14285 => x"2b8d0014",
    14286 => x"2b8e0010", 14287 => x"2b8f000c", 14288 => x"2b900008",
    14289 => x"379c0020", 14290 => x"c3a00000", 14291 => x"379cffd0",
    14292 => x"5b8b0010", 14293 => x"5b8c000c", 14294 => x"5b8d0008",
    14295 => x"5b9d0004", 14296 => x"780b0001", 14297 => x"396b8eec",
    14298 => x"31600000", 14299 => x"fbffffab", 14300 => x"3403ffed",
    14301 => x"44200023", 14302 => x"b9600800", 14303 => x"fbffffae",
    14304 => x"b8206000", 14305 => x"3403fffb", 14306 => x"5c20001e",
    14307 => x"378d0014", 14308 => x"b9601000", 14309 => x"34030010",
    14310 => x"b9a00800", 14311 => x"f800157a", 14312 => x"b9a00800",
    14313 => x"f80004e8", 14314 => x"78020001", 14315 => x"38428e88",
    14316 => x"5c2c0005", 14317 => x"34010001", 14318 => x"58410000",
    14319 => x"3403fffa", 14320 => x"e0000010", 14321 => x"2b830028",
    14322 => x"78010001", 14323 => x"38218e80", 14324 => x"58230000",
    14325 => x"2b83002c", 14326 => x"78010001", 14327 => x"38218e84",
    14328 => x"58230000", 14329 => x"2b830024", 14330 => x"78010001",
    14331 => x"38216f2c", 14332 => x"58230000", 14333 => x"34010002",
    14334 => x"58410000", 14335 => x"34030000", 14336 => x"b8600800",
    14337 => x"2b9d0004", 14338 => x"2b8b0010", 14339 => x"2b8c000c",
    14340 => x"2b8d0008", 14341 => x"379c0030", 14342 => x"c3a00000",
    14343 => x"379cffe0", 14344 => x"5b9b0008", 14345 => x"341b0020",
    14346 => x"b77cd800", 14347 => x"5b8b0020", 14348 => x"5b8c001c",
    14349 => x"5b8d0018", 14350 => x"5b8e0014", 14351 => x"5b8f0010",
    14352 => x"5b90000c", 14353 => x"5b9d0004", 14354 => x"780b0001",
    14355 => x"780c0001", 14356 => x"bb807800", 14357 => x"34020001",
    14358 => x"396b7020", 14359 => x"398c5650", 14360 => x"e0000012",
    14361 => x"bb808000", 14362 => x"379cffe4", 14363 => x"378e000b",
    14364 => x"01ce0003", 14365 => x"35a2002c", 14366 => x"3dce0003",
    14367 => x"34030014", 14368 => x"b9c00800", 14369 => x"f8001390",
    14370 => x"31c00013", 14371 => x"29a20020", 14372 => x"29630074",
    14373 => x"b9800800", 14374 => x"b9c02000", 14375 => x"fbfff991",
    14376 => x"34020000", 14377 => x"ba00e000", 14378 => x"b9600800",
    14379 => x"f80011ef", 14380 => x"b8206800", 14381 => x"5c20ffec",
    14382 => x"b9e0e000", 14383 => x"2b9d0004", 14384 => x"2b8b0020",
    14385 => x"2b8c001c", 14386 => x"2b8d0018", 14387 => x"2b8e0014",
    14388 => x"2b8f0010", 14389 => x"2b90000c", 14390 => x"2b9b0008",
    14391 => x"379c0020", 14392 => x"c3a00000", 14393 => x"379cffec",
    14394 => x"5b8b0014", 14395 => x"5b8c0010", 14396 => x"5b8d000c",
    14397 => x"5b8e0008", 14398 => x"5b9d0004", 14399 => x"780b0001",
    14400 => x"396b8e8c", 14401 => x"29610000", 14402 => x"5c200007",
    14403 => x"78010001", 14404 => x"38217020", 14405 => x"f80011b3",
    14406 => x"29610000", 14407 => x"34210001", 14408 => x"59610000",
    14409 => x"780b0001", 14410 => x"396b6f30", 14411 => x"780c0001",
    14412 => x"356d00f0", 14413 => x"398c7020", 14414 => x"e0000009",
    14415 => x"29620008", 14416 => x"2963000c", 14417 => x"29640010",
    14418 => x"296e0000", 14419 => x"b9800800", 14420 => x"f8001278",
    14421 => x"59c10000", 14422 => x"356b0018", 14423 => x"5d6dfff8",
    14424 => x"2b9d0004", 14425 => x"2b8b0014", 14426 => x"2b8c0010",
    14427 => x"2b8d000c", 14428 => x"2b8e0008", 14429 => x"379c0014",
    14430 => x"c3a00000", 14431 => x"379cfff4", 14432 => x"5b8b000c",
    14433 => x"5b8c0008", 14434 => x"5b9d0004", 14435 => x"34020000",
    14436 => x"b8206000", 14437 => x"f80004a7", 14438 => x"b8205800",
    14439 => x"4c200005", 14440 => x"78010001", 14441 => x"38215678",
    14442 => x"b9601000", 14443 => x"e0000004", 14444 => x"29820000",
    14445 => x"78010001", 14446 => x"382156a4", 14447 => x"fbfff949",
    14448 => x"b9600800", 14449 => x"2b9d0004", 14450 => x"2b8b000c",
    14451 => x"2b8c0008", 14452 => x"379c000c", 14453 => x"c3a00000",
    14454 => x"379cfffc", 14455 => x"5b9d0004", 14456 => x"78010001",
    14457 => x"38218e90", 14458 => x"58200000", 14459 => x"78020001",
    14460 => x"78010001", 14461 => x"38218ea4", 14462 => x"38428e94",
    14463 => x"3403ffff", 14464 => x"58230000", 14465 => x"58430000",
    14466 => x"58200008", 14467 => x"58400008", 14468 => x"58400004",
    14469 => x"58200004", 14470 => x"5840000c", 14471 => x"5820000c",
    14472 => x"34020000", 14473 => x"34010000", 14474 => x"f8000f66",
    14475 => x"2b9d0004", 14476 => x"379c0004", 14477 => x"c3a00000",
    14478 => x"379cfff4", 14479 => x"5b8b000c", 14480 => x"5b8c0008",
    14481 => x"5b9d0004", 14482 => x"b8206000", 14483 => x"34010000",
    14484 => x"f8001005", 14485 => x"b8205800", 14486 => x"34020000",
    14487 => x"5c200081", 14488 => x"fbfffacb", 14489 => x"78030001",
    14490 => x"38638e94", 14491 => x"28650008", 14492 => x"78020001",
    14493 => x"38428e90", 14494 => x"b8202000", 14495 => x"28420000",
    14496 => x"44ab0004", 14497 => x"34010001", 14498 => x"5ca1001d",
    14499 => x"e0000010", 14500 => x"34010001", 14501 => x"44810005",
    14502 => x"28610004", 14503 => x"34210001", 14504 => x"58610004",
    14505 => x"e0000002", 14506 => x"58600004", 14507 => x"78030001",
    14508 => x"38638e94", 14509 => x"28650004", 14510 => x"34010004",
    14511 => x"4c250010", 14512 => x"34010001", 14513 => x"58610008",
    14514 => x"e0000002", 14515 => x"44850003", 14516 => x"58600004",
    14517 => x"e000000a", 14518 => x"28650004", 14519 => x"34010004",
    14520 => x"34a50001", 14521 => x"58650004", 14522 => x"4c250005",
    14523 => x"34010002", 14524 => x"58610008", 14525 => x"3441fe0c",
    14526 => x"5861000c", 14527 => x"78030001", 14528 => x"38638ea4",
    14529 => x"28650008", 14530 => x"44a00004", 14531 => x"34010001",
    14532 => x"5ca1001c", 14533 => x"e000000f", 14534 => x"44850005",
    14535 => x"28610004", 14536 => x"34210001", 14537 => x"58610004",
    14538 => x"e0000002", 14539 => x"58600004", 14540 => x"78030001",
    14541 => x"38638ea4", 14542 => x"28640004", 14543 => x"34010004",
    14544 => x"4c240010", 14545 => x"34010001", 14546 => x"58610008",
    14547 => x"e0000002", 14548 => x"44800003", 14549 => x"58600004",
    14550 => x"e000000a", 14551 => x"28640004", 14552 => x"34010004",
    14553 => x"34840001", 14554 => x"58640004", 14555 => x"4c240005",
    14556 => x"34010002", 14557 => x"58610008", 14558 => x"3441fe0c",
    14559 => x"5861000c", 14560 => x"3401251b", 14561 => x"4c220030",
    14562 => x"78020001", 14563 => x"38428e94", 14564 => x"28440008",
    14565 => x"34010002", 14566 => x"3402ffff", 14567 => x"5c810031",
    14568 => x"78030001", 14569 => x"38638ea4", 14570 => x"28610008",
    14571 => x"5c24002d", 14572 => x"2862000c", 14573 => x"34011f3f",
    14574 => x"e0000002", 14575 => x"3442e0c0", 14576 => x"4841ffff",
    14577 => x"78030001", 14578 => x"38638ea4", 14579 => x"5862000c",
    14580 => x"78030001", 14581 => x"38638e94", 14582 => x"2863000c",
    14583 => x"34011f3f", 14584 => x"e0000002", 14585 => x"3463e0c0",
    14586 => x"4861ffff", 14587 => x"78040001", 14588 => x"38848e94",
    14589 => x"5883000c", 14590 => x"4c620003", 14591 => x"3444f060",
    14592 => x"e0000004", 14593 => x"34040000", 14594 => x"4c430002",
    14595 => x"34440fa0", 14596 => x"b4831800", 14597 => x"0062001f",
    14598 => x"b4431800", 14599 => x"14620001", 14600 => x"4c400003",
    14601 => x"34421f40", 14602 => x"e0000004", 14603 => x"34011f3f",
    14604 => x"4c220002", 14605 => x"3442e0c0", 14606 => x"59820000",
    14607 => x"34020001", 14608 => x"e0000008", 14609 => x"78010001",
    14610 => x"34420064", 14611 => x"38218e90", 14612 => x"58220000",
    14613 => x"34010000", 14614 => x"f8000eda", 14615 => x"34020000",
    14616 => x"b8400800", 14617 => x"2b9d0004", 14618 => x"2b8b000c",
    14619 => x"2b8c0008", 14620 => x"379c000c", 14621 => x"c3a00000",
    14622 => x"379cfff8", 14623 => x"5b8b0008", 14624 => x"5b9d0004",
    14625 => x"78020001", 14626 => x"b8205800", 14627 => x"b8400800",
    14628 => x"382156c4", 14629 => x"fbfff893", 14630 => x"e0000003",
    14631 => x"34010064", 14632 => x"fbfffe55", 14633 => x"34010000",
    14634 => x"fbfff9e1", 14635 => x"4420fffc", 14636 => x"34010003",
    14637 => x"34020000", 14638 => x"34030001", 14639 => x"f8000de6",
    14640 => x"78020001", 14641 => x"b8400800", 14642 => x"382156dc",
    14643 => x"fbfff885", 14644 => x"e0000003", 14645 => x"34010064",
    14646 => x"fbfffe47", 14647 => x"34010000", 14648 => x"f8000ea7",
    14649 => x"4420fffc", 14650 => x"78020001", 14651 => x"b8400800",
    14652 => x"38214cd8", 14653 => x"fbfff87b", 14654 => x"78020001",
    14655 => x"b8400800", 14656 => x"382156ec", 14657 => x"fbfff877",
    14658 => x"fbffff34", 14659 => x"b9600800", 14660 => x"fbffff4a",
    14661 => x"4420fffe", 14662 => x"2b9d0004", 14663 => x"2b8b0008",
    14664 => x"379c0008", 14665 => x"c3a00000", 14666 => x"379cfff0",
    14667 => x"5b8b000c", 14668 => x"5b8c0008", 14669 => x"5b9d0004",
    14670 => x"b8405800", 14671 => x"34020003", 14672 => x"5c220020",
    14673 => x"fbffff25", 14674 => x"b9600800", 14675 => x"fbffff3b",
    14676 => x"4420fffe", 14677 => x"4c200002", 14678 => x"e000001a",
    14679 => x"37810010", 14680 => x"34020000", 14681 => x"f80003b3",
    14682 => x"b8206000", 14683 => x"48010007", 14684 => x"29620000",
    14685 => x"2b810010", 14686 => x"3443ff38", 14687 => x"54610003",
    14688 => x"344200c8", 14689 => x"50410012", 14690 => x"34020001",
    14691 => x"b9600800", 14692 => x"f80003a8", 14693 => x"78030001",
    14694 => x"b8206000", 14695 => x"29620000", 14696 => x"38635714",
    14697 => x"4c200003", 14698 => x"78030001", 14699 => x"3863570c",
    14700 => x"78010001", 14701 => x"3821571c", 14702 => x"fbfff84a",
    14703 => x"e0000004", 14704 => x"b9600800", 14705 => x"fbfffeee",
    14706 => x"b8206000", 14707 => x"29610000", 14708 => x"fbffef83",
    14709 => x"b9800800", 14710 => x"2b9d0004", 14711 => x"2b8b000c",
    14712 => x"2b8c0008", 14713 => x"379c0010", 14714 => x"c3a00000",
    14715 => x"379cfffc", 14716 => x"5b9d0004", 14717 => x"34010800",
    14718 => x"34020001", 14719 => x"fbfffaf2", 14720 => x"34010400",
    14721 => x"34020000", 14722 => x"fbfffaef", 14723 => x"34011000",
    14724 => x"34020000", 14725 => x"fbfffaec", 14726 => x"2b9d0004",
    14727 => x"379c0004", 14728 => x"c3a00000", 14729 => x"78010001",
    14730 => x"38219254", 14731 => x"28210000", 14732 => x"78020001",
    14733 => x"3842923c", 14734 => x"58410000", 14735 => x"34020001",
    14736 => x"58220000", 14737 => x"34020006", 14738 => x"58220000",
    14739 => x"c3a00000", 14740 => x"78010001", 14741 => x"3821923c",
    14742 => x"28210000", 14743 => x"3402000e", 14744 => x"58220000",
    14745 => x"c3a00000", 14746 => x"78010001", 14747 => x"3821923c",
    14748 => x"28210000", 14749 => x"34020010", 14750 => x"58220000",
    14751 => x"c3a00000", 14752 => x"78010001", 14753 => x"3821923c",
    14754 => x"28210000", 14755 => x"34020020", 14756 => x"58220000",
    14757 => x"c3a00000", 14758 => x"379cffec", 14759 => x"5b8b0014",
    14760 => x"5b8c0010", 14761 => x"5b8d000c", 14762 => x"5b8e0008",
    14763 => x"5b9d0004", 14764 => x"780b0001", 14765 => x"396b923c",
    14766 => x"29610000", 14767 => x"780c0001", 14768 => x"398c4e54",
    14769 => x"2822000c", 14770 => x"780d0002", 14771 => x"b9800800",
    14772 => x"a04d1000", 14773 => x"fbfff803", 14774 => x"29610000",
    14775 => x"2822000c", 14776 => x"b9800800", 14777 => x"2042007f",
    14778 => x"fbfff7fe", 14779 => x"78010001", 14780 => x"382159c0",
    14781 => x"282e0000", 14782 => x"e0000005", 14783 => x"28420008",
    14784 => x"b9800800", 14785 => x"a04e1000", 14786 => x"fbfff7f6",
    14787 => x"29620000", 14788 => x"2841000c", 14789 => x"a02d0800",
    14790 => x"4420fff9", 14791 => x"34010000", 14792 => x"2b9d0004",
    14793 => x"2b8b0014", 14794 => x"2b8c0010", 14795 => x"2b8d000c",
    14796 => x"2b8e0008", 14797 => x"379c0014", 14798 => x"c3a00000",
    14799 => x"40230000", 14800 => x"78020001", 14801 => x"40240001",
    14802 => x"38429268", 14803 => x"28420000", 14804 => x"3c630008",
    14805 => x"b8831800", 14806 => x"58430010", 14807 => x"40240002",
    14808 => x"40230003", 14809 => x"3c840018", 14810 => x"3c630010",
    14811 => x"b8832000", 14812 => x"40230005", 14813 => x"b8832000",
    14814 => x"40230004", 14815 => x"3c630008", 14816 => x"b8830800",
    14817 => x"58410014", 14818 => x"c3a00000", 14819 => x"40230000",
    14820 => x"40240003", 14821 => x"78020001", 14822 => x"3c630018",
    14823 => x"38429268", 14824 => x"b8831800", 14825 => x"40240001",
    14826 => x"40210002", 14827 => x"28420000", 14828 => x"3c840010",
    14829 => x"3c210008", 14830 => x"b8641800", 14831 => x"b8611800",
    14832 => x"3401ff00", 14833 => x"58430018", 14834 => x"a0611800",
    14835 => x"34630001", 14836 => x"58410020", 14837 => x"3801ea60",
    14838 => x"5843001c", 14839 => x"58410024", 14840 => x"78030001",
    14841 => x"34210001", 14842 => x"386359c4", 14843 => x"58410028",
    14844 => x"34210001", 14845 => x"5841002c", 14846 => x"28610000",
    14847 => x"78030001", 14848 => x"386359c8", 14849 => x"58410030",
    14850 => x"38018cae", 14851 => x"58410034", 14852 => x"28610000",
    14853 => x"58410038", 14854 => x"34011f40", 14855 => x"5841003c",
    14856 => x"c3a00000", 14857 => x"379cfff4", 14858 => x"5b8b000c",
    14859 => x"5b8c0008", 14860 => x"5b9d0004", 14861 => x"780b0001",
    14862 => x"780c0001", 14863 => x"396b7350", 14864 => x"398c735c",
    14865 => x"e0000005", 14866 => x"29620000", 14867 => x"b9600800",
    14868 => x"356b000c", 14869 => x"d8400000", 14870 => x"558bfffc",
    14871 => x"2b9d0004", 14872 => x"2b8b000c", 14873 => x"2b8c0008",
    14874 => x"379c000c", 14875 => x"c3a00000", 14876 => x"379cfff0",
    14877 => x"5b8b0010", 14878 => x"5b8c000c", 14879 => x"5b8d0008",
    14880 => x"5b9d0004", 14881 => x"780b0001", 14882 => x"780d0001",
    14883 => x"340c0000", 14884 => x"396b7350", 14885 => x"39ad735c",
    14886 => x"e0000006", 14887 => x"29620000", 14888 => x"b9600800",
    14889 => x"356b000c", 14890 => x"d8400000", 14891 => x"b5816000",
    14892 => x"55abfffb", 14893 => x"69810000", 14894 => x"2b9d0004",
    14895 => x"2b8b0010", 14896 => x"2b8c000c", 14897 => x"2b8d0008",
    14898 => x"379c0010", 14899 => x"c3a00000", 14900 => x"379cffec",
    14901 => x"5b8b0014", 14902 => x"5b8c0010", 14903 => x"5b8d000c",
    14904 => x"5b8e0008", 14905 => x"5b9d0004", 14906 => x"780b0001",
    14907 => x"780d0001", 14908 => x"b8207000", 14909 => x"396b7350",
    14910 => x"39ad735c", 14911 => x"e000000c", 14912 => x"296c0008",
    14913 => x"e0000007", 14914 => x"b9c01000", 14915 => x"f800124e",
    14916 => x"5c200003", 14917 => x"29810004", 14918 => x"e0000007",
    14919 => x"358c0008", 14920 => x"29810000", 14921 => x"5c20fff9",
    14922 => x"356b000c", 14923 => x"55abfff5", 14924 => x"78018000",
    14925 => x"2b9d0004", 14926 => x"2b8b0014", 14927 => x"2b8c0010",
    14928 => x"2b8d000c", 14929 => x"2b8e0008", 14930 => x"379c0014",
    14931 => x"c3a00000", 14932 => x"b8201800", 14933 => x"5c200008",
    14934 => x"78010001", 14935 => x"78020001", 14936 => x"38217350",
    14937 => x"3842735c", 14938 => x"44220003", 14939 => x"28210008",
    14940 => x"c3a00000", 14941 => x"28620008", 14942 => x"34610008",
    14943 => x"5c400016", 14944 => x"78020001", 14945 => x"78040001",
    14946 => x"38427350", 14947 => x"3884735c", 14948 => x"e000000f",
    14949 => x"28410008", 14950 => x"e000000a", 14951 => x"5c230008",
    14952 => x"78030001", 14953 => x"3442000c", 14954 => x"3863735c",
    14955 => x"34010000", 14956 => x"50430009", 14957 => x"28410008",
    14958 => x"c3a00000", 14959 => x"34210008", 14960 => x"28250000",
    14961 => x"5ca0fff6", 14962 => x"3442000c", 14963 => x"5482fff2",
    14964 => x"34010000", 14965 => x"c3a00000", 14966 => x"379cffc8",
    14967 => x"5b8b0038", 14968 => x"5b8c0034", 14969 => x"5b8d0030",
    14970 => x"5b8e002c", 14971 => x"5b8f0028", 14972 => x"5b900024",
    14973 => x"5b910020", 14974 => x"5b92001c", 14975 => x"5b930018",
    14976 => x"5b940014", 14977 => x"5b950010", 14978 => x"5b96000c",
    14979 => x"5b970008", 14980 => x"5b9d0004", 14981 => x"b8207000",
    14982 => x"34010000", 14983 => x"b840b800", 14984 => x"78140001",
    14985 => x"fbffffcb", 14986 => x"78130001", 14987 => x"78120001",
    14988 => x"78110001", 14989 => x"78100001", 14990 => x"780f0001",
    14991 => x"b8206800", 14992 => x"34150000", 14993 => x"340b0000",
    14994 => x"3a945950", 14995 => x"3a734dfc", 14996 => x"3a525748",
    14997 => x"78168000", 14998 => x"3a315524", 14999 => x"3a104654",
    15000 => x"39ef551c", 15001 => x"e0000028", 15002 => x"3562000f",
    15003 => x"b5cb0800", 15004 => x"4ae20006", 15005 => x"78020001",
    15006 => x"38425740", 15007 => x"fbfff70b", 15008 => x"b5615800",
    15009 => x"e0000021", 15010 => x"29ac0004", 15011 => x"ba801800",
    15012 => x"46a00002", 15013 => x"ba601800", 15014 => x"29a40000",
    15015 => x"ba401000", 15016 => x"fbfff702", 15017 => x"b42b5800",
    15018 => x"5d960005", 15019 => x"b5cb0800", 15020 => x"b9e01000",
    15021 => x"fbfff6fd", 15022 => x"e000000e", 15023 => x"4d800006",
    15024 => x"b5cb0800", 15025 => x"ba001000", 15026 => x"fbfff6f8",
    15027 => x"c80c6000", 15028 => x"b5615800", 15029 => x"2184ffff",
    15030 => x"08842710", 15031 => x"15830010", 15032 => x"b5cb0800",
    15033 => x"00840010", 15034 => x"ba201000", 15035 => x"fbfff6ef",
    15036 => x"b42b5800", 15037 => x"b9a00800", 15038 => x"fbffff96",
    15039 => x"b8206800", 15040 => x"36b50001", 15041 => x"5da0ffd9",
    15042 => x"b9600800", 15043 => x"2b9d0004", 15044 => x"2b8b0038",
    15045 => x"2b8c0034", 15046 => x"2b8d0030", 15047 => x"2b8e002c",
    15048 => x"2b8f0028", 15049 => x"2b900024", 15050 => x"2b910020",
    15051 => x"2b92001c", 15052 => x"2b930018", 15053 => x"2b940014",
    15054 => x"2b950010", 15055 => x"2b96000c", 15056 => x"2b970008",
    15057 => x"379c0038", 15058 => x"c3a00000", 15059 => x"379cffa8",
    15060 => x"5b8b0008", 15061 => x"5b9d0004", 15062 => x"378b000c",
    15063 => x"b9600800", 15064 => x"34020050", 15065 => x"fbffff9d",
    15066 => x"78010001", 15067 => x"b9601000", 15068 => x"38214818",
    15069 => x"fbfff6db", 15070 => x"34010000", 15071 => x"2b9d0004",
    15072 => x"2b8b0008", 15073 => x"379c0058", 15074 => x"c3a00000",
    15075 => x"78010001", 15076 => x"38218f00", 15077 => x"28210000",
    15078 => x"28220008", 15079 => x"2821000c", 15080 => x"202100ff",
    15081 => x"c3a00000", 15082 => x"78010001", 15083 => x"78030001",
    15084 => x"386359cc", 15085 => x"38218f00", 15086 => x"28210000",
    15087 => x"28620000", 15088 => x"78040001", 15089 => x"388459d0",
    15090 => x"58220000", 15091 => x"58200014", 15092 => x"28830000",
    15093 => x"58200018", 15094 => x"58200010", 15095 => x"58230000",
    15096 => x"58220000", 15097 => x"5820001c", 15098 => x"c3a00000",
    15099 => x"78040001", 15100 => x"34050002", 15101 => x"38848f00",
    15102 => x"5c25000e", 15103 => x"28810000", 15104 => x"1444001f",
    15105 => x"20840007", 15106 => x"b4831800", 15107 => x"f4832000",
    15108 => x"00630003", 15109 => x"b4821000", 15110 => x"3c42001d",
    15111 => x"58200014", 15112 => x"58200018", 15113 => x"b8431800",
    15114 => x"58230010", 15115 => x"e0000006", 15116 => x"28810000",
    15117 => x"204200ff", 15118 => x"58230014", 15119 => x"58220018",
    15120 => x"58200010", 15121 => x"78010001", 15122 => x"38218f00",
    15123 => x"28210000", 15124 => x"28220000", 15125 => x"38420004",
    15126 => x"58220000", 15127 => x"34010000", 15128 => x"c3a00000",
    15129 => x"78050001", 15130 => x"38a58f00", 15131 => x"28a50000",
    15132 => x"202100ff", 15133 => x"00630003", 15134 => x"58a20014",
    15135 => x"58a10018", 15136 => x"58a30010", 15137 => x"34010003",
    15138 => x"5c810007", 15139 => x"28a20000", 15140 => x"3401fff3",
    15141 => x"a0410800", 15142 => x"38210008", 15143 => x"58a10000",
    15144 => x"c3a00000", 15145 => x"34010001", 15146 => x"5c810007",
    15147 => x"28a2001c", 15148 => x"3401ffe7", 15149 => x"a0410800",
    15150 => x"38210008", 15151 => x"58a1001c", 15152 => x"c3a00000",
    15153 => x"34010002", 15154 => x"5c810006", 15155 => x"28a2001c",
    15156 => x"3401ffe7", 15157 => x"a0410800", 15158 => x"38210010",
    15159 => x"58a1001c", 15160 => x"c3a00000", 15161 => x"379cffe0",
    15162 => x"5b8b0020", 15163 => x"5b8c001c", 15164 => x"5b8d0018",
    15165 => x"5b8e0014", 15166 => x"5b8f0010", 15167 => x"5b90000c",
    15168 => x"5b910008", 15169 => x"5b9d0004", 15170 => x"b8206000",
    15171 => x"78010001", 15172 => x"382159b4", 15173 => x"282f0000",
    15174 => x"780b0001", 15175 => x"b8406800", 15176 => x"396b8f00",
    15177 => x"fbffff9a", 15178 => x"b8208800", 15179 => x"29610000",
    15180 => x"b8408000", 15181 => x"282e0004", 15182 => x"a1cf7000",
    15183 => x"fbffff94", 15184 => x"5c31fff9", 15185 => x"5c50fff8",
    15186 => x"45800003", 15187 => x"59810000", 15188 => x"59820004",
    15189 => x"45a00003", 15190 => x"3dc10003", 15191 => x"59a10000",
    15192 => x"2b9d0004", 15193 => x"2b8b0020", 15194 => x"2b8c001c",
    15195 => x"2b8d0018", 15196 => x"2b8e0014", 15197 => x"2b8f0010",
    15198 => x"2b90000c", 15199 => x"2b910008", 15200 => x"379c0020",
    15201 => x"c3a00000", 15202 => x"78010001", 15203 => x"38218f00",
    15204 => x"28210000", 15205 => x"28210000", 15206 => x"20210004",
    15207 => x"64210000", 15208 => x"c3a00000", 15209 => x"78020001",
    15210 => x"38428f00", 15211 => x"28420000", 15212 => x"2843001c",
    15213 => x"44200003", 15214 => x"38630006", 15215 => x"e0000003",
    15216 => x"3401fff9", 15217 => x"a0611800", 15218 => x"5843001c",
    15219 => x"34010000", 15220 => x"c3a00000", 15221 => x"379cffe0",
    15222 => x"5b8b001c", 15223 => x"5b8c0018", 15224 => x"5b8d0014",
    15225 => x"5b8e0010", 15226 => x"5b8f000c", 15227 => x"5b900008",
    15228 => x"5b9d0004", 15229 => x"b8205800", 15230 => x"78010001",
    15231 => x"38218eb4", 15232 => x"b8406000", 15233 => x"40220000",
    15234 => x"b8607000", 15235 => x"b8807800", 15236 => x"b8a06800",
    15237 => x"3401ffff", 15238 => x"4440002b", 15239 => x"3d8c0001",
    15240 => x"b9600800", 15241 => x"fbfff8f6", 15242 => x"218200fe",
    15243 => x"b9600800", 15244 => x"fbfff93b", 15245 => x"01c20008",
    15246 => x"b9600800", 15247 => x"204200ff", 15248 => x"fbfff937",
    15249 => x"21c200ff", 15250 => x"b9600800", 15251 => x"fbfff934",
    15252 => x"b9600800", 15253 => x"fbfff8fe", 15254 => x"39820001",
    15255 => x"b9600800", 15256 => x"204200ff", 15257 => x"fbfff92e",
    15258 => x"340c0000", 15259 => x"35aeffff", 15260 => x"37900023",
    15261 => x"e0000009", 15262 => x"b9600800", 15263 => x"ba001000",
    15264 => x"34030000", 15265 => x"fbfff963", 15266 => x"43820023",
    15267 => x"b5ec0800", 15268 => x"358c0001", 15269 => x"30220000",
    15270 => x"55ccfff8", 15271 => x"b9600800", 15272 => x"ba001000",
    15273 => x"34030001", 15274 => x"fbfff95a", 15275 => x"43810023",
    15276 => x"b5ee7000", 15277 => x"31c10000", 15278 => x"b9600800",
    15279 => x"fbfff900", 15280 => x"b9a00800", 15281 => x"2b9d0004",
    15282 => x"2b8b001c", 15283 => x"2b8c0018", 15284 => x"2b8d0014",
    15285 => x"2b8e0010", 15286 => x"2b8f000c", 15287 => x"2b900008",
    15288 => x"379c0020", 15289 => x"c3a00000", 15290 => x"379cffe0",
    15291 => x"5b8b0020", 15292 => x"5b8c001c", 15293 => x"5b8d0018",
    15294 => x"5b8e0014", 15295 => x"5b8f0010", 15296 => x"5b90000c",
    15297 => x"5b910008", 15298 => x"5b9d0004", 15299 => x"b8205800",
    15300 => x"78010001", 15301 => x"38218eb4", 15302 => x"b8606800",
    15303 => x"40230000", 15304 => x"3c4f0001", 15305 => x"b8808000",
    15306 => x"b8a07000", 15307 => x"3401ffff", 15308 => x"21ef00ff",
    15309 => x"340c0000", 15310 => x"5c60001f", 15311 => x"e0000020",
    15312 => x"b9600800", 15313 => x"fbfff8ae", 15314 => x"b9e01000",
    15315 => x"b9600800", 15316 => x"fbfff8f3", 15317 => x"01a20008",
    15318 => x"b9600800", 15319 => x"204200ff", 15320 => x"fbfff8ef",
    15321 => x"21a200ff", 15322 => x"b9600800", 15323 => x"fbfff8ec",
    15324 => x"b60c1000", 15325 => x"40420000", 15326 => x"b9600800",
    15327 => x"35ad0001", 15328 => x"fbfff8e7", 15329 => x"b9600800",
    15330 => x"fbfff8cd", 15331 => x"b9600800", 15332 => x"fbfff89b",
    15333 => x"b9600800", 15334 => x"b9e01000", 15335 => x"fbfff8e0",
    15336 => x"b8208800", 15337 => x"b9600800", 15338 => x"fbfff8c5",
    15339 => x"5e20fff8", 15340 => x"358c0001", 15341 => x"55ccffe3",
    15342 => x"b9c00800", 15343 => x"2b9d0004", 15344 => x"2b8b0020",
    15345 => x"2b8c001c", 15346 => x"2b8d0018", 15347 => x"2b8e0014",
    15348 => x"2b8f0010", 15349 => x"2b90000c", 15350 => x"2b910008",
    15351 => x"379c0020", 15352 => x"c3a00000", 15353 => x"379cffec",
    15354 => x"5b8b0014", 15355 => x"5b8c0010", 15356 => x"5b8d000c",
    15357 => x"5b8e0008", 15358 => x"5b9d0004", 15359 => x"780d0001",
    15360 => x"780c0001", 15361 => x"39ad8eb8", 15362 => x"398c8ebc",
    15363 => x"780b0001", 15364 => x"59a10000", 15365 => x"59820000",
    15366 => x"34030001", 15367 => x"396b8eb4", 15368 => x"202100ff",
    15369 => x"204200ff", 15370 => x"31630000", 15371 => x"fbfff957",
    15372 => x"b8207000", 15373 => x"5c200006", 15374 => x"41a10003",
    15375 => x"41820003", 15376 => x"fbfff952", 15377 => x"5c2e0002",
    15378 => x"31600000", 15379 => x"2b9d0004", 15380 => x"2b8b0014",
    15381 => x"2b8c0010", 15382 => x"2b8d000c", 15383 => x"2b8e0008",
    15384 => x"379c0014", 15385 => x"c3a00000", 15386 => x"379cfff8",
    15387 => x"5b8b0008", 15388 => x"5b9d0004", 15389 => x"78010001",
    15390 => x"78020001", 15391 => x"38218eb8", 15392 => x"38428ebc",
    15393 => x"40420003", 15394 => x"780b0001", 15395 => x"40210003",
    15396 => x"396b70d8", 15397 => x"34031004", 15398 => x"b9602000",
    15399 => x"34050001", 15400 => x"31600000", 15401 => x"fbffff91",
    15402 => x"34030001", 15403 => x"3402ffff", 15404 => x"5c230002",
    15405 => x"41620000", 15406 => x"b8400800", 15407 => x"2b9d0004",
    15408 => x"2b8b0008", 15409 => x"379c0008", 15410 => x"c3a00000",
    15411 => x"379cffc4", 15412 => x"5b8b001c", 15413 => x"5b8c0018",
    15414 => x"5b8d0014", 15415 => x"5b8e0010", 15416 => x"5b8f000c",
    15417 => x"5b900008", 15418 => x"5b9d0004", 15419 => x"b8205800",
    15420 => x"206d00ff", 15421 => x"34010002", 15422 => x"204c00ff",
    15423 => x"3405fffc", 15424 => x"55a10087", 15425 => x"78040001",
    15426 => x"388470d8", 15427 => x"40820000", 15428 => x"340100ff",
    15429 => x"5c41000d", 15430 => x"78010001", 15431 => x"78020001",
    15432 => x"38218eb8", 15433 => x"38428ebc", 15434 => x"40420003",
    15435 => x"40210003", 15436 => x"34050001", 15437 => x"34031004",
    15438 => x"fbffff27", 15439 => x"34020001", 15440 => x"3405ffff",
    15441 => x"5c220076", 15442 => x"78010001", 15443 => x"382170d8",
    15444 => x"40230000", 15445 => x"340200ff", 15446 => x"5c620002",
    15447 => x"30200000", 15448 => x"5d800021", 15449 => x"78010001",
    15450 => x"382170d8", 15451 => x"40210000", 15452 => x"34050000",
    15453 => x"442c006a", 15454 => x"78010001", 15455 => x"78020001",
    15456 => x"38218eb8", 15457 => x"38428ebc", 15458 => x"09a3001d",
    15459 => x"40420003", 15460 => x"40210003", 15461 => x"3405001d",
    15462 => x"34631005", 15463 => x"b9602000", 15464 => x"fbffff0d",
    15465 => x"3402001d", 15466 => x"b9606000", 15467 => x"3405ffff",
    15468 => x"5c22005b", 15469 => x"3562001c", 15470 => x"34010000",
    15471 => x"e0000005", 15472 => x"41830000", 15473 => x"358c0001",
    15474 => x"b4230800", 15475 => x"202100ff", 15476 => x"5d82fffc",
    15477 => x"4162001c", 15478 => x"3405fffd", 15479 => x"5c410050",
    15480 => x"e000004a", 15481 => x"34010001", 15482 => x"5d810048",
    15483 => x"780f0001", 15484 => x"780e0001", 15485 => x"780d0001",
    15486 => x"340c0000", 15487 => x"39ef70d8", 15488 => x"39ce8eb8",
    15489 => x"39ad8ebc", 15490 => x"37900020", 15491 => x"e0000015",
    15492 => x"0983001d", 15493 => x"41a20003", 15494 => x"41c10003",
    15495 => x"34631005", 15496 => x"ba002000", 15497 => x"3405001d",
    15498 => x"fbfffeeb", 15499 => x"3402001d", 15500 => x"5c22003a",
    15501 => x"ba000800", 15502 => x"b9601000", 15503 => x"34030010",
    15504 => x"f8001084", 15505 => x"5c200005", 15506 => x"78010001",
    15507 => x"38215764", 15508 => x"fbfff524", 15509 => x"e0000005",
    15510 => x"358c0001", 15511 => x"218c00ff", 15512 => x"41e10000",
    15513 => x"542cffeb", 15514 => x"34010002", 15515 => x"3405fffe",
    15516 => x"5581002b", 15517 => x"3563001c", 15518 => x"b9600800",
    15519 => x"34020000", 15520 => x"e0000005", 15521 => x"40240000",
    15522 => x"34210001", 15523 => x"b4441000", 15524 => x"204200ff",
    15525 => x"5c23fffc", 15526 => x"780e0001", 15527 => x"780d0001",
    15528 => x"3162001c", 15529 => x"39ce8eb8", 15530 => x"39ad8ebc",
    15531 => x"0983001d", 15532 => x"41c10003", 15533 => x"41a20003",
    15534 => x"b9602000", 15535 => x"34631005", 15536 => x"3405001d",
    15537 => x"780b0001", 15538 => x"fbffff08", 15539 => x"396b70d8",
    15540 => x"41610000", 15541 => x"542c000d", 15542 => x"78010001",
    15543 => x"38215780", 15544 => x"fbfff500", 15545 => x"41610000",
    15546 => x"41a20003", 15547 => x"34031004", 15548 => x"34210001",
    15549 => x"31610000", 15550 => x"41c10003", 15551 => x"b9602000",
    15552 => x"34050001", 15553 => x"fbfffef9", 15554 => x"78010001",
    15555 => x"382170d8", 15556 => x"40250000", 15557 => x"e0000002",
    15558 => x"3405ffff", 15559 => x"b8a00800", 15560 => x"2b9d0004",
    15561 => x"2b8b001c", 15562 => x"2b8c0018", 15563 => x"2b8d0014",
    15564 => x"2b8e0010", 15565 => x"2b8f000c", 15566 => x"2b900008",
    15567 => x"379c003c", 15568 => x"c3a00000", 15569 => x"379cffcc",
    15570 => x"5b8b0014", 15571 => x"5b8c0010", 15572 => x"5b8d000c",
    15573 => x"5b8e0008", 15574 => x"5b9d0004", 15575 => x"340d0000",
    15576 => x"b8205800", 15577 => x"340c0001", 15578 => x"378e0018",
    15579 => x"e0000027", 15580 => x"b9c00800", 15581 => x"34020000",
    15582 => x"b9a01800", 15583 => x"fbffff54", 15584 => x"b8206000",
    15585 => x"4c010023", 15586 => x"b9c00800", 15587 => x"b9601000",
    15588 => x"34030010", 15589 => x"f800102f", 15590 => x"35ad0001",
    15591 => x"5c20001b", 15592 => x"2b81002c", 15593 => x"340c0001",
    15594 => x"00220018", 15595 => x"31610017", 15596 => x"31620014",
    15597 => x"00220010", 15598 => x"31620015", 15599 => x"00220008",
    15600 => x"2b810030", 15601 => x"31620016", 15602 => x"00220018",
    15603 => x"3161001b", 15604 => x"31620018", 15605 => x"00220010",
    15606 => x"31620019", 15607 => x"00220008", 15608 => x"2b810028",
    15609 => x"3162001a", 15610 => x"00220018", 15611 => x"31610013",
    15612 => x"31620010", 15613 => x"00220010", 15614 => x"31620011",
    15615 => x"00220008", 15616 => x"31620012", 15617 => x"e0000003",
    15618 => x"498dffda", 15619 => x"340c0000", 15620 => x"b9800800",
    15621 => x"2b9d0004", 15622 => x"2b8b0014", 15623 => x"2b8c0010",
    15624 => x"2b8d000c", 15625 => x"2b8e0008", 15626 => x"379c0034",
    15627 => x"c3a00000", 15628 => x"379cfff8", 15629 => x"5b8b0008",
    15630 => x"5b9d0004", 15631 => x"78030001", 15632 => x"b8205800",
    15633 => x"204200ff", 15634 => x"78010001", 15635 => x"38218eb8",
    15636 => x"38638ebc", 15637 => x"44400015", 15638 => x"29640000",
    15639 => x"78028000", 15640 => x"34050004", 15641 => x"b8821000",
    15642 => x"59620000", 15643 => x"40620003", 15644 => x"40210003",
    15645 => x"34031000", 15646 => x"b9602000", 15647 => x"fbfffe9b",
    15648 => x"7c210004", 15649 => x"78040001", 15650 => x"38845994",
    15651 => x"c8011000", 15652 => x"29630000", 15653 => x"28810000",
    15654 => x"38420001", 15655 => x"a0610800", 15656 => x"59610000",
    15657 => x"e0000013", 15658 => x"40620003", 15659 => x"40210003",
    15660 => x"34031000", 15661 => x"b9602000", 15662 => x"34050004",
    15663 => x"fbfffe46", 15664 => x"34030004", 15665 => x"3402ffff",
    15666 => x"5c23000a", 15667 => x"29610000", 15668 => x"34020000",
    15669 => x"4c200007", 15670 => x"78030001", 15671 => x"38635994",
    15672 => x"28620000", 15673 => x"a0220800", 15674 => x"59610000",
    15675 => x"34020001", 15676 => x"b8400800", 15677 => x"2b9d0004",
    15678 => x"2b8b0008", 15679 => x"379c0008", 15680 => x"c3a00000",
    15681 => x"379cfff8", 15682 => x"5b9d0004", 15683 => x"78010001",
    15684 => x"78020001", 15685 => x"38218eb8", 15686 => x"38428ebc",
    15687 => x"40420003", 15688 => x"40210003", 15689 => x"34031074",
    15690 => x"3784000a", 15691 => x"34050002", 15692 => x"0f80000a",
    15693 => x"fbfffe6d", 15694 => x"34030002", 15695 => x"3402ffff",
    15696 => x"5c230002", 15697 => x"2f82000a", 15698 => x"b8400800",
    15699 => x"2b9d0004", 15700 => x"379c0008", 15701 => x"c3a00000",
    15702 => x"379cffcc", 15703 => x"5b8b002c", 15704 => x"5b8c0028",
    15705 => x"5b8d0024", 15706 => x"5b8e0020", 15707 => x"5b8f001c",
    15708 => x"5b900018", 15709 => x"5b910014", 15710 => x"5b920010",
    15711 => x"5b93000c", 15712 => x"5b940008", 15713 => x"5b9d0004",
    15714 => x"78030001", 15715 => x"78020001", 15716 => x"38638eb8",
    15717 => x"b8208800", 15718 => x"38428ebc", 15719 => x"34010020",
    15720 => x"33810037", 15721 => x"40420003", 15722 => x"40610003",
    15723 => x"37840034", 15724 => x"34031074", 15725 => x"34050002",
    15726 => x"fbfffe07", 15727 => x"34020002", 15728 => x"340bffff",
    15729 => x"5c220051", 15730 => x"2f820034", 15731 => x"3801ffff",
    15732 => x"5c410002", 15733 => x"0f800034", 15734 => x"780d0001",
    15735 => x"780c0001", 15736 => x"340b0001", 15737 => x"39ad8eb8",
    15738 => x"398c8ebc", 15739 => x"37900037", 15740 => x"e0000023",
    15741 => x"41b40003", 15742 => x"41930003", 15743 => x"b9c00800",
    15744 => x"34721076", 15745 => x"f8000f64", 15746 => x"b8202800",
    15747 => x"b9c02000", 15748 => x"ba800800", 15749 => x"ba601000",
    15750 => x"ba401800", 15751 => x"fbfffe33", 15752 => x"b8207000",
    15753 => x"29e10000", 15754 => x"f8000f5b", 15755 => x"5dc10036",
    15756 => x"29e10000", 15757 => x"2f8e0034", 15758 => x"f8000f57",
    15759 => x"b5c11800", 15760 => x"41820003", 15761 => x"41a10003",
    15762 => x"2063ffff", 15763 => x"0f830034", 15764 => x"ba002000",
    15765 => x"34631076", 15766 => x"34050001", 15767 => x"fbfffe23",
    15768 => x"34020001", 15769 => x"5c220028", 15770 => x"2f810034",
    15771 => x"356b0001", 15772 => x"216b00ff", 15773 => x"34210001",
    15774 => x"0f810034", 15775 => x"3d6f0002", 15776 => x"2f830034",
    15777 => x"b62f7800", 15778 => x"29ee0000", 15779 => x"5dc0ffda",
    15780 => x"3401000a", 15781 => x"33810037", 15782 => x"41820003",
    15783 => x"41a10003", 15784 => x"34631075", 15785 => x"37840037",
    15786 => x"34050001", 15787 => x"fbfffe0f", 15788 => x"34020001",
    15789 => x"340bffff", 15790 => x"5c220014", 15791 => x"41a10003",
    15792 => x"41820003", 15793 => x"34031074", 15794 => x"37840034",
    15795 => x"34050002", 15796 => x"fbfffe06", 15797 => x"b8207000",
    15798 => x"34010002", 15799 => x"5dc1000b", 15800 => x"41a10003",
    15801 => x"41820003", 15802 => x"34031074", 15803 => x"37840032",
    15804 => x"34050002", 15805 => x"fbfffdb8", 15806 => x"e42e5800",
    15807 => x"356bffff", 15808 => x"e0000002", 15809 => x"340bffff",
    15810 => x"b9600800", 15811 => x"2b9d0004", 15812 => x"2b8b002c",
    15813 => x"2b8c0028", 15814 => x"2b8d0024", 15815 => x"2b8e0020",
    15816 => x"2b8f001c", 15817 => x"2b900018", 15818 => x"2b910014",
    15819 => x"2b920010", 15820 => x"2b93000c", 15821 => x"2b940008",
    15822 => x"379c0034", 15823 => x"c3a00000", 15824 => x"379cffe4",
    15825 => x"5b8b0018", 15826 => x"5b8c0014", 15827 => x"5b8d0010",
    15828 => x"5b8e000c", 15829 => x"5b8f0008", 15830 => x"5b9d0004",
    15831 => x"78010001", 15832 => x"78020001", 15833 => x"38218eb8",
    15834 => x"38428ebc", 15835 => x"40420003", 15836 => x"40210003",
    15837 => x"34031074", 15838 => x"3784001c", 15839 => x"34050002",
    15840 => x"fbfffd95", 15841 => x"34030002", 15842 => x"3402ffff",
    15843 => x"5c230025", 15844 => x"2f81001c", 15845 => x"3802fffd",
    15846 => x"3421ffff", 15847 => x"2021ffff", 15848 => x"50410005",
    15849 => x"78010001", 15850 => x"38214e80", 15851 => x"0f80001c",
    15852 => x"fbfff3cc", 15853 => x"780e0001", 15854 => x"780d0001",
    15855 => x"780c0001", 15856 => x"340b0000", 15857 => x"39ce8eb8",
    15858 => x"39ad8ebc", 15859 => x"378f001f", 15860 => x"398c4e7c",
    15861 => x"e000000e", 15862 => x"41a20003", 15863 => x"41c10003",
    15864 => x"35631076", 15865 => x"b9e02000", 15866 => x"34050001",
    15867 => x"fbfffd7a", 15868 => x"34020001", 15869 => x"5c22000a",
    15870 => x"4382001f", 15871 => x"b9800800", 15872 => x"356b0001",
    15873 => x"fbfff3b7", 15874 => x"216bffff", 15875 => x"2f81001c",
    15876 => x"542bfff2", 15877 => x"34020000", 15878 => x"e0000002",
    15879 => x"3402ffff", 15880 => x"b8400800", 15881 => x"2b9d0004",
    15882 => x"2b8b0018", 15883 => x"2b8c0014", 15884 => x"2b8d0010",
    15885 => x"2b8e000c", 15886 => x"2b8f0008", 15887 => x"379c001c",
    15888 => x"c3a00000", 15889 => x"379cffdc", 15890 => x"5b8b0024",
    15891 => x"5b8c0020", 15892 => x"5b8d001c", 15893 => x"5b8e0018",
    15894 => x"5b8f0014", 15895 => x"5b900010", 15896 => x"5b91000c",
    15897 => x"5b920008", 15898 => x"5b9d0004", 15899 => x"206300ff",
    15900 => x"b8208800", 15901 => x"205200ff", 15902 => x"5c600012",
    15903 => x"78040001", 15904 => x"78030001", 15905 => x"38848eb8",
    15906 => x"38638ebc", 15907 => x"40620003", 15908 => x"40810003",
    15909 => x"78040001", 15910 => x"34031074", 15911 => x"38848ec0",
    15912 => x"34050002", 15913 => x"fbfffd4c", 15914 => x"34020002",
    15915 => x"3403ffff", 15916 => x"5c22002b", 15917 => x"78030001",
    15918 => x"38638ec2", 15919 => x"0c610000", 15920 => x"78040001",
    15921 => x"38848ec2", 15922 => x"78030001", 15923 => x"38638ec0",
    15924 => x"2c820000", 15925 => x"2c610000", 15926 => x"34030000",
    15927 => x"3442fffe", 15928 => x"5041001f", 15929 => x"780d0001",
    15930 => x"780c0001", 15931 => x"340b0000", 15932 => x"b8807000",
    15933 => x"39ad8eb8", 15934 => x"398c8ebc", 15935 => x"3410000a",
    15936 => x"2dc30000", 15937 => x"3461fffe", 15938 => x"54320012",
    15939 => x"41820003", 15940 => x"41a10003", 15941 => x"34640001",
    15942 => x"b62b7800", 15943 => x"0dc40000", 15944 => x"34631074",
    15945 => x"b9e02000", 15946 => x"34050001", 15947 => x"fbfffd2a",
    15948 => x"34020001", 15949 => x"5c220009", 15950 => x"41e10000",
    15951 => x"356b0001", 15952 => x"216b00ff", 15953 => x"5c30ffef",
    15954 => x"b9601800", 15955 => x"e0000004", 15956 => x"3403fffd",
    15957 => x"e0000002", 15958 => x"3403ffff", 15959 => x"b8600800",
    15960 => x"2b9d0004", 15961 => x"2b8b0024", 15962 => x"2b8c0020",
    15963 => x"2b8d001c", 15964 => x"2b8e0018", 15965 => x"2b8f0014",
    15966 => x"2b900010", 15967 => x"2b91000c", 15968 => x"2b920008",
    15969 => x"379c0024", 15970 => x"c3a00000", 15971 => x"379cfffc",
    15972 => x"5b9d0004", 15973 => x"78010001", 15974 => x"38215798",
    15975 => x"fbfff351", 15976 => x"3401ffff", 15977 => x"2b9d0004",
    15978 => x"379c0004", 15979 => x"c3a00000", 15980 => x"379cfff8",
    15981 => x"5b8b0008", 15982 => x"5b9d0004", 15983 => x"78010001",
    15984 => x"b8405800", 15985 => x"78020001", 15986 => x"38425d78",
    15987 => x"382157bc", 15988 => x"fbfff344", 15989 => x"78020001",
    15990 => x"78010001", 15991 => x"38429188", 15992 => x"38219198",
    15993 => x"34460090", 15994 => x"34050022", 15995 => x"34040033",
    15996 => x"28220004", 15997 => x"204300ff", 15998 => x"7c670042",
    15999 => x"7c630028", 16000 => x"a0e31800", 16001 => x"5c60000b",
    16002 => x"28230000", 16003 => x"31650000", 16004 => x"31640001",
    16005 => x"31630002", 16006 => x"00430018", 16007 => x"31630003",
    16008 => x"00430010", 16009 => x"00420008", 16010 => x"31630004",
    16011 => x"31620005", 16012 => x"34210010", 16013 => x"5c26ffef",
    16014 => x"34010000", 16015 => x"2b9d0004", 16016 => x"2b8b0008",
    16017 => x"379c0008", 16018 => x"c3a00000", 16019 => x"379cffe8",
    16020 => x"5b8b0018", 16021 => x"5b8c0014", 16022 => x"5b8d0010",
    16023 => x"5b8e000c", 16024 => x"5b8f0008", 16025 => x"5b9d0004",
    16026 => x"780b0001", 16027 => x"b8207800", 16028 => x"b8407000",
    16029 => x"340d0008", 16030 => x"340c0001", 16031 => x"396b70dc",
    16032 => x"a18e1800", 16033 => x"29640008", 16034 => x"7c620000",
    16035 => x"b9e00800", 16036 => x"35adffff", 16037 => x"d8800000",
    16038 => x"3d8c0001", 16039 => x"5da0fff9", 16040 => x"2b9d0004",
    16041 => x"2b8b0018", 16042 => x"2b8c0014", 16043 => x"2b8d0010",
    16044 => x"2b8e000c", 16045 => x"2b8f0008", 16046 => x"379c0018",
    16047 => x"c3a00000", 16048 => x"379cffe8", 16049 => x"5b8b0018",
    16050 => x"5b8c0014", 16051 => x"5b8d0010", 16052 => x"5b8e000c",
    16053 => x"5b8f0008", 16054 => x"5b9d0004", 16055 => x"780b0001",
    16056 => x"b8207800", 16057 => x"340e0008", 16058 => x"340c0000",
    16059 => x"340d0001", 16060 => x"396b70dc", 16061 => x"29620004",
    16062 => x"b9e00800", 16063 => x"35ceffff", 16064 => x"d8400000",
    16065 => x"7c220000", 16066 => x"c8021000", 16067 => x"a1a21000",
    16068 => x"b9826000", 16069 => x"3dad0001", 16070 => x"5dc0fff7",
    16071 => x"34010064", 16072 => x"fbffe95b", 16073 => x"b9800800",
    16074 => x"2b9d0004", 16075 => x"2b8b0018", 16076 => x"2b8c0014",
    16077 => x"2b8d0010", 16078 => x"2b8e000c", 16079 => x"2b8f0008",
    16080 => x"379c0018", 16081 => x"c3a00000", 16082 => x"379cffc0",
    16083 => x"5b8b0040", 16084 => x"5b8c003c", 16085 => x"5b8d0038",
    16086 => x"5b8e0034", 16087 => x"5b8f0030", 16088 => x"5b90002c",
    16089 => x"5b910028", 16090 => x"5b920024", 16091 => x"5b930020",
    16092 => x"5b94001c", 16093 => x"5b950018", 16094 => x"5b960014",
    16095 => x"5b970010", 16096 => x"5b98000c", 16097 => x"5b990008",
    16098 => x"5b9d0004", 16099 => x"34020000", 16100 => x"b8206000",
    16101 => x"34030080", 16102 => x"34210008", 16103 => x"780d0001",
    16104 => x"f8000d47", 16105 => x"39ad70dc", 16106 => x"29a10000",
    16107 => x"340f0000", 16108 => x"44200061", 16109 => x"b9805800",
    16110 => x"34120000", 16111 => x"34110000", 16112 => x"78194000",
    16113 => x"34160001", 16114 => x"34180008", 16115 => x"596c0008",
    16116 => x"45e00022", 16117 => x"29610000", 16118 => x"78028000",
    16119 => x"34030000", 16120 => x"59610010", 16121 => x"29610004",
    16122 => x"59610014", 16123 => x"a0590800", 16124 => x"44200003",
    16125 => x"78024000", 16126 => x"34030000", 16127 => x"a0710800",
    16128 => x"a0522800", 16129 => x"b8a12800", 16130 => x"29640010",
    16131 => x"29610014", 16132 => x"5ca0000e", 16133 => x"a4603000",
    16134 => x"a0260800", 16135 => x"59610014", 16136 => x"00630001",
    16137 => x"3c41001f", 16138 => x"a4403800", 16139 => x"00420001",
    16140 => x"a0872000", 16141 => x"b8231800", 16142 => x"59640010",
    16143 => x"b8430800", 16144 => x"5c25ffeb", 16145 => x"e000003c",
    16146 => x"b8821000", 16147 => x"b8231800", 16148 => x"59620010",
    16149 => x"59630014", 16150 => x"35ee0001", 16151 => x"29a20000",
    16152 => x"3dce0004", 16153 => x"b9800800", 16154 => x"b58e7000",
    16155 => x"d8400000", 16156 => x"5c360031", 16157 => x"b9800800",
    16158 => x"340200f0", 16159 => x"fbffff74", 16160 => x"34140040",
    16161 => x"34130000", 16162 => x"34100001", 16163 => x"34120000",
    16164 => x"34110000", 16165 => x"29a20004", 16166 => x"b9800800",
    16167 => x"29d70004", 16168 => x"d8400000", 16169 => x"29a20004",
    16170 => x"b820a800", 16171 => x"b9800800", 16172 => x"a2f0b800",
    16173 => x"d8400000", 16174 => x"46a10008", 16175 => x"29a30008",
    16176 => x"baa01000", 16177 => x"7eb50000", 16178 => x"b9800800",
    16179 => x"d8600000", 16180 => x"5eb60011", 16181 => x"e0000007",
    16182 => x"29a30008", 16183 => x"b9800800", 16184 => x"bae01000",
    16185 => x"d8600000", 16186 => x"46e00009", 16187 => x"e000000a",
    16188 => x"29c10000", 16189 => x"b8330800", 16190 => x"59c10000",
    16191 => x"29c10004", 16192 => x"b8300800", 16193 => x"59c10004",
    16194 => x"e0000003", 16195 => x"ba539000", 16196 => x"ba308800",
    16197 => x"3e010001", 16198 => x"3e730001", 16199 => x"f6018000",
    16200 => x"3694ffff", 16201 => x"b6139800", 16202 => x"b8208000",
    16203 => x"5e80ffda", 16204 => x"e0000014", 16205 => x"b9e00800",
    16206 => x"2b9d0004", 16207 => x"2b8b0040", 16208 => x"2b8c003c",
    16209 => x"2b8d0038", 16210 => x"2b8e0034", 16211 => x"2b8f0030",
    16212 => x"2b90002c", 16213 => x"2b910028", 16214 => x"2b920024",
    16215 => x"2b930020", 16216 => x"2b94001c", 16217 => x"2b950018",
    16218 => x"2b960014", 16219 => x"2b970010", 16220 => x"2b98000c",
    16221 => x"2b990008", 16222 => x"379c0040", 16223 => x"c3a00000",
    16224 => x"35ef0001", 16225 => x"356b0010", 16226 => x"5df8ff91",
    16227 => x"e3ffffea", 16228 => x"379cfff0", 16229 => x"5b8b0010",
    16230 => x"5b8c000c", 16231 => x"5b8d0008", 16232 => x"5b9d0004",
    16233 => x"b8205800", 16234 => x"78010001", 16235 => x"382170dc",
    16236 => x"28220000", 16237 => x"29610000", 16238 => x"340c0000",
    16239 => x"340d0040", 16240 => x"d8400000", 16241 => x"29610000",
    16242 => x"34020055", 16243 => x"fbffff20", 16244 => x"29610008",
    16245 => x"2962000c", 16246 => x"b9801800", 16247 => x"358c0008",
    16248 => x"f8000b7c", 16249 => x"29610000", 16250 => x"fbffff19",
    16251 => x"5d8dfff9", 16252 => x"2b9d0004", 16253 => x"2b8b0010",
    16254 => x"2b8c000c", 16255 => x"2b8d0008", 16256 => x"379c0010",
    16257 => x"c3a00000", 16258 => x"28210000", 16259 => x"78020001",
    16260 => x"38429210", 16261 => x"28420000", 16262 => x"3c210008",
    16263 => x"3821000a", 16264 => x"58410000", 16265 => x"28410000",
    16266 => x"20230008", 16267 => x"5c60fffe", 16268 => x"20210001",
    16269 => x"18210001", 16270 => x"c3a00000", 16271 => x"28210000",
    16272 => x"78020001", 16273 => x"38429210", 16274 => x"28420000",
    16275 => x"3c210008", 16276 => x"38210009", 16277 => x"58410000",
    16278 => x"28410000", 16279 => x"20230008", 16280 => x"5c60fffe",
    16281 => x"20210001", 16282 => x"c3a00000", 16283 => x"28210000",
    16284 => x"78030001", 16285 => x"38639210", 16286 => x"3c210008",
    16287 => x"28630000", 16288 => x"7c420000", 16289 => x"38210008",
    16290 => x"b8221000", 16291 => x"58620000", 16292 => x"28610000",
    16293 => x"20210008", 16294 => x"5c20fffe", 16295 => x"c3a00000",
    16296 => x"78010001", 16297 => x"78030001", 16298 => x"38219210",
    16299 => x"386359d4", 16300 => x"28210000", 16301 => x"28620000",
    16302 => x"58220004", 16303 => x"c3a00000", 16304 => x"379cffc4",
    16305 => x"5b8b001c", 16306 => x"5b8c0018", 16307 => x"5b8d0014",
    16308 => x"5b8e0010", 16309 => x"5b8f000c", 16310 => x"5b900008",
    16311 => x"5b9d0004", 16312 => x"b8206000", 16313 => x"28210000",
    16314 => x"340bffff", 16315 => x"4420002a", 16316 => x"29820004",
    16317 => x"44400028", 16318 => x"fbffe819", 16319 => x"780e0001",
    16320 => x"b8206800", 16321 => x"340b0000", 16322 => x"3410001f",
    16323 => x"378f0020", 16324 => x"39ce57d8", 16325 => x"e000000b",
    16326 => x"fbffe811", 16327 => x"202400ff", 16328 => x"b56d1000",
    16329 => x"b5eb0800", 16330 => x"30240000", 16331 => x"b8401800",
    16332 => x"b9c00800", 16333 => x"b8802800", 16334 => x"fbfff1ea",
    16335 => x"356b0001", 16336 => x"29810004", 16337 => x"ee0b1800",
    16338 => x"358c0004", 16339 => x"7c220000", 16340 => x"a0621000",
    16341 => x"5c40fff1", 16342 => x"78010001", 16343 => x"b9602000",
    16344 => x"b9a01000", 16345 => x"b9e01800", 16346 => x"38219188",
    16347 => x"f80001cc", 16348 => x"b8206000", 16349 => x"b9601800",
    16350 => x"78010001", 16351 => x"fd8b5800", 16352 => x"382157fc",
    16353 => x"b9a01000", 16354 => x"b9802000", 16355 => x"fbfff1d5",
    16356 => x"c80b5800", 16357 => x"b9600800", 16358 => x"2b9d0004",
    16359 => x"2b8b001c", 16360 => x"2b8c0018", 16361 => x"2b8d0014",
    16362 => x"2b8e0010", 16363 => x"2b8f000c", 16364 => x"2b900008",
    16365 => x"379c003c", 16366 => x"c3a00000", 16367 => x"379cffc8",
    16368 => x"5b8b0018", 16369 => x"5b8c0014", 16370 => x"5b8d0010",
    16371 => x"5b8e000c", 16372 => x"5b8f0008", 16373 => x"5b9d0004",
    16374 => x"b8205800", 16375 => x"28210000", 16376 => x"3405ffff",
    16377 => x"4420002c", 16378 => x"29620004", 16379 => x"4440002a",
    16380 => x"fbffe7db", 16381 => x"b8207000", 16382 => x"29610004",
    16383 => x"fbffe7d8", 16384 => x"b8205800", 16385 => x"34010020",
    16386 => x"4c2b0002", 16387 => x"340b0020", 16388 => x"378d001c",
    16389 => x"78010001", 16390 => x"b9602000", 16391 => x"b9c01000",
    16392 => x"b9a01800", 16393 => x"38219188", 16394 => x"f8000189",
    16395 => x"b8206000", 16396 => x"78010001", 16397 => x"b9601800",
    16398 => x"3821581c", 16399 => x"b9c01000", 16400 => x"b9802000",
    16401 => x"fbfff1a7", 16402 => x"e98b5800", 16403 => x"ec0c0800",
    16404 => x"3405ffff", 16405 => x"b9615800", 16406 => x"5d60000f",
    16407 => x"b9a07800", 16408 => x"780d0001", 16409 => x"39ad57d8",
    16410 => x"b5eb0800", 16411 => x"40240000", 16412 => x"b56e1000",
    16413 => x"b9a00800", 16414 => x"b8401800", 16415 => x"b8802800",
    16416 => x"356b0001", 16417 => x"fbfff197", 16418 => x"498bfff8",
    16419 => x"fd8b2800", 16420 => x"c8052800", 16421 => x"b8a00800",
    16422 => x"2b9d0004", 16423 => x"2b8b0018", 16424 => x"2b8c0014",
    16425 => x"2b8d0010", 16426 => x"2b8e000c", 16427 => x"2b8f0008",
    16428 => x"379c0038", 16429 => x"c3a00000", 16430 => x"379cffe4",
    16431 => x"5b8b001c", 16432 => x"5b8c0018", 16433 => x"5b8d0014",
    16434 => x"5b8e0010", 16435 => x"5b8f000c", 16436 => x"5b900008",
    16437 => x"5b9d0004", 16438 => x"780d0001", 16439 => x"39ad9188",
    16440 => x"b9a00800", 16441 => x"780b0001", 16442 => x"780f0001",
    16443 => x"780e0001", 16444 => x"fbfffe96", 16445 => x"396b9198",
    16446 => x"340c0000", 16447 => x"39ef583c", 16448 => x"39ce5854",
    16449 => x"34100008", 16450 => x"29630000", 16451 => x"29640004",
    16452 => x"b8640800", 16453 => x"44200010", 16454 => x"b9801000",
    16455 => x"b9e00800", 16456 => x"fbfff170", 16457 => x"3d810004",
    16458 => x"34020000", 16459 => x"34210008", 16460 => x"b5a10800",
    16461 => x"f8000015", 16462 => x"2023ffff", 16463 => x"08632710",
    16464 => x"b8201000", 16465 => x"14420010", 16466 => x"14630010",
    16467 => x"b9c00800", 16468 => x"fbfff164", 16469 => x"358c0001",
    16470 => x"356b0010", 16471 => x"5d90ffeb", 16472 => x"34010000",
    16473 => x"2b9d0004", 16474 => x"2b8b001c", 16475 => x"2b8c0018",
    16476 => x"2b8d0014", 16477 => x"2b8e0010", 16478 => x"2b8f000c",
    16479 => x"2b900008", 16480 => x"379c001c", 16481 => x"c3a00000",
    16482 => x"379cffec", 16483 => x"5b8b0014", 16484 => x"5b8c0010",
    16485 => x"5b8d000c", 16486 => x"5b8e0008", 16487 => x"5b9d0004",
    16488 => x"402d000f", 16489 => x"b8206000", 16490 => x"34010028",
    16491 => x"b8407000", 16492 => x"45a10005", 16493 => x"34010042",
    16494 => x"45a10003", 16495 => x"34010010", 16496 => x"5da10034",
    16497 => x"21cb0002", 16498 => x"5d60000f", 16499 => x"b9800800",
    16500 => x"fbfffef0", 16501 => x"29810000", 16502 => x"34020044",
    16503 => x"21ce0001", 16504 => x"fbfffe1b", 16505 => x"34010000",
    16506 => x"5dcb002d", 16507 => x"780b0001", 16508 => x"396b70dc",
    16509 => x"29620004", 16510 => x"29810000", 16511 => x"d8400000",
    16512 => x"4420fffd", 16513 => x"b9800800", 16514 => x"fbfffee2",
    16515 => x"29810000", 16516 => x"780b0001", 16517 => x"340200be",
    16518 => x"396b8ec4", 16519 => x"fbfffe0c", 16520 => x"356e0008",
    16521 => x"e0000005", 16522 => x"29810000", 16523 => x"fbfffe25",
    16524 => x"31610000", 16525 => x"356b0001", 16526 => x"5d6efffc",
    16527 => x"78020001", 16528 => x"38428ec4", 16529 => x"40410001",
    16530 => x"40430000", 16531 => x"3c210008", 16532 => x"b8230800",
    16533 => x"34030028", 16534 => x"dc200800", 16535 => x"45a3000b",
    16536 => x"34030042", 16537 => x"45a30009", 16538 => x"34030010",
    16539 => x"5da3000b", 16540 => x"40420006", 16541 => x"3c21000f",
    16542 => x"3c42000c", 16543 => x"3421c000", 16544 => x"b8220800",
    16545 => x"e0000006", 16546 => x"3c21000c", 16547 => x"e0000004",
    16548 => x"78018000", 16549 => x"e0000002", 16550 => x"34010000",
    16551 => x"2b9d0004", 16552 => x"2b8b0014", 16553 => x"2b8c0010",
    16554 => x"2b8d000c", 16555 => x"2b8e0008", 16556 => x"379c0014",
    16557 => x"c3a00000", 16558 => x"379cfffc", 16559 => x"5b9d0004",
    16560 => x"34030000", 16561 => x"b8202000", 16562 => x"34090028",
    16563 => x"34080042", 16564 => x"34070010", 16565 => x"34060008",
    16566 => x"40850017", 16567 => x"44a90003", 16568 => x"44a80002",
    16569 => x"5ca70006", 16570 => x"3c630004", 16571 => x"34630008",
    16572 => x"b4230800", 16573 => x"fbffffa5", 16574 => x"e0000005",
    16575 => x"34630001", 16576 => x"34840010", 16577 => x"5c66fff5",
    16578 => x"78018000", 16579 => x"2b9d0004", 16580 => x"379c0004",
    16581 => x"c3a00000", 16582 => x"379cffe0", 16583 => x"5b8b0020",
    16584 => x"5b8c001c", 16585 => x"5b8d0018", 16586 => x"5b8e0014",
    16587 => x"5b8f0010", 16588 => x"5b90000c", 16589 => x"5b910008",
    16590 => x"5b9d0004", 16591 => x"b8205800", 16592 => x"b8408800",
    16593 => x"b8608000", 16594 => x"b8806000", 16595 => x"fbfffe91",
    16596 => x"29610000", 16597 => x"3402000f", 16598 => x"222e00ff",
    16599 => x"fbfffdbc", 16600 => x"29610000", 16601 => x"b9c01000",
    16602 => x"2231ff00", 16603 => x"fbfffdb8", 16604 => x"16310008",
    16605 => x"29610000", 16606 => x"ba201000", 16607 => x"340d0000",
    16608 => x"fbfffdb3", 16609 => x"e0000006", 16610 => x"b60d1000",
    16611 => x"29610000", 16612 => x"40420000", 16613 => x"35ad0001",
    16614 => x"fbfffdad", 16615 => x"498dfffb", 16616 => x"b9600800",
    16617 => x"fbfffe7b", 16618 => x"29610000", 16619 => x"340200aa",
    16620 => x"fbfffda7", 16621 => x"29610000", 16622 => x"fbfffdc2",
    16623 => x"b8207800", 16624 => x"5c2e0022", 16625 => x"29610000",
    16626 => x"fbfffdbe", 16627 => x"b8207000", 16628 => x"5c310020",
    16629 => x"29610000", 16630 => x"340d0000", 16631 => x"fbfffdb9",
    16632 => x"b8208800", 16633 => x"e0000007", 16634 => x"29610000",
    16635 => x"fbfffdb5", 16636 => x"b60d1000", 16637 => x"40420000",
    16638 => x"5c220018", 16639 => x"35ad0001", 16640 => x"498dfffa",
    16641 => x"b9600800", 16642 => x"fbfffe62", 16643 => x"29610000",
    16644 => x"34020055", 16645 => x"fbfffd8e", 16646 => x"29610000",
    16647 => x"b9e01000", 16648 => x"fbfffd8b", 16649 => x"29610000",
    16650 => x"b9c01000", 16651 => x"fbfffd88", 16652 => x"29610000",
    16653 => x"ba201000", 16654 => x"fbfffd85", 16655 => x"34012710",
    16656 => x"fbffe713", 16657 => x"e0000006", 16658 => x"340cffff",
    16659 => x"e0000004", 16660 => x"340cfffe", 16661 => x"e0000002",
    16662 => x"340cfffd", 16663 => x"b9800800", 16664 => x"2b9d0004",
    16665 => x"2b8b0020", 16666 => x"2b8c001c", 16667 => x"2b8d0018",
    16668 => x"2b8e0014", 16669 => x"2b8f0010", 16670 => x"2b90000c",
    16671 => x"2b910008", 16672 => x"379c0020", 16673 => x"c3a00000",
    16674 => x"379cffe4", 16675 => x"5b8b001c", 16676 => x"5b8c0018",
    16677 => x"5b8d0014", 16678 => x"5b8e0010", 16679 => x"5b8f000c",
    16680 => x"5b900008", 16681 => x"5b9d0004", 16682 => x"b8208000",
    16683 => x"2041001f", 16684 => x"b8405800", 16685 => x"b8607000",
    16686 => x"b8806000", 16687 => x"340d0000", 16688 => x"44200030",
    16689 => x"3441ffff", 16690 => x"b4240800", 16691 => x"1422001f",
    16692 => x"b8807800", 16693 => x"0042001b", 16694 => x"b4410800",
    16695 => x"1562001f", 16696 => x"14210005", 16697 => x"0042001b",
    16698 => x"b44b1000", 16699 => x"14420005", 16700 => x"4422000c",
    16701 => x"78010001", 16702 => x"382159d8", 16703 => x"28220000",
    16704 => x"a1621000", 16705 => x"4c400005", 16706 => x"3442ffff",
    16707 => x"3401ffe0", 16708 => x"b8411000", 16709 => x"34420001",
    16710 => x"340f0020", 16711 => x"c9e27800", 16712 => x"ba000800",
    16713 => x"b9601000", 16714 => x"b9c01800", 16715 => x"b9e02000",
    16716 => x"fbffff7a", 16717 => x"b8206800", 16718 => x"48010016",
    16719 => x"b5cf7000", 16720 => x"b56f5800", 16721 => x"c98f6000",
    16722 => x"e000000e", 16723 => x"b9802000", 16724 => x"4dec0002",
    16725 => x"34040020", 16726 => x"ba000800", 16727 => x"b9601000",
    16728 => x"b9c01800", 16729 => x"fbffff6d", 16730 => x"48010009",
    16731 => x"b5a16800", 16732 => x"35ce0020", 16733 => x"356b0020",
    16734 => x"358cffe0", 16735 => x"e0000002", 16736 => x"340f0020",
    16737 => x"4980fff2", 16738 => x"e0000002", 16739 => x"b8206800",
    16740 => x"b9a00800", 16741 => x"2b9d0004", 16742 => x"2b8b001c",
    16743 => x"2b8c0018", 16744 => x"2b8d0014", 16745 => x"2b8e0010",
    16746 => x"2b8f000c", 16747 => x"2b900008", 16748 => x"379c001c",
    16749 => x"c3a00000", 16750 => x"379cffec", 16751 => x"5b8b0014",
    16752 => x"5b8c0010", 16753 => x"5b8d000c", 16754 => x"5b8e0008",
    16755 => x"5b9d0004", 16756 => x"b8405800", 16757 => x"b8206000",
    16758 => x"b8607000", 16759 => x"b8806800", 16760 => x"fbfffdec",
    16761 => x"29810000", 16762 => x"340200f0", 16763 => x"fbfffd18",
    16764 => x"29810000", 16765 => x"216200ff", 16766 => x"fbfffd15",
    16767 => x"2162ff00", 16768 => x"29810000", 16769 => x"00420008",
    16770 => x"340b0000", 16771 => x"fbfffd10", 16772 => x"e0000006",
    16773 => x"29810000", 16774 => x"fbfffd2a", 16775 => x"b5cb1000",
    16776 => x"30410000", 16777 => x"356b0001", 16778 => x"49abfffb",
    16779 => x"b9a00800", 16780 => x"2b9d0004", 16781 => x"2b8b0014",
    16782 => x"2b8c0010", 16783 => x"2b8d000c", 16784 => x"2b8e0008",
    16785 => x"379c0014", 16786 => x"c3a00000", 16787 => x"379cfffc",
    16788 => x"5b9d0004", 16789 => x"34050000", 16790 => x"b8203000",
    16791 => x"34080043", 16792 => x"34070008", 16793 => x"40c90017",
    16794 => x"5d280006", 16795 => x"3ca50004", 16796 => x"34a50008",
    16797 => x"b4250800", 16798 => x"fbffffd0", 16799 => x"e0000005",
    16800 => x"34a50001", 16801 => x"34c60010", 16802 => x"5ca7fff7",
    16803 => x"3401ffff", 16804 => x"2b9d0004", 16805 => x"379c0004",
    16806 => x"c3a00000", 16807 => x"379cfffc", 16808 => x"5b9d0004",
    16809 => x"34050000", 16810 => x"b8203000", 16811 => x"34080043",
    16812 => x"34070008", 16813 => x"40c90017", 16814 => x"5d280006",
    16815 => x"3ca50004", 16816 => x"34a50008", 16817 => x"b4250800",
    16818 => x"fbffff70", 16819 => x"e0000005", 16820 => x"34a50001",
    16821 => x"34c60010", 16822 => x"5ca7fff7", 16823 => x"3401ffff",
    16824 => x"2b9d0004", 16825 => x"379c0004", 16826 => x"c3a00000",
    16827 => x"379cfff4", 16828 => x"5b8b000c", 16829 => x"5b8c0008",
    16830 => x"5b9d0004", 16831 => x"780b0001", 16832 => x"396b8ed4",
    16833 => x"29610000", 16834 => x"5c200009", 16835 => x"fbfff5b5",
    16836 => x"78020001", 16837 => x"342103e8", 16838 => x"38428ecc",
    16839 => x"58410000", 16840 => x"29610000", 16841 => x"34210001",
    16842 => x"59610000", 16843 => x"780b0001", 16844 => x"396b8ed0",
    16845 => x"296c0000", 16846 => x"fbfff5aa", 16847 => x"78020001",
    16848 => x"38428ecc", 16849 => x"28440000", 16850 => x"c8242800",
    16851 => x"34010000", 16852 => x"48050018", 16853 => x"21830001",
    16854 => x"78010001", 16855 => x"3c650002", 16856 => x"38215d8c",
    16857 => x"b4250800", 16858 => x"28210000", 16859 => x"b4242000",
    16860 => x"29610000", 16861 => x"58440000", 16862 => x"34020001",
    16863 => x"34210001", 16864 => x"59610000", 16865 => x"78010001",
    16866 => x"38219188", 16867 => x"44620003", 16868 => x"fbfffeca",
    16869 => x"e0000006", 16870 => x"34020002", 16871 => x"fbfffec7",
    16872 => x"78020001", 16873 => x"384270e8", 16874 => x"58410004",
    16875 => x"34010001", 16876 => x"2b9d0004", 16877 => x"2b8b000c",
    16878 => x"2b8c0008", 16879 => x"379c000c", 16880 => x"c3a00000",
    16881 => x"78010001", 16882 => x"38219240", 16883 => x"28220000",
    16884 => x"78010001", 16885 => x"3821926c", 16886 => x"58220000",
    16887 => x"340103c6", 16888 => x"58410004", 16889 => x"c3a00000",
    16890 => x"c3a00000", 16891 => x"379cfff8", 16892 => x"5b8b0008",
    16893 => x"5b9d0004", 16894 => x"b8205800", 16895 => x"3401000a",
    16896 => x"5d610003", 16897 => x"3401000d", 16898 => x"fbfffff9",
    16899 => x"78020001", 16900 => x"3842926c", 16901 => x"28420000",
    16902 => x"28410000", 16903 => x"20210001", 16904 => x"5c20fffe",
    16905 => x"584b0008", 16906 => x"2b9d0004", 16907 => x"2b8b0008",
    16908 => x"379c0008", 16909 => x"c3a00000", 16910 => x"379cfff4",
    16911 => x"5b8b000c", 16912 => x"5b8c0008", 16913 => x"5b9d0004",
    16914 => x"b8206000", 16915 => x"b8205800", 16916 => x"e0000004",
    16917 => x"b8400800", 16918 => x"356b0001", 16919 => x"fbffffe4",
    16920 => x"41620000", 16921 => x"5c40fffc", 16922 => x"c96c0800",
    16923 => x"2b9d0004", 16924 => x"2b8b000c", 16925 => x"2b8c0008",
    16926 => x"379c000c", 16927 => x"c3a00000", 16928 => x"78010001",
    16929 => x"3821926c", 16930 => x"28220000", 16931 => x"3401ffff",
    16932 => x"28430000", 16933 => x"20630002", 16934 => x"44600003",
    16935 => x"2841000c", 16936 => x"202100ff", 16937 => x"c3a00000",
    16938 => x"28250008", 16939 => x"28240000", 16940 => x"28260004",
    16941 => x"b4451800", 16942 => x"88642000", 16943 => x"5822001c",
    16944 => x"88461000", 16945 => x"b4821000", 16946 => x"2824000c",
    16947 => x"1442000c", 16948 => x"b4442000", 16949 => x"28220014",
    16950 => x"4c820005", 16951 => x"28240010", 16952 => x"44800008",
    16953 => x"4ca3000b", 16954 => x"e0000006", 16955 => x"28220018",
    16956 => x"4c440006", 16957 => x"28240010", 16958 => x"44800002",
    16959 => x"4c650005", 16960 => x"58230008", 16961 => x"e0000003",
    16962 => x"58230008", 16963 => x"b8801000", 16964 => x"58220020",
    16965 => x"b8400800", 16966 => x"c3a00000", 16967 => x"2822000c",
    16968 => x"58200008", 16969 => x"58220020", 16970 => x"c3a00000",
    16971 => x"379cfff8", 16972 => x"5b8b0008", 16973 => x"5b9d0004",
    16974 => x"b8205800", 16975 => x"58200014", 16976 => x"b8400800",
    16977 => x"f800093b", 16978 => x"2963000c", 16979 => x"29620000",
    16980 => x"4823000b", 16981 => x"29610004", 16982 => x"4c410003",
    16983 => x"34420001", 16984 => x"59620000", 16985 => x"29620000",
    16986 => x"5c410011", 16987 => x"34010001", 16988 => x"59610014",
    16989 => x"59610010", 16990 => x"e000000e", 16991 => x"29610008",
    16992 => x"4c220003", 16993 => x"3442ffff", 16994 => x"59620000",
    16995 => x"29620000", 16996 => x"5c410007", 16997 => x"34010001",
    16998 => x"59610014", 16999 => x"59600000", 17000 => x"59600010",
    17001 => x"3401ffff", 17002 => x"e0000002", 17003 => x"29610010",
    17004 => x"2b9d0004", 17005 => x"2b8b0008", 17006 => x"379c0008",
    17007 => x"c3a00000", 17008 => x"58200010", 17009 => x"58200000",
    17010 => x"58200014", 17011 => x"c3a00000", 17012 => x"78030001",
    17013 => x"3863924c", 17014 => x"28640000", 17015 => x"48810013",
    17016 => x"78030001", 17017 => x"38638ee8", 17018 => x"c8240800",
    17019 => x"44400007", 17020 => x"28620000", 17021 => x"34040001",
    17022 => x"bc810800", 17023 => x"28430028", 17024 => x"b8230800",
    17025 => x"e0000007", 17026 => x"28620000", 17027 => x"34040001",
    17028 => x"bc810800", 17029 => x"28430028", 17030 => x"a4200800",
    17031 => x"a0230800", 17032 => x"58410028", 17033 => x"c3a00000",
    17034 => x"78030001", 17035 => x"38638ee8", 17036 => x"44400007",
    17037 => x"28620000", 17038 => x"34040001", 17039 => x"bc810800",
    17040 => x"28430024", 17041 => x"b8230800", 17042 => x"e0000007",
    17043 => x"28620000", 17044 => x"34040001", 17045 => x"bc810800",
    17046 => x"28430024", 17047 => x"a4200800", 17048 => x"a0230800",
    17049 => x"58410024", 17050 => x"c3a00000", 17051 => x"379cfff0",
    17052 => x"5b8b0010", 17053 => x"5b8c000c", 17054 => x"5b8d0008",
    17055 => x"5b9d0004", 17056 => x"b8406800", 17057 => x"b8606000",
    17058 => x"34020000", 17059 => x"34030028", 17060 => x"b8205800",
    17061 => x"f800098a", 17062 => x"b9600800", 17063 => x"b9a01000",
    17064 => x"34030014", 17065 => x"f8000908", 17066 => x"596c0014",
    17067 => x"2b9d0004", 17068 => x"2b8b0010", 17069 => x"2b8c000c",
    17070 => x"2b8d0008", 17071 => x"379c0010", 17072 => x"c3a00000",
    17073 => x"b8201800", 17074 => x"e0000004", 17075 => x"28840000",
    17076 => x"34630008", 17077 => x"44820006", 17078 => x"28610004",
    17079 => x"b8602000", 17080 => x"5c20fffb", 17081 => x"78010001",
    17082 => x"38215870", 17083 => x"c3a00000", 17084 => x"78020001",
    17085 => x"38428ee8", 17086 => x"28420000", 17087 => x"b8201800",
    17088 => x"34010000", 17089 => x"28440008", 17090 => x"20840002",
    17091 => x"4480000c", 17092 => x"34040002", 17093 => x"58440008",
    17094 => x"78060001", 17095 => x"28420010", 17096 => x"38c659dc",
    17097 => x"28c40000", 17098 => x"3445ff9b", 17099 => x"54a40004",
    17100 => x"08420064", 17101 => x"34010001", 17102 => x"58620000",
    17103 => x"c3a00000", 17104 => x"379cfff0", 17105 => x"5b8b0010",
    17106 => x"5b8c000c", 17107 => x"5b8d0008", 17108 => x"5b9d0004",
    17109 => x"780b0001", 17110 => x"b8206000", 17111 => x"78010001",
    17112 => x"396b924c", 17113 => x"38219244", 17114 => x"28210000",
    17115 => x"296d0000", 17116 => x"b42d6800", 17117 => x"29810000",
    17118 => x"b9a01000", 17119 => x"f8000114", 17120 => x"29810004",
    17121 => x"29630000", 17122 => x"b9a01000", 17123 => x"f8000199",
    17124 => x"5980000c", 17125 => x"59800008", 17126 => x"2b9d0004",
    17127 => x"2b8b0010", 17128 => x"2b8c000c", 17129 => x"2b8d0008",
    17130 => x"379c0010", 17131 => x"c3a00000", 17132 => x"379cfff8",
    17133 => x"5b8b0008", 17134 => x"5b9d0004", 17135 => x"b8205800",
    17136 => x"28210000", 17137 => x"f800016c", 17138 => x"78010001",
    17139 => x"38218ee8", 17140 => x"28210000", 17141 => x"34020001",
    17142 => x"34030009", 17143 => x"58220004", 17144 => x"5963000c",
    17145 => x"78030001", 17146 => x"386359e0", 17147 => x"59620008",
    17148 => x"28620000", 17149 => x"5822004c", 17150 => x"2b9d0004",
    17151 => x"2b8b0008", 17152 => x"379c0008", 17153 => x"c3a00000",
    17154 => x"b8201000", 17155 => x"28210000", 17156 => x"2823004c",
    17157 => x"34010000", 17158 => x"44600016", 17159 => x"28430004",
    17160 => x"28630038", 17161 => x"44600013", 17162 => x"78030001",
    17163 => x"38638ee8", 17164 => x"28630000", 17165 => x"28640004",
    17166 => x"20840004", 17167 => x"4480000d", 17168 => x"28630004",
    17169 => x"20630008", 17170 => x"5c60000a", 17171 => x"2842000c",
    17172 => x"3403000a", 17173 => x"34010001", 17174 => x"54430006",
    17175 => x"78010001", 17176 => x"3c420002", 17177 => x"38215dbc",
    17178 => x"b4220800", 17179 => x"28210000", 17180 => x"c3a00000",
    17181 => x"379cfff0", 17182 => x"5b8b000c", 17183 => x"5b8c0008",
    17184 => x"5b9d0004", 17185 => x"2822000c", 17186 => x"b8205800",
    17187 => x"34010009", 17188 => x"3442ffff", 17189 => x"340c0000",
    17190 => x"544100a5", 17191 => x"78010001", 17192 => x"3c420002",
    17193 => x"38215d94", 17194 => x"b4220800", 17195 => x"28210000",
    17196 => x"c0200000", 17197 => x"78010001", 17198 => x"38218ee8",
    17199 => x"28210000", 17200 => x"340c0000", 17201 => x"28220004",
    17202 => x"20420008", 17203 => x"5c400098", 17204 => x"28230004",
    17205 => x"78028000", 17206 => x"b8621000", 17207 => x"58220004",
    17208 => x"3401000a", 17209 => x"e0000090", 17210 => x"78010001",
    17211 => x"38218ee8", 17212 => x"28210000", 17213 => x"78040001",
    17214 => x"38845994", 17215 => x"28230004", 17216 => x"28820000",
    17217 => x"a0621000", 17218 => x"58220004", 17219 => x"28220004",
    17220 => x"20420008", 17221 => x"5c400083", 17222 => x"28210004",
    17223 => x"340c0001", 17224 => x"20210004", 17225 => x"44220082",
    17226 => x"596c000c", 17227 => x"e0000080", 17228 => x"29610000",
    17229 => x"340c0000", 17230 => x"2821004c", 17231 => x"4420007c",
    17232 => x"fbffbd22", 17233 => x"29610004", 17234 => x"f8000151",
    17235 => x"fbffbd28", 17236 => x"34010008", 17237 => x"e0000074",
    17238 => x"78010001", 17239 => x"38218ee8", 17240 => x"28210000",
    17241 => x"34020002", 17242 => x"340c0000", 17243 => x"58220008",
    17244 => x"29610000", 17245 => x"2821004c", 17246 => x"4420006d",
    17247 => x"29610004", 17248 => x"28210038", 17249 => x"4420006a",
    17250 => x"78010001", 17251 => x"38218efc", 17252 => x"28210000",
    17253 => x"340300a2", 17254 => x"58230000", 17255 => x"34030003",
    17256 => x"58230010", 17257 => x"34030001", 17258 => x"5823001c",
    17259 => x"5962000c", 17260 => x"e000005e", 17261 => x"78010001",
    17262 => x"38218efc", 17263 => x"28210000", 17264 => x"340c0000",
    17265 => x"2822001c", 17266 => x"20420001", 17267 => x"44400058",
    17268 => x"34020002", 17269 => x"5822001c", 17270 => x"fbfff402",
    17271 => x"342107d0", 17272 => x"59610010", 17273 => x"34010003",
    17274 => x"e000004f", 17275 => x"fbfff3fd", 17276 => x"29620010",
    17277 => x"340c0000", 17278 => x"c8220800", 17279 => x"4801004c",
    17280 => x"34010007", 17281 => x"5961000c", 17282 => x"5960001c",
    17283 => x"e0000047", 17284 => x"37810010", 17285 => x"fbffff37",
    17286 => x"340c0000", 17287 => x"44200044", 17288 => x"78030001",
    17289 => x"386359e4", 17290 => x"28620000", 17291 => x"2b810010",
    17292 => x"f80007a4", 17293 => x"3802c34f", 17294 => x"e8221000",
    17295 => x"64210000", 17296 => x"b8410800", 17297 => x"44200005",
    17298 => x"34010064", 17299 => x"59610014", 17300 => x"3401ff9c",
    17301 => x"e0000003", 17302 => x"59600014", 17303 => x"34010064",
    17304 => x"59610018", 17305 => x"34010004", 17306 => x"e000002f",
    17307 => x"29610004", 17308 => x"340c0000", 17309 => x"f80001df",
    17310 => x"5c20002d", 17311 => x"37810010", 17312 => x"fbffff1c",
    17313 => x"442c002a", 17314 => x"78040001", 17315 => x"388459e4",
    17316 => x"2b810010", 17317 => x"28820000", 17318 => x"f800078a",
    17319 => x"29620014", 17320 => x"5b810010", 17321 => x"44220009",
    17322 => x"2961001c", 17323 => x"29620018", 17324 => x"b4410800",
    17325 => x"5961001c", 17326 => x"29610004", 17327 => x"2962001c",
    17328 => x"f80001aa", 17329 => x"e0000019", 17330 => x"29620014",
    17331 => x"340c0001", 17332 => x"5c220017", 17333 => x"2961001c",
    17334 => x"34217530", 17335 => x"5961001c", 17336 => x"29610004",
    17337 => x"2962001c", 17338 => x"f80001a0", 17339 => x"34010005",
    17340 => x"5961000c", 17341 => x"e000000e", 17342 => x"29610004",
    17343 => x"340c0000", 17344 => x"f80001bc", 17345 => x"5c20000a",
    17346 => x"34010006", 17347 => x"e0000006", 17348 => x"b9600800",
    17349 => x"fbffff3d", 17350 => x"340c0000", 17351 => x"5c200004",
    17352 => x"34010009", 17353 => x"5961000c", 17354 => x"340c0001",
    17355 => x"b9800800", 17356 => x"2b9d0004", 17357 => x"2b8b000c",
    17358 => x"2b8c0008", 17359 => x"379c0010", 17360 => x"c3a00000",
    17361 => x"78040001", 17362 => x"64630000", 17363 => x"38848ee8",
    17364 => x"28850000", 17365 => x"c8031800", 17366 => x"78048000",
    17367 => x"78060001", 17368 => x"a0641800", 17369 => x"38c659e8",
    17370 => x"b4641800", 17371 => x"28c40000", 17372 => x"3c210018",
    17373 => x"a0441000", 17374 => x"b8410800", 17375 => x"b8231800",
    17376 => x"58a3004c", 17377 => x"c3a00000", 17378 => x"78040001",
    17379 => x"64630000", 17380 => x"38848ee8", 17381 => x"28850000",
    17382 => x"c8031800", 17383 => x"78048000", 17384 => x"78060001",
    17385 => x"a0641800", 17386 => x"38c659e8", 17387 => x"b4641800",
    17388 => x"28c40000", 17389 => x"3c210018", 17390 => x"a0441000",
    17391 => x"b8410800", 17392 => x"b8231800", 17393 => x"58a3004c",
    17394 => x"c3a00000", 17395 => x"34030005", 17396 => x"5823002c",
    17397 => x"3803fffb", 17398 => x"58230030", 17399 => x"3403ff6a",
    17400 => x"5823001c", 17401 => x"3403fffe", 17402 => x"58230018",
    17403 => x"34030001", 17404 => x"58230028", 17405 => x"340300c8",
    17406 => x"58230048", 17407 => x"34032710", 17408 => x"58230040",
    17409 => x"34030064", 17410 => x"58230044", 17411 => x"5822000c",
    17412 => x"58200014", 17413 => x"c3a00000", 17414 => x"379cfff0",
    17415 => x"5b8b0010", 17416 => x"5b8c000c", 17417 => x"5b8d0008",
    17418 => x"5b9d0004", 17419 => x"b8205800", 17420 => x"2821000c",
    17421 => x"b8406800", 17422 => x"340c0000", 17423 => x"5c610047",
    17424 => x"34010022", 17425 => x"34030000", 17426 => x"fbffffbf",
    17427 => x"29620004", 17428 => x"34010025", 17429 => x"34030000",
    17430 => x"fbffffbb", 17431 => x"29610008", 17432 => x"4c200004",
    17433 => x"596d0004", 17434 => x"596d0008", 17435 => x"e000003b",
    17436 => x"4da10005", 17437 => x"29620000", 17438 => x"78010040",
    17439 => x"b4410800", 17440 => x"59610000", 17441 => x"29630000",
    17442 => x"78050001", 17443 => x"29620004", 17444 => x"38a559ec",
    17445 => x"28a10000", 17446 => x"b5a32000", 17447 => x"c8826000",
    17448 => x"482c0006", 17449 => x"78050001", 17450 => x"38a559f0",
    17451 => x"28a10000", 17452 => x"49810002", 17453 => x"e0000002",
    17454 => x"b8206000", 17455 => x"78050001", 17456 => x"38a559f4",
    17457 => x"28a10000", 17458 => x"4c240006", 17459 => x"4c220005",
    17460 => x"c8611800", 17461 => x"c8410800", 17462 => x"59630000",
    17463 => x"59610004", 17464 => x"29610004", 17465 => x"b9801000",
    17466 => x"596d0008", 17467 => x"34214000", 17468 => x"59610004",
    17469 => x"35610018", 17470 => x"fbfffdec", 17471 => x"78030001",
    17472 => x"38638ee8", 17473 => x"29620010", 17474 => x"b8206800",
    17475 => x"28610000", 17476 => x"34030000", 17477 => x"582d0040",
    17478 => x"34410001", 17479 => x"59610010", 17480 => x"34010026",
    17481 => x"fbffff88", 17482 => x"34010020", 17483 => x"b9a01000",
    17484 => x"34030000", 17485 => x"fbffff84", 17486 => x"b9801000",
    17487 => x"34010021", 17488 => x"34030001", 17489 => x"fbffff80",
    17490 => x"b9801000", 17491 => x"3561003c", 17492 => x"fbfffdf7",
    17493 => x"7c2c0000", 17494 => x"b9800800", 17495 => x"2b9d0004",
    17496 => x"2b8b0010", 17497 => x"2b8c000c", 17498 => x"2b8d0008",
    17499 => x"379c0010", 17500 => x"c3a00000", 17501 => x"379cfff8",
    17502 => x"5b8b0008", 17503 => x"5b9d0004", 17504 => x"b8205800",
    17505 => x"2821002c", 17506 => x"59600004", 17507 => x"59600000",
    17508 => x"59610024", 17509 => x"3401ffff", 17510 => x"59610008",
    17511 => x"59600010", 17512 => x"35610018", 17513 => x"fbfffdde",
    17514 => x"3561003c", 17515 => x"fbfffe05", 17516 => x"78020001",
    17517 => x"35610054", 17518 => x"34030010", 17519 => x"38425de8",
    17520 => x"fbfffe2b", 17521 => x"2961000c", 17522 => x"34020001",
    17523 => x"fbfffe01", 17524 => x"34010024", 17525 => x"34020001",
    17526 => x"34030001", 17527 => x"fbffff5a", 17528 => x"2b9d0004",
    17529 => x"2b8b0008", 17530 => x"379c0008", 17531 => x"c3a00000",
    17532 => x"379cfff8", 17533 => x"5b8b0008", 17534 => x"5b9d0004",
    17535 => x"b8205800", 17536 => x"34010005", 17537 => x"59610018",
    17538 => x"3801fffa", 17539 => x"5961001c", 17540 => x"34010001",
    17541 => x"59610014", 17542 => x"34017530", 17543 => x"59610010",
    17544 => x"3401fbb4", 17545 => x"59610008", 17546 => x"3401ffe2",
    17547 => x"59610004", 17548 => x"340104b0", 17549 => x"59610034",
    17550 => x"340103e8", 17551 => x"5961002c", 17552 => x"34010064",
    17553 => x"59610030", 17554 => x"78010001", 17555 => x"3821924c",
    17556 => x"28210000", 17557 => x"59630074", 17558 => x"59620070",
    17559 => x"c8611800", 17560 => x"59630080", 17561 => x"35610004",
    17562 => x"5960007c", 17563 => x"59600084", 17564 => x"fbfffdab",
    17565 => x"35610028", 17566 => x"fbfffdd2", 17567 => x"2b9d0004",
    17568 => x"2b8b0008", 17569 => x"379c0008", 17570 => x"c3a00000",
    17571 => x"379cfff8", 17572 => x"5b8b0008", 17573 => x"5b9d0004",
    17574 => x"b8205800", 17575 => x"58200044", 17576 => x"58200040",
    17577 => x"3401ffff", 17578 => x"59610048", 17579 => x"5961004c",
    17580 => x"59610050", 17581 => x"59610054", 17582 => x"34010001",
    17583 => x"59610084", 17584 => x"59600058", 17585 => x"35610004",
    17586 => x"5960005c", 17587 => x"59600060", 17588 => x"59600068",
    17589 => x"5960006c", 17590 => x"59600078", 17591 => x"fbfffd90",
    17592 => x"35610028", 17593 => x"fbfffdb7", 17594 => x"29610070",
    17595 => x"34020001", 17596 => x"fbfffdb8", 17597 => x"29610074",
    17598 => x"34020001", 17599 => x"fbfffdb5", 17600 => x"34010004",
    17601 => x"34020001", 17602 => x"34030001", 17603 => x"fbffff1f",
    17604 => x"2b9d0004", 17605 => x"2b8b0008", 17606 => x"379c0008",
    17607 => x"c3a00000", 17608 => x"379cfff8", 17609 => x"5b8b0008",
    17610 => x"5b9d0004", 17611 => x"b8205800", 17612 => x"28210074",
    17613 => x"34020000", 17614 => x"fbfffda6", 17615 => x"59600084",
    17616 => x"2b9d0004", 17617 => x"2b8b0008", 17618 => x"379c0008",
    17619 => x"c3a00000", 17620 => x"379cfff0", 17621 => x"5b8b0010",
    17622 => x"5b8c000c", 17623 => x"5b8d0008", 17624 => x"5b9d0004",
    17625 => x"28240084", 17626 => x"b8205800", 17627 => x"34010001",
    17628 => x"44800078", 17629 => x"29610070", 17630 => x"5c610002",
    17631 => x"59620048", 17632 => x"29610074", 17633 => x"5c610002",
    17634 => x"5962004c", 17635 => x"29610048", 17636 => x"48010009",
    17637 => x"29620050", 17638 => x"48020006", 17639 => x"4c220005",
    17640 => x"29630040", 17641 => x"78020040", 17642 => x"b4621000",
    17643 => x"59620040", 17644 => x"59610050", 17645 => x"2961004c",
    17646 => x"48010009", 17647 => x"29620054", 17648 => x"48020006",
    17649 => x"4c220005", 17650 => x"29630044", 17651 => x"78020040",
    17652 => x"b4621000", 17653 => x"59620044", 17654 => x"59610054",
    17655 => x"29630048", 17656 => x"34010000", 17657 => x"4803005b",
    17658 => x"2962004c", 17659 => x"48020059", 17660 => x"296c0040",
    17661 => x"29610038", 17662 => x"b46c1800", 17663 => x"296c0044",
    17664 => x"c8621000", 17665 => x"c84c6000", 17666 => x"44200006",
    17667 => x"218c3fff", 17668 => x"21812000", 17669 => x"44200003",
    17670 => x"3401c000", 17671 => x"b9816000", 17672 => x"b9801000",
    17673 => x"35610004", 17674 => x"fbfffd20", 17675 => x"29620080",
    17676 => x"78030001", 17677 => x"38638ee8", 17678 => x"2042000f",
    17679 => x"b8206800", 17680 => x"3c420010", 17681 => x"28610000",
    17682 => x"21a3ffff", 17683 => x"b8621000", 17684 => x"58220044",
    17685 => x"29630040", 17686 => x"29620048", 17687 => x"34010005",
    17688 => x"b4621000", 17689 => x"34030000", 17690 => x"fbfffec8",
    17691 => x"29630044", 17692 => x"2962004c", 17693 => x"34010002",
    17694 => x"b4621000", 17695 => x"34030000", 17696 => x"fbfffec2",
    17697 => x"34010001", 17698 => x"b9801000", 17699 => x"34030000",
    17700 => x"fbfffebe", 17701 => x"29620078", 17702 => x"34030000",
    17703 => x"34410001", 17704 => x"59610078", 17705 => x"34010006",
    17706 => x"fbfffeb8", 17707 => x"34010000", 17708 => x"b9a01000",
    17709 => x"34030001", 17710 => x"fbfffeb4", 17711 => x"78020001",
    17712 => x"3401ffff", 17713 => x"384259f8", 17714 => x"5961004c",
    17715 => x"59610048", 17716 => x"29630040", 17717 => x"28410000",
    17718 => x"4c23000a", 17719 => x"29620044", 17720 => x"4c220008",
    17721 => x"78040001", 17722 => x"388459fc", 17723 => x"28810000",
    17724 => x"b4611800", 17725 => x"b4410800", 17726 => x"59630040",
    17727 => x"59610044", 17728 => x"29610038", 17729 => x"4420000f",
    17730 => x"2961006c", 17731 => x"29620068", 17732 => x"4c220006",
    17733 => x"34210001", 17734 => x"5961006c", 17735 => x"29610040",
    17736 => x"3421ffff", 17737 => x"e0000006", 17738 => x"4c410006",
    17739 => x"3421ffff", 17740 => x"5961006c", 17741 => x"29610040",
    17742 => x"34210001", 17743 => x"59610040", 17744 => x"35610028",
    17745 => x"b9801000", 17746 => x"fbfffcf9", 17747 => x"7c210000",
    17748 => x"2b9d0004", 17749 => x"2b8b0010", 17750 => x"2b8c000c",
    17751 => x"2b8d0008", 17752 => x"379c0010", 17753 => x"c3a00000",
    17754 => x"379cfff0", 17755 => x"5b8b0008", 17756 => x"5b9d0004",
    17757 => x"b8205800", 17758 => x"1443001f", 17759 => x"3781000c",
    17760 => x"4802000b", 17761 => x"00440012", 17762 => x"3c63000e",
    17763 => x"3c42000e", 17764 => x"b8641800", 17765 => x"5b820010",
    17766 => x"34021f40", 17767 => x"5b83000c", 17768 => x"fbffc11e",
    17769 => x"2b820010", 17770 => x"e0000009", 17771 => x"0842c000",
    17772 => x"5b820010", 17773 => x"1442001f", 17774 => x"5b82000c",
    17775 => x"34021f40", 17776 => x"fbffc116", 17777 => x"2b820010",
    17778 => x"c8021000", 17779 => x"0041001f", 17780 => x"b4221000",
    17781 => x"14420001", 17782 => x"34010000", 17783 => x"59620068",
    17784 => x"2b9d0004", 17785 => x"2b8b0008", 17786 => x"379c0010",
    17787 => x"c3a00000", 17788 => x"28220068", 17789 => x"2821006c",
    17790 => x"fc410800", 17791 => x"c3a00000", 17792 => x"58220004",
    17793 => x"5820001c", 17794 => x"58230008", 17795 => x"5820000c",
    17796 => x"58200010", 17797 => x"58200000", 17798 => x"c3a00000",
    17799 => x"379cfffc", 17800 => x"5b9d0004", 17801 => x"34020001",
    17802 => x"58220000", 17803 => x"58200014", 17804 => x"5820001c",
    17805 => x"5820000c", 17806 => x"58200010", 17807 => x"28210004",
    17808 => x"fbfffce4", 17809 => x"78010001", 17810 => x"3821924c",
    17811 => x"28210000", 17812 => x"34020001", 17813 => x"fbfffcdf",
    17814 => x"2b9d0004", 17815 => x"379c0004", 17816 => x"c3a00000",
    17817 => x"379cffb0", 17818 => x"5b8b0010", 17819 => x"5b8c000c",
    17820 => x"5b8d0008", 17821 => x"5b9d0004", 17822 => x"b8205800",
    17823 => x"b8406000", 17824 => x"b8606800", 17825 => x"37810014",
    17826 => x"34020000", 17827 => x"34030040", 17828 => x"f800068b",
    17829 => x"3401c000", 17830 => x"78040001", 17831 => x"5b810020",
    17832 => x"3884924c", 17833 => x"34014000", 17834 => x"5b810044",
    17835 => x"28810000", 17836 => x"5da10005", 17837 => x"78030001",
    17838 => x"386371fc", 17839 => x"586c0000", 17840 => x"e0000027",
    17841 => x"3dad0005", 17842 => x"b56d5800", 17843 => x"29610000",
    17844 => x"44200023", 17845 => x"78030001", 17846 => x"386371fc",
    17847 => x"28610000", 17848 => x"29620010", 17849 => x"c9810800",
    17850 => x"20213fff", 17851 => x"1423000c", 17852 => x"5c400007",
    17853 => x"3c630002", 17854 => x"5961000c", 17855 => x"34010001",
    17856 => x"59630014", 17857 => x"59610010", 17858 => x"e0000015",
    17859 => x"2964000c", 17860 => x"34420001", 17861 => x"b4240800",
    17862 => x"29640014", 17863 => x"b4641800", 17864 => x"3c630002",
    17865 => x"37840050", 17866 => x"b4831800", 17867 => x"2863ffc4",
    17868 => x"59620010", 17869 => x"b4230800", 17870 => x"29630008",
    17871 => x"5961000c", 17872 => x"5c430007", 17873 => x"f8000532",
    17874 => x"59610018", 17875 => x"34010001", 17876 => x"5961001c",
    17877 => x"5960000c", 17878 => x"59600010", 17879 => x"34010000",
    17880 => x"2b9d0004", 17881 => x"2b8b0010", 17882 => x"2b8c000c",
    17883 => x"2b8d0008", 17884 => x"379c0050", 17885 => x"c3a00000",
    17886 => x"78030001", 17887 => x"38638ee8", 17888 => x"5c40000a",
    17889 => x"34040001", 17890 => x"28620000", 17891 => x"bc810800",
    17892 => x"202100ff", 17893 => x"28430020", 17894 => x"3c210010",
    17895 => x"a4200800", 17896 => x"a0230800", 17897 => x"e0000008",
    17898 => x"28620000", 17899 => x"34040001", 17900 => x"bc810800",
    17901 => x"28430020", 17902 => x"202100ff", 17903 => x"3c210010",
    17904 => x"b8230800", 17905 => x"58410020", 17906 => x"c3a00000",
    17907 => x"379cfff8", 17908 => x"5b8b0008", 17909 => x"5b9d0004",
    17910 => x"34020001", 17911 => x"44220009", 17912 => x"34020002",
    17913 => x"4422000c", 17914 => x"5c200017", 17915 => x"78010001",
    17916 => x"38218ee8", 17917 => x"282b0000", 17918 => x"356b0018",
    17919 => x"e000000a", 17920 => x"78010001", 17921 => x"38218ee8",
    17922 => x"282b0000", 17923 => x"356b0014", 17924 => x"e0000005",
    17925 => x"78010001", 17926 => x"38218ee8", 17927 => x"282b0000",
    17928 => x"356b001c", 17929 => x"340107d0", 17930 => x"fbfff173",
    17931 => x"78030001", 17932 => x"386359b4", 17933 => x"29620000",
    17934 => x"28610000", 17935 => x"a0410800", 17936 => x"e0000002",
    17937 => x"34010000", 17938 => x"2b9d0004", 17939 => x"2b8b0008",
    17940 => x"379c0008", 17941 => x"c3a00000", 17942 => x"379cfff8",
    17943 => x"5b8b0008", 17944 => x"5b9d0004", 17945 => x"b8201800",
    17946 => x"78010001", 17947 => x"b8405800", 17948 => x"38218fbc",
    17949 => x"44600007", 17950 => x"3461ffff", 17951 => x"08210090",
    17952 => x"78030001", 17953 => x"38638f04", 17954 => x"34210148",
    17955 => x"b4230800", 17956 => x"b9601000", 17957 => x"fbffff35",
    17958 => x"78010001", 17959 => x"38218f04", 17960 => x"582b0018",
    17961 => x"2b9d0004", 17962 => x"2b8b0008", 17963 => x"379c0008",
    17964 => x"c3a00000", 17965 => x"379cffec", 17966 => x"5b8b0014",
    17967 => x"5b8c0010", 17968 => x"5b8d000c", 17969 => x"5b8e0008",
    17970 => x"5b9d0004", 17971 => x"780c0001", 17972 => x"780d0001",
    17973 => x"b8207000", 17974 => x"340b0000", 17975 => x"398c924c",
    17976 => x"39ad8ed8", 17977 => x"e000000a", 17978 => x"29a10000",
    17979 => x"942b0800", 17980 => x"20210001", 17981 => x"44200005",
    17982 => x"35620013", 17983 => x"3c420005", 17984 => x"b5c20800",
    17985 => x"fbffff46", 17986 => x"356b0001", 17987 => x"29810000",
    17988 => x"482bfff6", 17989 => x"2b9d0004", 17990 => x"2b8b0014",
    17991 => x"2b8c0010", 17992 => x"2b8d000c", 17993 => x"2b8e0008",
    17994 => x"379c0014", 17995 => x"c3a00000", 17996 => x"379cffbc",
    17997 => x"5b8b0044", 17998 => x"5b8c0040", 17999 => x"5b8d003c",
    18000 => x"5b8e0038", 18001 => x"5b8f0034", 18002 => x"5b900030",
    18003 => x"5b91002c", 18004 => x"5b920028", 18005 => x"5b930024",
    18006 => x"5b940020", 18007 => x"5b95001c", 18008 => x"5b960018",
    18009 => x"5b970014", 18010 => x"5b980010", 18011 => x"5b99000c",
    18012 => x"5b9b0008", 18013 => x"5b9d0004", 18014 => x"781b0001",
    18015 => x"780b0001", 18016 => x"78190001", 18017 => x"780d0001",
    18018 => x"78110001", 18019 => x"78100001", 18020 => x"780c0001",
    18021 => x"78170001", 18022 => x"780f0001", 18023 => x"3b7b8ee8",
    18024 => x"396b8f04", 18025 => x"34140009", 18026 => x"3b395dfc",
    18027 => x"34180001", 18028 => x"34130003", 18029 => x"39ad8f9c",
    18030 => x"34120008", 18031 => x"3a318fbc", 18032 => x"3a108f20",
    18033 => x"398c924c", 18034 => x"3af79164", 18035 => x"39ef9244",
    18036 => x"e0000079", 18037 => x"2875007c", 18038 => x"780100ff",
    18039 => x"3821ffff", 18040 => x"02ae0018", 18041 => x"a2a1a800",
    18042 => x"29610004", 18043 => x"21ce007f", 18044 => x"3421ffff",
    18045 => x"54340050", 18046 => x"3c210002", 18047 => x"b7210800",
    18048 => x"28210000", 18049 => x"c0200000", 18050 => x"2961004c",
    18051 => x"58610040", 18052 => x"296100d4", 18053 => x"296200d0",
    18054 => x"b4410800", 18055 => x"0022001f", 18056 => x"b4410800",
    18057 => x"14210001", 18058 => x"34020001", 18059 => x"58610044",
    18060 => x"29810000", 18061 => x"fbfffbe7", 18062 => x"fbfff0ea",
    18063 => x"34210032", 18064 => x"59610008", 18065 => x"3401000a",
    18066 => x"e0000011", 18067 => x"29760008", 18068 => x"fbfff0e4",
    18069 => x"cac10800", 18070 => x"4c200037", 18071 => x"29610000",
    18072 => x"5c380003", 18073 => x"59780004", 18074 => x"e0000033",
    18075 => x"59730004", 18076 => x"e0000031", 18077 => x"29810000",
    18078 => x"34020000", 18079 => x"fbfffbd5", 18080 => x"b9a00800",
    18081 => x"fbfffc4b", 18082 => x"34010002", 18083 => x"59610004",
    18084 => x"e0000029", 18085 => x"b9a00800", 18086 => x"fbfffc5c",
    18087 => x"e0000012", 18088 => x"ba000800", 18089 => x"fbfffdb4",
    18090 => x"34010004", 18091 => x"e3fffff8", 18092 => x"29610068",
    18093 => x"44200020", 18094 => x"2961006c", 18095 => x"4420001e",
    18096 => x"29610000", 18097 => x"5c330009", 18098 => x"34010005",
    18099 => x"e3fffff0", 18100 => x"ba200800", 18101 => x"fbfffdee",
    18102 => x"34010006", 18103 => x"e3ffffec", 18104 => x"296100f0",
    18105 => x"44200014", 18106 => x"b9600800", 18107 => x"fbffff72",
    18108 => x"59720004", 18109 => x"e0000010", 18110 => x"29610000",
    18111 => x"5c380004", 18112 => x"b9a00800", 18113 => x"fbfffc41",
    18114 => x"44200007", 18115 => x"29610068", 18116 => x"44200005",
    18117 => x"29610000", 18118 => x"5c330007", 18119 => x"296100f0",
    18120 => x"5c200005", 18121 => x"29610010", 18122 => x"34210001",
    18123 => x"59610010", 18124 => x"59740004", 18125 => x"ba000800",
    18126 => x"baa01000", 18127 => x"b9c01800", 18128 => x"fbfffd36",
    18129 => x"29610068", 18130 => x"4420001b", 18131 => x"ba200800",
    18132 => x"baa01000", 18133 => x"b9c01800", 18134 => x"fbfffdfe",
    18135 => x"29610004", 18136 => x"5c320015", 18137 => x"29610000",
    18138 => x"34160000", 18139 => x"5c33000c", 18140 => x"e0000008",
    18141 => x"0ac10090", 18142 => x"baa01000", 18143 => x"b9c01800",
    18144 => x"34210148", 18145 => x"b5610800", 18146 => x"fbfffdf2",
    18147 => x"36d60001", 18148 => x"29e10000", 18149 => x"3421ffff",
    18150 => x"4836fff7", 18151 => x"29810000", 18152 => x"49c10005",
    18153 => x"bae00800", 18154 => x"baa01000", 18155 => x"b9c01800",
    18156 => x"fbfffead", 18157 => x"2b630000", 18158 => x"78020002",
    18159 => x"28610080", 18160 => x"a0220800", 18161 => x"4420ff84",
    18162 => x"29610014", 18163 => x"34210001", 18164 => x"59610014",
    18165 => x"34010001", 18166 => x"d0410000", 18167 => x"2b9d0004",
    18168 => x"2b8b0044", 18169 => x"2b8c0040", 18170 => x"2b8d003c",
    18171 => x"2b8e0038", 18172 => x"2b8f0034", 18173 => x"2b900030",
    18174 => x"2b91002c", 18175 => x"2b920028", 18176 => x"2b930024",
    18177 => x"2b940020", 18178 => x"2b95001c", 18179 => x"2b960018",
    18180 => x"2b970014", 18181 => x"2b980010", 18182 => x"2b99000c",
    18183 => x"2b9b0008", 18184 => x"379c0044", 18185 => x"c3a00000",
    18186 => x"78010001", 18187 => x"38218f00", 18188 => x"28220000",
    18189 => x"78030001", 18190 => x"78010001", 18191 => x"38218efc",
    18192 => x"38635a00", 18193 => x"58220000", 18194 => x"28610000",
    18195 => x"58410000", 18196 => x"c3a00000", 18197 => x"379cffd4",
    18198 => x"5b8b0028", 18199 => x"5b8c0024", 18200 => x"5b8d0020",
    18201 => x"5b8e001c", 18202 => x"5b8f0018", 18203 => x"5b900014",
    18204 => x"5b910010", 18205 => x"5b92000c", 18206 => x"5b930008",
    18207 => x"5b9d0004", 18208 => x"b8205800", 18209 => x"b8408000",
    18210 => x"b8609000", 18211 => x"fbffb94f", 18212 => x"78010001",
    18213 => x"3821927c", 18214 => x"28240000", 18215 => x"78010001",
    18216 => x"38218ee8", 18217 => x"58240000", 18218 => x"78010001",
    18219 => x"28850000", 18220 => x"38218f00", 18221 => x"28210000",
    18222 => x"78020001", 18223 => x"38428efc", 18224 => x"00a60010",
    18225 => x"58410000", 18226 => x"78020001", 18227 => x"3842924c",
    18228 => x"20c6003f", 18229 => x"00a50018", 18230 => x"58460000",
    18231 => x"78020001", 18232 => x"38429244", 18233 => x"20a50007",
    18234 => x"58450000", 18235 => x"78050001", 18236 => x"38a58f04",
    18237 => x"58ab0000", 18238 => x"58a00010", 18239 => x"58800040",
    18240 => x"58800044", 18241 => x"58800000", 18242 => x"58800028",
    18243 => x"58800024", 18244 => x"58800004", 18245 => x"78030001",
    18246 => x"58800020", 18247 => x"340203e8", 18248 => x"386359cc",
    18249 => x"58820048", 18250 => x"28620000", 18251 => x"5820001c",
    18252 => x"58220000", 18253 => x"34010004", 18254 => x"5d610004",
    18255 => x"34010007", 18256 => x"58a10004", 18257 => x"e0000006",
    18258 => x"34010009", 18259 => x"58a10004", 18260 => x"34010003",
    18261 => x"5d610002", 18262 => x"ba003000", 18263 => x"78010001",
    18264 => x"b8c01000", 18265 => x"38218f20", 18266 => x"780d0001",
    18267 => x"fbfffc98", 18268 => x"39ad924c", 18269 => x"29a30000",
    18270 => x"78010001", 18271 => x"38218fbc", 18272 => x"ba001000",
    18273 => x"780f0001", 18274 => x"780e0001", 18275 => x"fbfffd19",
    18276 => x"340c0000", 18277 => x"39ef9244", 18278 => x"39ce8f04",
    18279 => x"34130001", 18280 => x"e000000c", 18281 => x"09910090",
    18282 => x"29a40000", 18283 => x"ba001000", 18284 => x"36210148",
    18285 => x"34840001", 18286 => x"b48c1800", 18287 => x"b5c10800",
    18288 => x"b5d18800", 18289 => x"fbfffd0b", 18290 => x"358c0001",
    18291 => x"5a330140", 18292 => x"29e10000", 18293 => x"3421ffff",
    18294 => x"482cfff3", 18295 => x"34010002", 18296 => x"5d610006",
    18297 => x"78010001", 18298 => x"38218efc", 18299 => x"28210000",
    18300 => x"34020006", 18301 => x"5822001c", 18302 => x"780e0001",
    18303 => x"780d0001", 18304 => x"340c0000", 18305 => x"39ce924c",
    18306 => x"39ad8f04", 18307 => x"e0000008", 18308 => x"35810013",
    18309 => x"3c210005", 18310 => x"b9801000", 18311 => x"b5a10800",
    18312 => x"34030200", 18313 => x"fbfffdf7", 18314 => x"358c0001",
    18315 => x"29c20000", 18316 => x"484cfff8", 18317 => x"34010001",
    18318 => x"5d610017", 18319 => x"78010001", 18320 => x"38218ee8",
    18321 => x"28210000", 18322 => x"28210004", 18323 => x"20210002",
    18324 => x"44200021", 18325 => x"78010001", 18326 => x"78040001",
    18327 => x"38218f04", 18328 => x"38848f20", 18329 => x"58240098",
    18330 => x"78040001", 18331 => x"38848fbc", 18332 => x"5824009c",
    18333 => x"78010001", 18334 => x"38219244", 18335 => x"28240000",
    18336 => x"78010001", 18337 => x"38218f9c", 18338 => x"b4441000",
    18339 => x"ba401800", 18340 => x"fbfffb2c", 18341 => x"78010001",
    18342 => x"38218ee8", 18343 => x"28210000", 18344 => x"78020002",
    18345 => x"e0000003", 18346 => x"2823007c", 18347 => x"5b83002c",
    18348 => x"28230080", 18349 => x"a0621800", 18350 => x"4460fffc",
    18351 => x"34020001", 18352 => x"58220064", 18353 => x"28220028",
    18354 => x"38420001", 18355 => x"58220028", 18356 => x"fbffb8c7",
    18357 => x"2b9d0004", 18358 => x"2b8b0028", 18359 => x"2b8c0024",
    18360 => x"2b8d0020", 18361 => x"2b8e001c", 18362 => x"2b8f0018",
    18363 => x"2b900014", 18364 => x"2b910010", 18365 => x"2b92000c",
    18366 => x"2b930008", 18367 => x"379c002c", 18368 => x"c3a00000",
    18369 => x"379cfffc", 18370 => x"5b9d0004", 18371 => x"78020001",
    18372 => x"38428f04", 18373 => x"28430004", 18374 => x"64240000",
    18375 => x"7c630008", 18376 => x"b8831800", 18377 => x"5c600006",
    18378 => x"3421ffff", 18379 => x"08210090", 18380 => x"34210148",
    18381 => x"b4410800", 18382 => x"fbfffcd5", 18383 => x"2b9d0004",
    18384 => x"379c0004", 18385 => x"c3a00000", 18386 => x"379cfffc",
    18387 => x"5b9d0004", 18388 => x"44200008", 18389 => x"3421ffff",
    18390 => x"08210090", 18391 => x"78020001", 18392 => x"38428f04",
    18393 => x"34210148", 18394 => x"b4220800", 18395 => x"fbfffced",
    18396 => x"2b9d0004", 18397 => x"379c0004", 18398 => x"c3a00000",
    18399 => x"78020001", 18400 => x"b8201800", 18401 => x"38428f04",
    18402 => x"5c200004", 18403 => x"28410004", 18404 => x"64210008",
    18405 => x"c3a00000", 18406 => x"28450004", 18407 => x"34040008",
    18408 => x"34010000", 18409 => x"5ca40006", 18410 => x"3463ffff",
    18411 => x"08630090", 18412 => x"b4431000", 18413 => x"28410180",
    18414 => x"7c210000", 18415 => x"c3a00000", 18416 => x"379cffe8",
    18417 => x"5b8b0018", 18418 => x"5b8c0014", 18419 => x"5b8d0010",
    18420 => x"5b8e000c", 18421 => x"5b8f0008", 18422 => x"5b9d0004",
    18423 => x"3403ffff", 18424 => x"b8407800", 18425 => x"5c230016",
    18426 => x"34010000", 18427 => x"780c0001", 18428 => x"780d0001",
    18429 => x"fbfffe19", 18430 => x"340b0000", 18431 => x"398c9244",
    18432 => x"39ad8f04", 18433 => x"340e0004", 18434 => x"e0000009",
    18435 => x"09610090", 18436 => x"b5a10800", 18437 => x"28210140",
    18438 => x"5c2e0004", 18439 => x"35610001", 18440 => x"b9e01000",
    18441 => x"fbfffe0d", 18442 => x"356b0001", 18443 => x"29810000",
    18444 => x"3421ffff", 18445 => x"482bfff6", 18446 => x"e0000002",
    18447 => x"fbfffe07", 18448 => x"2b9d0004", 18449 => x"2b8b0018",
    18450 => x"2b8c0014", 18451 => x"2b8d0010", 18452 => x"2b8e000c",
    18453 => x"2b8f0008", 18454 => x"379c0018", 18455 => x"c3a00000",
    18456 => x"379cfff0", 18457 => x"5b8b0010", 18458 => x"5b8c000c",
    18459 => x"5b8d0008", 18460 => x"5b9d0004", 18461 => x"780b0001",
    18462 => x"b8406800", 18463 => x"b8606000", 18464 => x"396b8fbc",
    18465 => x"44200007", 18466 => x"342bffff", 18467 => x"096b0090",
    18468 => x"78010001", 18469 => x"38218f04", 18470 => x"356b0148",
    18471 => x"b5615800", 18472 => x"45a0000b", 18473 => x"2962006c",
    18474 => x"34041f40", 18475 => x"34030000", 18476 => x"3c420001",
    18477 => x"1441001f", 18478 => x"f80002ae", 18479 => x"3c210012",
    18480 => x"0044000e", 18481 => x"b8242000", 18482 => x"59a40000",
    18483 => x"4580000b", 18484 => x"29620068", 18485 => x"34030000",
    18486 => x"34041f40", 18487 => x"3c420001", 18488 => x"1441001f",
    18489 => x"f80002a3", 18490 => x"3c210012", 18491 => x"0042000e",
    18492 => x"b8221000", 18493 => x"59820000", 18494 => x"2b9d0004",
    18495 => x"2b8b0010", 18496 => x"2b8c000c", 18497 => x"2b8d0008",
    18498 => x"379c0010", 18499 => x"c3a00000", 18500 => x"379cfff0",
    18501 => x"5b8b0010", 18502 => x"5b8c000c", 18503 => x"5b8d0008",
    18504 => x"5b9d0004", 18505 => x"b8205800", 18506 => x"b8406800",
    18507 => x"78010001", 18508 => x"3d620005", 18509 => x"38218f04",
    18510 => x"b4220800", 18511 => x"28240278", 18512 => x"b8606000",
    18513 => x"4c800003", 18514 => x"34844000", 18515 => x"e0000004",
    18516 => x"34013fff", 18517 => x"4c240002", 18518 => x"3484c000",
    18519 => x"3c840001", 18520 => x"34010000", 18521 => x"20823ffe",
    18522 => x"34030000", 18523 => x"34041f40", 18524 => x"f8000280",
    18525 => x"3c210012", 18526 => x"0044000e", 18527 => x"b8242000",
    18528 => x"59a40000", 18529 => x"4580000d", 18530 => x"78010001",
    18531 => x"38218ed8", 18532 => x"35630013", 18533 => x"28220000",
    18534 => x"3c630005", 18535 => x"78010001", 18536 => x"38218f04",
    18537 => x"b4230800", 18538 => x"28210004", 18539 => x"94410800",
    18540 => x"20210001", 18541 => x"59810000", 18542 => x"3d6b0005",
    18543 => x"78020001", 18544 => x"38428f04", 18545 => x"b44b1000",
    18546 => x"2841027c", 18547 => x"2b9d0004", 18548 => x"2b8b0010",
    18549 => x"2b8c000c", 18550 => x"2b8d0008", 18551 => x"379c0010",
    18552 => x"c3a00000", 18553 => x"379cffec", 18554 => x"5b8b0014",
    18555 => x"5b8c0010", 18556 => x"5b9d000c", 18557 => x"780b0001",
    18558 => x"396b8f04", 18559 => x"29610000", 18560 => x"4c010014",
    18561 => x"296c0014", 18562 => x"29620004", 18563 => x"78010001",
    18564 => x"38215e24", 18565 => x"fbfffa2c", 18566 => x"29640000",
    18567 => x"b8201800", 18568 => x"296500a4", 18569 => x"29660068",
    18570 => x"296700f0", 18571 => x"29680054", 18572 => x"296200dc",
    18573 => x"29610010", 18574 => x"5b820004", 18575 => x"5b810008",
    18576 => x"78010001", 18577 => x"3821587c", 18578 => x"b9801000",
    18579 => x"fbffe925", 18580 => x"2b9d000c", 18581 => x"2b8b0014",
    18582 => x"2b8c0010", 18583 => x"379c0014", 18584 => x"c3a00000",
    18585 => x"379cfffc", 18586 => x"5b9d0004", 18587 => x"5c200004",
    18588 => x"78010001", 18589 => x"38218fbc", 18590 => x"e0000007",
    18591 => x"3421ffff", 18592 => x"08210090", 18593 => x"78020001",
    18594 => x"38428f04", 18595 => x"34210148", 18596 => x"b4220800",
    18597 => x"fbfffcd7", 18598 => x"2b9d0004", 18599 => x"379c0004",
    18600 => x"c3a00000", 18601 => x"379cfff0", 18602 => x"5b8b0010",
    18603 => x"5b8c000c", 18604 => x"5b8d0008", 18605 => x"5b9d0004",
    18606 => x"780d0001", 18607 => x"780b0001", 18608 => x"b8206000",
    18609 => x"39ad8f04", 18610 => x"396b8ed8", 18611 => x"4440000d",
    18612 => x"34020001", 18613 => x"fbfff9bf", 18614 => x"35810013",
    18615 => x"3c210005", 18616 => x"b5a10800", 18617 => x"fbfffcce",
    18618 => x"29610000", 18619 => x"34020001", 18620 => x"bc4c6000",
    18621 => x"b9816000", 18622 => x"596c0000", 18623 => x"e000000a",
    18624 => x"34030001", 18625 => x"29640000", 18626 => x"bc611800",
    18627 => x"a4601800", 18628 => x"a0641800", 18629 => x"59630000",
    18630 => x"29a30128", 18631 => x"44230002", 18632 => x"fbfff9ac",
    18633 => x"2b9d0004", 18634 => x"2b8b0010", 18635 => x"2b8c000c",
    18636 => x"2b8d0008", 18637 => x"379c0010", 18638 => x"c3a00000",
    18639 => x"08210090", 18640 => x"78020001", 18641 => x"38428f04",
    18642 => x"b4411000", 18643 => x"28410140", 18644 => x"28430140",
    18645 => x"34020004", 18646 => x"7c210001", 18647 => x"5c620002",
    18648 => x"38210002", 18649 => x"c3a00000", 18650 => x"4c200005",
    18651 => x"78010001", 18652 => x"38218f04", 18653 => x"28210054",
    18654 => x"c3a00000", 18655 => x"78020001", 18656 => x"38428f04",
    18657 => x"5c200003", 18658 => x"284100dc", 18659 => x"c3a00000",
    18660 => x"3421ffff", 18661 => x"08210090", 18662 => x"b4411000",
    18663 => x"2841016c", 18664 => x"c3a00000", 18665 => x"78030001",
    18666 => x"38638ee8", 18667 => x"4c200007", 18668 => x"78010001",
    18669 => x"38218f04", 18670 => x"58220054", 18671 => x"28610000",
    18672 => x"58220040", 18673 => x"c3a00000", 18674 => x"2024000f",
    18675 => x"28630000", 18676 => x"3c840010", 18677 => x"2045ffff",
    18678 => x"b8a42000", 18679 => x"58640044", 18680 => x"78030001",
    18681 => x"38638f04", 18682 => x"5c200003", 18683 => x"586200dc",
    18684 => x"c3a00000", 18685 => x"3421ffff", 18686 => x"08210090",
    18687 => x"b4611800", 18688 => x"5862016c", 18689 => x"c3a00000",
    18690 => x"379cffcc", 18691 => x"5b8b0034", 18692 => x"5b8c0030",
    18693 => x"5b8d002c", 18694 => x"5b8e0028", 18695 => x"5b8f0024",
    18696 => x"5b900020", 18697 => x"5b91001c", 18698 => x"5b920018",
    18699 => x"5b930014", 18700 => x"5b940010", 18701 => x"5b95000c",
    18702 => x"5b960008", 18703 => x"5b9d0004", 18704 => x"78010001",
    18705 => x"38218f04", 18706 => x"28220000", 18707 => x"34010001",
    18708 => x"34140000", 18709 => x"5c410005", 18710 => x"78010001",
    18711 => x"38218f9c", 18712 => x"fbfffa05", 18713 => x"b820a000",
    18714 => x"78110001", 18715 => x"780b0001", 18716 => x"780e0001",
    18717 => x"340d0000", 18718 => x"340c0001", 18719 => x"3a319244",
    18720 => x"396b8f04", 18721 => x"340f0001", 18722 => x"39ce8ee8",
    18723 => x"34120002", 18724 => x"34160003", 18725 => x"34150004",
    18726 => x"e0000047", 18727 => x"3593ffff", 18728 => x"0a700090",
    18729 => x"b5708000", 18730 => x"2a010140", 18731 => x"442f000f",
    18732 => x"29c10000", 18733 => x"bdec1000", 18734 => x"28210020",
    18735 => x"00210008", 18736 => x"202100ff", 18737 => x"a0220800",
    18738 => x"5c200008", 18739 => x"b9800800", 18740 => x"fbfffe9e",
    18741 => x"b9800800", 18742 => x"34020000", 18743 => x"fbfffca7",
    18744 => x"35ad0001", 18745 => x"5a0f0140", 18746 => x"0a610090",
    18747 => x"b5618000", 18748 => x"2a020140", 18749 => x"44520014",
    18750 => x"48520003", 18751 => x"5c4f002d", 18752 => x"e0000004",
    18753 => x"44560017", 18754 => x"5c55002a", 18755 => x"e000001e",
    18756 => x"296100f0", 18757 => x"44200027", 18758 => x"29c10000",
    18759 => x"bdec1000", 18760 => x"28210020", 18761 => x"00210008",
    18762 => x"202100ff", 18763 => x"a0220800", 18764 => x"44200020",
    18765 => x"b9800800", 18766 => x"fbfffe73", 18767 => x"5a120140",
    18768 => x"e000001b", 18769 => x"2a010180", 18770 => x"4420001a",
    18771 => x"29620018", 18772 => x"b9800800", 18773 => x"fbfffcc1",
    18774 => x"5a160140", 18775 => x"e0000014", 18776 => x"34210148",
    18777 => x"b5610800", 18778 => x"fbfffc22", 18779 => x"5c200011",
    18780 => x"b9800800", 18781 => x"34020001", 18782 => x"fbfffc80",
    18783 => x"5a150140", 18784 => x"e000000b", 18785 => x"296100f0",
    18786 => x"44200003", 18787 => x"2a010180", 18788 => x"5c200008",
    18789 => x"0a730090", 18790 => x"b9800800", 18791 => x"34020000",
    18792 => x"b5739800", 18793 => x"fbfffc75", 18794 => x"5a6f0140",
    18795 => x"35ad0001", 18796 => x"358c0001", 18797 => x"2a210000",
    18798 => x"482cffb9", 18799 => x"29630000", 18800 => x"78020001",
    18801 => x"38427204", 18802 => x"5843000c", 18803 => x"29630014",
    18804 => x"28410008", 18805 => x"7dad0000", 18806 => x"58430010",
    18807 => x"29630004", 18808 => x"34210002", 18809 => x"b5b4a000",
    18810 => x"58430014", 18811 => x"296300a4", 18812 => x"58410008",
    18813 => x"7e810000", 18814 => x"58430018", 18815 => x"29630068",
    18816 => x"5843001c", 18817 => x"296300f0", 18818 => x"58430020",
    18819 => x"29630054", 18820 => x"58430024", 18821 => x"296300dc",
    18822 => x"58430028", 18823 => x"29630010", 18824 => x"5843002c",
    18825 => x"2b9d0004", 18826 => x"2b8b0034", 18827 => x"2b8c0030",
    18828 => x"2b8d002c", 18829 => x"2b8e0028", 18830 => x"2b8f0024",
    18831 => x"2b900020", 18832 => x"2b91001c", 18833 => x"2b920018",
    18834 => x"2b930014", 18835 => x"2b940010", 18836 => x"2b95000c",
    18837 => x"2b960008", 18838 => x"379c0034", 18839 => x"c3a00000",
    18840 => x"379cfff8", 18841 => x"5b8b0008", 18842 => x"5b9d0004",
    18843 => x"fbffb6d7", 18844 => x"34020000", 18845 => x"3401ffff",
    18846 => x"fbffff4b", 18847 => x"34010001", 18848 => x"fbfffc53",
    18849 => x"380bffff", 18850 => x"b9601000", 18851 => x"3401ffff",
    18852 => x"fbffff45", 18853 => x"34010001", 18854 => x"fbfffc4d",
    18855 => x"34020000", 18856 => x"34010000", 18857 => x"fbffff40",
    18858 => x"34010000", 18859 => x"fbfffc48", 18860 => x"b9601000",
    18861 => x"34010000", 18862 => x"fbffff3b", 18863 => x"34010000",
    18864 => x"fbfffc43", 18865 => x"34010002", 18866 => x"fbfffc41",
    18867 => x"2b9d0004", 18868 => x"2b8b0008", 18869 => x"379c0008",
    18870 => x"c3a00000", 18871 => x"379cfff0", 18872 => x"5b8b0010",
    18873 => x"5b8c000c", 18874 => x"5b8d0008", 18875 => x"5b9d0004",
    18876 => x"78010001", 18877 => x"780b0001", 18878 => x"38215954",
    18879 => x"780c0001", 18880 => x"396bf800", 18881 => x"282d0000",
    18882 => x"398c5940", 18883 => x"e0000005", 18884 => x"b9800800",
    18885 => x"fbffe7f3", 18886 => x"340103e8", 18887 => x"fbffedb6",
    18888 => x"29610000", 18889 => x"5c2dfffb", 18890 => x"2b9d0004",
    18891 => x"2b8b0010", 18892 => x"2b8c000c", 18893 => x"2b8d0008",
    18894 => x"379c0010", 18895 => x"c3a00000", 18896 => x"c3a00000",
    18897 => x"379cfff8", 18898 => x"5b8b0008", 18899 => x"5b9d0004",
    18900 => x"28240014", 18901 => x"b8201800", 18902 => x"b8403000",
    18903 => x"44800015", 18904 => x"28250010", 18905 => x"20a50002",
    18906 => x"5ca00007", 18907 => x"b4862000", 18908 => x"b8800800",
    18909 => x"2b9d0004", 18910 => x"2b8b0008", 18911 => x"379c0008",
    18912 => x"c3a00000", 18913 => x"346b0030", 18914 => x"b4861000",
    18915 => x"b9600800", 18916 => x"34030040", 18917 => x"f80001cc",
    18918 => x"b9602000", 18919 => x"b8800800", 18920 => x"2b9d0004",
    18921 => x"2b8b0008", 18922 => x"379c0008", 18923 => x"c3a00000",
    18924 => x"28250010", 18925 => x"20a70004", 18926 => x"5ce4ffeb",
    18927 => x"2825001c", 18928 => x"34040000", 18929 => x"44a7ffeb",
    18930 => x"342b0030", 18931 => x"34040040", 18932 => x"b9601800",
    18933 => x"d8a00000", 18934 => x"b9602000", 18935 => x"e3fffff0",
    18936 => x"379cfff4", 18937 => x"5b8b0008", 18938 => x"5b9d0004",
    18939 => x"28220014", 18940 => x"b8205800", 18941 => x"44400013",
    18942 => x"2961000c", 18943 => x"b4411000", 18944 => x"28430000",
    18945 => x"78040001", 18946 => x"38845a04", 18947 => x"28820000",
    18948 => x"3401ffec", 18949 => x"5c620007", 18950 => x"78020001",
    18951 => x"38428edc", 18952 => x"28430000", 18953 => x"34010000",
    18954 => x"584b0000", 18955 => x"5963007c", 18956 => x"2b9d0004",
    18957 => x"2b8b0008", 18958 => x"379c000c", 18959 => x"c3a00000",
    18960 => x"28230010", 18961 => x"20630004", 18962 => x"5c62ffec",
    18963 => x"2825001c", 18964 => x"2822000c", 18965 => x"3783000c",
    18966 => x"34040004", 18967 => x"d8a00000", 18968 => x"2b83000c",
    18969 => x"e3ffffe8", 18970 => x"379cfff0", 18971 => x"5b8b0010",
    18972 => x"5b8c000c", 18973 => x"5b8d0008", 18974 => x"5b9d0004",
    18975 => x"b8205800", 18976 => x"44400047", 18977 => x"2822000c",
    18978 => x"58200080", 18979 => x"582000b0", 18980 => x"58220090",
    18981 => x"340c0000", 18982 => x"b9600800", 18983 => x"fbffffaa",
    18984 => x"59610028", 18985 => x"4022003f", 18986 => x"5c400006",
    18987 => x"78040001", 18988 => x"38845a04", 18989 => x"28230000",
    18990 => x"28820000", 18991 => x"4462005d", 18992 => x"34010000",
    18993 => x"45800030", 18994 => x"3583ffff", 18995 => x"346c0028",
    18996 => x"b58c0800", 18997 => x"b4210800", 18998 => x"b5610800",
    18999 => x"28220000", 19000 => x"5c40000f", 19001 => x"34010000",
    19002 => x"44620027", 19003 => x"34620027", 19004 => x"b4421000",
    19005 => x"b4421000", 19006 => x"b5621000", 19007 => x"e0000002",
    19008 => x"44610044", 19009 => x"28410000", 19010 => x"3463ffff",
    19011 => x"3442fffc", 19012 => x"4420fffc", 19013 => x"596300b0",
    19014 => x"346c0028", 19015 => x"346d0024", 19016 => x"b5ad6800",
    19017 => x"b5ad6800", 19018 => x"b56d6800", 19019 => x"29a20000",
    19020 => x"b9600800", 19021 => x"b58c6000", 19022 => x"fbffff83",
    19023 => x"b58c6000", 19024 => x"b56c1000", 19025 => x"29a40000",
    19026 => x"28430000", 19027 => x"296c00b0", 19028 => x"34840040",
    19029 => x"3463ffff", 19030 => x"59610028", 19031 => x"59a40000",
    19032 => x"58430000", 19033 => x"35830020", 19034 => x"b4631800",
    19035 => x"b4631800", 19036 => x"b5631800", 19037 => x"2824000c",
    19038 => x"28620000", 19039 => x"b4441000", 19040 => x"59620074",
    19041 => x"2b9d0004", 19042 => x"2b8b0010", 19043 => x"2b8c000c",
    19044 => x"2b8d0008", 19045 => x"379c0010", 19046 => x"c3a00000",
    19047 => x"28210028", 19048 => x"296300b0", 19049 => x"34050002",
    19050 => x"4024003f", 19051 => x"eca32800", 19052 => x"64840002",
    19053 => x"a0852000", 19054 => x"4482ffc5", 19055 => x"34620020",
    19056 => x"b4421000", 19057 => x"b4421000", 19058 => x"b5621000",
    19059 => x"28450000", 19060 => x"34640025", 19061 => x"28220004",
    19062 => x"b4842000", 19063 => x"b4842000", 19064 => x"b4a21000",
    19065 => x"b5642000", 19066 => x"58820000", 19067 => x"2824000c",
    19068 => x"34610021", 19069 => x"b4210800", 19070 => x"b4210800",
    19071 => x"b5610800", 19072 => x"b4852800", 19073 => x"346c0001",
    19074 => x"58250000", 19075 => x"e3ffffa3", 19076 => x"34010000",
    19077 => x"596000b0", 19078 => x"2b9d0004", 19079 => x"2b8b0010",
    19080 => x"2b8c000c", 19081 => x"2b8d0008", 19082 => x"379c0010",
    19083 => x"c3a00000", 19084 => x"35820024", 19085 => x"b4421000",
    19086 => x"b4421000", 19087 => x"b5621800", 19088 => x"2c250004",
    19089 => x"28640000", 19090 => x"35820028", 19091 => x"b4421000",
    19092 => x"b4421000", 19093 => x"b5621000", 19094 => x"34a5ffff",
    19095 => x"34840040", 19096 => x"58450000", 19097 => x"58640000",
    19098 => x"596c00b0", 19099 => x"e3ffffbe", 19100 => x"379cffec",
    19101 => x"5b8b0014", 19102 => x"5b8c0010", 19103 => x"5b8d000c",
    19104 => x"5b8e0008", 19105 => x"5b9d0004", 19106 => x"b8406000",
    19107 => x"34020001", 19108 => x"b8205800", 19109 => x"b8607000",
    19110 => x"b8806800", 19111 => x"fbffff73", 19112 => x"b9600800",
    19113 => x"34020000", 19114 => x"fbffff70", 19115 => x"b8202800",
    19116 => x"4420001e", 19117 => x"28a10018", 19118 => x"5c2cfffa",
    19119 => x"28a1001c", 19120 => x"5c2efff8", 19121 => x"28a10020",
    19122 => x"5c2dfff6", 19123 => x"296100b0", 19124 => x"59650028",
    19125 => x"28a2000c", 19126 => x"34210020", 19127 => x"b4210800",
    19128 => x"b4210800", 19129 => x"b5610800", 19130 => x"28230000",
    19131 => x"34010000", 19132 => x"b4431800", 19133 => x"59630074",
    19134 => x"28a30014", 19135 => x"59600078", 19136 => x"34630001",
    19137 => x"c8621000", 19138 => x"59620070", 19139 => x"2b9d0004",
    19140 => x"2b8b0014", 19141 => x"2b8c0010", 19142 => x"2b8d000c",
    19143 => x"2b8e0008", 19144 => x"379c0014", 19145 => x"c3a00000",
    19146 => x"3401fffe", 19147 => x"e3fffff8", 19148 => x"379cfff8",
    19149 => x"5b8b0008", 19150 => x"5b9d0004", 19151 => x"b8205800",
    19152 => x"fbffffcc", 19153 => x"4c200005", 19154 => x"2b9d0004",
    19155 => x"2b8b0008", 19156 => x"379c0008", 19157 => x"c3a00000",
    19158 => x"29610074", 19159 => x"59600028", 19160 => x"2b9d0004",
    19161 => x"2b8b0008", 19162 => x"379c0008", 19163 => x"c3a00000",
    19164 => x"2045ffff", 19165 => x"00460010", 19166 => x"2088ffff",
    19167 => x"00890010", 19168 => x"89053800", 19169 => x"89064000",
    19170 => x"89252800", 19171 => x"00ea0010", 19172 => x"89263000",
    19173 => x"b5052800", 19174 => x"b4aa2800", 19175 => x"50a80003",
    19176 => x"78080001", 19177 => x"b4c83000", 19178 => x"88431000",
    19179 => x"88812000", 19180 => x"00a10010", 19181 => x"3ca50010",
    19182 => x"b4c13000", 19183 => x"20e7ffff", 19184 => x"b4440800",
    19185 => x"b4260800", 19186 => x"b4a71000", 19187 => x"c3a00000",
    19188 => x"44600008", 19189 => x"34040020", 19190 => x"c8832000",
    19191 => x"48800006", 19192 => x"c8041000", 19193 => x"34030000",
    19194 => x"80221000", 19195 => x"b8600800", 19196 => x"c3a00000",
    19197 => x"bc242000", 19198 => x"80431000", 19199 => x"80231800",
    19200 => x"b8821000", 19201 => x"b8600800", 19202 => x"e3fffffa",
    19203 => x"379cfff8", 19204 => x"5b8b0008", 19205 => x"5b9d0004",
    19206 => x"44400022", 19207 => x"b8412000", 19208 => x"3403000f",
    19209 => x"5483000b", 19210 => x"78030001", 19211 => x"38635e7c",
    19212 => x"3c210004", 19213 => x"b4621000", 19214 => x"b4410800",
    19215 => x"40210000", 19216 => x"2b9d0004", 19217 => x"2b8b0008",
    19218 => x"379c0008", 19219 => x"c3a00000", 19220 => x"340b0000",
    19221 => x"4c200003", 19222 => x"c8010800", 19223 => x"340b0001",
    19224 => x"4c400003", 19225 => x"c8021000", 19226 => x"196b0001",
    19227 => x"90c01800", 19228 => x"20630002", 19229 => x"44600008",
    19230 => x"8c220800", 19231 => x"45600002", 19232 => x"c8010800",
    19233 => x"2b9d0004", 19234 => x"2b8b0008", 19235 => x"379c0008",
    19236 => x"c3a00000", 19237 => x"34030000", 19238 => x"f800004a",
    19239 => x"e3fffff8", 19240 => x"90000800", 19241 => x"20210001",
    19242 => x"3c210001", 19243 => x"d0010000", 19244 => x"90e00800",
    19245 => x"bba0f000", 19246 => x"342100a0", 19247 => x"c0200000",
    19248 => x"379cfff8", 19249 => x"5b8b0008", 19250 => x"5b9d0004",
    19251 => x"44400015", 19252 => x"340b0000", 19253 => x"4c200003",
    19254 => x"c8010800", 19255 => x"340b0001", 19256 => x"1443001f",
    19257 => x"90c02000", 19258 => x"98621000", 19259 => x"20840002",
    19260 => x"c8431000", 19261 => x"44800008", 19262 => x"c4220800",
    19263 => x"45600002", 19264 => x"c8010800", 19265 => x"2b9d0004",
    19266 => x"2b8b0008", 19267 => x"379c0008", 19268 => x"c3a00000",
    19269 => x"34030001", 19270 => x"f800002a", 19271 => x"e3fffff8",
    19272 => x"90000800", 19273 => x"20210001", 19274 => x"3c210001",
    19275 => x"d0010000", 19276 => x"90e00800", 19277 => x"bba0f000",
    19278 => x"342100a0", 19279 => x"c0200000", 19280 => x"379cfffc",
    19281 => x"5b9d0004", 19282 => x"44400006", 19283 => x"34030000",
    19284 => x"f800001c", 19285 => x"2b9d0004", 19286 => x"379c0004",
    19287 => x"c3a00000", 19288 => x"90000800", 19289 => x"20210001",
    19290 => x"3c210001", 19291 => x"d0010000", 19292 => x"90e00800",
    19293 => x"bba0f000", 19294 => x"342100a0", 19295 => x"c0200000",
    19296 => x"379cfffc", 19297 => x"5b9d0004", 19298 => x"44400006",
    19299 => x"34030001", 19300 => x"f800000c", 19301 => x"2b9d0004",
    19302 => x"379c0004", 19303 => x"c3a00000", 19304 => x"90000800",
    19305 => x"20210001", 19306 => x"3c210001", 19307 => x"d0010000",
    19308 => x"90e00800", 19309 => x"bba0f000", 19310 => x"342100a0",
    19311 => x"c0200000", 19312 => x"f4222000", 19313 => x"44800018",
    19314 => x"34040001", 19315 => x"4c40000b", 19316 => x"34050000",
    19317 => x"54410003", 19318 => x"c8220800", 19319 => x"b8a42800",
    19320 => x"00840001", 19321 => x"00420001", 19322 => x"5c80fffb",
    19323 => x"5c600002", 19324 => x"b8a00800", 19325 => x"c3a00000",
    19326 => x"3c420001", 19327 => x"3c840001", 19328 => x"f4222800",
    19329 => x"7c860000", 19330 => x"a0c52800", 19331 => x"44a00002",
    19332 => x"4c40fffa", 19333 => x"34050000", 19334 => x"4480fff5",
    19335 => x"34050000", 19336 => x"e3ffffed", 19337 => x"34040001",
    19338 => x"34050000", 19339 => x"e3ffffea", 19340 => x"1422001f",
    19341 => x"98410800", 19342 => x"c8220800", 19343 => x"c3a00000",
    19344 => x"34060003", 19345 => x"b8202000", 19346 => x"b8402800",
    19347 => x"50c3000c", 19348 => x"b8413000", 19349 => x"20c60003",
    19350 => x"5cc0000b", 19351 => x"34010003", 19352 => x"28860000",
    19353 => x"28a20000", 19354 => x"5cc20005", 19355 => x"3463fffc",
    19356 => x"34840004", 19357 => x"34a50004", 19358 => x"5461fffa",
    19359 => x"34010000", 19360 => x"4460000e", 19361 => x"40860000",
    19362 => x"40a10000", 19363 => x"3462ffff", 19364 => x"44c10006",
    19365 => x"e000000a", 19366 => x"40860000", 19367 => x"40a10000",
    19368 => x"3442ffff", 19369 => x"5cc10006", 19370 => x"34840001",
    19371 => x"34a50001", 19372 => x"5c40fffa", 19373 => x"34010000",
    19374 => x"c3a00000", 19375 => x"c8c10800", 19376 => x"c3a00000",
    19377 => x"3404000f", 19378 => x"b8203800", 19379 => x"b8403000",
    19380 => x"5083002d", 19381 => x"b8412000", 19382 => x"20840003",
    19383 => x"5c80002b", 19384 => x"b8402000", 19385 => x"b8202800",
    19386 => x"b8603000", 19387 => x"3407000f", 19388 => x"28880000",
    19389 => x"34c6fff0", 19390 => x"58a80000", 19391 => x"28880004",
    19392 => x"58a80004", 19393 => x"28880008", 19394 => x"58a80008",
    19395 => x"2888000c", 19396 => x"34840010", 19397 => x"58a8000c",
    19398 => x"34a50010", 19399 => x"54c7fff5", 19400 => x"3463fff0",
    19401 => x"00660004", 19402 => x"2063000f", 19403 => x"34c60001",
    19404 => x"3cc60004", 19405 => x"b4263800", 19406 => x"b4463000",
    19407 => x"34020003", 19408 => x"50430011", 19409 => x"34020000",
    19410 => x"34080003", 19411 => x"b4c22000", 19412 => x"28850000",
    19413 => x"b4e22000", 19414 => x"34420004", 19415 => x"58850000",
    19416 => x"c8622000", 19417 => x"5488fffa", 19418 => x"3463fffc",
    19419 => x"00620002", 19420 => x"20630003", 19421 => x"34420001",
    19422 => x"3c420002", 19423 => x"b4e23800", 19424 => x"b4c23000",
    19425 => x"44600008", 19426 => x"34020000", 19427 => x"b4c22000",
    19428 => x"40850000", 19429 => x"b4e22000", 19430 => x"34420001",
    19431 => x"30850000", 19432 => x"5c43fffb", 19433 => x"c3a00000",
    19434 => x"b8203800", 19435 => x"b8403000", 19436 => x"5041000c",
    19437 => x"b4432000", 19438 => x"5024000a", 19439 => x"4460003f",
    19440 => x"b4231000", 19441 => x"3484ffff", 19442 => x"40850000",
    19443 => x"3442ffff", 19444 => x"3463ffff", 19445 => x"30450000",
    19446 => x"5c60fffb", 19447 => x"c3a00000", 19448 => x"3404000f",
    19449 => x"5083002d", 19450 => x"b8412000", 19451 => x"20840003",
    19452 => x"5c80002b", 19453 => x"b8402000", 19454 => x"b8202800",
    19455 => x"b8603000", 19456 => x"3407000f", 19457 => x"28880000",
    19458 => x"34c6fff0", 19459 => x"58a80000", 19460 => x"28880004",
    19461 => x"58a80004", 19462 => x"28880008", 19463 => x"58a80008",
    19464 => x"2888000c", 19465 => x"34840010", 19466 => x"58a8000c",
    19467 => x"34a50010", 19468 => x"54c7fff5", 19469 => x"3463fff0",
    19470 => x"00660004", 19471 => x"2063000f", 19472 => x"34c60001",
    19473 => x"3cc60004", 19474 => x"b4263800", 19475 => x"b4463000",
    19476 => x"34020003", 19477 => x"50430011", 19478 => x"34020000",
    19479 => x"34080003", 19480 => x"b4c22000", 19481 => x"28850000",
    19482 => x"b4e22000", 19483 => x"34420004", 19484 => x"58850000",
    19485 => x"c8622000", 19486 => x"5488fffa", 19487 => x"3463fffc",
    19488 => x"00620002", 19489 => x"20630003", 19490 => x"34420001",
    19491 => x"3c420002", 19492 => x"b4e23800", 19493 => x"b4c23000",
    19494 => x"44600008", 19495 => x"34020000", 19496 => x"b4c22000",
    19497 => x"40850000", 19498 => x"b4e22000", 19499 => x"34420001",
    19500 => x"30850000", 19501 => x"5c43fffb", 19502 => x"c3a00000",
    19503 => x"20250003", 19504 => x"b8202000", 19505 => x"44a0000b",
    19506 => x"4460002c", 19507 => x"3463ffff", 19508 => x"204600ff",
    19509 => x"e0000003", 19510 => x"44600028", 19511 => x"3463ffff",
    19512 => x"30860000", 19513 => x"34840001", 19514 => x"20850003",
    19515 => x"5ca0fffb", 19516 => x"34050003", 19517 => x"50a3001a",
    19518 => x"204500ff", 19519 => x"3ca60008", 19520 => x"340a000f",
    19521 => x"b8c52800", 19522 => x"3ca60010", 19523 => x"b8804000",
    19524 => x"b8c53000", 19525 => x"b8603800", 19526 => x"b8802800",
    19527 => x"3409000f", 19528 => x"546a0017", 19529 => x"34040000",
    19530 => x"34070003", 19531 => x"b5042800", 19532 => x"34840004",
    19533 => x"58a60000", 19534 => x"c8642800", 19535 => x"54a7fffc",
    19536 => x"3463fffc", 19537 => x"00640002", 19538 => x"20630003",
    19539 => x"34840001", 19540 => x"3c840002", 19541 => x"b5044000",
    19542 => x"b9002000", 19543 => x"44600007", 19544 => x"204200ff",
    19545 => x"34050000", 19546 => x"b4853000", 19547 => x"30c20000",
    19548 => x"34a50001", 19549 => x"5c65fffd", 19550 => x"c3a00000",
    19551 => x"58a60000", 19552 => x"58a60004", 19553 => x"58a60008",
    19554 => x"58a6000c", 19555 => x"34e7fff0", 19556 => x"34a50010",
    19557 => x"54e9fffa", 19558 => x"3463fff0", 19559 => x"00680004",
    19560 => x"2063000f", 19561 => x"35080001", 19562 => x"3d080004",
    19563 => x"b4884000", 19564 => x"34040003", 19565 => x"5464ffdc",
    19566 => x"b9002000", 19567 => x"e3ffffe8", 19568 => x"78030001",
    19569 => x"38637200", 19570 => x"28670000", 19571 => x"b8204800",
    19572 => x"34030000", 19573 => x"34060001", 19574 => x"e0000009",
    19575 => x"40840000", 19576 => x"b4e44000", 19577 => x"41080001",
    19578 => x"21080003", 19579 => x"45060012", 19580 => x"c8a40800",
    19581 => x"5c200013", 19582 => x"44810012", 19583 => x"b5232800",
    19584 => x"40a50000", 19585 => x"b4432000", 19586 => x"34630001",
    19587 => x"b4e54000", 19588 => x"41080001", 19589 => x"21080003",
    19590 => x"5d06fff1", 19591 => x"40840000", 19592 => x"34a50020",
    19593 => x"b4e44000", 19594 => x"41080001", 19595 => x"21080003",
    19596 => x"5d06fff0", 19597 => x"34840020", 19598 => x"c8a40800",
    19599 => x"4420ffef", 19600 => x"c3a00000", 19601 => x"b8411800",
    19602 => x"20630003", 19603 => x"5c60001d", 19604 => x"b8202000",
    19605 => x"28430000", 19606 => x"28210000", 19607 => x"5c230018",
    19608 => x"78030001", 19609 => x"38635f7c", 19610 => x"28670000",
    19611 => x"78030001", 19612 => x"38635f80", 19613 => x"28660000",
    19614 => x"a4201800", 19615 => x"b4270800", 19616 => x"a0231800",
    19617 => x"a0661800", 19618 => x"34010000", 19619 => x"44600003",
    19620 => x"e000001c", 19621 => x"5c600019", 19622 => x"34840004",
    19623 => x"28810000", 19624 => x"34420004", 19625 => x"28480000",
    19626 => x"b4272800", 19627 => x"a4201800", 19628 => x"a0a31800",
    19629 => x"a0661800", 19630 => x"4428fff7", 19631 => x"b8800800",
    19632 => x"40230000", 19633 => x"5c600006", 19634 => x"e0000009",
    19635 => x"34210001", 19636 => x"40230000", 19637 => x"34420001",
    19638 => x"44600005", 19639 => x"40440000", 19640 => x"4464fffb",
    19641 => x"c8640800", 19642 => x"c3a00000", 19643 => x"40440000",
    19644 => x"c8640800", 19645 => x"c3a00000", 19646 => x"34010000",
    19647 => x"c3a00000", 19648 => x"c3a00000", 19649 => x"b8412800",
    19650 => x"20a50003", 19651 => x"b8403800", 19652 => x"b8202000",
    19653 => x"5ca00018", 19654 => x"78040001", 19655 => x"38845f7c",
    19656 => x"28430000", 19657 => x"28880000", 19658 => x"78040001",
    19659 => x"38845f80", 19660 => x"28870000", 19661 => x"a4603000",
    19662 => x"b4682000", 19663 => x"a0c43000", 19664 => x"a0c73000",
    19665 => x"b8202000", 19666 => x"5cc5000a", 19667 => x"58830000",
    19668 => x"34420004", 19669 => x"28430000", 19670 => x"34840004",
    19671 => x"a4603000", 19672 => x"b4682800", 19673 => x"a0c52800",
    19674 => x"a0a72800", 19675 => x"44a0fff8", 19676 => x"b8403800",
    19677 => x"34030000", 19678 => x"b4e32800", 19679 => x"40a50000",
    19680 => x"b4833000", 19681 => x"34630001", 19682 => x"30c50000",
    19683 => x"5ca0fffb", 19684 => x"c3a00000", 19685 => x"20220003",
    19686 => x"4440002c", 19687 => x"40230000", 19688 => x"34020000",
    19689 => x"44600027", 19690 => x"b8201000", 19691 => x"e0000003",
    19692 => x"40430000", 19693 => x"44600022", 19694 => x"34420001",
    19695 => x"20430003", 19696 => x"5c60fffc", 19697 => x"78040001",
    19698 => x"38845f7c", 19699 => x"28430000", 19700 => x"28860000",
    19701 => x"78040001", 19702 => x"38845f80", 19703 => x"28850000",
    19704 => x"a4602000", 19705 => x"b4661800", 19706 => x"a0641800",
    19707 => x"a0651800", 19708 => x"5c600011", 19709 => x"34420004",
    19710 => x"28430000", 19711 => x"b4662000", 19712 => x"a4601800",
    19713 => x"a0831800", 19714 => x"a0651800", 19715 => x"5c60000a",
    19716 => x"34420004", 19717 => x"28430000", 19718 => x"b4662000",
    19719 => x"a4601800", 19720 => x"a0831800", 19721 => x"a0651800",
    19722 => x"4460fff3", 19723 => x"e0000002", 19724 => x"34420001",
    19725 => x"40430000", 19726 => x"5c60fffe", 19727 => x"c8411000",
    19728 => x"b8400800", 19729 => x"c3a00000", 19730 => x"b8201000",
    19731 => x"e3ffffde", 19732 => x"34060000", 19733 => x"44600017",
    19734 => x"b8413800", 19735 => x"20e70003", 19736 => x"3464ffff",
    19737 => x"44e00015", 19738 => x"40230000", 19739 => x"40450000",
    19740 => x"5c65000f", 19741 => x"34060000", 19742 => x"4480000e",
    19743 => x"34210001", 19744 => x"34420001", 19745 => x"5c600004",
    19746 => x"e000000a", 19747 => x"44800033", 19748 => x"44600032",
    19749 => x"40230000", 19750 => x"40450000", 19751 => x"3484ffff",
    19752 => x"34210001", 19753 => x"34420001", 19754 => x"4465fff9",
    19755 => x"c8653000", 19756 => x"b8c00800", 19757 => x"c3a00000",
    19758 => x"b8202800", 19759 => x"34010003", 19760 => x"b8402000",
    19761 => x"50230028", 19762 => x"28a10000", 19763 => x"28420000",
    19764 => x"5c220025", 19765 => x"3463fffc", 19766 => x"b8e03000",
    19767 => x"4460fff5", 19768 => x"78020001", 19769 => x"38425f7c",
    19770 => x"28490000", 19771 => x"78020001", 19772 => x"38425f80",
    19773 => x"28480000", 19774 => x"a4201000", 19775 => x"b4290800",
    19776 => x"a0220800", 19777 => x"a0280800", 19778 => x"34070003",
    19779 => x"5c20ffe9", 19780 => x"34a50004", 19781 => x"34840004",
    19782 => x"54670006", 19783 => x"b8a00800", 19784 => x"b8801000",
    19785 => x"44600014", 19786 => x"3464ffff", 19787 => x"e3ffffcf",
    19788 => x"28a10000", 19789 => x"288a0000", 19790 => x"b4293000",
    19791 => x"a4201000", 19792 => x"a0c21000", 19793 => x"a0481000",
    19794 => x"5c2a0007", 19795 => x"3463fffc", 19796 => x"44600002",
    19797 => x"4440ffef", 19798 => x"34060000", 19799 => x"b8c00800",
    19800 => x"c3a00000", 19801 => x"b8801000", 19802 => x"b8a00800",
    19803 => x"3464ffff", 19804 => x"e3ffffbe", 19805 => x"40a30000",
    19806 => x"40850000", 19807 => x"c8653000", 19808 => x"e3ffffcc",
    19809 => x"b8412000", 19810 => x"20840003", 19811 => x"74650003",
    19812 => x"64840000", 19813 => x"b8403000", 19814 => x"a0852000",
    19815 => x"b8202800", 19816 => x"44800015", 19817 => x"78040001",
    19818 => x"38845f7c", 19819 => x"28890000", 19820 => x"78040001",
    19821 => x"38845f80", 19822 => x"28880000", 19823 => x"340a0003",
    19824 => x"e0000006", 19825 => x"58a40000", 19826 => x"3463fffc",
    19827 => x"34a50004", 19828 => x"34420004", 19829 => x"51430007",
    19830 => x"28440000", 19831 => x"a4803800", 19832 => x"b4893000",
    19833 => x"a0e63000", 19834 => x"a0c83000", 19835 => x"44c0fff6",
    19836 => x"b8403000", 19837 => x"44600014", 19838 => x"40c20000",
    19839 => x"3463ffff", 19840 => x"34a40001", 19841 => x"30a20000",
    19842 => x"44400009", 19843 => x"34c20001", 19844 => x"4460000e",
    19845 => x"40450000", 19846 => x"3463ffff", 19847 => x"34420001",
    19848 => x"30850000", 19849 => x"34840001", 19850 => x"5ca0fffa",
    19851 => x"34020000", 19852 => x"44600007", 19853 => x"b4822800",
    19854 => x"30a00000", 19855 => x"34420001", 19856 => x"5c62fffd",
    19857 => x"c3a00000", 19858 => x"c3a00000", 19859 => x"c3a00000",
    19860 => x"34030000", 19861 => x"4440000c", 19862 => x"40240000",
    19863 => x"4480000a", 19864 => x"3442ffff", 19865 => x"b8201800",
    19866 => x"e0000004", 19867 => x"40640000", 19868 => x"3442ffff",
    19869 => x"44800003", 19870 => x"34630001", 19871 => x"5c40fffc",
    19872 => x"c8611800", 19873 => x"b8600800", 19874 => x"c3a00000",
    19875 => x"57522043", 19876 => x"6f72653a", 19877 => x"20737461",
    19878 => x"7274696e", 19879 => x"67207570", 19880 => x"2e2e2e0a",
    19881 => x"00000000", 19882 => x"556e6162", 19883 => x"6c652074",
    19884 => x"6f206465", 19885 => x"7465726d", 19886 => x"696e6520",
    19887 => x"4d414320", 19888 => x"61646472", 19889 => x"6573730a",
    19890 => x"00000000", 19891 => x"4c6f6361", 19892 => x"6c204d41",
    19893 => x"43206164", 19894 => x"64726573", 19895 => x"733a2025",
    19896 => x"3032783a", 19897 => x"25303278", 19898 => x"3a253032",
    19899 => x"783a2530", 19900 => x"32783a25", 19901 => x"3032783a",
    19902 => x"25303278", 19903 => x"0a000000", 19904 => x"73706c6c",
    19905 => x"2d626800", 19906 => x"7368656c", 19907 => x"6c2b6775",
    19908 => x"69000000", 19909 => x"70747000", 19910 => x"75707469",
    19911 => x"6d650000", 19912 => x"63686563", 19913 => x"6b2d6c69",
    19914 => x"6e6b0000", 19915 => x"69646c65", 19916 => x"00000000",
    19917 => x"64696167", 19918 => x"2d66736d", 19919 => x"2d312d25",
    19920 => x"733a2025", 19921 => x"3039642e", 19922 => x"25303364",
    19923 => x"3a200000", 19924 => x"454e5445", 19925 => x"52202573",
    19926 => x"2c207061", 19927 => x"636b6574", 19928 => x"206c656e",
    19929 => x"2025690a", 19930 => x"00000000", 19931 => x"25733a20",
    19932 => x"7265656e", 19933 => x"74657220", 19934 => x"696e2025",
    19935 => x"69206d73", 19936 => x"0a000000", 19937 => x"4c454156",
    19938 => x"45202573", 19939 => x"20286e65", 19940 => x"78743a20",
    19941 => x"25336929", 19942 => x"0a0a0000", 19943 => x"52454356",
    19944 => x"20253032", 19945 => x"64206279", 19946 => x"74657320",
    19947 => x"61742025", 19948 => x"642e2530", 19949 => x"39642028",
    19950 => x"74797065", 19951 => x"2025782c", 19952 => x"20257329",
    19953 => x"0a000000", 19954 => x"66736d20", 19955 => x"666f7220",
    19956 => x"25733a20", 19957 => x"4572726f", 19958 => x"72202569",
    19959 => x"20696e20", 19960 => x"25730a00", 19961 => x"66736d3a",
    19962 => x"20556e6b", 19963 => x"6e6f776e", 19964 => x"20737461",
    19965 => x"74652066", 19966 => x"6f722070", 19967 => x"6f727420",
    19968 => x"25730a00", 19969 => x"70707369", 19970 => x"00000000",
    19971 => x"25732d25", 19972 => x"692d2573", 19973 => x"3a200000",
    19974 => x"25733a20", 19975 => x"6572726f", 19976 => x"72207061",
    19977 => x"7273696e", 19978 => x"67202225", 19979 => x"73220a00",
    19980 => x"64696167", 19981 => x"2d636f6e", 19982 => x"66696700",
    19983 => x"64696167", 19984 => x"2d657874", 19985 => x"656e7369",
    19986 => x"6f6e0000", 19987 => x"64696167", 19988 => x"2d626d63",
    19989 => x"00000000", 19990 => x"64696167", 19991 => x"2d736572",
    19992 => x"766f0000", 19993 => x"64696167", 19994 => x"2d667261",
    19995 => x"6d657300", 19996 => x"64696167", 19997 => x"2d74696d",
    19998 => x"65000000", 19999 => x"64696167", 20000 => x"2d66736d",
    20001 => x"00000000", 20002 => x"50505369", 20003 => x"20666f72",
    20004 => x"20575250", 20005 => x"432e2043", 20006 => x"6f6d6d69",
    20007 => x"74202573", 20008 => x"2c206275", 20009 => x"696c7420",
    20010 => x"6f6e2053", 20011 => x"65702032", 20012 => x"30203230",
    20013 => x"31360a00", 20014 => x"70707369", 20015 => x"2d763230",
    20016 => x"31342e30", 20017 => x"372d3139", 20018 => x"362d6763",
    20019 => x"39336437", 20020 => x"31300000", 20021 => x"50545020",
    20022 => x"73746172", 20023 => x"740a0000", 20024 => x"50545020",
    20025 => x"73746f70", 20026 => x"0a000000", 20027 => x"4c6f636b",
    20028 => x"696e6720", 20029 => x"504c4c00", 20030 => x"0a4c6f63",
    20031 => x"6b207469", 20032 => x"6d656f75", 20033 => x"742e0000",
    20034 => x"2e000000", 20035 => x"77723100", 20036 => x"25732573",
    20037 => x"25303278", 20038 => x"2d253032", 20039 => x"782d2530",
    20040 => x"32782d25", 20041 => x"3032782d", 20042 => x"25303278",
    20043 => x"2d253032", 20044 => x"782d2530", 20045 => x"32782d25",
    20046 => x"3032782d", 20047 => x"25303278", 20048 => x"2d253032",
    20049 => x"780a0000", 20050 => x"25732573", 20051 => x"25732028",
    20052 => x"73697a65", 20053 => x"20256929", 20054 => x"0a000000",
    20055 => x"25732573", 20056 => x"00000000", 20057 => x"25303278",
    20058 => x"00000000", 20059 => x"25735645", 20060 => x"5253494f",
    20061 => x"4e3a2075", 20062 => x"6e737570", 20063 => x"706f7274",
    20064 => x"65642028", 20065 => x"2569290a", 20066 => x"00000000",
    20067 => x"25735645", 20068 => x"5253494f", 20069 => x"4e3a2025",
    20070 => x"69202874", 20071 => x"79706520", 20072 => x"25692c20",
    20073 => x"6c656e20", 20074 => x"25692c20", 20075 => x"646f6d61",
    20076 => x"696e2025", 20077 => x"69290a00", 20078 => x"2573464c",
    20079 => x"4147533a", 20080 => x"20307825", 20081 => x"30347820",
    20082 => x"28636f72", 20083 => x"72656374", 20084 => x"696f6e20",
    20085 => x"2530386c", 20086 => x"75290a00", 20087 => x"504f5254",
    20088 => x"3a200000", 20089 => x"25735245", 20090 => x"53543a20",
    20091 => x"73657120", 20092 => x"25692c20", 20093 => x"6374726c",
    20094 => x"2025692c", 20095 => x"206c6f67", 20096 => x"2d696e74",
    20097 => x"65727661", 20098 => x"6c202569", 20099 => x"0a000000",
    20100 => x"25734d45", 20101 => x"53534147", 20102 => x"453a2028",
    20103 => x"45292053", 20104 => x"594e430a", 20105 => x"00000000",
    20106 => x"25732573", 20107 => x"256c752e", 20108 => x"25303969",
    20109 => x"0a000000", 20110 => x"4d53472d", 20111 => x"53594e43",
    20112 => x"3a200000", 20113 => x"25734d45", 20114 => x"53534147",
    20115 => x"453a2028", 20116 => x"45292044", 20117 => x"454c4159",
    20118 => x"5f524551", 20119 => x"0a000000", 20120 => x"4d53472d",
    20121 => x"44454c41", 20122 => x"595f5245", 20123 => x"513a2000",
    20124 => x"25734d45", 20125 => x"53534147", 20126 => x"453a2028",
    20127 => x"47292046", 20128 => x"4f4c4c4f", 20129 => x"575f5550",
    20130 => x"0a000000", 20131 => x"4d53472d", 20132 => x"464f4c4c",
    20133 => x"4f575f55", 20134 => x"503a2000", 20135 => x"25734d45",
    20136 => x"53534147", 20137 => x"453a2028", 20138 => x"47292044",
    20139 => x"454c4159", 20140 => x"5f524553", 20141 => x"500a0000",
    20142 => x"4d53472d", 20143 => x"44454c41", 20144 => x"595f5245",
    20145 => x"53503a20", 20146 => x"00000000", 20147 => x"25734d45",
    20148 => x"53534147", 20149 => x"453a2028", 20150 => x"47292041",
    20151 => x"4e4e4f55", 20152 => x"4e43450a", 20153 => x"00000000",
    20154 => x"4d53472d", 20155 => x"414e4e4f", 20156 => x"554e4345",
    20157 => x"3a207374", 20158 => x"616d7020", 20159 => x"00000000",
    20160 => x"25732573", 20161 => x"25303278", 20162 => x"2d253032",
    20163 => x"782d2530", 20164 => x"34780a00", 20165 => x"4d53472d",
    20166 => x"414e4e4f", 20167 => x"554e4345", 20168 => x"3a206772",
    20169 => x"616e646d", 20170 => x"61737465", 20171 => x"722d7175",
    20172 => x"616c6974", 20173 => x"79200000", 20174 => x"25734d53",
    20175 => x"472d414e", 20176 => x"4e4f554e", 20177 => x"43453a20",
    20178 => x"6772616e", 20179 => x"646d6173", 20180 => x"7465722d",
    20181 => x"7072696f", 20182 => x"20256920", 20183 => x"25690a00",
    20184 => x"25732573", 20185 => x"25303278", 20186 => x"2d253032",
    20187 => x"782d2530", 20188 => x"32782d25", 20189 => x"3032782d",
    20190 => x"25303278", 20191 => x"2d253032", 20192 => x"782d2530",
    20193 => x"32782d25", 20194 => x"3032780a", 20195 => x"00000000",
    20196 => x"4d53472d", 20197 => x"414e4e4f", 20198 => x"554e4345",
    20199 => x"3a206772", 20200 => x"616e646d", 20201 => x"61737465",
    20202 => x"722d6964", 20203 => x"20000000", 20204 => x"25734d45",
    20205 => x"53534147", 20206 => x"453a2028", 20207 => x"47292053",
    20208 => x"49474e41", 20209 => x"4c494e47", 20210 => x"0a000000",
    20211 => x"4d53472d", 20212 => x"5349474e", 20213 => x"414c494e",
    20214 => x"473a2074", 20215 => x"61726765", 20216 => x"742d706f",
    20217 => x"72742000", 20218 => x"2573544c", 20219 => x"563a2074",
    20220 => x"6f6f2073", 20221 => x"686f7274", 20222 => x"20282569",
    20223 => x"202d2025", 20224 => x"69203d20", 20225 => x"2569290a",
    20226 => x"00000000", 20227 => x"2573544c", 20228 => x"563a2074",
    20229 => x"79706520", 20230 => x"25303478", 20231 => x"206c656e",
    20232 => x"20256920", 20233 => x"6f756920", 20234 => x"25303278",
    20235 => x"3a253032", 20236 => x"783a2530", 20237 => x"32782073",
    20238 => x"75622025", 20239 => x"3032783a", 20240 => x"25303278",
    20241 => x"3a253032", 20242 => x"780a0000", 20243 => x"2573544c",
    20244 => x"563a2074", 20245 => x"6f6f2073", 20246 => x"686f7274",
    20247 => x"20286578", 20248 => x"70656374", 20249 => x"65642025",
    20250 => x"692c2074", 20251 => x"6f74616c", 20252 => x"20256929",
    20253 => x"0a000000", 20254 => x"544c563a", 20255 => x"20000000",
    20256 => x"746c762d", 20257 => x"636f6e74", 20258 => x"656e7400",
    20259 => x"44554d50", 20260 => x"3a200000", 20261 => x"7061796c",
    20262 => x"6f616400", 20263 => x"20696e76", 20264 => x"616c6964",
    20265 => x"00000000", 20266 => x"25735449", 20267 => x"4d453a20",
    20268 => x"28256c69", 20269 => x"202d2030", 20270 => x"78256c78",
    20271 => x"2920256c", 20272 => x"692e2530", 20273 => x"366c6925",
    20274 => x"730a0000", 20275 => x"2573564c", 20276 => x"414e2025",
    20277 => x"690a0000", 20278 => x"25734554", 20279 => x"483a2025",
    20280 => x"30347820", 20281 => x"28253032", 20282 => x"783a2530",
    20283 => x"32783a25", 20284 => x"3032783a", 20285 => x"25303278",
    20286 => x"3a253032", 20287 => x"783a2530", 20288 => x"3278202d",
    20289 => x"3e202530", 20290 => x"32783a25", 20291 => x"3032783a",
    20292 => x"25303278", 20293 => x"3a253032", 20294 => x"783a2530",
    20295 => x"32783a25", 20296 => x"30327829", 20297 => x"0a000000",
    20298 => x"25734950", 20299 => x"3a202569", 20300 => x"20282569",
    20301 => x"2e25692e", 20302 => x"25692e25", 20303 => x"69202d3e",
    20304 => x"2025692e", 20305 => x"25692e25", 20306 => x"692e2569",
    20307 => x"29206c65", 20308 => x"6e202569", 20309 => x"0a000000",
    20310 => x"25735544", 20311 => x"503a2028", 20312 => x"2569202d",
    20313 => x"3e202569", 20314 => x"29206c65", 20315 => x"6e202569",
    20316 => x"0a000000", 20317 => x"25733a20", 20318 => x"256c690a",
    20319 => x"00000000", 20320 => x"5761726e", 20321 => x"696e673a",
    20322 => x"2025733a", 20323 => x"2063616e", 20324 => x"206e6f74",
    20325 => x"2061646a", 20326 => x"75737420", 20327 => x"66726571",
    20328 => x"5f707062", 20329 => x"20256c69", 20330 => x"0a000000",
    20331 => x"25733a20", 20332 => x"25396c75", 20333 => x"2e253039",
    20334 => x"6c690a00", 20335 => x"25733a20", 20336 => x"736e743d",
    20337 => x"25642c20", 20338 => x"7365633d", 20339 => x"25642c20",
    20340 => x"6e736563", 20341 => x"3d25640a", 20342 => x"00000000",
    20343 => x"73656e64", 20344 => x"3a200000", 20345 => x"72656376",
    20346 => x"3a200000", 20347 => x"696e6974", 20348 => x"69616c69",
    20349 => x"7a696e67", 20350 => x"00000000", 20351 => x"6661756c",
    20352 => x"74790000", 20353 => x"64697361", 20354 => x"626c6564",
    20355 => x"00000000", 20356 => x"6c697374", 20357 => x"656e696e",
    20358 => x"67000000", 20359 => x"756e6361", 20360 => x"6c696272",
    20361 => x"61746564", 20362 => x"00000000", 20363 => x"736c6176",
    20364 => x"65000000", 20365 => x"756e6361", 20366 => x"6c696272",
    20367 => x"61746564", 20368 => x"2f77722d", 20369 => x"70726573",
    20370 => x"656e7400", 20371 => x"6d617374", 20372 => x"65722f77",
    20373 => x"722d6d2d", 20374 => x"6c6f636b", 20375 => x"00000000",
    20376 => x"756e6361", 20377 => x"6c696272", 20378 => x"61746564",
    20379 => x"2f77722d", 20380 => x"732d6c6f", 20381 => x"636b0000",
    20382 => x"756e6361", 20383 => x"6c696272", 20384 => x"61746564",
    20385 => x"2f77722d", 20386 => x"6c6f636b", 20387 => x"65640000",
    20388 => x"77722d63", 20389 => x"616c6962", 20390 => x"72617469",
    20391 => x"6f6e0000", 20392 => x"77722d63", 20393 => x"616c6962",
    20394 => x"72617465", 20395 => x"64000000", 20396 => x"77722d72",
    20397 => x"6573702d", 20398 => x"63616c69", 20399 => x"622d7265",
    20400 => x"71000000", 20401 => x"77722d6c", 20402 => x"696e6b2d",
    20403 => x"6f6e0000", 20404 => x"686f6f6b", 20405 => x"3a202573",
    20406 => x"0a000000", 20407 => x"5432206f", 20408 => x"72205433",
    20409 => x"20696e63", 20410 => x"6f727265", 20411 => x"63742c20",
    20412 => x"64697363", 20413 => x"61726469", 20414 => x"6e672074",
    20415 => x"75706c65", 20416 => x"0a000000", 20417 => x"48616e64",
    20418 => x"7368616b", 20419 => x"65206661", 20420 => x"696c7572",
    20421 => x"653a206e", 20422 => x"6f77206e", 20423 => x"6f6e2d77",
    20424 => x"72202573", 20425 => x"0a000000", 20426 => x"52657472",
    20427 => x"79206f6e", 20428 => x"2074696d", 20429 => x"656f7574",
    20430 => x"0a000000", 20431 => x"25733a20", 20432 => x"73756273",
    20433 => x"74617465", 20434 => x"2025690a", 20435 => x"00000000",
    20436 => x"54783d3e", 20437 => x"3e736361", 20438 => x"6c656450",
    20439 => x"69636f73", 20440 => x"65636f6e", 20441 => x"64732e6d",
    20442 => x"7362203d", 20443 => x"20307825", 20444 => x"780a0000",
    20445 => x"54783d3e", 20446 => x"3e736361", 20447 => x"6c656450",
    20448 => x"69636f73", 20449 => x"65636f6e", 20450 => x"64732e6c",
    20451 => x"7362203d", 20452 => x"20307825", 20453 => x"780a0000",
    20454 => x"52782066", 20455 => x"69786564", 20456 => x"2064656c",
    20457 => x"6179203d", 20458 => x"2025640a", 20459 => x"00000000",
    20460 => x"52783d3e", 20461 => x"3e736361", 20462 => x"6c656450",
    20463 => x"69636f73", 20464 => x"65636f6e", 20465 => x"64732e6d",
    20466 => x"7362203d", 20467 => x"20307825", 20468 => x"780a0000",
    20469 => x"52783d3e", 20470 => x"3e736361", 20471 => x"6c656450",
    20472 => x"69636f73", 20473 => x"65636f6e", 20474 => x"64732e6c",
    20475 => x"7362203d", 20476 => x"20307825", 20477 => x"780a0000",
    20478 => x"4552524f", 20479 => x"523a204e", 20480 => x"65772063",
    20481 => x"6c617373", 20482 => x"2025690a", 20483 => x"00000000",
    20484 => x"4255473a", 20485 => x"20547279", 20486 => x"696e6720",
    20487 => x"746f2073", 20488 => x"656e6420", 20489 => x"696e7661",
    20490 => x"6c696420", 20491 => x"77725f6d", 20492 => x"7367206d",
    20493 => x"6f64653d", 20494 => x"25782069", 20495 => x"643d2578",
    20496 => x"00000000", 20497 => x"68616e64", 20498 => x"6c652053",
    20499 => x"69676e61", 20500 => x"6c696e67", 20501 => x"206d7367",
    20502 => x"2c206661", 20503 => x"696c6564", 20504 => x"2c205468",
    20505 => x"69732069", 20506 => x"73206e6f", 20507 => x"74206f72",
    20508 => x"67616e69", 20509 => x"7a617469", 20510 => x"6f6e2065",
    20511 => x"7874656e", 20512 => x"73696f6e", 20513 => x"20544c56",
    20514 => x"203d2030", 20515 => x"7825780a", 20516 => x"00000000",
    20517 => x"68616e64", 20518 => x"6c652053", 20519 => x"69676e61",
    20520 => x"6c696e67", 20521 => x"206d7367", 20522 => x"2c206661",
    20523 => x"696c6564", 20524 => x"2c206e6f", 20525 => x"74204345",
    20526 => x"524e2773", 20527 => x"204f5549", 20528 => x"203d2030",
    20529 => x"7825780a", 20530 => x"00000000", 20531 => x"68616e64",
    20532 => x"6c652053", 20533 => x"69676e61", 20534 => x"6c696e67",
    20535 => x"206d7367", 20536 => x"2c206661", 20537 => x"696c6564",
    20538 => x"2c206e6f", 20539 => x"74205768", 20540 => x"69746520",
    20541 => x"52616262", 20542 => x"6974206d", 20543 => x"61676963",
    20544 => x"206e756d", 20545 => x"62657220", 20546 => x"3d203078",
    20547 => x"25780a00", 20548 => x"68616e64", 20549 => x"6c652053",
    20550 => x"69676e61", 20551 => x"6c696e67", 20552 => x"206d7367",
    20553 => x"2c206661", 20554 => x"696c6564", 20555 => x"2c206e6f",
    20556 => x"74207375", 20557 => x"70706f72", 20558 => x"74656420",
    20559 => x"76657273", 20560 => x"696f6e20", 20561 => x"6e756d62",
    20562 => x"6572203d", 20563 => x"20307825", 20564 => x"780a0000",
    20565 => x"25732825", 20566 => x"6429204d", 20567 => x"65737361",
    20568 => x"67652063", 20569 => x"616e2774", 20570 => x"20626520",
    20571 => x"73656e74", 20572 => x"0a000000", 20573 => x"53454e54",
    20574 => x"20253032", 20575 => x"64206279", 20576 => x"74657320",
    20577 => x"61742025", 20578 => x"642e2530", 20579 => x"39642028",
    20580 => x"2573290a", 20581 => x"00000000", 20582 => x"556e696e",
    20583 => x"69746961", 20584 => x"6c697a65", 20585 => x"64000000",
    20586 => x"20287761", 20587 => x"69742066", 20588 => x"6f722068",
    20589 => x"77290000", 20590 => x"4552524f", 20591 => x"523a2025",
    20592 => x"733a2054", 20593 => x"696d6573", 20594 => x"74616d70",
    20595 => x"73496e63", 20596 => x"6f727265", 20597 => x"63743a20",
    20598 => x"25642025", 20599 => x"64202564", 20600 => x"2025640a",
    20601 => x"00000000", 20602 => x"2573203d", 20603 => x"2025643a",
    20604 => x"25643a25", 20605 => x"640a0000", 20606 => x"73657276",
    20607 => x"6f3a7431", 20608 => x"00000000", 20609 => x"73657276",
    20610 => x"6f3a7432", 20611 => x"00000000", 20612 => x"73657276",
    20613 => x"6f3a7433", 20614 => x"00000000", 20615 => x"73657276",
    20616 => x"6f3a7434", 20617 => x"00000000", 20618 => x"2d3e6d64",
    20619 => x"656c6179", 20620 => x"00000000", 20621 => x"504c4c20",
    20622 => x"4f75744f", 20623 => x"664c6f63", 20624 => x"6b2c2073",
    20625 => x"686f756c", 20626 => x"64207265", 20627 => x"73746172",
    20628 => x"74207379", 20629 => x"6e630a00", 20630 => x"73657276",
    20631 => x"6f3a6275", 20632 => x"73790a00", 20633 => x"6f666673",
    20634 => x"65745f68", 20635 => x"773a2025", 20636 => x"6c692e25",
    20637 => x"30396c69", 20638 => x"20282b25", 20639 => x"6c69290a",
    20640 => x"00000000", 20641 => x"77725f73", 20642 => x"6572766f",
    20643 => x"20737461", 20644 => x"74653a20", 20645 => x"25732573",
    20646 => x"0a000000", 20647 => x"6f6c6473", 20648 => x"65747020",
    20649 => x"25692c20", 20650 => x"6f666673", 20651 => x"65742025",
    20652 => x"693a2530", 20653 => x"34690a00", 20654 => x"61646a75",
    20655 => x"73742070", 20656 => x"68617365", 20657 => x"2025690a",
    20658 => x"00000000", 20659 => x"53594e43", 20660 => x"5f4e5345",
    20661 => x"43000000", 20662 => x"53594e43", 20663 => x"5f534543",
    20664 => x"00000000", 20665 => x"53594e43", 20666 => x"5f504841",
    20667 => x"53450000", 20668 => x"54524143", 20669 => x"4b5f5048",
    20670 => x"41534500", 20671 => x"57414954", 20672 => x"5f4f4646",
    20673 => x"5345545f", 20674 => x"53544142", 20675 => x"4c450000",
    20676 => x"7072652d", 20677 => x"6d617374", 20678 => x"65720000",
    20679 => x"70617373", 20680 => x"69766500", 20681 => x"25733a20",
    20682 => x"63616e27", 20683 => x"7420696e", 20684 => x"69742065",
    20685 => x"7874656e", 20686 => x"73696f6e", 20687 => x"0a000000",
    20688 => x"636c6f63", 20689 => x"6b20636c", 20690 => x"61737320",
    20691 => x"3d202564", 20692 => x"0a000000", 20693 => x"636c6f63",
    20694 => x"6b206163", 20695 => x"63757261", 20696 => x"6379203d",
    20697 => x"2025640a", 20698 => x"00000000", 20699 => x"70705f73",
    20700 => x"6c617665", 20701 => x"203a2044", 20702 => x"656c6179",
    20703 => x"20526573", 20704 => x"7020646f", 20705 => x"65736e27",
    20706 => x"74206d61", 20707 => x"74636820", 20708 => x"44656c61",
    20709 => x"79205265", 20710 => x"710a0000", 20711 => x"4e657720",
    20712 => x"666f7265", 20713 => x"69676e20", 20714 => x"4d617374",
    20715 => x"65722025", 20716 => x"69206164", 20717 => x"6465640a",
    20718 => x"00000000", 20719 => x"4552524f", 20720 => x"523a2025",
    20721 => x"733a2046", 20722 => x"6f6c6c6f", 20723 => x"77207570",
    20724 => x"206d6573", 20725 => x"73616765", 20726 => x"20697320",
    20727 => x"6e6f7420", 20728 => x"66726f6d", 20729 => x"20637572",
    20730 => x"72656e74", 20731 => x"20706172", 20732 => x"656e740a",
    20733 => x"00000000", 20734 => x"4552524f", 20735 => x"523a2025",
    20736 => x"733a2053", 20737 => x"6c617665", 20738 => x"20776173",
    20739 => x"206e6f74", 20740 => x"20776169", 20741 => x"74696e67",
    20742 => x"20612066", 20743 => x"6f6c6c6f", 20744 => x"77207570",
    20745 => x"206d6573", 20746 => x"73616765", 20747 => x"0a000000",
    20748 => x"4552524f", 20749 => x"523a2025", 20750 => x"733a2053",
    20751 => x"65717565", 20752 => x"6e636549", 20753 => x"44202564",
    20754 => x"20646f65", 20755 => x"736e2774", 20756 => x"206d6174",
    20757 => x"6368206c", 20758 => x"61737420", 20759 => x"53796e63",
    20760 => x"206d6573", 20761 => x"73616765", 20762 => x"2025640a",
    20763 => x"00000000", 20764 => x"416e6e6f", 20765 => x"756e6365",
    20766 => x"206d6573", 20767 => x"73616765", 20768 => x"2066726f",
    20769 => x"6d20616e", 20770 => x"6f746865", 20771 => x"7220666f",
    20772 => x"72656967", 20773 => x"6e206d61", 20774 => x"73746572",
    20775 => x"0a000000", 20776 => x"25733a25", 20777 => x"693a2045",
    20778 => x"72726f72", 20779 => x"20310a00", 20780 => x"25733a25",
    20781 => x"693a2045", 20782 => x"72726f72", 20783 => x"20320a00",
    20784 => x"42657374", 20785 => x"20666f72", 20786 => x"6569676e",
    20787 => x"206d6173", 20788 => x"74657220", 20789 => x"69732025",
    20790 => x"692f2569", 20791 => x"0a000000", 20792 => x"25733a20",
    20793 => x"6572726f", 20794 => x"720a0000", 20795 => x"25733a20",
    20796 => x"70617373", 20797 => x"6976650a", 20798 => x"00000000",
    20799 => x"25733a20", 20800 => x"6d617374", 20801 => x"65720a00",
    20802 => x"4e657720", 20803 => x"55544320", 20804 => x"6f666673",
    20805 => x"65743a20", 20806 => x"25690a00", 20807 => x"25733a20",
    20808 => x"736c6176", 20809 => x"650a0000", 20810 => x"73796e63",
    20811 => x"00000000", 20812 => x"64656c61", 20813 => x"795f7265",
    20814 => x"71000000", 20815 => x"7064656c", 20816 => x"61795f72",
    20817 => x"65710000", 20818 => x"7064656c", 20819 => x"61795f72",
    20820 => x"65737000", 20821 => x"64656c61", 20822 => x"795f7265",
    20823 => x"73700000", 20824 => x"7064656c", 20825 => x"61795f72",
    20826 => x"6573705f", 20827 => x"666f6c6c", 20828 => x"6f775f75",
    20829 => x"70000000", 20830 => x"616e6e6f", 20831 => x"756e6365",
    20832 => x"00000000", 20833 => x"7369676e", 20834 => x"616c696e",
    20835 => x"67000000", 20836 => x"6d616e61", 20837 => x"67656d65",
    20838 => x"6e740000", 20839 => x"4552524f", 20840 => x"523a2042",
    20841 => x"55473a20", 20842 => x"25732064", 20843 => x"6f65736e",
    20844 => x"27742073", 20845 => x"7570706f", 20846 => x"7274206e",
    20847 => x"65676174", 20848 => x"69766573", 20849 => x"0a000000",
    20850 => x"4552524f", 20851 => x"523a204e", 20852 => x"65676174",
    20853 => x"69766520", 20854 => x"76616c75", 20855 => x"65206361",
    20856 => x"6e6e6f74", 20857 => x"20626520", 20858 => x"636f6e76",
    20859 => x"65727465", 20860 => x"6420696e", 20861 => x"746f2074",
    20862 => x"696d6573", 20863 => x"74616d70", 20864 => x"0a000000",
    20865 => x"4552524f", 20866 => x"523a2074", 20867 => x"6f5f5469",
    20868 => x"6d65496e", 20869 => x"7465726e", 20870 => x"616c3a20",
    20871 => x"7365636f", 20872 => x"6e647320", 20873 => x"6669656c",
    20874 => x"64206973", 20875 => x"20686967", 20876 => x"68657220",
    20877 => x"7468616e", 20878 => x"20736967", 20879 => x"6e656420",
    20880 => x"696e7465", 20881 => x"67657220", 20882 => x"28333262",
    20883 => x"69747329", 20884 => x"0a000000", 20885 => x"2d000000",
    20886 => x"25732564", 20887 => x"2e253039", 20888 => x"64000000",
    20889 => x"6572726f", 20890 => x"7220696e", 20891 => x"20745f6f",
    20892 => x"70732d3e", 20893 => x"73657276", 20894 => x"6f5f696e",
    20895 => x"69740000", 20896 => x"496e6974", 20897 => x"69616c69",
    20898 => x"7a65643a", 20899 => x"206f6273", 20900 => x"5f647269",
    20901 => x"66742025", 20902 => x"6c6c690a", 20903 => x"00000000",
    20904 => x"636f7272", 20905 => x"65637469", 20906 => x"6f6e2066",
    20907 => x"69656c64", 20908 => x"20313a20", 20909 => x"25730a00",
    20910 => x"64697363", 20911 => x"61726420", 20912 => x"54332f54",
    20913 => x"343a2077", 20914 => x"65206d69", 20915 => x"73732054",
    20916 => x"312f5432", 20917 => x"0a000000", 20918 => x"636f7272",
    20919 => x"65637469", 20920 => x"6f6e2066", 20921 => x"69656c64",
    20922 => x"20323a20", 20923 => x"25730a00", 20924 => x"54313a20",
    20925 => x"25730a00", 20926 => x"54323a20", 20927 => x"25730a00",
    20928 => x"54333a20", 20929 => x"25730a00", 20930 => x"54343a20",
    20931 => x"25730a00", 20932 => x"4d617374", 20933 => x"65722074",
    20934 => x"6f20736c", 20935 => x"6176653a", 20936 => x"2025730a",
    20937 => x"00000000", 20938 => x"536c6176", 20939 => x"6520746f",
    20940 => x"206d6173", 20941 => x"7465723a", 20942 => x"2025730a",
    20943 => x"00000000", 20944 => x"6d65616e", 20945 => x"50617468",
    20946 => x"44656c61", 20947 => x"793a2025", 20948 => x"730a0000",
    20949 => x"73657276", 20950 => x"6f206162", 20951 => x"6f727465",
    20952 => x"642c2064", 20953 => x"656c6179", 20954 => x"20677265",
    20955 => x"61746572", 20956 => x"20746861", 20957 => x"6e203120",
    20958 => x"7365636f", 20959 => x"6e640a00", 20960 => x"73657276",
    20961 => x"6f206162", 20962 => x"6f727465", 20963 => x"642c2064",
    20964 => x"656c6179", 20965 => x"20256420", 20966 => x"6f722025",
    20967 => x"64206772", 20968 => x"65617465", 20969 => x"72207468",
    20970 => x"616e2063", 20971 => x"6f6e6669", 20972 => x"67757265",
    20973 => x"64206d61", 20974 => x"78696d75", 20975 => x"6d202564",
    20976 => x"0a000000", 20977 => x"5472696d", 20978 => x"20746f6f",
    20979 => x"2d6c6f6e", 20980 => x"67206d70", 20981 => x"643a2025",
    20982 => x"690a0000", 20983 => x"41667465", 20984 => x"72206176",
    20985 => x"67282569", 20986 => x"292c206d", 20987 => x"65616e50",
    20988 => x"61746844", 20989 => x"656c6179", 20990 => x"3a202569",
    20991 => x"0a000000", 20992 => x"4f666673", 20993 => x"65742066",
    20994 => x"726f6d20", 20995 => x"6d617374", 20996 => x"65723a20",
    20997 => x"20202020", 20998 => x"25730a00", 20999 => x"73657276",
    21000 => x"6f206162", 21001 => x"6f727465", 21002 => x"642c206f",
    21003 => x"66667365", 21004 => x"74206772", 21005 => x"65617465",
    21006 => x"72207468", 21007 => x"616e2031", 21008 => x"20736563",
    21009 => x"6f6e640a", 21010 => x"00000000", 21011 => x"73657276",
    21012 => x"6f206162", 21013 => x"6f727465", 21014 => x"642c206f",
    21015 => x"66667365", 21016 => x"74206772", 21017 => x"65617465",
    21018 => x"72207468", 21019 => x"616e2063", 21020 => x"6f6e6669",
    21021 => x"67757265", 21022 => x"64206d61", 21023 => x"78696d75",
    21024 => x"6d202564", 21025 => x"0a000000", 21026 => x"4f627365",
    21027 => x"72766564", 21028 => x"20647269", 21029 => x"66743a20",
    21030 => x"2539690a", 21031 => x"00000000", 21032 => x"74696d65",
    21033 => x"6f757420", 21034 => x"65787069", 21035 => x"7265643a",
    21036 => x"2025730a", 21037 => x"00000000", 21038 => x"50505f54",
    21039 => x"4f5f4445", 21040 => x"4c415952", 21041 => x"45510000",
    21042 => x"50505f54", 21043 => x"4f5f5359", 21044 => x"4e430000",
    21045 => x"50505f54", 21046 => x"4f5f414e", 21047 => x"4e5f5245",
    21048 => x"43454950", 21049 => x"54000000", 21050 => x"50505f54",
    21051 => x"4f5f414e", 21052 => x"4e5f494e", 21053 => x"54455256",
    21054 => x"414c0000", 21055 => x"50505f54", 21056 => x"4f5f4641",
    21057 => x"554c5459", 21058 => x"00000000", 21059 => x"50505f54",
    21060 => x"4f5f4558", 21061 => x"545f3000", 21062 => x"50505f54",
    21063 => x"4f5f4558", 21064 => x"545f3100", 21065 => x"50505f54",
    21066 => x"4f5f4558", 21067 => x"545f3200", 21068 => x"536c6176",
    21069 => x"65204f6e", 21070 => x"6c792c20", 21071 => x"636c6f63",
    21072 => x"6b20636c", 21073 => x"61737320", 21074 => x"73657420",
    21075 => x"746f2032", 21076 => x"35350a00", 21077 => x"25750000",
    21078 => x"25752575", 21079 => x"00000000", 21080 => x"6c6e6b3a",
    21081 => x"25642072", 21082 => x"783a2564", 21083 => x"2074783a",
    21084 => x"25642000", 21085 => x"6c6f636b", 21086 => x"3a256420",
    21087 => x"00000000", 21088 => x"7074703a", 21089 => x"25732000",
    21090 => x"73763a25", 21091 => x"64200000", 21092 => x"73733a27",
    21093 => x"25732720", 21094 => x"00000000", 21095 => x"6175783a",
    21096 => x"25782000", 21097 => x"7365633a", 21098 => x"2564206e",
    21099 => x"7365633a", 21100 => x"25642000", 21101 => x"6d753a25",
    21102 => x"73200000", 21103 => x"646d733a", 21104 => x"25732000",
    21105 => x"6474786d", 21106 => x"3a256420", 21107 => x"6472786d",
    21108 => x"3a256420", 21109 => x"00000000", 21110 => x"64747873",
    21111 => x"3a256420", 21112 => x"64727873", 21113 => x"3a256420",
    21114 => x"00000000", 21115 => x"6173796d", 21116 => x"3a256420",
    21117 => x"00000000", 21118 => x"63727474", 21119 => x"3a257320",
    21120 => x"00000000", 21121 => x"636b6f3a", 21122 => x"25642000",
    21123 => x"73657470", 21124 => x"3a256420", 21125 => x"00000000",
    21126 => x"75636e74", 21127 => x"3a256420", 21128 => x"00000000",
    21129 => x"68643a25", 21130 => x"64206d64", 21131 => x"3a256420",
    21132 => x"61643a25", 21133 => x"64200000", 21134 => x"70636200",
    21135 => x"74656d70", 21136 => x"3a202564", 21137 => x"2e253034",
    21138 => x"64204300", 21139 => x"0a0a5054", 21140 => x"50207374",
    21141 => x"61747573", 21142 => x"3a200000", 21143 => x"25730000",
    21144 => x"0a0a5379", 21145 => x"6e632069", 21146 => x"6e666f20",
    21147 => x"6e6f7420", 21148 => x"76616c69", 21149 => x"640a0a00",
    21150 => x"0a0a5379", 21151 => x"6e636872", 21152 => x"6f6e697a",
    21153 => x"6174696f", 21154 => x"6e207374", 21155 => x"61747573",
    21156 => x"3a0a0a00", 21157 => x"57522050", 21158 => x"54502043",
    21159 => x"6f726520", 21160 => x"53796e63", 21161 => x"204d6f6e",
    21162 => x"69746f72", 21163 => x"20762031", 21164 => x"2e300000",
    21165 => x"45736320", 21166 => x"3d206578", 21167 => x"69740000",
    21168 => x"0a0a5441", 21169 => x"49205469", 21170 => x"6d653a20",
    21171 => x"20202020", 21172 => x"20202020", 21173 => x"20202020",
    21174 => x"20202020", 21175 => x"20000000", 21176 => x"0a0a4c69",
    21177 => x"6e6b2073", 21178 => x"74617475", 21179 => x"733a0000",
    21180 => x"25733a20", 21181 => x"00000000", 21182 => x"77727531",
    21183 => x"00000000", 21184 => x"4c696e6b", 21185 => x"20757020",
    21186 => x"20200000", 21187 => x"4c696e6b", 21188 => x"20646f77",
    21189 => x"6e200000", 21190 => x"2852583a", 21191 => x"2025642c",
    21192 => x"2054583a", 21193 => x"20256429", 21194 => x"2c206d6f",
    21195 => x"64653a20", 21196 => x"00000000", 21197 => x"5752204f",
    21198 => x"66660000", 21199 => x"436c6f63", 21200 => x"6b206f66",
    21201 => x"66736574", 21202 => x"3a202020", 21203 => x"20202020",
    21204 => x"20202020", 21205 => x"20202020", 21206 => x"20200000",
    21207 => x"2532692e", 21208 => x"25303969", 21209 => x"20730000",
    21210 => x"25396920", 21211 => x"6e730000", 21212 => x"0a4f6e65",
    21213 => x"2d776179", 21214 => x"2064656c", 21215 => x"61792061",
    21216 => x"76657261", 21217 => x"6765643a", 21218 => x"20202020",
    21219 => x"20202000", 21220 => x"0a4f6273", 21221 => x"65727665",
    21222 => x"64206472", 21223 => x"6966743a", 21224 => x"20202020",
    21225 => x"20202020", 21226 => x"20202020", 21227 => x"20202000",
    21228 => x"5752204d", 21229 => x"61737465", 21230 => x"72202000",
    21231 => x"57522053", 21232 => x"6c617665", 21233 => x"20202000",
    21234 => x"57522055", 21235 => x"6e6b6e6f", 21236 => x"776e2020",
    21237 => x"20000000", 21238 => x"4c6f636b", 21239 => x"65642020",
    21240 => x"00000000", 21241 => x"4e6f4c6f", 21242 => x"636b2020",
    21243 => x"00000000", 21244 => x"43616c69", 21245 => x"62726174",
    21246 => x"65642020", 21247 => x"00000000", 21248 => x"556e6361",
    21249 => x"6c696272", 21250 => x"61746564", 21251 => x"20200000",
    21252 => x"0a495076", 21253 => x"343a2000", 21254 => x"424f4f54",
    21255 => x"50207275", 21256 => x"6e6e696e", 21257 => x"67000000",
    21258 => x"25732028", 21259 => x"66726f6d", 21260 => x"20626f6f",
    21261 => x"74702900", 21262 => x"25732028", 21263 => x"73746174",
    21264 => x"69632061", 21265 => x"73736967", 21266 => x"6e6d656e",
    21267 => x"74290000", 21268 => x"53657276", 21269 => x"6f207374",
    21270 => x"6174653a", 21271 => x"20202020", 21272 => x"20202020",
    21273 => x"20202020", 21274 => x"20202000", 21275 => x"50686173",
    21276 => x"65207472", 21277 => x"61636b69", 21278 => x"6e673a20",
    21279 => x"20202020", 21280 => x"20202020", 21281 => x"20202000",
    21282 => x"4f4e0a00", 21283 => x"4f46460a", 21284 => x"00000000",
    21285 => x"41757820", 21286 => x"636c6f63", 21287 => x"6b207374",
    21288 => x"61747573", 21289 => x"3a202020", 21290 => x"20202020",
    21291 => x"20202000", 21292 => x"656e6162", 21293 => x"6c656400",
    21294 => x"2c206c6f", 21295 => x"636b6564", 21296 => x"00000000",
    21297 => x"0a54696d", 21298 => x"696e6720", 21299 => x"70617261",
    21300 => x"6d657465", 21301 => x"72733a0a", 21302 => x"0a000000",
    21303 => x"526f756e", 21304 => x"642d7472", 21305 => x"69702074",
    21306 => x"696d6520", 21307 => x"286d7529", 21308 => x"3a202020",
    21309 => x"20000000", 21310 => x"25732070", 21311 => x"730a0000",
    21312 => x"4d617374", 21313 => x"65722d73", 21314 => x"6c617665",
    21315 => x"2064656c", 21316 => x"61793a20", 21317 => x"20202020",
    21318 => x"20000000", 21319 => x"4d617374", 21320 => x"65722050",
    21321 => x"48592064", 21322 => x"656c6179", 21323 => x"733a2020",
    21324 => x"20202020", 21325 => x"20000000", 21326 => x"54583a20",
    21327 => x"25642070", 21328 => x"732c2052", 21329 => x"583a2025",
    21330 => x"64207073", 21331 => x"0a000000", 21332 => x"536c6176",
    21333 => x"65205048", 21334 => x"59206465", 21335 => x"6c617973",
    21336 => x"3a202020", 21337 => x"20202020", 21338 => x"20000000",
    21339 => x"546f7461", 21340 => x"6c206c69", 21341 => x"6e6b2061",
    21342 => x"73796d6d", 21343 => x"65747279", 21344 => x"3a202020",
    21345 => x"20000000", 21346 => x"25396420", 21347 => x"70730a00",
    21348 => x"4361626c", 21349 => x"65207274", 21350 => x"74206465",
    21351 => x"6c61793a", 21352 => x"20202020", 21353 => x"20202020",
    21354 => x"20000000", 21355 => x"436c6f63", 21356 => x"6b206f66",
    21357 => x"66736574", 21358 => x"3a202020", 21359 => x"20202020",
    21360 => x"20202020", 21361 => x"20000000", 21362 => x"50686173",
    21363 => x"65207365", 21364 => x"74706f69", 21365 => x"6e743a20",
    21366 => x"20202020", 21367 => x"20202020", 21368 => x"20000000",
    21369 => x"536b6577", 21370 => x"3a202020", 21371 => x"20202020",
    21372 => x"20202020", 21373 => x"20202020", 21374 => x"20202020",
    21375 => x"20000000", 21376 => x"55706461", 21377 => x"74652063",
    21378 => x"6f756e74", 21379 => x"65723a20", 21380 => x"20202020",
    21381 => x"20202020", 21382 => x"20000000", 21383 => x"2539640a",
    21384 => x"00000000", 21385 => x"2d2d0000", 21386 => x"756e6b6e",
    21387 => x"6f776e00", 21388 => x"73746174", 21389 => x"73000000",
    21390 => x"1b5b3125", 21391 => x"63000000", 21392 => x"436f6d6d",
    21393 => x"616e6420", 21394 => x"22257322", 21395 => x"3a206572",
    21396 => x"726f7220", 21397 => x"25640a00", 21398 => x"556e7265",
    21399 => x"636f676e", 21400 => x"697a6564", 21401 => x"20636f6d",
    21402 => x"6d616e64", 21403 => x"20222573", 21404 => x"222e0a00",
    21405 => x"77726323", 21406 => x"20000000", 21407 => x"25630000",
    21408 => x"456d7074", 21409 => x"7920696e", 21410 => x"69742073",
    21411 => x"63726970", 21412 => x"742e2e2e", 21413 => x"0a000000",
    21414 => x"65786563", 21415 => x"7574696e", 21416 => x"673a2025",
    21417 => x"730a0000", 21418 => x"57522043", 21419 => x"6f726520",
    21420 => x"6275696c", 21421 => x"643a2025", 21422 => x"7325730a",
    21423 => x"00000000", 21424 => x"2028756e", 21425 => x"73757070",
    21426 => x"6f727465", 21427 => x"64206465", 21428 => x"76656c6f",
    21429 => x"70657220", 21430 => x"6275696c", 21431 => x"64290000",
    21432 => x"4275696c", 21433 => x"743a2025", 21434 => x"73202573",
    21435 => x"20627920", 21436 => x"25730a00", 21437 => x"4275696c",
    21438 => x"7420666f", 21439 => x"72202564", 21440 => x"206b4220",
    21441 => x"52414d2c", 21442 => x"20737461", 21443 => x"636b2069",
    21444 => x"73202564", 21445 => x"20627974", 21446 => x"65730a00",
    21447 => x"5741524e", 21448 => x"494e473a", 21449 => x"20686172",
    21450 => x"64776172", 21451 => x"65207361", 21452 => x"79732025",
    21453 => x"696b4220", 21454 => x"3c3d2052", 21455 => x"414d203c",
    21456 => x"2025696b", 21457 => x"420a0000", 21458 => x"76657200",
    21459 => x"73746172", 21460 => x"74000000", 21461 => x"73746f70",
    21462 => x"00000000", 21463 => x"676d0000", 21464 => x"6d6f6465",
    21465 => x"00000000", 21466 => x"6772616e", 21467 => x"646d6173",
    21468 => x"74657200", 21469 => x"41766169", 21470 => x"6c61626c",
    21471 => x"6520636f", 21472 => x"6d6d616e", 21473 => x"64733a0a",
    21474 => x"00000000", 21475 => x"20202573", 21476 => x"0a000000",
    21477 => x"68656c70", 21478 => x"00000000", 21479 => x"25303278",
    21480 => x"3a253032", 21481 => x"783a2530", 21482 => x"32783a25",
    21483 => x"3032783a", 21484 => x"25303278", 21485 => x"3a253032",
    21486 => x"78000000", 21487 => x"67657400", 21488 => x"67657470",
    21489 => x"00000000", 21490 => x"73657400", 21491 => x"73657470",
    21492 => x"00000000", 21493 => x"4d41432d", 21494 => x"61646472",
    21495 => x"6573733a", 21496 => x"2025730a", 21497 => x"00000000",
    21498 => x"6d616300", 21499 => x"72657365", 21500 => x"74000000",
    21501 => x"20697465", 21502 => x"72617469", 21503 => x"6f6e7320",
    21504 => x"20202020", 21505 => x"7365636f", 21506 => x"6e64732e",
    21507 => x"6d696372", 21508 => x"6f732020", 21509 => x"20206e61",
    21510 => x"6d650a00", 21511 => x"20202539", 21512 => x"6c692020",
    21513 => x"2025396c", 21514 => x"692e2530", 21515 => x"366c6920",
    21516 => x"2025730a", 21517 => x"00000000", 21518 => x"70730000",
    21519 => x"55736167", 21520 => x"653a2072", 21521 => x"65667265",
    21522 => x"7368203c", 21523 => x"7365636f", 21524 => x"6e64733e",
    21525 => x"0a000000", 21526 => x"72656672", 21527 => x"65736800",
    21528 => x"73746174", 21529 => x"69737469", 21530 => x"6373206e",
    21531 => x"6f77206f", 21532 => x"66660a00", 21533 => x"62747300",
    21534 => x"6f666600", 21535 => x"73746174", 21536 => x"00000000",
    21537 => x"57726f6e", 21538 => x"67207061", 21539 => x"72616d65",
    21540 => x"7465720a", 21541 => x"00000000", 21542 => x"65726173",
    21543 => x"65000000", 21544 => x"436f756c", 21545 => x"64206e6f",
    21546 => x"74206572", 21547 => x"61736520", 21548 => x"44420a00",
    21549 => x"61646400", 21550 => x"53465020", 21551 => x"44422069",
    21552 => x"73206675", 21553 => x"6c6c0a00", 21554 => x"49324320",
    21555 => x"6572726f", 21556 => x"720a0000", 21557 => x"53465020",
    21558 => x"64617461", 21559 => x"62617365", 21560 => x"20657272",
    21561 => x"6f722028", 21562 => x"2564290a", 21563 => x"00000000",
    21564 => x"25642053", 21565 => x"46507320", 21566 => x"696e2044",
    21567 => x"420a0000", 21568 => x"73686f77", 21569 => x"00000000",
    21570 => x"53465020", 21571 => x"64617461", 21572 => x"62617365",
    21573 => x"20656d70", 21574 => x"74790a00", 21575 => x"25643a20",
    21576 => x"504e3a00", 21577 => x"20645478", 21578 => x"3a202538",
    21579 => x"64206452", 21580 => x"783a2025", 21581 => x"38642061",
    21582 => x"6c706861", 21583 => x"3a202538", 21584 => x"640a0000",
    21585 => x"6d617463", 21586 => x"68000000", 21587 => x"4e6f2053",
    21588 => x"46502e0a", 21589 => x"00000000", 21590 => x"53465020",
    21591 => x"72656164", 21592 => x"20657272", 21593 => x"6f720a00",
    21594 => x"436f756c", 21595 => x"64206e6f", 21596 => x"74206d61",
    21597 => x"74636820", 21598 => x"746f2044", 21599 => x"420a0000",
    21600 => x"53465020", 21601 => x"6d617463", 21602 => x"6865642c",
    21603 => x"20645478", 21604 => x"3d256420", 21605 => x"6452783d",
    21606 => x"25642061", 21607 => x"6c706861", 21608 => x"3d25640a",
    21609 => x"00000000", 21610 => x"656e6100", 21611 => x"73667000",
    21612 => x"696e6974", 21613 => x"00000000", 21614 => x"636c0000",
    21615 => x"73707300", 21616 => x"67707300", 21617 => x"25642025",
    21618 => x"640a0000", 21619 => x"73646163", 21620 => x"00000000",
    21621 => x"67646163", 21622 => x"00000000", 21623 => x"63686563",
    21624 => x"6b76636f", 21625 => x"00000000", 21626 => x"706c6c00",
    21627 => x"666f7263", 21628 => x"65000000", 21629 => x"466f756e",
    21630 => x"64207068", 21631 => x"61736520", 21632 => x"7472616e",
    21633 => x"73697469", 21634 => x"6f6e2069", 21635 => x"6e204545",
    21636 => x"50524f4d", 21637 => x"3a202564", 21638 => x"70730a00",
    21639 => x"4d656173", 21640 => x"7572696e", 21641 => x"67207432",
    21642 => x"2f743420", 21643 => x"70686173", 21644 => x"65207472",
    21645 => x"616e7369", 21646 => x"74696f6e", 21647 => x"2e2e2e0a",
    21648 => x"00000000", 21649 => x"63616c69", 21650 => x"62726174",
    21651 => x"696f6e00", 21652 => x"73657473", 21653 => x"65630000",
    21654 => x"7365746e", 21655 => x"73656300", 21656 => x"72617700",
    21657 => x"2573202b", 21658 => x"2564206e", 21659 => x"616e6f73",
    21660 => x"65636f6e", 21661 => x"64732e0a", 21662 => x"00000000",
    21663 => x"74696d65", 21664 => x"00000000", 21665 => x"67756900",
    21666 => x"73646200", 21667 => x"4f4e0000", 21668 => x"4f464600",
    21669 => x"656e6162", 21670 => x"6c650000", 21671 => x"64697361",
    21672 => x"626c6500", 21673 => x"70686173", 21674 => x"65207472",
    21675 => x"61636b69", 21676 => x"6e672025", 21677 => x"730a0000",
    21678 => x"70747261", 21679 => x"636b0000", 21680 => x"63616c63",
    21681 => x"00000000", 21682 => x"63683100", 21683 => x"63683200",
    21684 => x"70636e00", 21685 => x"25642e25", 21686 => x"642e2564",
    21687 => x"2e256400", 21688 => x"49502d61", 21689 => x"64647265",
    21690 => x"73733a20", 21691 => x"696e2074", 21692 => x"7261696e",
    21693 => x"696e670a", 21694 => x"00000000", 21695 => x"49502d61",
    21696 => x"64647265", 21697 => x"73733a20", 21698 => x"25732028",
    21699 => x"66726f6d", 21700 => x"20626f6f", 21701 => x"7470290a",
    21702 => x"00000000", 21703 => x"49502d61", 21704 => x"64647265",
    21705 => x"73733a20", 21706 => x"25732028", 21707 => x"73746174",
    21708 => x"69632061", 21709 => x"73736967", 21710 => x"6e6d656e",
    21711 => x"74290a00", 21712 => x"69700000", 21713 => x"50505349",
    21714 => x"20766572", 21715 => x"626f7369", 21716 => x"74793a20",
    21717 => x"2530386c", 21718 => x"780a0000", 21719 => x"76657262",
    21720 => x"6f736500", 21721 => x"436f756c", 21722 => x"64206e6f",
    21723 => x"74206572", 21724 => x"61736520", 21725 => x"696e6974",
    21726 => x"20736372", 21727 => x"6970740a", 21728 => x"00000000",
    21729 => x"436f756c", 21730 => x"64206e6f", 21731 => x"74206164",
    21732 => x"64207468", 21733 => x"6520636f", 21734 => x"6d6d616e",
    21735 => x"640a0000", 21736 => x"4f4b2e0a", 21737 => x"00000000",
    21738 => x"626f6f74", 21739 => x"00000000", 21740 => x"25732c20",
    21741 => x"25732025", 21742 => x"642c2025", 21743 => x"642c2025",
    21744 => x"3032643a", 21745 => x"25303264", 21746 => x"3a253032",
    21747 => x"64000000", 21748 => x"25732025", 21749 => x"32642025",
    21750 => x"3032643a", 21751 => x"25303264", 21752 => x"3a253032",
    21753 => x"64000000", 21754 => x"2534642d", 21755 => x"25303264",
    21756 => x"2d253032", 21757 => x"642d2530", 21758 => x"32643a25",
    21759 => x"3032643a", 21760 => x"25303264", 21761 => x"00000000",
    21762 => x"1b5b3025", 21763 => x"643b3325", 21764 => x"646d0000",
    21765 => x"1b5b6d00", 21766 => x"1b5b2564", 21767 => x"3b256466",
    21768 => x"00000000", 21769 => x"1b5b324a", 21770 => x"1b5b313b",
    21771 => x"31480000", 21772 => x"53756e00", 21773 => x"4d6f6e00",
    21774 => x"54756500", 21775 => x"57656400", 21776 => x"54687500",
    21777 => x"46726900", 21778 => x"53617400", 21779 => x"4a616e00",
    21780 => x"46656200", 21781 => x"4d617200", 21782 => x"41707200",
    21783 => x"4d617900", 21784 => x"4a756e00", 21785 => x"4a756c00",
    21786 => x"41756700", 21787 => x"53657000", 21788 => x"4f637400",
    21789 => x"4e6f7600", 21790 => x"44656300", 21791 => x"4c6f6f70",
    21792 => x"73207065", 21793 => x"72206a69", 21794 => x"6666793a",
    21795 => x"2025690a", 21796 => x"00000000", 21797 => x"25733a20",
    21798 => x"6e6f2073", 21799 => x"6f636b65", 21800 => x"7420736c",
    21801 => x"6f747320", 21802 => x"6c656674", 21803 => x"0a000000",
    21804 => x"77723000", 21805 => x"6e65742d", 21806 => x"62680000",
    21807 => x"69707634", 21808 => x"00000000", 21809 => x"61727000",
    21810 => x"44697363", 21811 => x"6f766572", 21812 => x"65642049",
    21813 => x"50206164", 21814 => x"64726573", 21815 => x"73202825",
    21816 => x"642e2564", 21817 => x"2e25642e", 21818 => x"25642921",
    21819 => x"0a000000", 21820 => x"534e4d50", 21821 => x"3a205346",
    21822 => x"50207570", 21823 => x"64617465", 21824 => x"6420696e",
    21825 => x"206d656d", 21826 => x"6f72792c", 21827 => x"20726573",
    21828 => x"74617274", 21829 => x"20505450", 21830 => x"0a000000",
    21831 => x"494e5641", 21832 => x"4c494400", 21833 => x"25642e25",
    21834 => x"30346400", 21835 => x"736e6d70", 21836 => x"00000000",
    21837 => x"53657020", 21838 => x"32302032", 21839 => x"30313620",
    21840 => x"31373a33", 21841 => x"303a3136", 21842 => x"00000000",
    21843 => x"30313233", 21844 => x"34353637", 21845 => x"38396162",
    21846 => x"63646566", 21847 => x"00000000", 21848 => x"49443a20",
    21849 => x"25780a00", 21850 => x"6e6f2070", 21851 => x"66696c74",
    21852 => x"65722072", 21853 => x"756c652d", 21854 => x"73657421",
    21855 => x"0a000000", 21856 => x"7066696c", 21857 => x"7465723a",
    21858 => x"2077726f", 21859 => x"6e67206d", 21860 => x"61676963",
    21861 => x"206e756d", 21862 => x"62657220", 21863 => x"28676f74",
    21864 => x"20307825", 21865 => x"78290a00", 21866 => x"7066696c",
    21867 => x"7465723a", 21868 => x"2077726f", 21869 => x"6e672072",
    21870 => x"756c652d", 21871 => x"7365742c", 21872 => x"2063616e",
    21873 => x"27742061", 21874 => x"70706c79", 21875 => x"0a000000",
    21876 => x"696e7661", 21877 => x"6c696420", 21878 => x"64657363",
    21879 => x"72697074", 21880 => x"6f722040", 21881 => x"2578203d",
    21882 => x"2025780a", 21883 => x"00000000", 21884 => x"5761726e",
    21885 => x"696e673a", 21886 => x"20747820", 21887 => x"6e6f7420",
    21888 => x"7465726d", 21889 => x"696e6174", 21890 => x"65642069",
    21891 => x"6e66696e", 21892 => x"69746520", 21893 => x"6d63723d",
    21894 => x"30782578", 21895 => x"0a000000", 21896 => x"5761726e",
    21897 => x"696e673a", 21898 => x"20747820", 21899 => x"74696d65",
    21900 => x"7374616d", 21901 => x"70206e65", 21902 => x"76657220",
    21903 => x"62656361", 21904 => x"6d652061", 21905 => x"7661696c",
    21906 => x"61626c65", 21907 => x"0a000000", 21908 => x"64657620",
    21909 => x"20307825", 21910 => x"30386c78", 21911 => x"20402025",
    21912 => x"30366c78", 21913 => x"2c202573", 21914 => x"0a000000",
    21915 => x"66706761", 21916 => x"2d617265", 21917 => x"61000000",
    21918 => x"4572726f", 21919 => x"72202564", 21920 => x"20776869",
    21921 => x"6c652072", 21922 => x"65616469", 21923 => x"6e672074",
    21924 => x"32347020", 21925 => x"66726f6d", 21926 => x"2073746f",
    21927 => x"72616765", 21928 => x"0a000000", 21929 => x"74323470",
    21930 => x"20726561", 21931 => x"64206672", 21932 => x"6f6d2073",
    21933 => x"746f7261", 21934 => x"67653a20", 21935 => x"25642070",
    21936 => x"730a0000", 21937 => x"57616974", 21938 => x"696e6720",
    21939 => x"666f7220", 21940 => x"6c696e6b", 21941 => x"2e2e2e0a",
    21942 => x"00000000", 21943 => x"4c6f636b", 21944 => x"696e6720",
    21945 => x"504c4c2e", 21946 => x"2e2e0a00", 21947 => x"43616c69",
    21948 => x"62726174", 21949 => x"696e6720", 21950 => x"52582074",
    21951 => x"696d6573", 21952 => x"74616d70", 21953 => x"65722e2e",
    21954 => x"2e0a0000", 21955 => x"4661696c", 21956 => x"65640000",
    21957 => x"53756363", 21958 => x"65737300", 21959 => x"57726f74",
    21960 => x"65206e65", 21961 => x"77207432", 21962 => x"34702076",
    21963 => x"616c7565", 21964 => x"3a202564", 21965 => x"20707320",
    21966 => x"28257329", 21967 => x"0a000000", 21968 => x"20454e4f",
    21969 => x"53504300", 21970 => x"25732573", 21971 => x"3a000000",
    21972 => x"74656d70", 21973 => x"00000000", 21974 => x"74656d70",
    21975 => x"65726174", 21976 => x"75726500", 21977 => x"55706461",
    21978 => x"74652065", 21979 => x"78697374", 21980 => x"696e6720",
    21981 => x"53465020", 21982 => x"656e7472", 21983 => x"790a0000",
    21984 => x"41646469", 21985 => x"6e67206e", 21986 => x"65772053",
    21987 => x"46502065", 21988 => x"6e747279", 21989 => x"0a000000",
    21990 => x"43616e27", 21991 => x"74207361", 21992 => x"76652070",
    21993 => x"65727369", 21994 => x"7374656e", 21995 => x"74204d41",
    21996 => x"43206164", 21997 => x"64726573", 21998 => x"730a0000",
    21999 => x"25733a20", 22000 => x"5573696e", 22001 => x"67205731",
    22002 => x"20736572", 22003 => x"69616c20", 22004 => x"6e756d62",
    22005 => x"65720a00", 22006 => x"6f666673", 22007 => x"65742025",
    22008 => x"34692028", 22009 => x"30782530", 22010 => x"3378293a",
    22011 => x"20253369", 22012 => x"20283078", 22013 => x"25303278",
    22014 => x"290a0000", 22015 => x"77726974", 22016 => x"65283078",
    22017 => x"25782c20", 22018 => x"2569293a", 22019 => x"20726573",
    22020 => x"756c7420", 22021 => x"3d202569", 22022 => x"0a000000",
    22023 => x"72656164", 22024 => x"28307825", 22025 => x"782c2025",
    22026 => x"69293a20", 22027 => x"72657375", 22028 => x"6c74203d",
    22029 => x"2025690a", 22030 => x"00000000", 22031 => x"64657669",
    22032 => x"63652025", 22033 => x"693a2025", 22034 => x"30387825",
    22035 => x"3038780a", 22036 => x"00000000", 22037 => x"74656d70",
    22038 => x"3a202564", 22039 => x"2e253034", 22040 => x"640a0000",
    22041 => x"77310000", 22042 => x"77317200", 22043 => x"77317700",
    22044 => x"3c756e6b", 22045 => x"6e6f776e", 22046 => x"3e000000",
    22047 => x"736f6674", 22048 => x"706c6c3a", 22049 => x"20697271",
    22050 => x"73202564", 22051 => x"20736571", 22052 => x"20257320",
    22053 => x"6d6f6465", 22054 => x"20256420", 22055 => x"616c6967",
    22056 => x"6e6d656e", 22057 => x"745f7374", 22058 => x"61746520",
    22059 => x"25642048", 22060 => x"4c256420", 22061 => x"4d4c2564",
    22062 => x"2048593d", 22063 => x"2564204d", 22064 => x"593d2564",
    22065 => x"2044656c", 22066 => x"436e743d", 22067 => x"25640a00",
    22068 => x"73746172", 22069 => x"742d6578", 22070 => x"74000000",
    22071 => x"77616974", 22072 => x"2d657874", 22073 => x"00000000",
    22074 => x"73746172", 22075 => x"742d6865", 22076 => x"6c706572",
    22077 => x"00000000", 22078 => x"77616974", 22079 => x"2d68656c",
    22080 => x"70657200", 22081 => x"73746172", 22082 => x"742d6d61",
    22083 => x"696e0000", 22084 => x"77616974", 22085 => x"2d6d6169",
    22086 => x"6e000000", 22087 => x"72656164", 22088 => x"79000000",
    22089 => x"636c6561", 22090 => x"722d6461", 22091 => x"63730000",
    22092 => x"77616974", 22093 => x"2d636c65", 22094 => x"61722d64",
    22095 => x"61637300", 22096 => x"53746163", 22097 => x"6b206f76",
    22098 => x"6572666c", 22099 => x"6f77210a", 22100 => x"00000000",
    22101 => x"badc0ffe", 22102 => x"3b9aca00", 22103 => x"000f4240",
    22104 => x"00080030", 22105 => x"d4a51000", 22106 => x"3b9ac9ff",
    22107 => x"c4653600", 22108 => x"7ffffffe", 22109 => x"80000001",
    22110 => x"fff06000", 22111 => x"0007d000", 22112 => x"41c64e6d",
    22113 => x"00010043", 22114 => x"00010044", 22115 => x"00015180",
    22116 => x"83aa7e80", 22117 => x"7fffffff", 22118 => x"00062000",
    22119 => x"005ee000", 22120 => x"01000001", 22121 => x"11223344",
    22122 => x"e0001fff", 22123 => x"111ee000", 22124 => x"01554000",
    22125 => x"0fffffff", 22126 => x"059682f0", 22127 => x"0ee6b27f",
    22128 => x"0003ffff", 22129 => x"c0a80001", 22130 => x"4b002f40",
    22131 => x"01312d02", 22132 => x"01312d0a", 22133 => x"003d0137",
    22134 => x"8000001f", 22135 => x"009895b6", 22136 => x"c4000001",
    22137 => x"000186a0", 22138 => x"00ffffff", 22139 => x"fffdb610",
    22140 => x"000249f0", 22141 => x"05f5e100", 22142 => x"0bebc200",
    22143 => x"fa0a1f00", 22144 => x"01312d03", 22145 => x"5344422d",
    22146 => x"011b1900", 22147 => x"00000000", 22148 => x"70705f64",
    22149 => x"6961675f", 22150 => x"70617273", 22151 => x"65000000",
    22152 => x"00000000", 22153 => x"00013830", 22154 => x"0001383c",
    22155 => x"0001384c", 22156 => x"00013858", 22157 => x"00013864",
    22158 => x"00013870", 22159 => x"0001387c", 22160 => x"0000150c",
    22161 => x"0000157c", 22162 => x"00001834", 22163 => x"00001834",
    22164 => x"00001834", 22165 => x"00001834", 22166 => x"00001834",
    22167 => x"00001834", 22168 => x"000015f8", 22169 => x"00001668",
    22170 => x"00001834", 22171 => x"000016fc", 22172 => x"00001808",
    22173 => x"77727063", 22174 => x"5f74696d", 22175 => x"655f6164",
    22176 => x"6a757374", 22177 => x"5f6f6666", 22178 => x"73657400",
    22179 => x"77725f73", 22180 => x"31000000", 22181 => x"77727063",
    22182 => x"5f74696d", 22183 => x"655f6164", 22184 => x"6a757374",
    22185 => x"00000000", 22186 => x"77727063", 22187 => x"5f74696d",
    22188 => x"655f7365", 22189 => x"74000000", 22190 => x"77727063",
    22191 => x"5f74696d", 22192 => x"655f6765", 22193 => x"74000000",
    22194 => x"77727063", 22195 => x"5f6e6574", 22196 => x"5f73656e",
    22197 => x"64000000", 22198 => x"77725f75", 22199 => x"6e706163",
    22200 => x"6b5f616e", 22201 => x"6e6f756e", 22202 => x"63650000",
    22203 => x"77725f73", 22204 => x"6572766f", 22205 => x"5f757064",
    22206 => x"61746500", 22207 => x"77725f70", 22208 => x"61636b5f",
    22209 => x"616e6e6f", 22210 => x"756e6365", 22211 => x"00000000",
    22212 => x"77725f68", 22213 => x"616e646c", 22214 => x"655f666f",
    22215 => x"6c6c6f77", 22216 => x"75700000", 22217 => x"77725f68",
    22218 => x"616e646c", 22219 => x"655f616e", 22220 => x"6e6f756e",
    22221 => x"63650000", 22222 => x"77725f65", 22223 => x"78656375",
    22224 => x"74655f73", 22225 => x"6c617665", 22226 => x"00000000",
    22227 => x"77725f68", 22228 => x"616e646c", 22229 => x"655f7265",
    22230 => x"73700000", 22231 => x"77725f6e", 22232 => x"65775f73",
    22233 => x"6c617665", 22234 => x"00000000", 22235 => x"77725f6d",
    22236 => x"61737465", 22237 => x"725f6d73", 22238 => x"67000000",
    22239 => x"77725f6c", 22240 => x"69737465", 22241 => x"6e696e67",
    22242 => x"00000000", 22243 => x"77725f6f", 22244 => x"70656e00",
    22245 => x"77725f69", 22246 => x"6e697400", 22247 => x"00002e0c",
    22248 => x"00002e34", 22249 => x"00002e54", 22250 => x"00002ec4",
    22251 => x"00002ee4", 22252 => x"00002f00", 22253 => x"00002f20",
    22254 => x"00002fac", 22255 => x"00002fcc", 22256 => x"77725f63",
    22257 => x"616c6962", 22258 => x"72617469", 22259 => x"6f6e0000",
    22260 => x"00004450", 22261 => x"00004438", 22262 => x"00004478",
    22263 => x"00004584", 22264 => x"000044cc", 22265 => x"00014198",
    22266 => x"000142cc", 22267 => x"000142d8", 22268 => x"000142e4",
    22269 => x"000142f0", 22270 => x"000142fc", 22271 => x"70705f69",
    22272 => x"6e697469", 22273 => x"616c697a", 22274 => x"696e6700",
    22275 => x"73745f63", 22276 => x"6f6d5f73", 22277 => x"6c617665",
    22278 => x"5f68616e", 22279 => x"646c655f", 22280 => x"666f6c6c",
    22281 => x"6f777570", 22282 => x"00000000", 22283 => x"626d635f",
    22284 => x"64617461", 22285 => x"7365745f", 22286 => x"636d7000",
    22287 => x"626d635f", 22288 => x"73746174", 22289 => x"655f6465",
    22290 => x"63697369", 22291 => x"6f6e0000", 22292 => x"63466965",
    22293 => x"6c645f74", 22294 => x"6f5f5469", 22295 => x"6d65496e",
    22296 => x"7465726e", 22297 => x"616c0000", 22298 => x"00014e28",
    22299 => x"00014f68", 22300 => x"00014314", 22301 => x"00013e2c",
    22302 => x"0000001f", 22303 => x"0000001c", 22304 => x"0000001f",
    22305 => x"0000001e", 22306 => x"0000001f", 22307 => x"0000001e",
    22308 => x"0000001f", 22309 => x"0000001f", 22310 => x"0000001e",
    22311 => x"0000001f", 22312 => x"0000001e", 22313 => x"0000001f",
    22314 => x"0000001f", 22315 => x"0000001d", 22316 => x"0000001f",
    22317 => x"0000001e", 22318 => x"0000001f", 22319 => x"0000001e",
    22320 => x"0000001f", 22321 => x"0000001f", 22322 => x"0000001e",
    22323 => x"0000001f", 22324 => x"0000001e", 22325 => x"0000001f",
    22326 => x"00015430", 22327 => x"00015434", 22328 => x"00015438",
    22329 => x"0001543c", 22330 => x"00015440", 22331 => x"00015444",
    22332 => x"00015448", 22333 => x"0001544c", 22334 => x"00015450",
    22335 => x"00015454", 22336 => x"00015458", 22337 => x"0001545c",
    22338 => x"00015460", 22339 => x"00015464", 22340 => x"00015468",
    22341 => x"0001546c", 22342 => x"00015470", 22343 => x"00015474",
    22344 => x"00015478", 22345 => x"70747064", 22346 => x"5f6e6574",
    22347 => x"69665f63", 22348 => x"72656174", 22349 => x"655f736f",
    22350 => x"636b6574", 22351 => x"00000000", 22352 => x"0000b6f8",
    22353 => x"0000b708", 22354 => x"0000b76c", 22355 => x"0000b76c",
    22356 => x"0000b718", 22357 => x"0000b76c", 22358 => x"0000b76c",
    22359 => x"30ff0201", 22360 => x"fa040670", 22361 => x"75626c69",
    22362 => x"63fdff02", 22363 => x"f90201fc", 22364 => x"0201fb30",
    22365 => x"ff30ff06", 22366 => x"6765745f", 22367 => x"70657273",
    22368 => x"69737465", 22369 => x"6e745f6d", 22370 => x"61630000",
    22371 => x"000000c8", 22372 => x"000039d0", 22373 => x"00010d30",
    22374 => x"00010db4", 22375 => x"00010dec", 22376 => x"00010e6c",
    22377 => x"00010ef8", 22378 => x"00010f10", 22379 => x"00010e10",
    22380 => x"00010d58", 22381 => x"00010cb4", 22382 => x"00010ce8",
    22383 => x"00000000", 22384 => x"00000000", 22385 => x"00000000",
    22386 => x"00000000", 22387 => x"00000001", 22388 => x"00000001",
    22389 => x"00000001", 22390 => x"00000001", 22391 => x"00000000",
    22392 => x"00000000", 22393 => x"00000000", 22394 => x"0000ece8",
    22395 => x"0000ece8", 22396 => x"00000000", 22397 => x"0000d9d0",
    22398 => x"00000000", 22399 => x"00011a74", 22400 => x"00011a94",
    22401 => x"00011aa0", 22402 => x"00011ab0", 22403 => x"00011ad0",
    22404 => x"00011ae0", 22405 => x"00011b34", 22406 => x"00011af8",
    22407 => x"00011a08", 22408 => x"00011a4c", 22409 => x"00000001",
    22410 => x"000158d0", 22411 => x"00000002", 22412 => x"000158dc",
    22413 => x"00000003", 22414 => x"000158e8", 22415 => x"00000004",
    22416 => x"000158f8", 22417 => x"00000005", 22418 => x"00015904",
    22419 => x"00000006", 22420 => x"00015910", 22421 => x"00000007",
    22422 => x"00013e04", 22423 => x"00000008", 22424 => x"0001591c",
    22425 => x"00000009", 22426 => x"00015924", 22427 => x"0000000a",
    22428 => x"00015930", 22429 => x"00000000", 22430 => x"00000000",
    22431 => x"00000000", 22432 => x"00000000", 22433 => x"00000000",
    22434 => x"00000000", 22435 => x"00010000", 22436 => x"00000000",
    22437 => x"00000000", 22438 => x"00000000", 22439 => x"00020100",
    22440 => x"00000000", 22441 => x"00000000", 22442 => x"00000000",
    22443 => x"00030101", 22444 => x"00000000", 22445 => x"00000000",
    22446 => x"00000000", 22447 => x"00040201", 22448 => x"01000000",
    22449 => x"00000000", 22450 => x"00000000", 22451 => x"00050201",
    22452 => x"01010000", 22453 => x"00000000", 22454 => x"00000000",
    22455 => x"00060302", 22456 => x"01010100", 22457 => x"00000000",
    22458 => x"00000000", 22459 => x"00070302", 22460 => x"01010101",
    22461 => x"00000000", 22462 => x"00000000", 22463 => x"00080402",
    22464 => x"02010101", 22465 => x"01000000", 22466 => x"00000000",
    22467 => x"00090403", 22468 => x"02010101", 22469 => x"01010000",
    22470 => x"00000000", 22471 => x"000a0503", 22472 => x"02020101",
    22473 => x"01010100", 22474 => x"00000000", 22475 => x"000b0503",
    22476 => x"02020101", 22477 => x"01010101", 22478 => x"00000000",
    22479 => x"000c0604", 22480 => x"03020201", 22481 => x"01010101",
    22482 => x"01000000", 22483 => x"000d0604", 22484 => x"03020201",
    22485 => x"01010101", 22486 => x"01010000", 22487 => x"000e0704",
    22488 => x"03020202", 22489 => x"01010101", 22490 => x"01010100",
    22491 => x"000f0705", 22492 => x"03030202", 22493 => x"01010101",
    22494 => x"01010101", 22495 => x"fefefeff", 22496 => x"80808080",
    22497 => x"00202020", 22498 => x"20202020", 22499 => x"20202828",
    22500 => x"28282820", 22501 => x"20202020", 22502 => x"20202020",
    22503 => x"20202020", 22504 => x"20202020", 22505 => x"20881010",
    22506 => x"10101010", 22507 => x"10101010", 22508 => x"10101010",
    22509 => x"10040404", 22510 => x"04040404", 22511 => x"04040410",
    22512 => x"10101010", 22513 => x"10104141", 22514 => x"41414141",
    22515 => x"01010101", 22516 => x"01010101", 22517 => x"01010101",
    22518 => x"01010101", 22519 => x"01010101", 22520 => x"10101010",
    22521 => x"10104242", 22522 => x"42424242", 22523 => x"02020202",
    22524 => x"02020202", 22525 => x"02020202", 22526 => x"02020202",
    22527 => x"02020202", 22528 => x"10101010", 22529 => x"20000000",
    22530 => x"00000000", 22531 => x"00000000", 22532 => x"00000000",
    22533 => x"00000000", 22534 => x"00000000", 22535 => x"00000000",
    22536 => x"00000000", 22537 => x"00000000", 22538 => x"00000000",
    22539 => x"00000000", 22540 => x"00000000", 22541 => x"00000000",
    22542 => x"00000000", 22543 => x"00000000", 22544 => x"00000000",
    22545 => x"00000000", 22546 => x"00000000", 22547 => x"00000000",
    22548 => x"00000000", 22549 => x"00000000", 22550 => x"00000000",
    22551 => x"00000000", 22552 => x"00000000", 22553 => x"00000000",
    22554 => x"00000000", 22555 => x"00000000", 22556 => x"00000000",
    22557 => x"00000000", 22558 => x"00000000", 22559 => x"00000000",
    22560 => x"00000000", 22561 => x"00000000", 22562 => x"00017238",
    22563 => x"00017258", 22564 => x"00017268", 22565 => x"00017278",
    22566 => x"000003e8", 22567 => x"00000001", 22568 => x"00000955",
    22569 => x"ffffffff", 22570 => x"00000000", 22571 => x"00000000",
    22572 => x"00000000", 22573 => x"00000000", 22574 => x"00000000",
    22575 => x"00000000", 22576 => x"00000000", 22577 => x"00000000",
    22578 => x"0001641c", 22579 => x"0001653c", 22580 => x"00016520",
    22581 => x"00017558", 22582 => x"000175d8", 22583 => x"00000000",
    22584 => x"00000000", 22585 => x"00000000", 22586 => x"00000000",
    22587 => x"00000000", 22588 => x"00000000", 22589 => x"00000000",
    22590 => x"00000000", 22591 => x"00000000", 22592 => x"00000000",
    22593 => x"00000000", 22594 => x"00000000", 22595 => x"00000000",
    22596 => x"00000000", 22597 => x"00000000", 22598 => x"00000000",
    22599 => x"00000000", 22600 => x"00000000", 22601 => x"00000000",
    22602 => x"00000000", 22603 => x"00000000", 22604 => x"00000000",
    22605 => x"00000000", 22606 => x"00000000", 22607 => x"00000000",
    22608 => x"00000000", 22609 => x"00000000", 22610 => x"00000000",
    22611 => x"00000000", 22612 => x"00000000", 22613 => x"00000000",
    22614 => x"00000000", 22615 => x"00000000", 22616 => x"00000000",
    22617 => x"00000000", 22618 => x"00000000", 22619 => x"00000000",
    22620 => x"00000000", 22621 => x"00000000", 22622 => x"00000000",
    22623 => x"00000000", 22624 => x"00000000", 22625 => x"00000000",
    22626 => x"00000000", 22627 => x"00000000", 22628 => x"00000000",
    22629 => x"00000000", 22630 => x"00000000", 22631 => x"00000000",
    22632 => x"00000000", 22633 => x"00000000", 22634 => x"00000000",
    22635 => x"00000000", 22636 => x"00000000", 22637 => x"00000000",
    22638 => x"00000000", 22639 => x"00000000", 22640 => x"00000000",
    22641 => x"00000000", 22642 => x"00000000", 22643 => x"00000000",
    22644 => x"00000000", 22645 => x"00000000", 22646 => x"00000000",
    22647 => x"00000000", 22648 => x"00000000", 22649 => x"00000000",
    22650 => x"00000000", 22651 => x"00000000", 22652 => x"00000000",
    22653 => x"00000000", 22654 => x"00000000", 22655 => x"00000000",
    22656 => x"00000000", 22657 => x"00000000", 22658 => x"00000000",
    22659 => x"00000000", 22660 => x"00000000", 22661 => x"00000000",
    22662 => x"00000000", 22663 => x"00000000", 22664 => x"00000000",
    22665 => x"00000000", 22666 => x"00000000", 22667 => x"00000000",
    22668 => x"00000000", 22669 => x"00000000", 22670 => x"00000000",
    22671 => x"00000000", 22672 => x"00000000", 22673 => x"00000000",
    22674 => x"00000000", 22675 => x"00000000", 22676 => x"00000000",
    22677 => x"00000000", 22678 => x"00000000", 22679 => x"00000000",
    22680 => x"00000000", 22681 => x"00000000", 22682 => x"00000000",
    22683 => x"00000000", 22684 => x"00000000", 22685 => x"00000000",
    22686 => x"00000000", 22687 => x"00000000", 22688 => x"00000000",
    22689 => x"00000000", 22690 => x"00000000", 22691 => x"00000000",
    22692 => x"00000000", 22693 => x"00000000", 22694 => x"00000000",
    22695 => x"00000000", 22696 => x"00000000", 22697 => x"00000000",
    22698 => x"00000000", 22699 => x"00000000", 22700 => x"00000000",
    22701 => x"00000000", 22702 => x"00000000", 22703 => x"00000000",
    22704 => x"00000000", 22705 => x"00000000", 22706 => x"00000000",
    22707 => x"00000000", 22708 => x"00000000", 22709 => x"00000000",
    22710 => x"00000000", 22711 => x"00000000", 22712 => x"00000000",
    22713 => x"00000000", 22714 => x"00000000", 22715 => x"00000000",
    22716 => x"00000000", 22717 => x"00000000", 22718 => x"00000000",
    22719 => x"00000000", 22720 => x"00000000", 22721 => x"00000000",
    22722 => x"00000000", 22723 => x"00000000", 22724 => x"00000000",
    22725 => x"00000000", 22726 => x"00000000", 22727 => x"00000000",
    22728 => x"00000000", 22729 => x"00000000", 22730 => x"00000000",
    22731 => x"00000000", 22732 => x"00000000", 22733 => x"00000000",
    22734 => x"00000000", 22735 => x"00000000", 22736 => x"00000000",
    22737 => x"00000000", 22738 => x"00000000", 22739 => x"00000000",
    22740 => x"00000000", 22741 => x"00000000", 22742 => x"00000000",
    22743 => x"00000000", 22744 => x"00000000", 22745 => x"00000000",
    22746 => x"00000000", 22747 => x"00000000", 22748 => x"00016464",
    22749 => x"00000000", 22750 => x"00000000", 22751 => x"00000000",
    22752 => x"00000000", 22753 => x"00000000", 22754 => x"00000000",
    22755 => x"00000000", 22756 => x"00000000", 22757 => x"00000000",
    22758 => x"00000000", 22759 => x"00000000", 22760 => x"00000000",
    22761 => x"00000000", 22762 => x"00000000", 22763 => x"00000000",
    22764 => x"00000000", 22765 => x"00000000", 22766 => x"00000000",
    22767 => x"00000000", 22768 => x"00000000", 22769 => x"00000000",
    22770 => x"00000000", 22771 => x"00000000", 22772 => x"00000000",
    22773 => x"00000000", 22774 => x"0001390c", 22775 => x"0001390c",
    22776 => x"00000000", 22777 => x"00000001", 22778 => x"00000000",
    22779 => x"00000000", 22780 => x"00000000", 22781 => x"00000000",
    22782 => x"00000000", 22783 => x"00000000", 22784 => x"00000000",
    22785 => x"00000000", 22786 => x"00000000", 22787 => x"00000000",
    22788 => x"00000000", 22789 => x"00000000", 22790 => x"00000000",
    22791 => x"000160a8", 22792 => x"00017658", 22793 => x"00000000",
    22794 => x"00017698", 22795 => x"000176b4", 22796 => x"000176e4",
    22797 => x"00017704", 22798 => x"00000000", 22799 => x"00000000",
    22800 => x"00000000", 22801 => x"00000000", 22802 => x"00000000",
    22803 => x"00000000", 22804 => x"00000000", 22805 => x"00000000",
    22806 => x"00000000", 22807 => x"00017728", 22808 => x"000003e8",
    22809 => x"00000000", 22810 => x"00000000", 22811 => x"00000000",
    22812 => x"00000000", 22813 => x"00016478", 22814 => x"000164e4",
    22815 => x"00000000", 22816 => x"00000000", 22817 => x"00000000",
    22818 => x"00000000", 22819 => x"00000000", 22820 => x"00000000",
    22821 => x"00000000", 22822 => x"00000000", 22823 => x"00000000",
    22824 => x"00000000", 22825 => x"00000000", 22826 => x"00000000",
    22827 => x"00000000", 22828 => x"00000000", 22829 => x"00000000",
    22830 => x"00000000", 22831 => x"00000000", 22832 => x"00000000",
    22833 => x"00000000", 22834 => x"00000000", 22835 => x"00000000",
    22836 => x"00000000", 22837 => x"00000000", 22838 => x"00000000",
    22839 => x"00000000", 22840 => x"00000000", 22841 => x"00000a88",
    22842 => x"00000abc", 22843 => x"00000b3c", 22844 => x"00000b44",
    22845 => x"00000b9c", 22846 => x"00000bc8", 22847 => x"00000c20",
    22848 => x"00000c44", 22849 => x"00000d08", 22850 => x"00000d10",
    22851 => x"00000d18", 22852 => x"00000d7c", 22853 => x"00000d98",
    22854 => x"00000b68", 22855 => x"00000000", 22856 => x"00001cbc",
    22857 => x"00001c40", 22858 => x"00001be4", 22859 => x"00001b8c",
    22860 => x"00000000", 22861 => x"00000000", 22862 => x"00001b5c",
    22863 => x"00001f48", 22864 => x"00001f28", 22865 => x"00001e58",
    22866 => x"00001d3c", 22867 => x"00000000", 22868 => x"00000000",
    22869 => x"00000000", 22870 => x"00000000", 22871 => x"00000000",
    22872 => x"00000000", 22873 => x"00000000", 22874 => x"00000000",
    22875 => x"00000000", 22876 => x"00000000", 22877 => x"00000000",
    22878 => x"00000200", 22879 => x"00000000", 22880 => x"00017838",
    22881 => x"00000001", 22882 => x"00013dec", 22883 => x"00004778",
    22884 => x"00000002", 22885 => x"00013dfc", 22886 => x"00004944",
    22887 => x"00000003", 22888 => x"00013e04", 22889 => x"00004a00",
    22890 => x"00000004", 22891 => x"00013e10", 22892 => x"00004a10",
    22893 => x"00000006", 22894 => x"00014314", 22895 => x"00004bbc",
    22896 => x"00000008", 22897 => x"00013e1c", 22898 => x"00004efc",
    22899 => x"00000009", 22900 => x"00013e2c", 22901 => x"00004f70",
    22902 => x"00000064", 22903 => x"00013e34", 22904 => x"00002844",
    22905 => x"00000066", 22906 => x"00013e4c", 22907 => x"000029bc",
    22908 => x"00000065", 22909 => x"00013e60", 22910 => x"00002ae8",
    22911 => x"00000067", 22912 => x"00013e78", 22913 => x"00002bec",
    22914 => x"00000068", 22915 => x"00013e90", 22916 => x"00002d18",
    22917 => x"00000069", 22918 => x"00013ea0", 22919 => x"00003034",
    22920 => x"0000006a", 22921 => x"00013eb0", 22922 => x"00003148",
    22923 => x"0000006b", 22924 => x"00013ec4", 22925 => x"000032cc",
    22926 => x"00000000", 22927 => x"00000000", 22928 => x"00000000",
    22929 => x"00000001", 22930 => x"00013dec", 22931 => x"00004778",
    22932 => x"00000002", 22933 => x"00013dfc", 22934 => x"00004944",
    22935 => x"00000003", 22936 => x"00013e04", 22937 => x"00004a00",
    22938 => x"00000004", 22939 => x"00013e10", 22940 => x"00004a10",
    22941 => x"00000005", 22942 => x"00014310", 22943 => x"00004b28",
    22944 => x"00000006", 22945 => x"00014314", 22946 => x"00004bbc",
    22947 => x"00000007", 22948 => x"0001431c", 22949 => x"00004e38",
    22950 => x"00000008", 22951 => x"00013e1c", 22952 => x"00004efc",
    22953 => x"00000009", 22954 => x"00013e2c", 22955 => x"00004f70",
    22956 => x"00000000", 22957 => x"00000000", 22958 => x"00000000",
    22959 => x"00002248", 22960 => x"00002168", 22961 => x"00000000",
    22962 => x"00002120", 22963 => x"000025e0", 22964 => x"00002598",
    22965 => x"000024ac", 22966 => x"00002090", 22967 => x"00002004",
    22968 => x"00002434", 22969 => x"000023bc", 22970 => x"00002354",
    22971 => x"000022e8", 22972 => x"00000001", 22973 => x"00014528",
    22974 => x"00014530", 22975 => x"0001453c", 22976 => x"00014548",
    22977 => x"00000000", 22978 => x"00000000", 22979 => x"00000000",
    22980 => x"00000000", 22981 => x"0001456c", 22982 => x"00014554",
    22983 => x"00014560", 22984 => x"00014578", 22985 => x"00014584",
    22986 => x"00014590", 22987 => x"00000000", 22988 => x"00000000",
    22989 => x"000148b8", 22990 => x"000148c8", 22991 => x"000148d4",
    22992 => x"000148e8", 22993 => x"000148fc", 22994 => x"0001490c",
    22995 => x"00014918", 22996 => x"00014924", 22997 => x"bbfef060",
    22998 => x"00000000", 22999 => x"00000000", 23000 => x"00000000",
    23001 => x"00000000", 23002 => x"00000000", 23003 => x"00000000",
    23004 => x"00000000", 23005 => x"00000000", 23006 => x"00000000",
    23007 => x"00000000", 23008 => x"00000000", 23009 => x"00000000",
    23010 => x"00000001", 23011 => x"00000000", 23012 => x"000a03e8",
    23013 => x"00060100", 23014 => x"80800000", 23015 => x"00000000",
    23016 => x"000160a8", 23017 => x"00000000", 23018 => x"00000000",
    23019 => x"00000000", 23020 => x"00000000", 23021 => x"00000000",
    23022 => x"00000000", 23023 => x"00000000", 23024 => x"00000000",
    23025 => x"00000000", 23026 => x"00000000", 23027 => x"00000200",
    23028 => x"00000000", 23029 => x"00017d64", 23030 => x"00000000",
    23031 => x"00000000", 23032 => x"00000000", 23033 => x"00000000",
    23034 => x"00000000", 23035 => x"00000000", 23036 => x"00000000",
    23037 => x"00000000", 23038 => x"00000000", 23039 => x"00000000",
    23040 => x"00000060", 23041 => x"00000000", 23042 => x"00017f64",
    23043 => x"00000000", 23044 => x"00000000", 23045 => x"00000000",
    23046 => x"00000000", 23047 => x"00000000", 23048 => x"00000000",
    23049 => x"00000000", 23050 => x"00000000", 23051 => x"00000000",
    23052 => x"00000000", 23053 => x"00000080", 23054 => x"00000000",
    23055 => x"00017fc4", 23056 => x"00000000", 23057 => x"00000000",
    23058 => x"00000000", 23059 => x"00000000", 23060 => x"00000000",
    23061 => x"00000000", 23062 => x"00000000", 23063 => x"00000000",
    23064 => x"00000000", 23065 => x"00000000", 23066 => x"00000080",
    23067 => x"00000000", 23068 => x"00018048", 23069 => x"63757465",
    23070 => x"70636e00", 23071 => x"00000000", 23072 => x"00000000",
    23073 => x"00000000", 23074 => x"00000000", 23075 => x"00000000",
    23076 => x"00000000", 23077 => x"00016958", 23078 => x"0000bc48",
    23079 => x"00016964", 23080 => x"09000000", 23081 => x"000169c8",
    23082 => x"0000bc48", 23083 => x"000169d4", 23084 => x"09000000",
    23085 => x"00016a24", 23086 => x"0000ba38", 23087 => x"00016a30",
    23088 => x"0a000000", 23089 => x"00016a6c", 23090 => x"0000bc48",
    23091 => x"00016a78", 23092 => x"09000000", 23093 => x"00016b40",
    23094 => x"0000bc48", 23095 => x"00016b4c", 23096 => x"09000000",
    23097 => x"00016cb4", 23098 => x"0000bc48", 23099 => x"00016cc0",
    23100 => x"09000000", 23101 => x"00016d4c", 23102 => x"0000bc48",
    23103 => x"00016d58", 23104 => x"09000000", 23105 => x"00016dd0",
    23106 => x"0000ba38", 23107 => x"00016ddc", 23108 => x"0a000000",
    23109 => x"00000000", 23110 => x"00000000", 23111 => x"00000000",
    23112 => x"00000000", 23113 => x"00000000", 23114 => x"00000000",
    23115 => x"00000000", 23116 => x"00000000", 23117 => x"00000000",
    23118 => x"00000000", 23119 => x"00000000", 23120 => x"00000000",
    23121 => x"00000000", 23122 => x"00000000", 23123 => x"00000100",
    23124 => x"00000000", 23125 => x"000180f0", 23126 => x"2b060104",
    23127 => x"01606501", 23128 => x"01000000", 23129 => x"00016e40",
    23130 => x"0000c1c4", 23131 => x"00000000", 23132 => x"00016874",
    23133 => x"02040020", 23134 => x"00016e44", 23135 => x"0000c198",
    23136 => x"00000000", 23137 => x"00016088", 23138 => x"02040004",
    23139 => x"00016e48", 23140 => x"0000c198", 23141 => x"00000000",
    23142 => x"00016094", 23143 => x"02040004", 23144 => x"00016e4c",
    23145 => x"0000c198", 23146 => x"00000000", 23147 => x"00016e50",
    23148 => x"02040004", 23149 => x"00000000", 23150 => x"00000000",
    23151 => x"00000000", 23152 => x"00000000", 23153 => x"00000000",
    23154 => x"2b060104", 23155 => x"01606501", 23156 => x"02000000",
    23157 => x"00016e54", 23158 => x"0000c55c", 23159 => x"00000000",
    23160 => x"00000004", 23161 => x"02460001", 23162 => x"00016e58",
    23163 => x"0000c55c", 23164 => x"00000000", 23165 => x"00000005",
    23166 => x"02040001", 23167 => x"00016e5c", 23168 => x"0000c55c",
    23169 => x"00000000", 23170 => x"00000002", 23171 => x"02430001",
    23172 => x"00000000", 23173 => x"00000000", 23174 => x"00000000",
    23175 => x"00000000", 23176 => x"00000000", 23177 => x"2b060104",
    23178 => x"01606501", 23179 => x"03010000", 23180 => x"00016e60",
    23181 => x"0000c42c", 23182 => x"00000000", 23183 => x"00000000",
    23184 => x"01040001", 23185 => x"00016e64", 23186 => x"0000c42c",
    23187 => x"00000000", 23188 => x"00000000", 23189 => x"01040001",
    23190 => x"00000000", 23191 => x"00000000", 23192 => x"00000000",
    23193 => x"00000000", 23194 => x"00000000", 23195 => x"2b060104",
    23196 => x"01606501", 23197 => x"04000000", 23198 => x"00016e68",
    23199 => x"0000c1c4", 23200 => x"00000000", 23201 => x"00017210",
    23202 => x"02020004", 23203 => x"00016e6c", 23204 => x"0000c1c4",
    23205 => x"00000000", 23206 => x"00017214", 23207 => x"02410004",
    23208 => x"00016e70", 23209 => x"0000c1c4", 23210 => x"00000000",
    23211 => x"00017218", 23212 => x"02020004", 23213 => x"00016e74",
    23214 => x"0000c1c4", 23215 => x"00000000", 23216 => x"0001721c",
    23217 => x"02020004", 23218 => x"00016e78", 23219 => x"0000c1c4",
    23220 => x"00000000", 23221 => x"00017220", 23222 => x"02410004",
    23223 => x"00016e7c", 23224 => x"0000c1c4", 23225 => x"00000000",
    23226 => x"00017224", 23227 => x"02410004", 23228 => x"00016e80",
    23229 => x"0000c1c4", 23230 => x"00000000", 23231 => x"00017228",
    23232 => x"02020004", 23233 => x"00016e84", 23234 => x"0000c1c4",
    23235 => x"00000000", 23236 => x"0001722c", 23237 => x"02020004",
    23238 => x"00016e88", 23239 => x"0000c1c4", 23240 => x"00000000",
    23241 => x"00017230", 23242 => x"02410004", 23243 => x"00000000",
    23244 => x"00000000", 23245 => x"00000000", 23246 => x"00000000",
    23247 => x"00000000", 23248 => x"2b060104", 23249 => x"01606501",
    23250 => x"05000000", 23251 => x"00016e8c", 23252 => x"0000c198",
    23253 => x"00000000", 23254 => x"000180cc", 23255 => x"02021404",
    23256 => x"00016e90", 23257 => x"0000c10c", 23258 => x"00000000",
    23259 => x"000180cc", 23260 => x"0202e808", 23261 => x"00016e94",
    23262 => x"0000c10c", 23263 => x"00000000", 23264 => x"000180cc",
    23265 => x"0202e008", 23266 => x"00016e98", 23267 => x"0000c198",
    23268 => x"00000000", 23269 => x"000180cc", 23270 => x"0246a008",
    23271 => x"00016e9c", 23272 => x"0000c198", 23273 => x"00000000",
    23274 => x"000180cc", 23275 => x"0241b804", 23276 => x"00016ea0",
    23277 => x"0000c00c", 23278 => x"00000000", 23279 => x"00000001",
    23280 => x"02460001", 23281 => x"00016ea4", 23282 => x"0000c198",
    23283 => x"00000000", 23284 => x"000180cc", 23285 => x"02021804",
    23286 => x"00016ea8", 23287 => x"0000c198", 23288 => x"00000000",
    23289 => x"000180cc", 23290 => x"02021c04", 23291 => x"00016eac",
    23292 => x"0000c198", 23293 => x"00000000", 23294 => x"000180cc",
    23295 => x"02022004", 23296 => x"00016eb0", 23297 => x"0000c198",
    23298 => x"00000000", 23299 => x"000180cc", 23300 => x"02022404",
    23301 => x"00016eb4", 23302 => x"0000c198", 23303 => x"00000000",
    23304 => x"000180cc", 23305 => x"0241f004", 23306 => x"00016eb8",
    23307 => x"0000c198", 23308 => x"00000000", 23309 => x"000180cc",
    23310 => x"0241f404", 23311 => x"00016ebc", 23312 => x"0000c198",
    23313 => x"00000000", 23314 => x"000180cc", 23315 => x"0241f804",
    23316 => x"00016ec0", 23317 => x"0000c00c", 23318 => x"00000000",
    23319 => x"00000002", 23320 => x"02460001", 23321 => x"00016ec4",
    23322 => x"0000c1c4", 23323 => x"00000000", 23324 => x"00016414",
    23325 => x"02410004", 23326 => x"00016ec8", 23327 => x"0000c1c4",
    23328 => x"00000000", 23329 => x"00016418", 23330 => x"02410004",
    23331 => x"00016ecc", 23332 => x"0000c198", 23333 => x"00000000",
    23334 => x"000180cc", 23335 => x"02022804", 23336 => x"00000000",
    23337 => x"00000000", 23338 => x"00000000", 23339 => x"00000000",
    23340 => x"00000000", 23341 => x"2b060104", 23342 => x"01606501",
    23343 => x"06000000", 23344 => x"00016ed0", 23345 => x"0000c1c4",
    23346 => x"0000c24c", 23347 => x"000181f0", 23348 => x"02020004",
    23349 => x"00016ed4", 23350 => x"0000c1c4", 23351 => x"0000c2ac",
    23352 => x"000181f4", 23353 => x"02020004", 23354 => x"00016ed8",
    23355 => x"0000c1c4", 23356 => x"0000ba14", 23357 => x"000180d0",
    23358 => x"02040010", 23359 => x"00016edc", 23360 => x"0000c1c4",
    23361 => x"0000ba14", 23362 => x"000180e4", 23363 => x"02020004",
    23364 => x"00016ee0", 23365 => x"0000c1c4", 23366 => x"0000ba14",
    23367 => x"000180e8", 23368 => x"02020004", 23369 => x"00016ee4",
    23370 => x"0000c1c4", 23371 => x"0000ba14", 23372 => x"000180e0",
    23373 => x"02020004", 23374 => x"00000000", 23375 => x"00000000",
    23376 => x"00000000", 23377 => x"00000000", 23378 => x"00000000",
    23379 => x"2b060104", 23380 => x"01606501", 23381 => x"07000000",
    23382 => x"00016ee8", 23383 => x"0000c1ec", 23384 => x"00000000",
    23385 => x"00000001", 23386 => x"02020001", 23387 => x"00016eec",
    23388 => x"0000c1c4", 23389 => x"00000000", 23390 => x"00018eec",
    23391 => x"02040010", 23392 => x"00016ef0", 23393 => x"0000c1c4",
    23394 => x"00000000", 23395 => x"00018e88", 23396 => x"02020004",
    23397 => x"00016ef4", 23398 => x"0000c1c4", 23399 => x"00000000",
    23400 => x"00019234", 23401 => x"02410004", 23402 => x"00016ef8",
    23403 => x"0000c1c4", 23404 => x"00000000", 23405 => x"00019238",
    23406 => x"02410004", 23407 => x"00000000", 23408 => x"00000000",
    23409 => x"00000000", 23410 => x"00000000", 23411 => x"00000000",
    23412 => x"2b060104", 23413 => x"01606501", 23414 => x"08010000",
    23415 => x"00016efc", 23416 => x"0000bedc", 23417 => x"00000000",
    23418 => x"00000000", 23419 => x"01040001", 23420 => x"00016f00",
    23421 => x"0000bedc", 23422 => x"00000000", 23423 => x"00000000",
    23424 => x"01020001", 23425 => x"00016f04", 23426 => x"0000bedc",
    23427 => x"00000000", 23428 => x"00000000", 23429 => x"01020001",
    23430 => x"00016f08", 23431 => x"0000bedc", 23432 => x"00000000",
    23433 => x"00000000", 23434 => x"01020001", 23435 => x"00000000",
    23436 => x"00000000", 23437 => x"00000000", 23438 => x"00000000",
    23439 => x"00000000", 23440 => x"01000000", 23441 => x"02000000",
    23442 => x"03000000", 23443 => x"04000000", 23444 => x"00015534",
    23445 => x"01000000", 23446 => x"02000000", 23447 => x"03000000",
    23448 => x"02000000", 23449 => x"03000000", 23450 => x"01000000",
    23451 => x"02000000", 23452 => x"03000000", 23453 => x"04000000",
    23454 => x"05000000", 23455 => x"06000000", 23456 => x"07000000",
    23457 => x"08000000", 23458 => x"09000000", 23459 => x"05000000",
    23460 => x"08000000", 23461 => x"09000000", 23462 => x"0a000000",
    23463 => x"0c000000", 23464 => x"0d000000", 23465 => x"0e000000",
    23466 => x"0f000000", 23467 => x"10000000", 23468 => x"11000000",
    23469 => x"12000000", 23470 => x"13000000", 23471 => x"14000000",
    23472 => x"16000000", 23473 => x"17000000", 23474 => x"18000000",
    23475 => x"1a000000", 23476 => x"01000000", 23477 => x"02000000",
    23478 => x"03000000", 23479 => x"04000000", 23480 => x"05000000",
    23481 => x"06000000", 23482 => x"01000000", 23483 => x"02000000",
    23484 => x"03000000", 23485 => x"04000000", 23486 => x"05000000",
    23487 => x"02000000", 23488 => x"03000000", 23489 => x"04000000",
    23490 => x"05000000", 23491 => x"000170f8", 23492 => x"000171fc",
    23493 => x"00000000", 23494 => x"00000000", 23495 => x"00000004",
    23496 => x"00000008", 23497 => x"00000100", 23498 => x"00000200",
    23499 => x"046362a0", 23500 => x"00019274", 23501 => x"00000000",
    23502 => x"00000000", 23503 => x"0000ce42", 23504 => x"ab28633a",
    23505 => x"00000000", 23506 => x"00018ee0", 23507 => x"00000000",
    23508 => x"00000000", 23509 => x"0000ce42", 23510 => x"650c2d4f",
    23511 => x"00000000", 23512 => x"0001927c", 23513 => x"00000000",
    23514 => x"00000000", 23515 => x"0000ce42", 23516 => x"65158dc0",
    23517 => x"00000000", 23518 => x"00018f00", 23519 => x"00000000",
    23520 => x"00000000", 23521 => x"0000ce42", 23522 => x"de0d8ced",
    23523 => x"00000000", 23524 => x"00019278", 23525 => x"00000000",
    23526 => x"00000000", 23527 => x"0000ce42", 23528 => x"ff07fc47",
    23529 => x"00000000", 23530 => x"00019240", 23531 => x"00000000",
    23532 => x"00000000", 23533 => x"0000ce42", 23534 => x"e2d13d04",
    23535 => x"00000000", 23536 => x"00019210", 23537 => x"00000000",
    23538 => x"00000000", 23539 => x"0000ce42", 23540 => x"779c5443",
    23541 => x"00000000", 23542 => x"00019270", 23543 => x"00000000",
    23544 => x"00000000", 23545 => x"00000651", 23546 => x"68202b22",
    23547 => x"00000000", 23548 => x"00019268", 23549 => x"00000000",
    23550 => x"00000000", 23551 => x"00001103", 23552 => x"c0413599",
    23553 => x"00000000", 23554 => x"00019254", 23555 => x"00000000",
    23556 => x"00000000", 23557 => x"00001103", 23558 => x"f0f43591",
    23559 => x"00000000", 23560 => x"0001566c", 23561 => x"00000000",
    23562 => x"00000001", 23563 => x"00030000", 23564 => x"00000004",
    23565 => x"00000000", 23566 => x"00000000", 23567 => x"00000000",
    23568 => x"00000000", 23569 => x"00000000", 23570 => x"00000000",
    23571 => x"00000000", 23572 => x"00000000", 23573 => x"00000000",
    23574 => x"00000000", 23575 => x"00000000", 23576 => x"00000000",
    23577 => x"00000000", 23578 => x"00000000", 23579 => x"00000000",
    23580 => x"00000000", 23581 => x"00000000", 23582 => x"00000000",
    23583 => x"00000000", 23584 => x"00000000", 23585 => x"00000000",
    23586 => x"00000000", 23587 => x"00000000", 23588 => x"00000000",
    23589 => x"00000000", 23590 => x"00000000", 23591 => x"00000000",
    23592 => x"00000000", 23593 => x"00000000", 23594 => x"00000000",
    23595 => x"00000000", 23596 => x"00000000", 23597 => x"00000000",
    23598 => x"00000000", 23599 => x"00000000", 23600 => x"00000000",
    23601 => x"00000000", 23602 => x"00000000", 23603 => x"00000000",
    23604 => x"00000000", 23605 => x"00000000", 23606 => x"ff000000",
    23607 => x"0000fe08", 23608 => x"0000fe3c", 23609 => x"0000fe6c",
    23610 => x"00014a38", 23611 => x"80000000", 23612 => x"00000000",
    23613 => x"00000000", 23614 => x"44332211", 23615 => x"00000000",
    23616 => x"04000000", 23617 => x"138046e2", 23618 => x"01000000",
    23619 => x"9000cfea", 23620 => x"01000000", 23621 => x"108157f3",
    23622 => x"01000000", 23623 => x"0be0ffff", 23624 => x"01000000",
    23625 => x"88e0ffff", 23626 => x"01000000", 23627 => x"08e1ffff",
    23628 => x"01000000", 23629 => x"1b0020e0", 23630 => x"01000000",
    23631 => x"9800c0eb", 23632 => x"01000000", 23633 => x"6b2130e0",
    23634 => x"01000000", 23635 => x"69610de0", 23636 => x"01000000",
    23637 => x"10a38900", 23638 => x"04000000", 23639 => x"6b0320f0",
    23640 => x"01000000", 23641 => x"bb0d8001", 23642 => x"04000000",
    23643 => x"33e31ef1", 23644 => x"01000000", 23645 => x"31c35ff9",
    23646 => x"01000000", 23647 => x"2b0300e1", 23648 => x"01000000",
    23649 => x"33e31ef1", 23650 => x"01000000", 23651 => x"43c300e1",
    23652 => x"01000000", 23653 => x"79411400", 23654 => x"04000000",
    23655 => x"cb250060", 23656 => x"00000000", 23657 => x"d3250260",
    23658 => x"00000000", 23659 => x"50ea8101", 23660 => x"04000000",
    23661 => x"81c88001", 23662 => x"04000000", 23663 => x"802fc100",
    23664 => x"04000000", 23665 => x"5b090080", 23666 => x"01000000",
    23667 => x"59092080", 23668 => x"01000000", 23669 => x"c06ac100",
    23670 => x"04000000", 23671 => x"63097afd", 23672 => x"01000000",
    23673 => x"f88a8101", 23674 => x"04000000", 23675 => x"f48a8101",
    23676 => x"04000000", 23677 => x"00000000", 23678 => x"08000000",
    23679 => x"ffffffff", 23680 => x"00015f84", 23681 => x"5b1157a7",
    23682 => x"00000003", 23683 => x"00000000", 23684 => x"00000000",
    23685 => x"00000000", 23686 => x"00000000", 23687 => x"00000000",
    23688 => x"00000000", 23689 => x"00000000", 23690 => x"00000000",
    23691 => x"00000000", 23692 => x"00000000", 23693 => x"00000000",
    23694 => x"77727063", 23695 => x"2d76332e", 23696 => x"302d3131",
    23697 => x"2d673038", 23698 => x"34376234", 23699 => x"392d6469",
    23700 => x"72747900", 23701 => x"00000000", 23702 => x"53657020",
    23703 => x"32302032", 23704 => x"30313600", 23705 => x"00000000",
    23706 => x"31373a33", 23707 => x"303a3137", 23708 => x"00000000",
    23709 => x"00000000", 23710 => x"686f6e67", 23711 => x"6d696e67",
    23712 => x"00000000", 23713 => x"00000000", 23714 => x"00000000",
    23715 => x"00000000", 23716 => x"00000000", 23717 => x"00000000",
    23718 => x"00014f48", 23719 => x"000088b0", 23720 => x"00013714",
    23721 => x"00008970", 23722 => x"00014f60", 23723 => x"000089d0",
    23724 => x"00014f94", 23725 => x"00008a6c", 23726 => x"00014fe8",
    23727 => x"00008b84", 23728 => x"00015038", 23729 => x"00008c94",
    23730 => x"00015058", 23731 => x"00008d74", 23732 => x"0001507c",
    23733 => x"00008dd4", 23734 => x"000151ac", 23735 => x"00008ed8",
    23736 => x"000151e8", 23737 => x"00009270", 23738 => x"00015244",
    23739 => x"000094d8", 23740 => x"0001527c", 23741 => x"000095b0",
    23742 => x"00015284", 23743 => x"00009710", 23744 => x"00015288",
    23745 => x"00009728", 23746 => x"000152b8", 23747 => x"00009744",
    23748 => x"000152d0", 23749 => x"000097f0", 23750 => x"00015340",
    23751 => x"00009948", 23752 => x"0001535c", 23753 => x"00009a38",
    23754 => x"000151b0", 23755 => x"00009a80", 23756 => x"00015750",
    23757 => x"0000eb4c", 23758 => x"00015864", 23759 => x"000100b8",
    23760 => x"00015868", 23761 => x"0000ffbc", 23762 => x"0001586c",
    23763 => x"0000fec0", 23764 => x"000106ec", 23765 => x"00000000",
    23766 => x"000170e8", 23767 => x"0001372c", 23768 => x"00000000",
    23769 => x"00000214", 23770 => x"00000000", 23771 => x"00000000",
    23772 => x"00000000", 23773 => x"00000000", 23774 => x"00013700",
    23775 => x"00000000", 23776 => x"00000000", 23777 => x"00012408",
    23778 => x"00000000", 23779 => x"00000000", 23780 => x"00000000",
    23781 => x"00013708", 23782 => x"00000000", 23783 => x"00008804",
    23784 => x"000004f8", 23785 => x"00000000", 23786 => x"00000000",
    23787 => x"00000000", 23788 => x"00013714", 23789 => x"00000000",
    23790 => x"00000000", 23791 => x"00001118", 23792 => x"00000000",
    23793 => x"00000000", 23794 => x"00000000", 23795 => x"00013718",
    23796 => x"00000000", 23797 => x"000004d4", 23798 => x"00000468",
    23799 => x"00000000", 23800 => x"00000000", 23801 => x"00000000",
    23802 => x"00013720", 23803 => x"00000000", 23804 => x"00000000",
    23805 => x"00000378", 23806 => x"00000000", 23807 => x"00000000",
    23808 => x"00000000", 23809 => x"00014e30", 23810 => x"00000000",
    23811 => x"00000000", 23812 => x"000076a8", 23813 => x"00000000",
    23814 => x"00000000", 23815 => x"00000000", 23816 => x"000154b4",
    23817 => x"00019258", 23818 => x"00000000", 23819 => x"0000a1bc",
    23820 => x"00000000", 23821 => x"00000000", 23822 => x"00000000",
    23823 => x"000154bc", 23824 => x"00019258", 23825 => x"0000a92c",
    23826 => x"0000a9dc", 23827 => x"00000000", 23828 => x"00000000",
    23829 => x"00000000", 23830 => x"000154c4", 23831 => x"00019258",
    23832 => x"0000aee8", 23833 => x"0000ad5c", 23834 => x"00000000",
    23835 => x"00000000", 23836 => x"00000000", 23837 => x"0001552c",
    23838 => x"00019258", 23839 => x"0000c608", 23840 => x"0000b630",
    23841 => x"00000000", 23842 => x"00000000", 23843 => x"00000000",
    23844 => x"00015758", 23845 => x"00000000", 23846 => x"0000e824",
    23847 => x"0000e870", 23848 => x"00000000", 23849 => x"00000000",
    23850 => x"00000000", 23851 => x"00000000", 23852 => x"00000000",
    23853 => x"00000000", 23854 => x"00000000", 23855 => x"00000000",
    23856 => x"00000000", 23857 => x"00000000", 23858 => x"00000000",
    23859 => x"00000000", 23860 => x"00000000", 23861 => x"00000000",
    23862 => x"00000000", 23863 => x"00000000", 23864 => x"00000000",
    23865 => x"00000000", 23866 => x"00000000", 23867 => x"00000000",
    23868 => x"00000000", 23869 => x"00000000", 23870 => x"00000000",
    23871 => x"00000000", 23872 => x"00000000", 23873 => x"00000000",
    23874 => x"00000000", 23875 => x"00000000", 23876 => x"00000000",
    23877 => x"00000000", 23878 => x"00000000", 23879 => x"00000000",
    23880 => x"00000000", 23881 => x"00000000", 23882 => x"00000000",
    23883 => x"00000000", 23884 => x"00000000", 23885 => x"00000000",
    23886 => x"00000000", 23887 => x"00000000", 23888 => x"00000000",
    23889 => x"00000000", 23890 => x"00000000", 23891 => x"00000000",
    23892 => x"00000000", 23893 => x"00000000", 23894 => x"00000000",
    23895 => x"00000000", 23896 => x"00000000", 23897 => x"00000000",
    23898 => x"00000000", 23899 => x"00000000", 23900 => x"00000000",
    23901 => x"00000000", 23902 => x"00000000", 23903 => x"00000000",
    23904 => x"00000000", 23905 => x"00000000", 23906 => x"00000000",
    23907 => x"00000000", 23908 => x"00000000", 23909 => x"00000000",
    23910 => x"00000000", 23911 => x"00000000", 23912 => x"00000000",
    23913 => x"00000000", 23914 => x"00000000", 23915 => x"00000000",
    23916 => x"00000000", 23917 => x"00000000", 23918 => x"00000000",
    23919 => x"00000000", 23920 => x"00000000", 23921 => x"00000000",
    23922 => x"00000000", 23923 => x"00000000", 23924 => x"00000000",
    23925 => x"00000000", 23926 => x"00000000", 23927 => x"00000000",
    23928 => x"00000000", 23929 => x"00000000", 23930 => x"00000000",
    23931 => x"00000000", 23932 => x"00000000", 23933 => x"00000000",
    23934 => x"00000000", 23935 => x"00000000", 23936 => x"00000000",
    23937 => x"00000000", 23938 => x"00000000", 23939 => x"00000000",
    23940 => x"00000000", 23941 => x"00000000", 23942 => x"00000000",
    23943 => x"00000000", 23944 => x"00000000", 23945 => x"00000000",
    23946 => x"00000000", 23947 => x"00000000", 23948 => x"00000000",
    23949 => x"00000000", 23950 => x"00000000", 23951 => x"00000000",
    23952 => x"00000000", 23953 => x"00000000", 23954 => x"00000000",
    23955 => x"00000000", 23956 => x"00000000", 23957 => x"00000000",
    23958 => x"00000000", 23959 => x"00000000", 23960 => x"00000000",
    23961 => x"00000000", 23962 => x"00000000", 23963 => x"00000000",
    23964 => x"00000000", 23965 => x"00000000", 23966 => x"00000000",
    23967 => x"00000000", 23968 => x"00000000", 23969 => x"00000000",
    23970 => x"00000000", 23971 => x"00000000", 23972 => x"00000000",
    23973 => x"00000000", 23974 => x"00000000", 23975 => x"00000000",
    23976 => x"00000000", 23977 => x"00000000", 23978 => x"00000000",
    23979 => x"00000000", 23980 => x"00000000", 23981 => x"00000000",
    23982 => x"00000000", 23983 => x"00000000", 23984 => x"00000000",
    23985 => x"00000000", 23986 => x"00000000", 23987 => x"00000000",
    23988 => x"00000000", 23989 => x"00000000", 23990 => x"00000000",
    23991 => x"00000000", 23992 => x"00000000", 23993 => x"00000000",
    23994 => x"00000000", 23995 => x"00000000", 23996 => x"00000000",
    23997 => x"00000000", 23998 => x"00000000", 23999 => x"00000000",
    24000 => x"00000000", 24001 => x"00000000", 24002 => x"00000000",
    24003 => x"00000000", 24004 => x"00000000", 24005 => x"00000000",
    24006 => x"00000000", 24007 => x"00000000", 24008 => x"00000000",
    24009 => x"00000000", 24010 => x"00000000", 24011 => x"00000000",
    24012 => x"00000000", 24013 => x"00000000", 24014 => x"00000000",
    24015 => x"00000000", 24016 => x"00000000", 24017 => x"00000000",
    24018 => x"00000000", 24019 => x"00000000", 24020 => x"00000000",
    24021 => x"00000000", 24022 => x"00000000", 24023 => x"00000000",
    24024 => x"00000000", 24025 => x"00000000", 24026 => x"00000000",
    24027 => x"00000000", 24028 => x"00000000", 24029 => x"00000000",
    24030 => x"00000000", 24031 => x"00000000", 24032 => x"00000000",
    24033 => x"00000000", 24034 => x"00000000", 24035 => x"00000000",
    24036 => x"00000000", 24037 => x"00000000", 24038 => x"00000000",
    24039 => x"00000000", 24040 => x"00000000", 24041 => x"00000000",
    24042 => x"00000000", 24043 => x"00000000", 24044 => x"00000000",
    24045 => x"00000000", 24046 => x"00000000", 24047 => x"00000000",
    24048 => x"00000000", 24049 => x"00000000", 24050 => x"00000000",
    24051 => x"00000000", 24052 => x"00000000", 24053 => x"00000000",
    24054 => x"00000000", 24055 => x"00000000", 24056 => x"00000000",
    24057 => x"00000000", 24058 => x"00000000", 24059 => x"00000000",
    24060 => x"00000000", 24061 => x"00000000", 24062 => x"00000000",
    24063 => x"00000000", 24064 => x"00000000", 24065 => x"00000000",
    24066 => x"00000000", 24067 => x"00000000", 24068 => x"00000000",
    24069 => x"00000000", 24070 => x"00000000", 24071 => x"00000000",
    24072 => x"00000000", 24073 => x"00000000", 24074 => x"00000000",
    24075 => x"00000000", 24076 => x"00000000", 24077 => x"00000000",
    24078 => x"00000000", 24079 => x"00000000", 24080 => x"00000000",
    24081 => x"00000000", 24082 => x"00000000", 24083 => x"00000000",
    24084 => x"00000000", 24085 => x"00000000", 24086 => x"00000000",
    24087 => x"00000000", 24088 => x"00000000", 24089 => x"00000000",
    24090 => x"00000000", 24091 => x"00000000", 24092 => x"00000000",
    24093 => x"00000000", 24094 => x"00000000", 24095 => x"00000000",
    24096 => x"00000000", 24097 => x"00000000", 24098 => x"00000000",
    24099 => x"00000000", 24100 => x"00000000", 24101 => x"00000000",
    24102 => x"00000000", 24103 => x"00000000", 24104 => x"00000000",
    24105 => x"00000000", 24106 => x"00000000", 24107 => x"00000000",
    24108 => x"00000000", 24109 => x"00000000", 24110 => x"00000000",
    24111 => x"00000000", 24112 => x"00000000", 24113 => x"00000000",
    24114 => x"00000000", 24115 => x"00000000", 24116 => x"00000000",
    24117 => x"00000000", 24118 => x"00000000", 24119 => x"00000000",
    24120 => x"00000000", 24121 => x"00000000", 24122 => x"00000000",
    24123 => x"00000000", 24124 => x"00000000", 24125 => x"00000000",
    24126 => x"00000000", 24127 => x"00000000", 24128 => x"00000000",
    24129 => x"00000000", 24130 => x"00000000", 24131 => x"00000000",
    24132 => x"00000000", 24133 => x"00000000", 24134 => x"00000000",
    24135 => x"00000000", 24136 => x"00000000", 24137 => x"00000000",
    24138 => x"00000000", 24139 => x"00000000", 24140 => x"00000000",
    24141 => x"00000000", 24142 => x"00000000", 24143 => x"00000000",
    24144 => x"00000000", 24145 => x"00000000", 24146 => x"00000000",
    24147 => x"00000000", 24148 => x"00000000", 24149 => x"00000000",
    24150 => x"00000000", 24151 => x"00000000", 24152 => x"00000000",
    24153 => x"00000000", 24154 => x"00000000", 24155 => x"00000000",
    24156 => x"00000000", 24157 => x"00000000", 24158 => x"00000000",
    24159 => x"00000000", 24160 => x"00000000", 24161 => x"00000000",
    24162 => x"00000000", 24163 => x"00000000", 24164 => x"00000000",
    24165 => x"00000000", 24166 => x"00000000", 24167 => x"00000000",
    24168 => x"00000000", 24169 => x"00000000", 24170 => x"00000000",
    24171 => x"00000000", 24172 => x"00000000", 24173 => x"00000000",
    24174 => x"00000000", 24175 => x"00000000", 24176 => x"00000000",
    24177 => x"00000000", 24178 => x"00000000", 24179 => x"00000000",
    24180 => x"00000000", 24181 => x"00000000", 24182 => x"00000000",
    24183 => x"00000000", 24184 => x"00000000", 24185 => x"00000000",
    24186 => x"00000000", 24187 => x"00000000", 24188 => x"00000000",
    24189 => x"00000000", 24190 => x"00000000", 24191 => x"00000000",
    24192 => x"00000000", 24193 => x"00000000", 24194 => x"00000000",
    24195 => x"00000000", 24196 => x"00000000", 24197 => x"00000000",
    24198 => x"00000000", 24199 => x"00000000", 24200 => x"00000000",
    24201 => x"00000000", 24202 => x"00000000", 24203 => x"00000000",
    24204 => x"00000000", 24205 => x"00000000", 24206 => x"00000000",
    24207 => x"00000000", 24208 => x"00000000", 24209 => x"00000000",
    24210 => x"00000000", 24211 => x"00000000", 24212 => x"00000000",
    24213 => x"00000000", 24214 => x"00000000", 24215 => x"00000000",
    24216 => x"00000000", 24217 => x"00000000", 24218 => x"00000000",
    24219 => x"00000000", 24220 => x"00000000", 24221 => x"00000000",
    24222 => x"00000000", 24223 => x"00000000", 24224 => x"00000000",
    24225 => x"00000000", 24226 => x"00000000", 24227 => x"00000000",
    24228 => x"00000000", 24229 => x"00000000", 24230 => x"00000000",
    24231 => x"00000000", 24232 => x"00000000", 24233 => x"00000000",
    24234 => x"00000000", 24235 => x"00000000", 24236 => x"00000000",
    24237 => x"00000000", 24238 => x"00000000", 24239 => x"00000000",
    24240 => x"00000000", 24241 => x"00000000", 24242 => x"00000000",
    24243 => x"00000000", 24244 => x"00000000", 24245 => x"00000000",
    24246 => x"00000000", 24247 => x"00000000", 24248 => x"00000000",
    24249 => x"00000000", 24250 => x"00000000", 24251 => x"00000000",
    24252 => x"00000000", 24253 => x"00000000", 24254 => x"00000000",
    24255 => x"00000000", 24256 => x"00000000", 24257 => x"00000000",
    24258 => x"00000000", 24259 => x"00000000", 24260 => x"00000000",
    24261 => x"00000000", 24262 => x"00000000", 24263 => x"00000000",
    24264 => x"00000000", 24265 => x"00000000", 24266 => x"00000000",
    24267 => x"00000000", 24268 => x"00000000", 24269 => x"00000000",
    24270 => x"00000000", 24271 => x"00000000", 24272 => x"00000000",
    24273 => x"00000000", 24274 => x"00000000", 24275 => x"00000000",
    24276 => x"00000000", 24277 => x"00000000", 24278 => x"00000000",
    24279 => x"00000000", 24280 => x"00000000", 24281 => x"00000000",
    24282 => x"00000000", 24283 => x"00000000", 24284 => x"00000000",
    24285 => x"00000000", 24286 => x"00000000", 24287 => x"00000000",
    24288 => x"00000000", 24289 => x"00000000", 24290 => x"00000000",
    24291 => x"00000000", 24292 => x"00000000", 24293 => x"00000000",
    24294 => x"00000000", 24295 => x"00000000", 24296 => x"00000000",
    24297 => x"00000000", 24298 => x"00000000", 24299 => x"00000000",
    24300 => x"00000000", 24301 => x"00000000", 24302 => x"00000000",
    24303 => x"00000000", 24304 => x"00000000", 24305 => x"00000000",
    24306 => x"00000000", 24307 => x"00000000", 24308 => x"00000000",
    24309 => x"00000000", 24310 => x"00000000", 24311 => x"00000000",
    24312 => x"00000000", 24313 => x"00000000", 24314 => x"00000000",
    24315 => x"00000000", 24316 => x"00000000", 24317 => x"00000000",
    24318 => x"00000000", 24319 => x"00000000", 24320 => x"00000000",
    24321 => x"00000000", 24322 => x"00000000", 24323 => x"00000000",
    24324 => x"00000000", 24325 => x"00000000", 24326 => x"00000000",
    24327 => x"00000000", 24328 => x"00000000", 24329 => x"00000000",
    24330 => x"00000000", 24331 => x"00000000", 24332 => x"00000000",
    24333 => x"00000000", 24334 => x"00000000", 24335 => x"00000000",
    24336 => x"00000000", 24337 => x"00000000", 24338 => x"00000000",
    24339 => x"00000000", 24340 => x"00000000", 24341 => x"00000000",
    24342 => x"00000000", 24343 => x"00000000", 24344 => x"00000000",
    24345 => x"00000000", 24346 => x"00000000", 24347 => x"00000000",
    24348 => x"00000000", 24349 => x"00000000", 24350 => x"00000000",
    24351 => x"00000000", 24352 => x"00000000", 24353 => x"00000000",
    24354 => x"00000000", 24355 => x"00000000", 24356 => x"00000000",
    24357 => x"00000000", 24358 => x"00000000", 24359 => x"00000000",
    24360 => x"00000000", 24361 => x"00000000", 24362 => x"00000000",
    24363 => x"00000000", 24364 => x"00000000", 24365 => x"00000000",
    24366 => x"00000000", 24367 => x"00000000", 24368 => x"00000000",
    24369 => x"00000000", 24370 => x"00000000", 24371 => x"00000000",
    24372 => x"00000000", 24373 => x"00000000", 24374 => x"00000000",
    24375 => x"00000000", 24376 => x"00000000", 24377 => x"00000000",
    24378 => x"00000000", 24379 => x"00000000", 24380 => x"00000000",
    24381 => x"00000000", 24382 => x"00000000", 24383 => x"00000000",
    24384 => x"00000000", 24385 => x"00000000", 24386 => x"00000000",
    24387 => x"00000000", 24388 => x"00000000", 24389 => x"00000000",
    24390 => x"00000000", 24391 => x"00000000", 24392 => x"00000000",
    24393 => x"00000000", 24394 => x"00000000", 24395 => x"00000000",
    24396 => x"00000000", 24397 => x"00000000", 24398 => x"00000000",
    24399 => x"00000000", 24400 => x"00000000", 24401 => x"00000000",
    24402 => x"00000000", 24403 => x"00000000", 24404 => x"00000000",
    24405 => x"00000000", 24406 => x"00000000", 24407 => x"00000000",
    24408 => x"00000000", 24409 => x"00000000", 24410 => x"00000000",
    24411 => x"00000000", 24412 => x"00000000", 24413 => x"00000000",
    24414 => x"00000000", 24415 => x"00000000", 24416 => x"00000000",
    24417 => x"00000000", 24418 => x"00000000", 24419 => x"00000000",
    24420 => x"00000000", 24421 => x"00000000", 24422 => x"00000000",
    24423 => x"00000000", 24424 => x"00000000", 24425 => x"00000000",
    24426 => x"00000000", 24427 => x"00000000", 24428 => x"00000000",
    24429 => x"00000000", 24430 => x"00000000", 24431 => x"00000000",
    24432 => x"00000000", 24433 => x"00000000", 24434 => x"00000000",
    24435 => x"00000000", 24436 => x"00000000", 24437 => x"00000000",
    24438 => x"00000000", 24439 => x"00000000", 24440 => x"00000000",
    24441 => x"00000000", 24442 => x"00000000", 24443 => x"00000000",
    24444 => x"00000000", 24445 => x"00000000", 24446 => x"00000000",
    24447 => x"00000000", 24448 => x"00000000", 24449 => x"00000000",
    24450 => x"00000000", 24451 => x"00000000", 24452 => x"00000000",
    24453 => x"00000000", 24454 => x"00000000", 24455 => x"00000000",
    24456 => x"00000000", 24457 => x"00000000", 24458 => x"00000000",
    24459 => x"00000000", 24460 => x"00000000", 24461 => x"00000000",
    24462 => x"00000000", 24463 => x"00000000", 24464 => x"00000000",
    24465 => x"00000000", 24466 => x"00000000", 24467 => x"00000000",
    24468 => x"00000000", 24469 => x"00000000", 24470 => x"00000000",
    24471 => x"00000000", 24472 => x"00000000", 24473 => x"00000000",
    24474 => x"00000000", 24475 => x"00000000", 24476 => x"00000000",
    24477 => x"00000000", 24478 => x"00000000", 24479 => x"00000000",
    24480 => x"00000000", 24481 => x"00000000", 24482 => x"00000000",
    24483 => x"00000000", 24484 => x"00000000", 24485 => x"00000000",
    24486 => x"00000000", 24487 => x"00000000", 24488 => x"00000000",
    24489 => x"00000000", 24490 => x"00000000", 24491 => x"00000000",
    24492 => x"00000000", 24493 => x"00000000", 24494 => x"00000000",
    24495 => x"00000000", 24496 => x"00000000", 24497 => x"00000000",
    24498 => x"00000000", 24499 => x"00000000", 24500 => x"00000000",
    24501 => x"00000000", 24502 => x"00000000", 24503 => x"00000000",
    24504 => x"00000000", 24505 => x"00000000", 24506 => x"00000000",
    24507 => x"00000000", 24508 => x"00000000", 24509 => x"00000000",
    24510 => x"00000000", 24511 => x"00000000", 24512 => x"00000000",
    24513 => x"00000000", 24514 => x"00000000", 24515 => x"00000000",
    24516 => x"00000000", 24517 => x"00000000", 24518 => x"00000000",
    24519 => x"00000000", 24520 => x"00000000", 24521 => x"00000000",
    24522 => x"00000000", 24523 => x"00000000", 24524 => x"00000000",
    24525 => x"00000000", 24526 => x"00000000", 24527 => x"00000000",
    24528 => x"00000000", 24529 => x"00000000", 24530 => x"00000000",
    24531 => x"00000000", 24532 => x"00000000", 24533 => x"00000000",
    24534 => x"00000000", 24535 => x"00000000", 24536 => x"00000000",
    24537 => x"00000000", 24538 => x"00000000", 24539 => x"00000000",
    24540 => x"00000000", 24541 => x"00000000", 24542 => x"00000000",
    24543 => x"00000000", 24544 => x"00000000", 24545 => x"00000000",
    24546 => x"00000000", 24547 => x"00000000", 24548 => x"00000000",
    24549 => x"00000000", 24550 => x"00000000", 24551 => x"00000000",
    24552 => x"00000000", 24553 => x"00000000", 24554 => x"00000000",
    24555 => x"00000000", 24556 => x"00000000", 24557 => x"00000000",
    24558 => x"00000000", 24559 => x"00000000", 24560 => x"00000000",
    24561 => x"00000000", 24562 => x"00000000", 24563 => x"00000000",
    24564 => x"00000000", 24565 => x"00000000", 24566 => x"00000000",
    24567 => x"00000000", 24568 => x"00000000", 24569 => x"00000000",
    24570 => x"00000000", 24571 => x"00000000", 24572 => x"00000000",
    24573 => x"00000000", 24574 => x"00000000", 24575 => x"00000000",
    24576 => x"00000000", 24577 => x"00000000", 24578 => x"00000000",
    24579 => x"00000000", 24580 => x"00000000", 24581 => x"00000000",
    24582 => x"00000000", 24583 => x"00000000", 24584 => x"00000000",
    24585 => x"00000000", 24586 => x"00000000", 24587 => x"00000000",
    24588 => x"00000000", 24589 => x"00000000", 24590 => x"00000000",
    24591 => x"00000000", 24592 => x"00000000", 24593 => x"00000000",
    24594 => x"00000000", 24595 => x"00000000", 24596 => x"00000000",
    24597 => x"00000000", 24598 => x"00000000", 24599 => x"00000000",
    24600 => x"00000000", 24601 => x"00000000", 24602 => x"00000000",
    24603 => x"00000000", 24604 => x"00000000", 24605 => x"00000000",
    24606 => x"00000000", 24607 => x"00000000", 24608 => x"00000000",
    24609 => x"00000000", 24610 => x"00000000", 24611 => x"00000000",
    24612 => x"00000000", 24613 => x"00000000", 24614 => x"00000000",
    24615 => x"00000000", 24616 => x"00000000", 24617 => x"00000000",
    24618 => x"00000000", 24619 => x"00000000", 24620 => x"00000000",
    24621 => x"00000000", 24622 => x"00000000", 24623 => x"00000000",
    24624 => x"00000000", 24625 => x"00000000", 24626 => x"00000000",
    24627 => x"00000000", 24628 => x"00000000", 24629 => x"00000000",
    24630 => x"00000000", 24631 => x"00000000", 24632 => x"00000000",
    24633 => x"00000000", 24634 => x"00000000", 24635 => x"00000000",
    24636 => x"00000000", 24637 => x"00000000", 24638 => x"00000000",
    24639 => x"00000000", 24640 => x"00000000", 24641 => x"00000000",
    24642 => x"00000000", 24643 => x"00000000", 24644 => x"00000000",
    24645 => x"00000000", 24646 => x"00000000", 24647 => x"00000000",
    24648 => x"00000000", 24649 => x"00000000", 24650 => x"00000000",
    24651 => x"00000000", 24652 => x"00000000", 24653 => x"00000000",
    24654 => x"00000000", 24655 => x"00000000", 24656 => x"00000000",
    24657 => x"00000000", 24658 => x"00000000", 24659 => x"00000000",
    24660 => x"00000000", 24661 => x"00000000", 24662 => x"00000000",
    24663 => x"00000000", 24664 => x"00000000", 24665 => x"00000000",
    24666 => x"00000000", 24667 => x"00000000", 24668 => x"00000000",
    24669 => x"00000000", 24670 => x"00000000", 24671 => x"00000000",
    24672 => x"00000000", 24673 => x"00000000", 24674 => x"00000000",
    24675 => x"00000000", 24676 => x"00000000", 24677 => x"00000000",
    24678 => x"00000000", 24679 => x"00000000", 24680 => x"00000000",
    24681 => x"00000000", 24682 => x"00000000", 24683 => x"00000000",
    24684 => x"00000000", 24685 => x"00000000", 24686 => x"00000000",
    24687 => x"00000000", 24688 => x"00000000", 24689 => x"00000000",
    24690 => x"00000000", 24691 => x"00000000", 24692 => x"00000000",
    24693 => x"00000000", 24694 => x"00000000", 24695 => x"00000000",
    24696 => x"00000000", 24697 => x"00000000", 24698 => x"00000000",
    24699 => x"00000000", 24700 => x"00000000", 24701 => x"00000000",
    24702 => x"00000000", 24703 => x"00000000", 24704 => x"00000000",
    24705 => x"00000000", 24706 => x"00000000", 24707 => x"00000000",
    24708 => x"00000000", 24709 => x"00000000", 24710 => x"00000000",
    24711 => x"00000000", 24712 => x"00000000", 24713 => x"00000000",
    24714 => x"00000000", 24715 => x"00000000", 24716 => x"00000000",
    24717 => x"00000000", 24718 => x"00000000", 24719 => x"00000000",
    24720 => x"00000000", 24721 => x"00000000", 24722 => x"00000000",
    24723 => x"00000000", 24724 => x"00000000", 24725 => x"00000000",
    24726 => x"00000000", 24727 => x"00000000", 24728 => x"00000000",
    24729 => x"00000000", 24730 => x"00000000", 24731 => x"00000000",
    24732 => x"00000000", 24733 => x"00000000", 24734 => x"00000000",
    24735 => x"00000000", 24736 => x"00000000", 24737 => x"00000000",
    24738 => x"00000000", 24739 => x"00000000", 24740 => x"00000000",
    24741 => x"00000000", 24742 => x"00000000", 24743 => x"00000000",
    24744 => x"00000000", 24745 => x"00000000", 24746 => x"00000000",
    24747 => x"00000000", 24748 => x"00000000", 24749 => x"00000000",
    24750 => x"00000000", 24751 => x"00000000", 24752 => x"00000000",
    24753 => x"00000000", 24754 => x"00000000", 24755 => x"00000000",
    24756 => x"00000000", 24757 => x"00000000", 24758 => x"00000000",
    24759 => x"00000000", 24760 => x"00000000", 24761 => x"00000000",
    24762 => x"00000000", 24763 => x"00000000", 24764 => x"00000000",
    24765 => x"00000000", 24766 => x"00000000", 24767 => x"00000000",
    24768 => x"00000000", 24769 => x"00000000", 24770 => x"00000000",
    24771 => x"00000000", 24772 => x"00000000", 24773 => x"00000000",
    24774 => x"00000000", 24775 => x"00000000", 24776 => x"00000000",
    24777 => x"00000000", 24778 => x"00000000", 24779 => x"00000000",
    24780 => x"00000000", 24781 => x"00000000", 24782 => x"00000000",
    24783 => x"00000000", 24784 => x"00000000", 24785 => x"00000000",
    24786 => x"00000000", 24787 => x"00000000", 24788 => x"00000000",
    24789 => x"00000000", 24790 => x"00000000", 24791 => x"00000000",
    24792 => x"00000000", 24793 => x"00000000", 24794 => x"00000000",
    24795 => x"00000000", 24796 => x"00000000", 24797 => x"00000000",
    24798 => x"00000000", 24799 => x"00000000", 24800 => x"00000000",
    24801 => x"00000000", 24802 => x"00000000", 24803 => x"00000000",
    24804 => x"00000000", 24805 => x"00000000", 24806 => x"00000000",
    24807 => x"00000000", 24808 => x"00000000", 24809 => x"00000000",
    24810 => x"00000000", 24811 => x"00000000", 24812 => x"00000000",
    24813 => x"00000000", 24814 => x"00000000", 24815 => x"00000000",
    24816 => x"00000000", 24817 => x"00000000", 24818 => x"00000000",
    24819 => x"00000000", 24820 => x"00000000", 24821 => x"00000000",
    24822 => x"00000000", 24823 => x"00000000", 24824 => x"00000000",
    24825 => x"00000000", 24826 => x"00000000", 24827 => x"00000000",
    24828 => x"00000000", 24829 => x"00000000", 24830 => x"00000000",
    24831 => x"00000000", 24832 => x"00000000", 24833 => x"00000000",
    24834 => x"00000000", 24835 => x"00000000", 24836 => x"00000000",
    24837 => x"00000000", 24838 => x"00000000", 24839 => x"00000000",
    24840 => x"00000000", 24841 => x"00000000", 24842 => x"00000000",
    24843 => x"00000000", 24844 => x"00000000", 24845 => x"00000000",
    24846 => x"00000000", 24847 => x"00000000", 24848 => x"00000000",
    24849 => x"00000000", 24850 => x"00000000", 24851 => x"00000000",
    24852 => x"00000000", 24853 => x"00000000", 24854 => x"00000000",
    24855 => x"00000000", 24856 => x"00000000", 24857 => x"00000000",
    24858 => x"00000000", 24859 => x"00000000", 24860 => x"00000000",
    24861 => x"00000000", 24862 => x"00000000", 24863 => x"00000000",
    24864 => x"00000000", 24865 => x"00000000", 24866 => x"00000000",
    24867 => x"00000000", 24868 => x"00000000", 24869 => x"00000000",
    24870 => x"00000000", 24871 => x"00000000", 24872 => x"00000000",
    24873 => x"00000000", 24874 => x"00000000", 24875 => x"00000000",
    24876 => x"00000000", 24877 => x"00000000", 24878 => x"00000000",
    24879 => x"00000000", 24880 => x"00000000", 24881 => x"00000000",
    24882 => x"00000000", 24883 => x"00000000", 24884 => x"00000000",
    24885 => x"00000000", 24886 => x"00000000", 24887 => x"00000000",
    24888 => x"00000000", 24889 => x"00000000", 24890 => x"00000000",
    24891 => x"00000000", 24892 => x"00000000", 24893 => x"00000000",
    24894 => x"00000000", 24895 => x"00000000", 24896 => x"00000000",
    24897 => x"00000000", 24898 => x"00000000", 24899 => x"00000000",
    24900 => x"00000000", 24901 => x"00000000", 24902 => x"00000000",
    24903 => x"00000000", 24904 => x"00000000", 24905 => x"00000000",
    24906 => x"00000000", 24907 => x"00000000", 24908 => x"00000000",
    24909 => x"00000000", 24910 => x"00000000", 24911 => x"00000000",
    24912 => x"00000000", 24913 => x"00000000", 24914 => x"00000000",
    24915 => x"00000000", 24916 => x"00000000", 24917 => x"00000000",
    24918 => x"00000000", 24919 => x"00000000", 24920 => x"00000000",
    24921 => x"00000000", 24922 => x"00000000", 24923 => x"00000000",
    24924 => x"00000000", 24925 => x"00000000", 24926 => x"00000000",
    24927 => x"00000000", 24928 => x"00000000", 24929 => x"00000000",
    24930 => x"00000000", 24931 => x"00000000", 24932 => x"00000000",
    24933 => x"00000000", 24934 => x"00000000", 24935 => x"00000000",
    24936 => x"00000000", 24937 => x"00000000", 24938 => x"00000000",
    24939 => x"00000000", 24940 => x"00000000", 24941 => x"00000000",
    24942 => x"00000000", 24943 => x"00000000", 24944 => x"00000000",
    24945 => x"00000000", 24946 => x"00000000", 24947 => x"00000000",
    24948 => x"00000000", 24949 => x"00000000", 24950 => x"00000000",
    24951 => x"00000000", 24952 => x"00000000", 24953 => x"00000000",
    24954 => x"00000000", 24955 => x"00000000", 24956 => x"00000000",
    24957 => x"00000000", 24958 => x"00000000", 24959 => x"00000000",
    24960 => x"00000000", 24961 => x"00000000", 24962 => x"00000000",
    24963 => x"00000000", 24964 => x"00000000", 24965 => x"00000000",
    24966 => x"00000000", 24967 => x"00000000", 24968 => x"00000000",
    24969 => x"00000000", 24970 => x"00000000", 24971 => x"00000000",
    24972 => x"00000000", 24973 => x"00000000", 24974 => x"00000000",
    24975 => x"00000000", 24976 => x"00000000", 24977 => x"00000000",
    24978 => x"00000000", 24979 => x"00000000", 24980 => x"00000000",
    24981 => x"00000000", 24982 => x"00000000", 24983 => x"00000000",
    24984 => x"00000000", 24985 => x"00000000", 24986 => x"00000000",
    24987 => x"00000000", 24988 => x"00000000", 24989 => x"00000000",
    24990 => x"00000000", 24991 => x"00000000", 24992 => x"00000000",
    24993 => x"00000000", 24994 => x"00000000", 24995 => x"00000000",
    24996 => x"00000000", 24997 => x"00000000", 24998 => x"00000000",
    24999 => x"00000000", 25000 => x"00000000", 25001 => x"00000000",
    25002 => x"00000000", 25003 => x"00000000", 25004 => x"00000000",
    25005 => x"00000000", 25006 => x"00000000", 25007 => x"00000000",
    25008 => x"00000000", 25009 => x"00000000", 25010 => x"00000000",
    25011 => x"00000000", 25012 => x"00000000", 25013 => x"00000000",
    25014 => x"00000000", 25015 => x"00000000", 25016 => x"00000000",
    25017 => x"00000000", 25018 => x"00000000", 25019 => x"00000000",
    25020 => x"00000000", 25021 => x"00000000", 25022 => x"00000000",
    25023 => x"00000000", 25024 => x"00000000", 25025 => x"00000000",
    25026 => x"00000000", 25027 => x"00000000", 25028 => x"00000000",
    25029 => x"00000000", 25030 => x"00000000", 25031 => x"00000000",
    25032 => x"00000000", 25033 => x"00000000", 25034 => x"00000000",
    25035 => x"00000000", 25036 => x"00000000", 25037 => x"00000000",
    25038 => x"00000000", 25039 => x"00000000", 25040 => x"00000000",
    25041 => x"00000000", 25042 => x"00000000", 25043 => x"00000000",
    25044 => x"00000000", 25045 => x"00000000", 25046 => x"00000000",
    25047 => x"00000000", 25048 => x"00000000", 25049 => x"00000000",
    25050 => x"00000000", 25051 => x"00000000", 25052 => x"00000000",
    25053 => x"00000000", 25054 => x"00000000", 25055 => x"00000000",
    25056 => x"00000000", 25057 => x"00000000", 25058 => x"00000000",
    25059 => x"00000000", 25060 => x"00000000", 25061 => x"00000000",
    25062 => x"00000000", 25063 => x"00000000", 25064 => x"00000000",
    25065 => x"00000000", 25066 => x"00000000", 25067 => x"00000000",
    25068 => x"00000000", 25069 => x"00000000", 25070 => x"00000000",
    25071 => x"00000000", 25072 => x"00000000", 25073 => x"00000000",
    25074 => x"00000000", 25075 => x"00000000", 25076 => x"00000000",
    25077 => x"00000000", 25078 => x"00000000", 25079 => x"00000000",
    25080 => x"00000000", 25081 => x"00000000", 25082 => x"00000000",
    25083 => x"00000000", 25084 => x"00000000", 25085 => x"00000000",
    25086 => x"00000000", 25087 => x"00000000", 25088 => x"00000000",
    25089 => x"00000000", 25090 => x"00000000", 25091 => x"00000000",
    25092 => x"00000000", 25093 => x"00000000", 25094 => x"00000000",
    25095 => x"00000000", 25096 => x"00000000", 25097 => x"00000000",
    25098 => x"00000000", 25099 => x"00000000", 25100 => x"00000000",
    25101 => x"00000000", 25102 => x"00000000", 25103 => x"00000000",
    25104 => x"00000000", 25105 => x"00000000", 25106 => x"00000000",
    25107 => x"00000000", 25108 => x"00000000", 25109 => x"00000000",
    25110 => x"00000000", 25111 => x"00000000", 25112 => x"00000000",
    25113 => x"00000000", 25114 => x"00000000", 25115 => x"00000000",
    25116 => x"00000000", 25117 => x"00000000", 25118 => x"00000000",
    25119 => x"00000000", 25120 => x"00000000", 25121 => x"00000000",
    25122 => x"00000000", 25123 => x"00000000", 25124 => x"00000000",
    25125 => x"00000000", 25126 => x"00000000", 25127 => x"00000000",
    25128 => x"00000000", 25129 => x"00000000", 25130 => x"00000000",
    25131 => x"00000000", 25132 => x"00000000", 25133 => x"00000000",
    25134 => x"00000000", 25135 => x"00000000", 25136 => x"00000000",
    25137 => x"00000000", 25138 => x"00000000", 25139 => x"00000000",
    25140 => x"00000000", 25141 => x"00000000", 25142 => x"00000000",
    25143 => x"00000000", 25144 => x"00000000", 25145 => x"00000000",
    25146 => x"00000000", 25147 => x"00000000", 25148 => x"00000000",
    25149 => x"00000000", 25150 => x"00000000", 25151 => x"00000000",
    25152 => x"00000000", 25153 => x"00000000", 25154 => x"00000000",
    25155 => x"00000000", 25156 => x"00000000", 25157 => x"00000000",
    25158 => x"00000000", 25159 => x"00000000", 25160 => x"00000000",
    25161 => x"00000000", 25162 => x"00000000", 25163 => x"00000000",
    25164 => x"00000000", 25165 => x"00000000", 25166 => x"00000000",
    25167 => x"00000000", 25168 => x"00000000", 25169 => x"00000000",
    25170 => x"00000000", 25171 => x"00000000", 25172 => x"00000000",
    25173 => x"00000000", 25174 => x"00000000", 25175 => x"00000000",
    25176 => x"00000000", 25177 => x"00000000", 25178 => x"00000000",
    25179 => x"00000000", 25180 => x"00000000", 25181 => x"00000000",
    25182 => x"00000000", 25183 => x"00000000", 25184 => x"00000000",
    25185 => x"00000000", 25186 => x"00000000", 25187 => x"00000000",
    25188 => x"00000000", 25189 => x"00000000", 25190 => x"00000000",
    25191 => x"00000000", 25192 => x"00000000", 25193 => x"00000000",
    25194 => x"00000000", 25195 => x"00000000", 25196 => x"00000000",
    25197 => x"00000000", 25198 => x"00000000", 25199 => x"00000000",
    25200 => x"00000000", 25201 => x"00000000", 25202 => x"00000000",
    25203 => x"00000000", 25204 => x"00000000", 25205 => x"00000000",
    25206 => x"00000000", 25207 => x"00000000", 25208 => x"00000000",
    25209 => x"00000000", 25210 => x"00000000", 25211 => x"00000000",
    25212 => x"00000000", 25213 => x"00000000", 25214 => x"00000000",
    25215 => x"00000000", 25216 => x"00000000", 25217 => x"00000000",
    25218 => x"00000000", 25219 => x"00000000", 25220 => x"00000000",
    25221 => x"00000000", 25222 => x"00000000", 25223 => x"00000000",
    25224 => x"00000000", 25225 => x"00000000", 25226 => x"00000000",
    25227 => x"00000000", 25228 => x"00000000", 25229 => x"00000000",
    25230 => x"00000000", 25231 => x"00000000", 25232 => x"00000000",
    25233 => x"00000000", 25234 => x"00000000", 25235 => x"00000000",
    25236 => x"00000000", 25237 => x"00000000", 25238 => x"00000000",
    25239 => x"00000000", 25240 => x"00000000", 25241 => x"00000000",
    25242 => x"00000000", 25243 => x"00000000", 25244 => x"00000000",
    25245 => x"00000000", 25246 => x"00000000", 25247 => x"00000000",
    25248 => x"00000000", 25249 => x"00000000", 25250 => x"00000000",
    25251 => x"00000000", 25252 => x"00000000", 25253 => x"00000000",
    25254 => x"00000000", 25255 => x"00000000", 25256 => x"00000000",
    25257 => x"00000000", 25258 => x"00000000", 25259 => x"00000000",
    25260 => x"00000000", 25261 => x"00000000", 25262 => x"00000000",
    25263 => x"00000000", 25264 => x"00000000", 25265 => x"00000000",
    25266 => x"00000000", 25267 => x"00000000", 25268 => x"00000000",
    25269 => x"00000000", 25270 => x"00000000", 25271 => x"00000000",
    25272 => x"00000000", 25273 => x"00000000", 25274 => x"00000000",
    25275 => x"00000000", 25276 => x"00000000", 25277 => x"00000000",
    25278 => x"00000000", 25279 => x"00000000", 25280 => x"00000000",
    25281 => x"00000000", 25282 => x"00000000", 25283 => x"00000000",
    25284 => x"00000000", 25285 => x"00000000", 25286 => x"00000000",
    25287 => x"00000000", 25288 => x"00000000", 25289 => x"00000000",
    25290 => x"00000000", 25291 => x"00000000", 25292 => x"00000000",
    25293 => x"00000000", 25294 => x"00000000", 25295 => x"00000000",
    25296 => x"00000000", 25297 => x"00000000", 25298 => x"00000000",
    25299 => x"00000000", 25300 => x"00000000", 25301 => x"00000000",
    25302 => x"00000000", 25303 => x"00000000", 25304 => x"00000000",
    25305 => x"00000000", 25306 => x"00000000", 25307 => x"00000000",
    25308 => x"00000000", 25309 => x"00000000", 25310 => x"00000000",
    25311 => x"00000000", 25312 => x"00000000", 25313 => x"00000000",
    25314 => x"00000000", 25315 => x"00000000", 25316 => x"00000000",
    25317 => x"00000000", 25318 => x"00000000", 25319 => x"00000000",
    25320 => x"00000000", 25321 => x"00000000", 25322 => x"00000000",
    25323 => x"00000000", 25324 => x"00000000", 25325 => x"00000000",
    25326 => x"00000000", 25327 => x"00000000", 25328 => x"00000000",
    25329 => x"00000000", 25330 => x"00000000", 25331 => x"00000000",
    25332 => x"00000000", 25333 => x"00000000", 25334 => x"00000000",
    25335 => x"00000000", 25336 => x"00000000", 25337 => x"00000000",
    25338 => x"00000000", 25339 => x"00000000", 25340 => x"00000000",
    25341 => x"00000000", 25342 => x"00000000", 25343 => x"00000000",
    25344 => x"00000000", 25345 => x"00000000", 25346 => x"00000000",
    25347 => x"00000000", 25348 => x"00000000", 25349 => x"00000000",
    25350 => x"00000000", 25351 => x"00000000", 25352 => x"00000000",
    25353 => x"00000000", 25354 => x"00000000", 25355 => x"00000000",
    25356 => x"00000000", 25357 => x"00000000", 25358 => x"00000000",
    25359 => x"00000000", 25360 => x"00000000", 25361 => x"00000000",
    25362 => x"00000000", 25363 => x"00000000", 25364 => x"00000000",
    25365 => x"00000000", 25366 => x"00000000", 25367 => x"00000000",
    25368 => x"00000000", 25369 => x"00000000", 25370 => x"00000000",
    25371 => x"00000000", 25372 => x"00000000", 25373 => x"00000000",
    25374 => x"00000000", 25375 => x"00000000", 25376 => x"00000000",
    25377 => x"00000000", 25378 => x"00000000", 25379 => x"00000000",
    25380 => x"00000000", 25381 => x"00000000", 25382 => x"00000000",
    25383 => x"00000000", 25384 => x"00000000", 25385 => x"00000000",
    25386 => x"00000000", 25387 => x"00000000", 25388 => x"00000000",
    25389 => x"00000000", 25390 => x"00000000", 25391 => x"00000000",
    25392 => x"00000000", 25393 => x"00000000", 25394 => x"00000000",
    25395 => x"00000000", 25396 => x"00000000", 25397 => x"00000000",
    25398 => x"00000000", 25399 => x"00000000", 25400 => x"00000000",
    25401 => x"00000000", 25402 => x"00000000", 25403 => x"00000000",
    25404 => x"00000000", 25405 => x"00000000", 25406 => x"00000000",
    25407 => x"00000000", 25408 => x"00000000", 25409 => x"00000000",
    25410 => x"00000000", 25411 => x"00000000", 25412 => x"00000000",
    25413 => x"00000000", 25414 => x"00000000", 25415 => x"00000000",
    25416 => x"00000000", 25417 => x"00000000", 25418 => x"00000000",
    25419 => x"00000000", 25420 => x"00000000", 25421 => x"00000000",
    25422 => x"00000000", 25423 => x"00000000", 25424 => x"00000000",
    25425 => x"00000000", 25426 => x"00000000", 25427 => x"00000000",
    25428 => x"00000000", 25429 => x"00000000", 25430 => x"00000000",
    25431 => x"00000000", 25432 => x"00000000", 25433 => x"00000000",
    25434 => x"00000000", 25435 => x"00000000", 25436 => x"00000000",
    25437 => x"00000000", 25438 => x"00000000", 25439 => x"00000000",
    25440 => x"00000000", 25441 => x"00000000", 25442 => x"00000000",
    25443 => x"00000000", 25444 => x"00000000", 25445 => x"00000000",
    25446 => x"00000000", 25447 => x"00000000", 25448 => x"00000000",
    25449 => x"00000000", 25450 => x"00000000", 25451 => x"00000000",
    25452 => x"00000000", 25453 => x"00000000", 25454 => x"00000000",
    25455 => x"00000000", 25456 => x"00000000", 25457 => x"00000000",
    25458 => x"00000000", 25459 => x"00000000", 25460 => x"00000000",
    25461 => x"00000000", 25462 => x"00000000", 25463 => x"00000000",
    25464 => x"00000000", 25465 => x"00000000", 25466 => x"00000000",
    25467 => x"00000000", 25468 => x"00000000", 25469 => x"00000000",
    25470 => x"00000000", 25471 => x"00000000", 25472 => x"00000000",
    25473 => x"00000000", 25474 => x"00000000", 25475 => x"00000000",
    25476 => x"00000000", 25477 => x"00000000", 25478 => x"00000000",
    25479 => x"00000000", 25480 => x"00000000", 25481 => x"00000000",
    25482 => x"00000000", 25483 => x"00000000", 25484 => x"00000000",
    25485 => x"00000000", 25486 => x"00000000", 25487 => x"00000000",
    25488 => x"00000000", 25489 => x"00000000", 25490 => x"00000000",
    25491 => x"00000000", 25492 => x"00000000", 25493 => x"00000000",
    25494 => x"00000000", 25495 => x"00000000", 25496 => x"00000000",
    25497 => x"00000000", 25498 => x"00000000", 25499 => x"00000000",
    25500 => x"00000000", 25501 => x"00000000", 25502 => x"00000000",
    25503 => x"00000000", 25504 => x"00000000", 25505 => x"00000000",
    25506 => x"00000000", 25507 => x"00000000", 25508 => x"00000000",
    25509 => x"00000000", 25510 => x"00000000", 25511 => x"00000000",
    25512 => x"00000000", 25513 => x"00000000", 25514 => x"00000000",
    25515 => x"00000000", 25516 => x"00000000", 25517 => x"00000000",
    25518 => x"00000000", 25519 => x"00000000", 25520 => x"00000000",
    25521 => x"00000000", 25522 => x"00000000", 25523 => x"00000000",
    25524 => x"00000000", 25525 => x"00000000", 25526 => x"00000000",
    25527 => x"00000000", 25528 => x"00000000", 25529 => x"00000000",
    25530 => x"00000000", 25531 => x"00000000", 25532 => x"00000000",
    25533 => x"00000000", 25534 => x"00000000", 25535 => x"00000000",
    25536 => x"00000000", 25537 => x"00000000", 25538 => x"00000000",
    25539 => x"00000000", 25540 => x"00000000", 25541 => x"00000000",
    25542 => x"00000000", 25543 => x"00000000", 25544 => x"00000000",
    25545 => x"00000000", 25546 => x"00000000", 25547 => x"00000000",
    25548 => x"00000000", 25549 => x"00000000", 25550 => x"00000000",
    25551 => x"00000000", 25552 => x"00000000", 25553 => x"00000000",
    25554 => x"00000000", 25555 => x"00000000", 25556 => x"00000000",
    25557 => x"00000000", 25558 => x"00000000", 25559 => x"00000000",
    25560 => x"00000000", 25561 => x"00000000", 25562 => x"00000000",
    25563 => x"00000000", 25564 => x"00000000", 25565 => x"00000000",
    25566 => x"00000000", 25567 => x"00000000", 25568 => x"00000000",
    25569 => x"00000000", 25570 => x"00000000", 25571 => x"00000000",
    25572 => x"00000000", 25573 => x"00000000", 25574 => x"00000000",
    25575 => x"00000000", 25576 => x"00000000", 25577 => x"00000000",
    25578 => x"00000000", 25579 => x"00000000", 25580 => x"00000000",
    25581 => x"00000000", 25582 => x"00000000", 25583 => x"00000000",
    25584 => x"00000000", 25585 => x"00000000", 25586 => x"00000000",
    25587 => x"00000000", 25588 => x"00000000", 25589 => x"00000000",
    25590 => x"00000000", 25591 => x"00000000", 25592 => x"00000000",
    25593 => x"00000000", 25594 => x"00000000", 25595 => x"00000000",
    25596 => x"00000000", 25597 => x"00000000", 25598 => x"00000000",
    25599 => x"00000000", 25600 => x"00000000", 25601 => x"00000000",
    25602 => x"00000000", 25603 => x"00000000", 25604 => x"00000000",
    25605 => x"00000000", 25606 => x"00000000", 25607 => x"00000000",
    25608 => x"00000000", 25609 => x"00000000", 25610 => x"00000000",
    25611 => x"00000000", 25612 => x"00000000", 25613 => x"00000000",
    25614 => x"00000000", 25615 => x"00000000", 25616 => x"00000000",
    25617 => x"00000000", 25618 => x"00000000", 25619 => x"00000000",
    25620 => x"00000000", 25621 => x"00000000", 25622 => x"00000000",
    25623 => x"00000000", 25624 => x"00000000", 25625 => x"00000000",
    25626 => x"00000000", 25627 => x"00000000", 25628 => x"00000000",
    25629 => x"00000000", 25630 => x"00000000", 25631 => x"00000000",
    25632 => x"00000000", 25633 => x"00000000", 25634 => x"00000000",
    25635 => x"00000000", 25636 => x"00000000", 25637 => x"00000000",
    25638 => x"00000000", 25639 => x"00000000", 25640 => x"00000000",
    25641 => x"00000000", 25642 => x"00000000", 25643 => x"00000000",
    25644 => x"00000000", 25645 => x"00000000", 25646 => x"00000000",
    25647 => x"00000000", 25648 => x"00000000", 25649 => x"00000000",
    25650 => x"00000000", 25651 => x"00000000", 25652 => x"00000000",
    25653 => x"00000000", 25654 => x"00000000", 25655 => x"00000000",
    25656 => x"00000000", 25657 => x"00000000", 25658 => x"00000000",
    25659 => x"00000000", 25660 => x"00000000", 25661 => x"00000000",
    25662 => x"00000000", 25663 => x"00000000", 25664 => x"00000000",
    25665 => x"00000000", 25666 => x"00000000", 25667 => x"00000000",
    25668 => x"00000000", 25669 => x"00000000", 25670 => x"00000000",
    25671 => x"00000000", 25672 => x"00000000", 25673 => x"00000000",
    25674 => x"00000000", 25675 => x"00000000", 25676 => x"00000000",
    25677 => x"00000000", 25678 => x"00000000", 25679 => x"00000000",
    25680 => x"00000000", 25681 => x"00000000", 25682 => x"00000000",
    25683 => x"00000000", 25684 => x"00000000", 25685 => x"00000000",
    25686 => x"00000000", 25687 => x"00000000", 25688 => x"00000000",
    25689 => x"00000000", 25690 => x"00000000", 25691 => x"00000000",
    25692 => x"00000000", 25693 => x"00000000", 25694 => x"00000000",
    25695 => x"00000000", 25696 => x"00000000", 25697 => x"00000000",
    25698 => x"00000000", 25699 => x"00000000", 25700 => x"00000000",
    25701 => x"00000000", 25702 => x"00000000", 25703 => x"00000000",
    25704 => x"00000000", 25705 => x"00000000", 25706 => x"00000000",
    25707 => x"00000000", 25708 => x"00000000", 25709 => x"00000000",
    25710 => x"00000000", 25711 => x"00000000", 25712 => x"00000000",
    25713 => x"00000000", 25714 => x"00000000", 25715 => x"00000000",
    25716 => x"00000000", 25717 => x"00000000", 25718 => x"00000000",
    25719 => x"00000000", 25720 => x"00000000", 25721 => x"00000000",
    25722 => x"00000000", 25723 => x"00000000", 25724 => x"00000000",
    25725 => x"00000000", 25726 => x"00000000", 25727 => x"00000000",
    25728 => x"00000000", 25729 => x"00000000", 25730 => x"00000000",
    25731 => x"00000000", 25732 => x"00000000", 25733 => x"00000000",
    25734 => x"00000000", 25735 => x"00000000", 25736 => x"00000000",
    25737 => x"00000000", 25738 => x"00000000", 25739 => x"00000000",
    25740 => x"00000000", 25741 => x"00000000", 25742 => x"00000000",
    25743 => x"00000000", 25744 => x"00000000", 25745 => x"00000000",
    25746 => x"00000000", 25747 => x"00000000", 25748 => x"00000000",
    25749 => x"00000000", 25750 => x"00000000", 25751 => x"00000000",
    25752 => x"00000000", 25753 => x"00000000", 25754 => x"00000000",
    25755 => x"00000000", 25756 => x"00000000", 25757 => x"00000000",
    25758 => x"00000000", 25759 => x"00000000", 25760 => x"00000000",
    25761 => x"00000000", 25762 => x"00000000", 25763 => x"00000000",
    25764 => x"00000000", 25765 => x"00000000", 25766 => x"00000000",
    25767 => x"00000000", 25768 => x"00000000", 25769 => x"00000000",
    25770 => x"00000000", 25771 => x"00000000", 25772 => x"00000000",
    25773 => x"00000000", 25774 => x"00000000", 25775 => x"00000000",
    25776 => x"00000000", 25777 => x"00000000", 25778 => x"00000000",
    25779 => x"00000000", 25780 => x"00000000", 25781 => x"00000000",
    25782 => x"00000000", 25783 => x"00000000", 25784 => x"00000000",
    25785 => x"00000000", 25786 => x"00000000", 25787 => x"00000000",
    25788 => x"00000000", 25789 => x"00000000", 25790 => x"00000000",
    25791 => x"00000000", 25792 => x"00000000", 25793 => x"00000000",
    25794 => x"00000000", 25795 => x"00000000", 25796 => x"00000000",
    25797 => x"00000000", 25798 => x"00000000", 25799 => x"00000000",
    25800 => x"00000000", 25801 => x"00000000", 25802 => x"00000000",
    25803 => x"00000000", 25804 => x"00000000", 25805 => x"00000000",
    25806 => x"00000000", 25807 => x"00000000", 25808 => x"00000000",
    25809 => x"00000000", 25810 => x"00000000", 25811 => x"00000000",
    25812 => x"00000000", 25813 => x"00000000", 25814 => x"00000000",
    25815 => x"00000000", 25816 => x"00000000", 25817 => x"00000000",
    25818 => x"00000000", 25819 => x"00000000", 25820 => x"00000000",
    25821 => x"00000000", 25822 => x"00000000", 25823 => x"00000000",
    25824 => x"00000000", 25825 => x"00000000", 25826 => x"00000000",
    25827 => x"00000000", 25828 => x"00000000", 25829 => x"00000000",
    25830 => x"00000000", 25831 => x"00000000", 25832 => x"00000000",
    25833 => x"00000000", 25834 => x"00000000", 25835 => x"00000000",
    25836 => x"00000000", 25837 => x"00000000", 25838 => x"00000000",
    25839 => x"00000000", 25840 => x"00000000", 25841 => x"00000000",
    25842 => x"00000000", 25843 => x"00000000", 25844 => x"00000000",
    25845 => x"00000000", 25846 => x"00000000", 25847 => x"00000000",
    25848 => x"00000000", 25849 => x"00000000", 25850 => x"00000000",
    25851 => x"00000000", 25852 => x"00000000", 25853 => x"00000000",
    25854 => x"00000000", 25855 => x"00000000", 25856 => x"00000000",
    25857 => x"00000000", 25858 => x"00000000", 25859 => x"00000000",
    25860 => x"00000000", 25861 => x"00000000", 25862 => x"00000000",
    25863 => x"00000000", 25864 => x"00000000", 25865 => x"00000000",
    25866 => x"00000000", 25867 => x"00000000", 25868 => x"00000000",
    25869 => x"00000000", 25870 => x"00000000", 25871 => x"00000000",
    25872 => x"00000000", 25873 => x"00000000", 25874 => x"00000000",
    25875 => x"00000000", 25876 => x"00000000", 25877 => x"00000000",
    25878 => x"00000000", 25879 => x"00000000", 25880 => x"00000000",
    25881 => x"00000000", 25882 => x"00000000", 25883 => x"00000000",
    25884 => x"00000000", 25885 => x"00000000", 25886 => x"00000000",
    25887 => x"00000000", 25888 => x"00000000", 25889 => x"00000000",
    25890 => x"00000000", 25891 => x"00000000", 25892 => x"00000000",
    25893 => x"00000000", 25894 => x"00000000", 25895 => x"00000000",
    25896 => x"00000000", 25897 => x"00000000", 25898 => x"00000000",
    25899 => x"00000000", 25900 => x"00000000", 25901 => x"00000000",
    25902 => x"00000000", 25903 => x"00000000", 25904 => x"00000000",
    25905 => x"00000000", 25906 => x"00000000", 25907 => x"00000000",
    25908 => x"00000000", 25909 => x"00000000", 25910 => x"00000000",
    25911 => x"00000000", 25912 => x"00000000", 25913 => x"00000000",
    25914 => x"00000000", 25915 => x"00000000", 25916 => x"00000000",
    25917 => x"00000000", 25918 => x"00000000", 25919 => x"00000000",
    25920 => x"00000000", 25921 => x"00000000", 25922 => x"00000000",
    25923 => x"00000000", 25924 => x"00000000", 25925 => x"00000000",
    25926 => x"00000000", 25927 => x"00000000", 25928 => x"00000000",
    25929 => x"00000000", 25930 => x"00000000", 25931 => x"00000000",
    25932 => x"00000000", 25933 => x"00000000", 25934 => x"00000000",
    25935 => x"00000000", 25936 => x"00000000", 25937 => x"00000000",
    25938 => x"00000000", 25939 => x"00000000", 25940 => x"00000000",
    25941 => x"00000000", 25942 => x"00000000", 25943 => x"00000000",
    25944 => x"00000000", 25945 => x"00000000", 25946 => x"00000000",
    25947 => x"00000000", 25948 => x"00000000", 25949 => x"00000000",
    25950 => x"00000000", 25951 => x"00000000", 25952 => x"00000000",
    25953 => x"00000000", 25954 => x"00000000", 25955 => x"00000000",
    25956 => x"00000000", 25957 => x"00000000", 25958 => x"00000000",
    25959 => x"00000000", 25960 => x"00000000", 25961 => x"00000000",
    25962 => x"00000000", 25963 => x"00000000", 25964 => x"00000000",
    25965 => x"00000000", 25966 => x"00000000", 25967 => x"00000000",
    25968 => x"00000000", 25969 => x"00000000", 25970 => x"00000000",
    25971 => x"00000000", 25972 => x"00000000", 25973 => x"00000000",
    25974 => x"00000000", 25975 => x"00000000", 25976 => x"00000000",
    25977 => x"00000000", 25978 => x"00000000", 25979 => x"00000000",
    25980 => x"00000000", 25981 => x"00000000", 25982 => x"00000000",
    25983 => x"00000000", 25984 => x"00000000", 25985 => x"00000000",
    25986 => x"00000000", 25987 => x"00000000", 25988 => x"00000000",
    25989 => x"00000000", 25990 => x"00000000", 25991 => x"00000000",
    25992 => x"00000000", 25993 => x"00000000", 25994 => x"00000000",
    25995 => x"00000000", 25996 => x"00000000", 25997 => x"00000000",
    25998 => x"00000000", 25999 => x"00000000", 26000 => x"00000000",
    26001 => x"00000000", 26002 => x"00000000", 26003 => x"00000000",
    26004 => x"00000000", 26005 => x"00000000", 26006 => x"00000000",
    26007 => x"00000000", 26008 => x"00000000", 26009 => x"00000000",
    26010 => x"00000000", 26011 => x"00000000", 26012 => x"00000000",
    26013 => x"00000000", 26014 => x"00000000", 26015 => x"00000000",
    26016 => x"00000000", 26017 => x"00000000", 26018 => x"00000000",
    26019 => x"00000000", 26020 => x"00000000", 26021 => x"00000000",
    26022 => x"00000000", 26023 => x"00000000", 26024 => x"00000000",
    26025 => x"00000000", 26026 => x"00000000", 26027 => x"00000000",
    26028 => x"00000000", 26029 => x"00000000", 26030 => x"00000000",
    26031 => x"00000000", 26032 => x"00000000", 26033 => x"00000000",
    26034 => x"00000000", 26035 => x"00000000", 26036 => x"00000000",
    26037 => x"00000000", 26038 => x"00000000", 26039 => x"00000000",
    26040 => x"00000000", 26041 => x"00000000", 26042 => x"00000000",
    26043 => x"00000000", 26044 => x"00000000", 26045 => x"00000000",
    26046 => x"00000000", 26047 => x"00000000", 26048 => x"00000000",
    26049 => x"00000000", 26050 => x"00000000", 26051 => x"00000000",
    26052 => x"00000000", 26053 => x"00000000", 26054 => x"00000000",
    26055 => x"00000000", 26056 => x"00000000", 26057 => x"00000000",
    26058 => x"00000000", 26059 => x"00000000", 26060 => x"00000000",
    26061 => x"00000000", 26062 => x"00000000", 26063 => x"00000000",
    26064 => x"00000000", 26065 => x"00000000", 26066 => x"00000000",
    26067 => x"00000000", 26068 => x"00000000", 26069 => x"00000000",
    26070 => x"00000000", 26071 => x"00000000", 26072 => x"00000000",
    26073 => x"00000000", 26074 => x"00000000", 26075 => x"00000000",
    26076 => x"00000000", 26077 => x"00000000", 26078 => x"00000000",
    26079 => x"00000000", 26080 => x"00000000", 26081 => x"00000000",
    26082 => x"00000000", 26083 => x"00000000", 26084 => x"00000000",
    26085 => x"00000000", 26086 => x"00000000", 26087 => x"00000000",
    26088 => x"00000000", 26089 => x"00000000", 26090 => x"00000000",
    26091 => x"00000000", 26092 => x"00000000", 26093 => x"00000000",
    26094 => x"00000000", 26095 => x"00000000", 26096 => x"00000000",
    26097 => x"00000000", 26098 => x"00000000", 26099 => x"00000000",
    26100 => x"00000000", 26101 => x"00000000", 26102 => x"00000000",
    26103 => x"00000000", 26104 => x"00000000", 26105 => x"00000000",
    26106 => x"00000000", 26107 => x"00000000", 26108 => x"00000000",
    26109 => x"00000000", 26110 => x"00000000", 26111 => x"00000000",
    26112 => x"00000000", 26113 => x"00000000", 26114 => x"00000000",
    26115 => x"00000000", 26116 => x"00000000", 26117 => x"00000000",
    26118 => x"00000000", 26119 => x"00000000", 26120 => x"00000000",
    26121 => x"00000000", 26122 => x"00000000", 26123 => x"00000000",
    26124 => x"00000000", 26125 => x"00000000", 26126 => x"00000000",
    26127 => x"00000000", 26128 => x"00000000", 26129 => x"00000000",
    26130 => x"00000000", 26131 => x"00000000", 26132 => x"00000000",
    26133 => x"00000000", 26134 => x"00000000", 26135 => x"00000000",
    26136 => x"00000000", 26137 => x"00000000", 26138 => x"00000000",
    26139 => x"00000000", 26140 => x"00000000", 26141 => x"00000000",
    26142 => x"00000000", 26143 => x"00000000", 26144 => x"00000000",
    26145 => x"00000000", 26146 => x"00000000", 26147 => x"00000000",
    26148 => x"00000000", 26149 => x"00000000", 26150 => x"00000000",
    26151 => x"00000000", 26152 => x"00000000", 26153 => x"00000000",
    26154 => x"00000000", 26155 => x"00000000", 26156 => x"00000000",
    26157 => x"00000000", 26158 => x"00000000", 26159 => x"00000000",
    26160 => x"00000000", 26161 => x"00000000", 26162 => x"00000000",
    26163 => x"00000000", 26164 => x"00000000", 26165 => x"00000000",
    26166 => x"00000000", 26167 => x"00000000", 26168 => x"00000000",
    26169 => x"00000000", 26170 => x"00000000", 26171 => x"00000000",
    26172 => x"00000000", 26173 => x"00000000", 26174 => x"00000000",
    26175 => x"00000000", 26176 => x"00000000", 26177 => x"00000000",
    26178 => x"00000000", 26179 => x"00000000", 26180 => x"00000000",
    26181 => x"00000000", 26182 => x"00000000", 26183 => x"00000000",
    26184 => x"00000000", 26185 => x"00000000", 26186 => x"00000000",
    26187 => x"00000000", 26188 => x"00000000", 26189 => x"00000000",
    26190 => x"00000000", 26191 => x"00000000", 26192 => x"00000000",
    26193 => x"00000000", 26194 => x"00000000", 26195 => x"00000000",
    26196 => x"00000000", 26197 => x"00000000", 26198 => x"00000000",
    26199 => x"00000000", 26200 => x"00000000", 26201 => x"00000000",
    26202 => x"00000000", 26203 => x"00000000", 26204 => x"00000000",
    26205 => x"00000000", 26206 => x"00000000", 26207 => x"00000000",
    26208 => x"00000000", 26209 => x"00000000", 26210 => x"00000000",
    26211 => x"00000000", 26212 => x"00000000", 26213 => x"00000000",
    26214 => x"00000000", 26215 => x"00000000", 26216 => x"00000000",
    26217 => x"00000000", 26218 => x"00000000", 26219 => x"00000000",
    26220 => x"00000000", 26221 => x"00000000", 26222 => x"00000000",
    26223 => x"00000000", 26224 => x"00000000", 26225 => x"00000000",
    26226 => x"00000000", 26227 => x"00000000", 26228 => x"00000000",
    26229 => x"00000000", 26230 => x"00000000", 26231 => x"00000000",
    26232 => x"00000000", 26233 => x"00000000", 26234 => x"00000000",
    26235 => x"00000000", 26236 => x"00000000", 26237 => x"00000000",
    26238 => x"00000000", 26239 => x"00000000", 26240 => x"00000000",
    26241 => x"00000000", 26242 => x"00000000", 26243 => x"00000000",
    26244 => x"00000000", 26245 => x"00000000", 26246 => x"00000000",
    26247 => x"00000000", 26248 => x"00000000", 26249 => x"00000000",
    26250 => x"00000000", 26251 => x"00000000", 26252 => x"00000000",
    26253 => x"00000000", 26254 => x"00000000", 26255 => x"00000000",
    26256 => x"00000000", 26257 => x"00000000", 26258 => x"00000000",
    26259 => x"00000000", 26260 => x"00000000", 26261 => x"00000000",
    26262 => x"00000000", 26263 => x"00000000", 26264 => x"00000000",
    26265 => x"00000000", 26266 => x"00000000", 26267 => x"00000000",
    26268 => x"00000000", 26269 => x"00000000", 26270 => x"00000000",
    26271 => x"00000000", 26272 => x"00000000", 26273 => x"00000000",
    26274 => x"00000000", 26275 => x"00000000", 26276 => x"00000000",
    26277 => x"00000000", 26278 => x"00000000", 26279 => x"00000000",
    26280 => x"00000000", 26281 => x"00000000", 26282 => x"00000000",
    26283 => x"00000000", 26284 => x"00000000", 26285 => x"00000000",
    26286 => x"00000000", 26287 => x"00000000", 26288 => x"00000000",
    26289 => x"00000000", 26290 => x"00000000", 26291 => x"00000000",
    26292 => x"00000000", 26293 => x"00000000", 26294 => x"00000000",
    26295 => x"00000000", 26296 => x"00000000", 26297 => x"00000000",
    26298 => x"00000000", 26299 => x"00000000", 26300 => x"00000000",
    26301 => x"00000000", 26302 => x"00000000", 26303 => x"00000000",
    26304 => x"00000000", 26305 => x"00000000", 26306 => x"00000000",
    26307 => x"00000000", 26308 => x"00000000", 26309 => x"00000000",
    26310 => x"00000000", 26311 => x"00000000", 26312 => x"00000000",
    26313 => x"00000000", 26314 => x"00000000", 26315 => x"00000000",
    26316 => x"00000000", 26317 => x"00000000", 26318 => x"00000000",
    26319 => x"00000000", 26320 => x"00000000", 26321 => x"00000000",
    26322 => x"00000000", 26323 => x"00000000", 26324 => x"00000000",
    26325 => x"00000000", 26326 => x"00000000", 26327 => x"00000000",
    26328 => x"00000000", 26329 => x"00000000", 26330 => x"00000000",
    26331 => x"00000000", 26332 => x"00000000", 26333 => x"00000000",
    26334 => x"00000000", 26335 => x"00000000", 26336 => x"00000000",
    26337 => x"00000000", 26338 => x"00000000", 26339 => x"00000000",
    26340 => x"00000000", 26341 => x"00000000", 26342 => x"00000000",
    26343 => x"00000000", 26344 => x"00000000", 26345 => x"00000000",
    26346 => x"00000000", 26347 => x"00000000", 26348 => x"00000000",
    26349 => x"00000000", 26350 => x"00000000", 26351 => x"00000000",
    26352 => x"00000000", 26353 => x"00000000", 26354 => x"00000000",
    26355 => x"00000000", 26356 => x"00000000", 26357 => x"00000000",
    26358 => x"00000000", 26359 => x"00000000", 26360 => x"00000000",
    26361 => x"00000000", 26362 => x"00000000", 26363 => x"00000000",
    26364 => x"00000000", 26365 => x"00000000", 26366 => x"00000000",
    26367 => x"00000000", 26368 => x"00000000", 26369 => x"00000000",
    26370 => x"00000000", 26371 => x"00000000", 26372 => x"00000000",
    26373 => x"00000000", 26374 => x"00000000", 26375 => x"00000000",
    26376 => x"00000000", 26377 => x"00000000", 26378 => x"00000000",
    26379 => x"00000000", 26380 => x"00000000", 26381 => x"00000000",
    26382 => x"00000000", 26383 => x"00000000", 26384 => x"00000000",
    26385 => x"00000000", 26386 => x"00000000", 26387 => x"00000000",
    26388 => x"00000000", 26389 => x"00000000", 26390 => x"00000000",
    26391 => x"00000000", 26392 => x"00000000", 26393 => x"00000000",
    26394 => x"00000000", 26395 => x"00000000", 26396 => x"00000000",
    26397 => x"00000000", 26398 => x"00000000", 26399 => x"00000000",
    26400 => x"00000000", 26401 => x"00000000", 26402 => x"00000000",
    26403 => x"00000000", 26404 => x"00000000", 26405 => x"00000000",
    26406 => x"00000000", 26407 => x"00000000", 26408 => x"00000000",
    26409 => x"00000000", 26410 => x"00000000", 26411 => x"00000000",
    26412 => x"00000000", 26413 => x"00000000", 26414 => x"00000000",
    26415 => x"00000000", 26416 => x"00000000", 26417 => x"00000000",
    26418 => x"00000000", 26419 => x"00000000", 26420 => x"00000000",
    26421 => x"00000000", 26422 => x"00000000", 26423 => x"00000000",
    26424 => x"00000000", 26425 => x"00000000", 26426 => x"00000000",
    26427 => x"00000000", 26428 => x"00000000", 26429 => x"00000000",
    26430 => x"00000000", 26431 => x"00000000", 26432 => x"00000000",
    26433 => x"00000000", 26434 => x"00000000", 26435 => x"00000000",
    26436 => x"00000000", 26437 => x"00000000", 26438 => x"00000000",
    26439 => x"00000000", 26440 => x"00000000", 26441 => x"00000000",
    26442 => x"00000000", 26443 => x"00000000", 26444 => x"00000000",
    26445 => x"00000000", 26446 => x"00000000", 26447 => x"00000000",
    26448 => x"00000000", 26449 => x"00000000", 26450 => x"00000000",
    26451 => x"00000000", 26452 => x"00000000", 26453 => x"00000000",
    26454 => x"00000000", 26455 => x"00000000", 26456 => x"00000000",
    26457 => x"00000000", 26458 => x"00000000", 26459 => x"00000000",
    26460 => x"00000000", 26461 => x"00000000", 26462 => x"00000000",
    26463 => x"00000000", 26464 => x"00000000", 26465 => x"00000000",
    26466 => x"00000000", 26467 => x"00000000", 26468 => x"00000000",
    26469 => x"00000000", 26470 => x"00000000", 26471 => x"00000000",
    26472 => x"00000000", 26473 => x"00000000", 26474 => x"00000000",
    26475 => x"00000000", 26476 => x"00000000", 26477 => x"00000000",
    26478 => x"00000000", 26479 => x"00000000", 26480 => x"00000000",
    26481 => x"00000000", 26482 => x"00000000", 26483 => x"00000000",
    26484 => x"00000000", 26485 => x"00000000", 26486 => x"00000000",
    26487 => x"00000000", 26488 => x"00000000", 26489 => x"00000000",
    26490 => x"00000000", 26491 => x"00000000", 26492 => x"00000000",
    26493 => x"00000000", 26494 => x"00000000", 26495 => x"00000000",
    26496 => x"00000000", 26497 => x"00000000", 26498 => x"00000000",
    26499 => x"00000000", 26500 => x"00000000", 26501 => x"00000000",
    26502 => x"00000000", 26503 => x"00000000", 26504 => x"00000000",
    26505 => x"00000000", 26506 => x"00000000", 26507 => x"00000000",
    26508 => x"00000000", 26509 => x"00000000", 26510 => x"00000000",
    26511 => x"00000000", 26512 => x"00000000", 26513 => x"00000000",
    26514 => x"00000000", 26515 => x"00000000", 26516 => x"00000000",
    26517 => x"00000000", 26518 => x"00000000", 26519 => x"00000000",
    26520 => x"00000000", 26521 => x"00000000", 26522 => x"00000000",
    26523 => x"00000000", 26524 => x"00000000", 26525 => x"00000000",
    26526 => x"00000000", 26527 => x"00000000", 26528 => x"00000000",
    26529 => x"00000000", 26530 => x"00000000", 26531 => x"00000000",
    26532 => x"00000000", 26533 => x"00000000", 26534 => x"00000000",
    26535 => x"00000000", 26536 => x"00000000", 26537 => x"00000000",
    26538 => x"00000000", 26539 => x"00000000", 26540 => x"00000000",
    26541 => x"00000000", 26542 => x"00000000", 26543 => x"00000000",
    26544 => x"00000000", 26545 => x"00000000", 26546 => x"00000000",
    26547 => x"00000000", 26548 => x"00000000", 26549 => x"00000000",
    26550 => x"00000000", 26551 => x"00000000", 26552 => x"00000000",
    26553 => x"00000000", 26554 => x"00000000", 26555 => x"00000000",
    26556 => x"00000000", 26557 => x"00000000", 26558 => x"00000000",
    26559 => x"00000000", 26560 => x"00000000", 26561 => x"00000000",
    26562 => x"00000000", 26563 => x"00000000", 26564 => x"00000000",
    26565 => x"00000000", 26566 => x"00000000", 26567 => x"00000000",
    26568 => x"00000000", 26569 => x"00000000", 26570 => x"00000000",
    26571 => x"00000000", 26572 => x"00000000", 26573 => x"00000000",
    26574 => x"00000000", 26575 => x"00000000", 26576 => x"00000000",
    26577 => x"00000000", 26578 => x"00000000", 26579 => x"00000000",
    26580 => x"00000000", 26581 => x"00000000", 26582 => x"00000000",
    26583 => x"00000000", 26584 => x"00000000", 26585 => x"00000000",
    26586 => x"00000000", 26587 => x"00000000", 26588 => x"00000000",
    26589 => x"00000000", 26590 => x"00000000", 26591 => x"00000000",
    26592 => x"00000000", 26593 => x"00000000", 26594 => x"00000000",
    26595 => x"00000000", 26596 => x"00000000", 26597 => x"00000000",
    26598 => x"00000000", 26599 => x"00000000", 26600 => x"00000000",
    26601 => x"00000000", 26602 => x"00000000", 26603 => x"00000000",
    26604 => x"00000000", 26605 => x"00000000", 26606 => x"00000000",
    26607 => x"00000000", 26608 => x"00000000", 26609 => x"00000000",
    26610 => x"00000000", 26611 => x"00000000", 26612 => x"00000000",
    26613 => x"00000000", 26614 => x"00000000", 26615 => x"00000000",
    26616 => x"00000000", 26617 => x"00000000", 26618 => x"00000000",
    26619 => x"00000000", 26620 => x"00000000", 26621 => x"00000000",
    26622 => x"00000000", 26623 => x"00000000", 26624 => x"00000000",
    26625 => x"00000000", 26626 => x"00000000", 26627 => x"00000000",
    26628 => x"00000000", 26629 => x"00000000", 26630 => x"00000000",
    26631 => x"00000000", 26632 => x"00000000", 26633 => x"00000000",
    26634 => x"00000000", 26635 => x"00000000", 26636 => x"00000000",
    26637 => x"00000000", 26638 => x"00000000", 26639 => x"00000000",
    26640 => x"00000000", 26641 => x"00000000", 26642 => x"00000000",
    26643 => x"00000000", 26644 => x"00000000", 26645 => x"00000000",
    26646 => x"00000000", 26647 => x"00000000", 26648 => x"00000000",
    26649 => x"00000000", 26650 => x"00000000", 26651 => x"00000000",
    26652 => x"00000000", 26653 => x"00000000", 26654 => x"00000000",
    26655 => x"00000000", 26656 => x"00000000", 26657 => x"00000000",
    26658 => x"00000000", 26659 => x"00000000", 26660 => x"00000000",
    26661 => x"00000000", 26662 => x"00000000", 26663 => x"00000000",
    26664 => x"00000000", 26665 => x"00000000", 26666 => x"00000000",
    26667 => x"00000000", 26668 => x"00000000", 26669 => x"00000000",
    26670 => x"00000000", 26671 => x"00000000", 26672 => x"00000000",
    26673 => x"00000000", 26674 => x"00000000", 26675 => x"00000000",
    26676 => x"00000000", 26677 => x"00000000", 26678 => x"00000000",
    26679 => x"00000000", 26680 => x"00000000", 26681 => x"00000000",
    26682 => x"00000000", 26683 => x"00000000", 26684 => x"00000000",
    26685 => x"00000000", 26686 => x"00000000", 26687 => x"00000000",
    26688 => x"00000000", 26689 => x"00000000", 26690 => x"00000000",
    26691 => x"00000000", 26692 => x"00000000", 26693 => x"00000000",
    26694 => x"00000000", 26695 => x"00000000", 26696 => x"00000000",
    26697 => x"00000000", 26698 => x"00000000", 26699 => x"00000000",
    26700 => x"00000000", 26701 => x"00000000", 26702 => x"00000000",
    26703 => x"00000000", 26704 => x"00000000", 26705 => x"00000000",
    26706 => x"00000000", 26707 => x"00000000", 26708 => x"00000000",
    26709 => x"00000000", 26710 => x"00000000", 26711 => x"00000000",
    26712 => x"00000000", 26713 => x"00000000", 26714 => x"00000000",
    26715 => x"00000000", 26716 => x"00000000", 26717 => x"00000000",
    26718 => x"00000000", 26719 => x"00000000", 26720 => x"00000000",
    26721 => x"00000000", 26722 => x"00000000", 26723 => x"00000000",
    26724 => x"00000000", 26725 => x"00000000", 26726 => x"00000000",
    26727 => x"00000000", 26728 => x"00000000", 26729 => x"00000000",
    26730 => x"00000000", 26731 => x"00000000", 26732 => x"00000000",
    26733 => x"00000000", 26734 => x"00000000", 26735 => x"00000000",
    26736 => x"00000000", 26737 => x"00000000", 26738 => x"00000000",
    26739 => x"00000000", 26740 => x"00000000", 26741 => x"00000000",
    26742 => x"00000000", 26743 => x"00000000", 26744 => x"00000000",
    26745 => x"00000000", 26746 => x"00000000", 26747 => x"00000000",
    26748 => x"00000000", 26749 => x"00000000", 26750 => x"00000000",
    26751 => x"00000000", 26752 => x"00000000", 26753 => x"00000000",
    26754 => x"00000000", 26755 => x"00000000", 26756 => x"00000000",
    26757 => x"00000000", 26758 => x"00000000", 26759 => x"00000000",
    26760 => x"00000000", 26761 => x"00000000", 26762 => x"00000000",
    26763 => x"00000000", 26764 => x"00000000", 26765 => x"00000000",
    26766 => x"00000000", 26767 => x"00000000", 26768 => x"00000000",
    26769 => x"00000000", 26770 => x"00000000", 26771 => x"00000000",
    26772 => x"00000000", 26773 => x"00000000", 26774 => x"00000000",
    26775 => x"00000000", 26776 => x"00000000", 26777 => x"00000000",
    26778 => x"00000000", 26779 => x"00000000", 26780 => x"00000000",
    26781 => x"00000000", 26782 => x"00000000", 26783 => x"00000000",
    26784 => x"00000000", 26785 => x"00000000", 26786 => x"00000000",
    26787 => x"00000000", 26788 => x"00000000", 26789 => x"00000000",
    26790 => x"00000000", 26791 => x"00000000", 26792 => x"00000000",
    26793 => x"00000000", 26794 => x"00000000", 26795 => x"00000000",
    26796 => x"00000000", 26797 => x"00000000", 26798 => x"00000000",
    26799 => x"00000000", 26800 => x"00000000", 26801 => x"00000000",
    26802 => x"00000000", 26803 => x"00000000", 26804 => x"00000000",
    26805 => x"00000000", 26806 => x"00000000", 26807 => x"00000000",
    26808 => x"00000000", 26809 => x"00000000", 26810 => x"00000000",
    26811 => x"00000000", 26812 => x"00000000", 26813 => x"00000000",
    26814 => x"00000000", 26815 => x"00000000", 26816 => x"00000000",
    26817 => x"00000000", 26818 => x"00000000", 26819 => x"00000000",
    26820 => x"00000000", 26821 => x"00000000", 26822 => x"00000000",
    26823 => x"00000000", 26824 => x"00000000", 26825 => x"00000000",
    26826 => x"00000000", 26827 => x"00000000", 26828 => x"00000000",
    26829 => x"00000000", 26830 => x"00000000", 26831 => x"00000000",
    26832 => x"00000000", 26833 => x"00000000", 26834 => x"00000000",
    26835 => x"00000000", 26836 => x"00000000", 26837 => x"00000000",
    26838 => x"00000000", 26839 => x"00000000", 26840 => x"00000000",
    26841 => x"00000000", 26842 => x"00000000", 26843 => x"00000000",
    26844 => x"00000000", 26845 => x"00000000", 26846 => x"00000000",
    26847 => x"00000000", 26848 => x"00000000", 26849 => x"00000000",
    26850 => x"00000000", 26851 => x"00000000", 26852 => x"00000000",
    26853 => x"00000000", 26854 => x"00000000", 26855 => x"00000000",
    26856 => x"00000000", 26857 => x"00000000", 26858 => x"00000000",
    26859 => x"00000000", 26860 => x"00000000", 26861 => x"00000000",
    26862 => x"00000000", 26863 => x"00000000", 26864 => x"00000000",
    26865 => x"00000000", 26866 => x"00000000", 26867 => x"00000000",
    26868 => x"00000000", 26869 => x"00000000", 26870 => x"00000000",
    26871 => x"00000000", 26872 => x"00000000", 26873 => x"00000000",
    26874 => x"00000000", 26875 => x"00000000", 26876 => x"00000000",
    26877 => x"00000000", 26878 => x"00000000", 26879 => x"00000000",
    26880 => x"00000000", 26881 => x"00000000", 26882 => x"00000000",
    26883 => x"00000000", 26884 => x"00000000", 26885 => x"00000000",
    26886 => x"00000000", 26887 => x"00000000", 26888 => x"00000000",
    26889 => x"00000000", 26890 => x"00000000", 26891 => x"00000000",
    26892 => x"00000000", 26893 => x"00000000", 26894 => x"00000000",
    26895 => x"00000000", 26896 => x"00000000", 26897 => x"00000000",
    26898 => x"00000000", 26899 => x"00000000", 26900 => x"00000000",
    26901 => x"00000000", 26902 => x"00000000", 26903 => x"00000000",
    26904 => x"00000000", 26905 => x"00000000", 26906 => x"00000000",
    26907 => x"00000000", 26908 => x"00000000", 26909 => x"00000000",
    26910 => x"00000000", 26911 => x"00000000", 26912 => x"00000000",
    26913 => x"00000000", 26914 => x"00000000", 26915 => x"00000000",
    26916 => x"00000000", 26917 => x"00000000", 26918 => x"00000000",
    26919 => x"00000000", 26920 => x"00000000", 26921 => x"00000000",
    26922 => x"00000000", 26923 => x"00000000", 26924 => x"00000000",
    26925 => x"00000000", 26926 => x"00000000", 26927 => x"00000000",
    26928 => x"00000000", 26929 => x"00000000", 26930 => x"00000000",
    26931 => x"00000000", 26932 => x"00000000", 26933 => x"00000000",
    26934 => x"00000000", 26935 => x"00000000", 26936 => x"00000000",
    26937 => x"00000000", 26938 => x"00000000", 26939 => x"00000000",
    26940 => x"00000000", 26941 => x"00000000", 26942 => x"00000000",
    26943 => x"00000000", 26944 => x"00000000", 26945 => x"00000000",
    26946 => x"00000000", 26947 => x"00000000", 26948 => x"00000000",
    26949 => x"00000000", 26950 => x"00000000", 26951 => x"00000000",
    26952 => x"00000000", 26953 => x"00000000", 26954 => x"00000000",
    26955 => x"00000000", 26956 => x"00000000", 26957 => x"00000000",
    26958 => x"00000000", 26959 => x"00000000", 26960 => x"00000000",
    26961 => x"00000000", 26962 => x"00000000", 26963 => x"00000000",
    26964 => x"00000000", 26965 => x"00000000", 26966 => x"00000000",
    26967 => x"00000000", 26968 => x"00000000", 26969 => x"00000000",
    26970 => x"00000000", 26971 => x"00000000", 26972 => x"00000000",
    26973 => x"00000000", 26974 => x"00000000", 26975 => x"00000000",
    26976 => x"00000000", 26977 => x"00000000", 26978 => x"00000000",
    26979 => x"00000000", 26980 => x"00000000", 26981 => x"00000000",
    26982 => x"00000000", 26983 => x"00000000", 26984 => x"00000000",
    26985 => x"00000000", 26986 => x"00000000", 26987 => x"00000000",
    26988 => x"00000000", 26989 => x"00000000", 26990 => x"00000000",
    26991 => x"00000000", 26992 => x"00000000", 26993 => x"00000000",
    26994 => x"00000000", 26995 => x"00000000", 26996 => x"00000000",
    26997 => x"00000000", 26998 => x"00000000", 26999 => x"00000000",
    27000 => x"00000000", 27001 => x"00000000", 27002 => x"00000000",
    27003 => x"00000000", 27004 => x"00000000", 27005 => x"00000000",
    27006 => x"00000000", 27007 => x"00000000", 27008 => x"00000000",
    27009 => x"00000000", 27010 => x"00000000", 27011 => x"00000000",
    27012 => x"00000000", 27013 => x"00000000", 27014 => x"00000000",
    27015 => x"00000000", 27016 => x"00000000", 27017 => x"00000000",
    27018 => x"00000000", 27019 => x"00000000", 27020 => x"00000000",
    27021 => x"00000000", 27022 => x"00000000", 27023 => x"00000000",
    27024 => x"00000000", 27025 => x"00000000", 27026 => x"00000000",
    27027 => x"00000000", 27028 => x"00000000", 27029 => x"00000000",
    27030 => x"00000000", 27031 => x"00000000", 27032 => x"00000000",
    27033 => x"00000000", 27034 => x"00000000", 27035 => x"00000000",
    27036 => x"00000000", 27037 => x"00000000", 27038 => x"00000000",
    27039 => x"00000000", 27040 => x"00000000", 27041 => x"00000000",
    27042 => x"00000000", 27043 => x"00000000", 27044 => x"00000000",
    27045 => x"00000000", 27046 => x"00000000", 27047 => x"00000000",
    27048 => x"00000000", 27049 => x"00000000", 27050 => x"00000000",
    27051 => x"00000000", 27052 => x"00000000", 27053 => x"00000000",
    27054 => x"00000000", 27055 => x"00000000", 27056 => x"00000000",
    27057 => x"00000000", 27058 => x"00000000", 27059 => x"00000000",
    27060 => x"00000000", 27061 => x"00000000", 27062 => x"00000000",
    27063 => x"00000000", 27064 => x"00000000", 27065 => x"00000000",
    27066 => x"00000000", 27067 => x"00000000", 27068 => x"00000000",
    27069 => x"00000000", 27070 => x"00000000", 27071 => x"00000000",
    27072 => x"00000000", 27073 => x"00000000", 27074 => x"00000000",
    27075 => x"00000000", 27076 => x"00000000", 27077 => x"00000000",
    27078 => x"00000000", 27079 => x"00000000", 27080 => x"00000000",
    27081 => x"00000000", 27082 => x"00000000", 27083 => x"00000000",
    27084 => x"00000000", 27085 => x"00000000", 27086 => x"00000000",
    27087 => x"00000000", 27088 => x"00000000", 27089 => x"00000000",
    27090 => x"00000000", 27091 => x"00000000", 27092 => x"00000000",
    27093 => x"00000000", 27094 => x"00000000", 27095 => x"00000000",
    27096 => x"00000000", 27097 => x"00000000", 27098 => x"00000000",
    27099 => x"00000000", 27100 => x"00000000", 27101 => x"00000000",
    27102 => x"00000000", 27103 => x"00000000", 27104 => x"00000000",
    27105 => x"00000000", 27106 => x"00000000", 27107 => x"00000000",
    27108 => x"00000000", 27109 => x"00000000", 27110 => x"00000000",
    27111 => x"00000000", 27112 => x"00000000", 27113 => x"00000000",
    27114 => x"00000000", 27115 => x"00000000", 27116 => x"00000000",
    27117 => x"00000000", 27118 => x"00000000", 27119 => x"00000000",
    27120 => x"00000000", 27121 => x"00000000", 27122 => x"00000000",
    27123 => x"00000000", 27124 => x"00000000", 27125 => x"00000000",
    27126 => x"00000000", 27127 => x"00000000", 27128 => x"00000000",
    27129 => x"00000000", 27130 => x"00000000", 27131 => x"00000000",
    27132 => x"00000000", 27133 => x"00000000", 27134 => x"00000000",
    27135 => x"00000000", 27136 => x"00000000", 27137 => x"00000000",
    27138 => x"00000000", 27139 => x"00000000", 27140 => x"00000000",
    27141 => x"00000000", 27142 => x"00000000", 27143 => x"00000000",
    27144 => x"00000000", 27145 => x"00000000", 27146 => x"00000000",
    27147 => x"00000000", 27148 => x"00000000", 27149 => x"00000000",
    27150 => x"00000000", 27151 => x"00000000", 27152 => x"00000000",
    27153 => x"00000000", 27154 => x"00000000", 27155 => x"00000000",
    27156 => x"00000000", 27157 => x"00000000", 27158 => x"00000000",
    27159 => x"00000000", 27160 => x"00000000", 27161 => x"00000000",
    27162 => x"00000000", 27163 => x"00000000", 27164 => x"00000000",
    27165 => x"00000000", 27166 => x"00000000", 27167 => x"00000000",
    27168 => x"00000000", 27169 => x"00000000", 27170 => x"00000000",
    27171 => x"00000000", 27172 => x"00000000", 27173 => x"00000000",
    27174 => x"00000000", 27175 => x"00000000", 27176 => x"00000000",
    27177 => x"00000000", 27178 => x"00000000", 27179 => x"00000000",
    27180 => x"00000000", 27181 => x"00000000", 27182 => x"00000000",
    27183 => x"00000000", 27184 => x"00000000", 27185 => x"00000000",
    27186 => x"00000000", 27187 => x"00000000", 27188 => x"00000000",
    27189 => x"00000000", 27190 => x"00000000", 27191 => x"00000000",
    27192 => x"00000000", 27193 => x"00000000", 27194 => x"00000000",
    27195 => x"00000000", 27196 => x"00000000", 27197 => x"00000000",
    27198 => x"00000000", 27199 => x"00000000", 27200 => x"00000000",
    27201 => x"00000000", 27202 => x"00000000", 27203 => x"00000000",
    27204 => x"00000000", 27205 => x"00000000", 27206 => x"00000000",
    27207 => x"00000000", 27208 => x"00000000", 27209 => x"00000000",
    27210 => x"00000000", 27211 => x"00000000", 27212 => x"00000000",
    27213 => x"00000000", 27214 => x"00000000", 27215 => x"00000000",
    27216 => x"00000000", 27217 => x"00000000", 27218 => x"00000000",
    27219 => x"00000000", 27220 => x"00000000", 27221 => x"00000000",
    27222 => x"00000000", 27223 => x"00000000", 27224 => x"00000000",
    27225 => x"00000000", 27226 => x"00000000", 27227 => x"00000000",
    27228 => x"00000000", 27229 => x"00000000", 27230 => x"00000000",
    27231 => x"00000000", 27232 => x"00000000", 27233 => x"00000000",
    27234 => x"00000000", 27235 => x"00000000", 27236 => x"00000000",
    27237 => x"00000000", 27238 => x"00000000", 27239 => x"00000000",
    27240 => x"00000000", 27241 => x"00000000", 27242 => x"00000000",
    27243 => x"00000000", 27244 => x"00000000", 27245 => x"00000000",
    27246 => x"00000000", 27247 => x"00000000", 27248 => x"00000000",
    27249 => x"00000000", 27250 => x"00000000", 27251 => x"00000000",
    27252 => x"00000000", 27253 => x"00000000", 27254 => x"00000000",
    27255 => x"00000000", 27256 => x"00000000", 27257 => x"00000000",
    27258 => x"00000000", 27259 => x"00000000", 27260 => x"00000000",
    27261 => x"00000000", 27262 => x"00000000", 27263 => x"00000000",
    27264 => x"00000000", 27265 => x"00000000", 27266 => x"00000000",
    27267 => x"00000000", 27268 => x"00000000", 27269 => x"00000000",
    27270 => x"00000000", 27271 => x"00000000", 27272 => x"00000000",
    27273 => x"00000000", 27274 => x"00000000", 27275 => x"00000000",
    27276 => x"00000000", 27277 => x"00000000", 27278 => x"00000000",
    27279 => x"00000000", 27280 => x"00000000", 27281 => x"00000000",
    27282 => x"00000000", 27283 => x"00000000", 27284 => x"00000000",
    27285 => x"00000000", 27286 => x"00000000", 27287 => x"00000000",
    27288 => x"00000000", 27289 => x"00000000", 27290 => x"00000000",
    27291 => x"00000000", 27292 => x"00000000", 27293 => x"00000000",
    27294 => x"00000000", 27295 => x"00000000", 27296 => x"00000000",
    27297 => x"00000000", 27298 => x"00000000", 27299 => x"00000000",
    27300 => x"00000000", 27301 => x"00000000", 27302 => x"00000000",
    27303 => x"00000000", 27304 => x"00000000", 27305 => x"00000000",
    27306 => x"00000000", 27307 => x"00000000", 27308 => x"00000000",
    27309 => x"00000000", 27310 => x"00000000", 27311 => x"00000000",
    27312 => x"00000000", 27313 => x"00000000", 27314 => x"00000000",
    27315 => x"00000000", 27316 => x"00000000", 27317 => x"00000000",
    27318 => x"00000000", 27319 => x"00000000", 27320 => x"00000000",
    27321 => x"00000000", 27322 => x"00000000", 27323 => x"00000000",
    27324 => x"00000000", 27325 => x"00000000", 27326 => x"00000000",
    27327 => x"00000000", 27328 => x"00000000", 27329 => x"00000000",
    27330 => x"00000000", 27331 => x"00000000", 27332 => x"00000000",
    27333 => x"00000000", 27334 => x"00000000", 27335 => x"00000000",
    27336 => x"00000000", 27337 => x"00000000", 27338 => x"00000000",
    27339 => x"00000000", 27340 => x"00000000", 27341 => x"00000000",
    27342 => x"00000000", 27343 => x"00000000", 27344 => x"00000000",
    27345 => x"00000000", 27346 => x"00000000", 27347 => x"00000000",
    27348 => x"00000000", 27349 => x"00000000", 27350 => x"00000000",
    27351 => x"00000000", 27352 => x"00000000", 27353 => x"00000000",
    27354 => x"00000000", 27355 => x"00000000", 27356 => x"00000000",
    27357 => x"00000000", 27358 => x"00000000", 27359 => x"00000000",
    27360 => x"00000000", 27361 => x"00000000", 27362 => x"00000000",
    27363 => x"00000000", 27364 => x"00000000", 27365 => x"00000000",
    27366 => x"00000000", 27367 => x"00000000", 27368 => x"00000000",
    27369 => x"00000000", 27370 => x"00000000", 27371 => x"00000000",
    27372 => x"00000000", 27373 => x"00000000", 27374 => x"00000000",
    27375 => x"00000000", 27376 => x"00000000", 27377 => x"00000000",
    27378 => x"00000000", 27379 => x"00000000", 27380 => x"00000000",
    27381 => x"00000000", 27382 => x"00000000", 27383 => x"00000000",
    27384 => x"00000000", 27385 => x"00000000", 27386 => x"00000000",
    27387 => x"00000000", 27388 => x"00000000", 27389 => x"00000000",
    27390 => x"00000000", 27391 => x"00000000", 27392 => x"00000000",
    27393 => x"00000000", 27394 => x"00000000", 27395 => x"00000000",
    27396 => x"00000000", 27397 => x"00000000", 27398 => x"00000000",
    27399 => x"00000000", 27400 => x"00000000", 27401 => x"00000000",
    27402 => x"00000000", 27403 => x"00000000", 27404 => x"00000000",
    27405 => x"00000000", 27406 => x"00000000", 27407 => x"00000000",
    27408 => x"00000000", 27409 => x"00000000", 27410 => x"00000000",
    27411 => x"00000000", 27412 => x"00000000", 27413 => x"00000000",
    27414 => x"00000000", 27415 => x"00000000", 27416 => x"00000000",
    27417 => x"00000000", 27418 => x"00000000", 27419 => x"00000000",
    27420 => x"00000000", 27421 => x"00000000", 27422 => x"00000000",
    27423 => x"00000000", 27424 => x"00000000", 27425 => x"00000000",
    27426 => x"00000000", 27427 => x"00000000", 27428 => x"00000000",
    27429 => x"00000000", 27430 => x"00000000", 27431 => x"00000000",
    27432 => x"00000000", 27433 => x"00000000", 27434 => x"00000000",
    27435 => x"00000000", 27436 => x"00000000", 27437 => x"00000000",
    27438 => x"00000000", 27439 => x"00000000", 27440 => x"00000000",
    27441 => x"00000000", 27442 => x"00000000", 27443 => x"00000000",
    27444 => x"00000000", 27445 => x"00000000", 27446 => x"00000000",
    27447 => x"00000000", 27448 => x"00000000", 27449 => x"00000000",
    27450 => x"00000000", 27451 => x"00000000", 27452 => x"00000000",
    27453 => x"00000000", 27454 => x"00000000", 27455 => x"00000000",
    27456 => x"00000000", 27457 => x"00000000", 27458 => x"00000000",
    27459 => x"00000000", 27460 => x"00000000", 27461 => x"00000000",
    27462 => x"00000000", 27463 => x"00000000", 27464 => x"00000000",
    27465 => x"00000000", 27466 => x"00000000", 27467 => x"00000000",
    27468 => x"00000000", 27469 => x"00000000", 27470 => x"00000000",
    27471 => x"00000000", 27472 => x"00000000", 27473 => x"00000000",
    27474 => x"00000000", 27475 => x"00000000", 27476 => x"00000000",
    27477 => x"00000000", 27478 => x"00000000", 27479 => x"00000000",
    27480 => x"00000000", 27481 => x"00000000", 27482 => x"00000000",
    27483 => x"00000000", 27484 => x"00000000", 27485 => x"00000000",
    27486 => x"00000000", 27487 => x"00000000", 27488 => x"00000000",
    27489 => x"00000000", 27490 => x"00000000", 27491 => x"00000000",
    27492 => x"00000000", 27493 => x"00000000", 27494 => x"00000000",
    27495 => x"00000000", 27496 => x"00000000", 27497 => x"00000000",
    27498 => x"00000000", 27499 => x"00000000", 27500 => x"00000000",
    27501 => x"00000000", 27502 => x"00000000", 27503 => x"00000000",
    27504 => x"00000000", 27505 => x"00000000", 27506 => x"00000000",
    27507 => x"00000000", 27508 => x"00000000", 27509 => x"00000000",
    27510 => x"00000000", 27511 => x"00000000", 27512 => x"00000000",
    27513 => x"00000000", 27514 => x"00000000", 27515 => x"00000000",
    27516 => x"00000000", 27517 => x"00000000", 27518 => x"00000000",
    27519 => x"00000000", 27520 => x"00000000", 27521 => x"00000000",
    27522 => x"00000000", 27523 => x"00000000", 27524 => x"00000000",
    27525 => x"00000000", 27526 => x"00000000", 27527 => x"00000000",
    27528 => x"00000000", 27529 => x"00000000", 27530 => x"00000000",
    27531 => x"00000000", 27532 => x"00000000", 27533 => x"00000000",
    27534 => x"00000000", 27535 => x"00000000", 27536 => x"00000000",
    27537 => x"00000000", 27538 => x"00000000", 27539 => x"00000000",
    27540 => x"00000000", 27541 => x"00000000", 27542 => x"00000000",
    27543 => x"00000000", 27544 => x"00000000", 27545 => x"00000000",
    27546 => x"00000000", 27547 => x"00000000", 27548 => x"00000000",
    27549 => x"00000000", 27550 => x"00000000", 27551 => x"00000000",
    27552 => x"00000000", 27553 => x"00000000", 27554 => x"00000000",
    27555 => x"00000000", 27556 => x"00000000", 27557 => x"00000000",
    27558 => x"00000000", 27559 => x"00000000", 27560 => x"00000000",
    27561 => x"00000000", 27562 => x"00000000", 27563 => x"00000000",
    27564 => x"00000000", 27565 => x"00000000", 27566 => x"00000000",
    27567 => x"00000000", 27568 => x"00000000", 27569 => x"00000000",
    27570 => x"00000000", 27571 => x"00000000", 27572 => x"00000000",
    27573 => x"00000000", 27574 => x"00000000", 27575 => x"00000000",
    27576 => x"00000000", 27577 => x"00000000", 27578 => x"00000000",
    27579 => x"00000000", 27580 => x"00000000", 27581 => x"00000000",
    27582 => x"00000000", 27583 => x"00000000", 27584 => x"00000000",
    27585 => x"00000000", 27586 => x"00000000", 27587 => x"00000000",
    27588 => x"00000000", 27589 => x"00000000", 27590 => x"00000000",
    27591 => x"00000000", 27592 => x"00000000", 27593 => x"00000000",
    27594 => x"00000000", 27595 => x"00000000", 27596 => x"00000000",
    27597 => x"00000000", 27598 => x"00000000", 27599 => x"00000000",
    27600 => x"00000000", 27601 => x"00000000", 27602 => x"00000000",
    27603 => x"00000000", 27604 => x"00000000", 27605 => x"00000000",
    27606 => x"00000000", 27607 => x"00000000", 27608 => x"00000000",
    27609 => x"00000000", 27610 => x"00000000", 27611 => x"00000000",
    27612 => x"00000000", 27613 => x"00000000", 27614 => x"00000000",
    27615 => x"00000000", 27616 => x"00000000", 27617 => x"00000000",
    27618 => x"00000000", 27619 => x"00000000", 27620 => x"00000000",
    27621 => x"00000000", 27622 => x"00000000", 27623 => x"00000000",
    27624 => x"00000000", 27625 => x"00000000", 27626 => x"00000000",
    27627 => x"00000000", 27628 => x"00000000", 27629 => x"00000000",
    27630 => x"00000000", 27631 => x"00000000", 27632 => x"00000000",
    27633 => x"00000000", 27634 => x"00000000", 27635 => x"00000000",
    27636 => x"00000000", 27637 => x"00000000", 27638 => x"00000000",
    27639 => x"00000000", 27640 => x"00000000", 27641 => x"00000000",
    27642 => x"00000000", 27643 => x"00000000", 27644 => x"00000000",
    27645 => x"00000000", 27646 => x"00000000", 27647 => x"00000000",
    27648 => x"00000000", 27649 => x"00000000", 27650 => x"00000000",
    27651 => x"00000000", 27652 => x"00000000", 27653 => x"00000000",
    27654 => x"00000000", 27655 => x"00000000", 27656 => x"00000000",
    27657 => x"00000000", 27658 => x"00000000", 27659 => x"00000000",
    27660 => x"00000000", 27661 => x"00000000", 27662 => x"00000000",
    27663 => x"00000000", 27664 => x"00000000", 27665 => x"00000000",
    27666 => x"00000000", 27667 => x"00000000", 27668 => x"00000000",
    27669 => x"00000000", 27670 => x"00000000", 27671 => x"00000000",
    27672 => x"00000000", 27673 => x"00000000", 27674 => x"00000000",
    27675 => x"00000000", 27676 => x"00000000", 27677 => x"00000000",
    27678 => x"00000000", 27679 => x"00000000", 27680 => x"00000000",
    27681 => x"00000000", 27682 => x"00000000", 27683 => x"00000000",
    27684 => x"00000000", 27685 => x"00000000", 27686 => x"00000000",
    27687 => x"00000000", 27688 => x"00000000", 27689 => x"00000000",
    27690 => x"00000000", 27691 => x"00000000", 27692 => x"00000000",
    27693 => x"00000000", 27694 => x"00000000", 27695 => x"00000000",
    27696 => x"00000000", 27697 => x"00000000", 27698 => x"00000000",
    27699 => x"00000000", 27700 => x"00000000", 27701 => x"00000000",
    27702 => x"00000000", 27703 => x"00000000", 27704 => x"00000000",
    27705 => x"00000000", 27706 => x"00000000", 27707 => x"00000000",
    27708 => x"00000000", 27709 => x"00000000", 27710 => x"00000000",
    27711 => x"00000000", 27712 => x"00000000", 27713 => x"00000000",
    27714 => x"00000000", 27715 => x"00000000", 27716 => x"00000000",
    27717 => x"00000000", 27718 => x"00000000", 27719 => x"00000000",
    27720 => x"00000000", 27721 => x"00000000", 27722 => x"00000000",
    27723 => x"00000000", 27724 => x"00000000", 27725 => x"00000000",
    27726 => x"00000000", 27727 => x"00000000", 27728 => x"00000000",
    27729 => x"00000000", 27730 => x"00000000", 27731 => x"00000000",
    27732 => x"00000000", 27733 => x"00000000", 27734 => x"00000000",
    27735 => x"00000000", 27736 => x"00000000", 27737 => x"00000000",
    27738 => x"00000000", 27739 => x"00000000", 27740 => x"00000000",
    27741 => x"00000000", 27742 => x"00000000", 27743 => x"00000000",
    27744 => x"00000000", 27745 => x"00000000", 27746 => x"00000000",
    27747 => x"00000000", 27748 => x"00000000", 27749 => x"00000000",
    27750 => x"00000000", 27751 => x"00000000", 27752 => x"00000000",
    27753 => x"00000000", 27754 => x"00000000", 27755 => x"00000000",
    27756 => x"00000000", 27757 => x"00000000", 27758 => x"00000000",
    27759 => x"00000000", 27760 => x"00000000", 27761 => x"00000000",
    27762 => x"00000000", 27763 => x"00000000", 27764 => x"00000000",
    27765 => x"00000000", 27766 => x"00000000", 27767 => x"00000000",
    27768 => x"00000000", 27769 => x"00000000", 27770 => x"00000000",
    27771 => x"00000000", 27772 => x"00000000", 27773 => x"00000000",
    27774 => x"00000000", 27775 => x"00000000", 27776 => x"00000000",
    27777 => x"00000000", 27778 => x"00000000", 27779 => x"00000000",
    27780 => x"00000000", 27781 => x"00000000", 27782 => x"00000000",
    27783 => x"00000000", 27784 => x"00000000", 27785 => x"00000000",
    27786 => x"00000000", 27787 => x"00000000", 27788 => x"00000000",
    27789 => x"00000000", 27790 => x"00000000", 27791 => x"00000000",
    27792 => x"00000000", 27793 => x"00000000", 27794 => x"00000000",
    27795 => x"00000000", 27796 => x"00000000", 27797 => x"00000000",
    27798 => x"00000000", 27799 => x"00000000", 27800 => x"00000000",
    27801 => x"00000000", 27802 => x"00000000", 27803 => x"00000000",
    27804 => x"00000000", 27805 => x"00000000", 27806 => x"00000000",
    27807 => x"00000000", 27808 => x"00000000", 27809 => x"00000000",
    27810 => x"00000000", 27811 => x"00000000", 27812 => x"00000000",
    27813 => x"00000000", 27814 => x"00000000", 27815 => x"00000000",
    27816 => x"00000000", 27817 => x"00000000", 27818 => x"00000000",
    27819 => x"00000000", 27820 => x"00000000", 27821 => x"00000000",
    27822 => x"00000000", 27823 => x"00000000", 27824 => x"00000000",
    27825 => x"00000000", 27826 => x"00000000", 27827 => x"00000000",
    27828 => x"00000000", 27829 => x"00000000", 27830 => x"00000000",
    27831 => x"00000000", 27832 => x"00000000", 27833 => x"00000000",
    27834 => x"00000000", 27835 => x"00000000", 27836 => x"00000000",
    27837 => x"00000000", 27838 => x"00000000", 27839 => x"00000000",
    27840 => x"00000000", 27841 => x"00000000", 27842 => x"00000000",
    27843 => x"00000000", 27844 => x"00000000", 27845 => x"00000000",
    27846 => x"00000000", 27847 => x"00000000", 27848 => x"00000000",
    27849 => x"00000000", 27850 => x"00000000", 27851 => x"00000000",
    27852 => x"00000000", 27853 => x"00000000", 27854 => x"00000000",
    27855 => x"00000000", 27856 => x"00000000", 27857 => x"00000000",
    27858 => x"00000000", 27859 => x"00000000", 27860 => x"00000000",
    27861 => x"00000000", 27862 => x"00000000", 27863 => x"00000000",
    27864 => x"00000000", 27865 => x"00000000", 27866 => x"00000000",
    27867 => x"00000000", 27868 => x"00000000", 27869 => x"00000000",
    27870 => x"00000000", 27871 => x"00000000", 27872 => x"00000000",
    27873 => x"00000000", 27874 => x"00000000", 27875 => x"00000000",
    27876 => x"00000000", 27877 => x"00000000", 27878 => x"00000000",
    27879 => x"00000000", 27880 => x"00000000", 27881 => x"00000000",
    27882 => x"00000000", 27883 => x"00000000", 27884 => x"00000000",
    27885 => x"00000000", 27886 => x"00000000", 27887 => x"00000000",
    27888 => x"00000000", 27889 => x"00000000", 27890 => x"00000000",
    27891 => x"00000000", 27892 => x"00000000", 27893 => x"00000000",
    27894 => x"00000000", 27895 => x"00000000", 27896 => x"00000000",
    27897 => x"00000000", 27898 => x"00000000", 27899 => x"00000000",
    27900 => x"00000000", 27901 => x"00000000", 27902 => x"00000000",
    27903 => x"00000000", 27904 => x"00000000", 27905 => x"00000000",
    27906 => x"00000000", 27907 => x"00000000", 27908 => x"00000000",
    27909 => x"00000000", 27910 => x"00000000", 27911 => x"00000000",
    27912 => x"00000000", 27913 => x"00000000", 27914 => x"00000000",
    27915 => x"00000000", 27916 => x"00000000", 27917 => x"00000000",
    27918 => x"00000000", 27919 => x"00000000", 27920 => x"00000000",
    27921 => x"00000000", 27922 => x"00000000", 27923 => x"00000000",
    27924 => x"00000000", 27925 => x"00000000", 27926 => x"00000000",
    27927 => x"00000000", 27928 => x"00000000", 27929 => x"00000000",
    27930 => x"00000000", 27931 => x"00000000", 27932 => x"00000000",
    27933 => x"00000000", 27934 => x"00000000", 27935 => x"00000000",
    27936 => x"00000000", 27937 => x"00000000", 27938 => x"00000000",
    27939 => x"00000000", 27940 => x"00000000", 27941 => x"00000000",
    27942 => x"00000000", 27943 => x"00000000", 27944 => x"00000000",
    27945 => x"00000000", 27946 => x"00000000", 27947 => x"00000000",
    27948 => x"00000000", 27949 => x"00000000", 27950 => x"00000000",
    27951 => x"00000000", 27952 => x"00000000", 27953 => x"00000000",
    27954 => x"00000000", 27955 => x"00000000", 27956 => x"00000000",
    27957 => x"00000000", 27958 => x"00000000", 27959 => x"00000000",
    27960 => x"00000000", 27961 => x"00000000", 27962 => x"00000000",
    27963 => x"00000000", 27964 => x"00000000", 27965 => x"00000000",
    27966 => x"00000000", 27967 => x"00000000", 27968 => x"00000000",
    27969 => x"00000000", 27970 => x"00000000", 27971 => x"00000000",
    27972 => x"00000000", 27973 => x"00000000", 27974 => x"00000000",
    27975 => x"00000000", 27976 => x"00000000", 27977 => x"00000000",
    27978 => x"00000000", 27979 => x"00000000", 27980 => x"00000000",
    27981 => x"00000000", 27982 => x"00000000", 27983 => x"00000000",
    27984 => x"00000000", 27985 => x"00000000", 27986 => x"00000000",
    27987 => x"00000000", 27988 => x"00000000", 27989 => x"00000000",
    27990 => x"00000000", 27991 => x"00000000", 27992 => x"00000000",
    27993 => x"00000000", 27994 => x"00000000", 27995 => x"00000000",
    27996 => x"00000000", 27997 => x"00000000", 27998 => x"00000000",
    27999 => x"00000000", 28000 => x"00000000", 28001 => x"00000000",
    28002 => x"00000000", 28003 => x"00000000", 28004 => x"00000000",
    28005 => x"00000000", 28006 => x"00000000", 28007 => x"00000000",
    28008 => x"00000000", 28009 => x"00000000", 28010 => x"00000000",
    28011 => x"00000000", 28012 => x"00000000", 28013 => x"00000000",
    28014 => x"00000000", 28015 => x"00000000", 28016 => x"00000000",
    28017 => x"00000000", 28018 => x"00000000", 28019 => x"00000000",
    28020 => x"00000000", 28021 => x"00000000", 28022 => x"00000000",
    28023 => x"00000000", 28024 => x"00000000", 28025 => x"00000000",
    28026 => x"00000000", 28027 => x"00000000", 28028 => x"00000000",
    28029 => x"00000000", 28030 => x"00000000", 28031 => x"00000000",
    28032 => x"00000000", 28033 => x"00000000", 28034 => x"00000000",
    28035 => x"00000000", 28036 => x"00000000", 28037 => x"00000000",
    28038 => x"00000000", 28039 => x"00000000", 28040 => x"00000000",
    28041 => x"00000000", 28042 => x"00000000", 28043 => x"00000000",
    28044 => x"00000000", 28045 => x"00000000", 28046 => x"00000000",
    28047 => x"00000000", 28048 => x"00000000", 28049 => x"00000000",
    28050 => x"00000000", 28051 => x"00000000", 28052 => x"00000000",
    28053 => x"00000000", 28054 => x"00000000", 28055 => x"00000000",
    28056 => x"00000000", 28057 => x"00000000", 28058 => x"00000000",
    28059 => x"00000000", 28060 => x"00000000", 28061 => x"00000000",
    28062 => x"00000000", 28063 => x"00000000", 28064 => x"00000000",
    28065 => x"00000000", 28066 => x"00000000", 28067 => x"00000000",
    28068 => x"00000000", 28069 => x"00000000", 28070 => x"00000000",
    28071 => x"00000000", 28072 => x"00000000", 28073 => x"00000000",
    28074 => x"00000000", 28075 => x"00000000", 28076 => x"00000000",
    28077 => x"00000000", 28078 => x"00000000", 28079 => x"00000000",
    28080 => x"00000000", 28081 => x"00000000", 28082 => x"00000000",
    28083 => x"00000000", 28084 => x"00000000", 28085 => x"00000000",
    28086 => x"00000000", 28087 => x"00000000", 28088 => x"00000000",
    28089 => x"00000000", 28090 => x"00000000", 28091 => x"00000000",
    28092 => x"00000000", 28093 => x"00000000", 28094 => x"00000000",
    28095 => x"00000000", 28096 => x"00000000", 28097 => x"00000000",
    28098 => x"00000000", 28099 => x"00000000", 28100 => x"00000000",
    28101 => x"00000000", 28102 => x"00000000", 28103 => x"00000000",
    28104 => x"00000000", 28105 => x"00000000", 28106 => x"00000000",
    28107 => x"00000000", 28108 => x"00000000", 28109 => x"00000000",
    28110 => x"00000000", 28111 => x"00000000", 28112 => x"00000000",
    28113 => x"00000000", 28114 => x"00000000", 28115 => x"00000000",
    28116 => x"00000000", 28117 => x"00000000", 28118 => x"00000000",
    28119 => x"00000000", 28120 => x"00000000", 28121 => x"00000000",
    28122 => x"00000000", 28123 => x"00000000", 28124 => x"00000000",
    28125 => x"00000000", 28126 => x"00000000", 28127 => x"00000000",
    28128 => x"00000000", 28129 => x"00000000", 28130 => x"00000000",
    28131 => x"00000000", 28132 => x"00000000", 28133 => x"00000000",
    28134 => x"00000000", 28135 => x"00000000", 28136 => x"00000000",
    28137 => x"00000000", 28138 => x"00000000", 28139 => x"00000000",
    28140 => x"00000000", 28141 => x"00000000", 28142 => x"00000000",
    28143 => x"00000000", 28144 => x"00000000", 28145 => x"00000000",
    28146 => x"00000000", 28147 => x"00000000", 28148 => x"00000000",
    28149 => x"00000000", 28150 => x"00000000", 28151 => x"00000000",
    28152 => x"00000000", 28153 => x"00000000", 28154 => x"00000000",
    28155 => x"00000000", 28156 => x"00000000", 28157 => x"00000000",
    28158 => x"00000000", 28159 => x"00000000", 28160 => x"00000000",
    28161 => x"00000000", 28162 => x"00000000", 28163 => x"00000000",
    28164 => x"00000000", 28165 => x"00000000", 28166 => x"00000000",
    28167 => x"00000000", 28168 => x"00000000", 28169 => x"00000000",
    28170 => x"00000000", 28171 => x"00000000", 28172 => x"00000000",
    28173 => x"00000000", 28174 => x"00000000", 28175 => x"00000000",
    28176 => x"00000000", 28177 => x"00000000", 28178 => x"00000000",
    28179 => x"00000000", 28180 => x"00000000", 28181 => x"00000000",
    28182 => x"00000000", 28183 => x"00000000", 28184 => x"00000000",
    28185 => x"00000000", 28186 => x"00000000", 28187 => x"00000000",
    28188 => x"00000000", 28189 => x"00000000", 28190 => x"00000000",
    28191 => x"00000000", 28192 => x"00000000", 28193 => x"00000000",
    28194 => x"00000000", 28195 => x"00000000", 28196 => x"00000000",
    28197 => x"00000000", 28198 => x"00000000", 28199 => x"00000000",
    28200 => x"00000000", 28201 => x"00000000", 28202 => x"00000000",
    28203 => x"00000000", 28204 => x"00000000", 28205 => x"00000000",
    28206 => x"00000000", 28207 => x"00000000", 28208 => x"00000000",
    28209 => x"00000000", 28210 => x"00000000", 28211 => x"00000000",
    28212 => x"00000000", 28213 => x"00000000", 28214 => x"00000000",
    28215 => x"00000000", 28216 => x"00000000", 28217 => x"00000000",
    28218 => x"00000000", 28219 => x"00000000", 28220 => x"00000000",
    28221 => x"00000000", 28222 => x"00000000", 28223 => x"00000000",
    28224 => x"00000000", 28225 => x"00000000", 28226 => x"00000000",
    28227 => x"00000000", 28228 => x"00000000", 28229 => x"00000000",
    28230 => x"00000000", 28231 => x"00000000", 28232 => x"00000000",
    28233 => x"00000000", 28234 => x"00000000", 28235 => x"00000000",
    28236 => x"00000000", 28237 => x"00000000", 28238 => x"00000000",
    28239 => x"00000000", 28240 => x"00000000", 28241 => x"00000000",
    28242 => x"00000000", 28243 => x"00000000", 28244 => x"00000000",
    28245 => x"00000000", 28246 => x"00000000", 28247 => x"00000000",
    28248 => x"00000000", 28249 => x"00000000", 28250 => x"00000000",
    28251 => x"00000000", 28252 => x"00000000", 28253 => x"00000000",
    28254 => x"00000000", 28255 => x"00000000", 28256 => x"00000000",
    28257 => x"00000000", 28258 => x"00000000", 28259 => x"00000000",
    28260 => x"00000000", 28261 => x"00000000", 28262 => x"00000000",
    28263 => x"00000000", 28264 => x"00000000", 28265 => x"00000000",
    28266 => x"00000000", 28267 => x"00000000", 28268 => x"00000000",
    28269 => x"00000000", 28270 => x"00000000", 28271 => x"00000000",
    28272 => x"00000000", 28273 => x"00000000", 28274 => x"00000000",
    28275 => x"00000000", 28276 => x"00000000", 28277 => x"00000000",
    28278 => x"00000000", 28279 => x"00000000", 28280 => x"00000000",
    28281 => x"00000000", 28282 => x"00000000", 28283 => x"00000000",
    28284 => x"00000000", 28285 => x"00000000", 28286 => x"00000000",
    28287 => x"00000000", 28288 => x"00000000", 28289 => x"00000000",
    28290 => x"00000000", 28291 => x"00000000", 28292 => x"00000000",
    28293 => x"00000000", 28294 => x"00000000", 28295 => x"00000000",
    28296 => x"00000000", 28297 => x"00000000", 28298 => x"00000000",
    28299 => x"00000000", 28300 => x"00000000", 28301 => x"00000000",
    28302 => x"00000000", 28303 => x"00000000", 28304 => x"00000000",
    28305 => x"00000000", 28306 => x"00000000", 28307 => x"00000000",
    28308 => x"00000000", 28309 => x"00000000", 28310 => x"00000000",
    28311 => x"00000000", 28312 => x"00000000", 28313 => x"00000000",
    28314 => x"00000000", 28315 => x"00000000", 28316 => x"00000000",
    28317 => x"00000000", 28318 => x"00000000", 28319 => x"00000000",
    28320 => x"00000000", 28321 => x"00000000", 28322 => x"00000000",
    28323 => x"00000000", 28324 => x"00000000", 28325 => x"00000000",
    28326 => x"00000000", 28327 => x"00000000", 28328 => x"00000000",
    28329 => x"00000000", 28330 => x"00000000", 28331 => x"00000000",
    28332 => x"00000000", 28333 => x"00000000", 28334 => x"00000000",
    28335 => x"00000000", 28336 => x"00000000", 28337 => x"00000000",
    28338 => x"00000000", 28339 => x"00000000", 28340 => x"00000000",
    28341 => x"00000000", 28342 => x"00000000", 28343 => x"00000000",
    28344 => x"00000000", 28345 => x"00000000", 28346 => x"00000000",
    28347 => x"00000000", 28348 => x"00000000", 28349 => x"00000000",
    28350 => x"00000000", 28351 => x"00000000", 28352 => x"00000000",
    28353 => x"00000000", 28354 => x"00000000", 28355 => x"00000000",
    28356 => x"00000000", 28357 => x"00000000", 28358 => x"00000000",
    28359 => x"00000000", 28360 => x"00000000", 28361 => x"00000000",
    28362 => x"00000000", 28363 => x"00000000", 28364 => x"00000000",
    28365 => x"00000000", 28366 => x"00000000", 28367 => x"00000000",
    28368 => x"00000000", 28369 => x"00000000", 28370 => x"00000000",
    28371 => x"00000000", 28372 => x"00000000", 28373 => x"00000000",
    28374 => x"00000000", 28375 => x"00000000", 28376 => x"00000000",
    28377 => x"00000000", 28378 => x"00000000", 28379 => x"00000000",
    28380 => x"00000000", 28381 => x"00000000", 28382 => x"00000000",
    28383 => x"00000000", 28384 => x"00000000", 28385 => x"00000000",
    28386 => x"00000000", 28387 => x"00000000", 28388 => x"00000000",
    28389 => x"00000000", 28390 => x"00000000", 28391 => x"00000000",
    28392 => x"00000000", 28393 => x"00000000", 28394 => x"00000000",
    28395 => x"00000000", 28396 => x"00000000", 28397 => x"00000000",
    28398 => x"00000000", 28399 => x"00000000", 28400 => x"00000000",
    28401 => x"00000000", 28402 => x"00000000", 28403 => x"00000000",
    28404 => x"00000000", 28405 => x"00000000", 28406 => x"00000000",
    28407 => x"00000000", 28408 => x"00000000", 28409 => x"00000000",
    28410 => x"00000000", 28411 => x"00000000", 28412 => x"00000000",
    28413 => x"00000000", 28414 => x"00000000", 28415 => x"00000000",
    28416 => x"00000000", 28417 => x"00000000", 28418 => x"00000000",
    28419 => x"00000000", 28420 => x"00000000", 28421 => x"00000000",
    28422 => x"00000000", 28423 => x"00000000", 28424 => x"00000000",
    28425 => x"00000000", 28426 => x"00000000", 28427 => x"00000000",
    28428 => x"00000000", 28429 => x"00000000", 28430 => x"00000000",
    28431 => x"00000000", 28432 => x"00000000", 28433 => x"00000000",
    28434 => x"00000000", 28435 => x"00000000", 28436 => x"00000000",
    28437 => x"00000000", 28438 => x"00000000", 28439 => x"00000000",
    28440 => x"00000000", 28441 => x"00000000", 28442 => x"00000000",
    28443 => x"00000000", 28444 => x"00000000", 28445 => x"00000000",
    28446 => x"00000000", 28447 => x"00000000", 28448 => x"00000000",
    28449 => x"00000000", 28450 => x"00000000", 28451 => x"00000000",
    28452 => x"00000000", 28453 => x"00000000", 28454 => x"00000000",
    28455 => x"00000000", 28456 => x"00000000", 28457 => x"00000000",
    28458 => x"00000000", 28459 => x"00000000", 28460 => x"00000000",
    28461 => x"00000000", 28462 => x"00000000", 28463 => x"00000000",
    28464 => x"00000000", 28465 => x"00000000", 28466 => x"00000000",
    28467 => x"00000000", 28468 => x"00000000", 28469 => x"00000000",
    28470 => x"00000000", 28471 => x"00000000", 28472 => x"00000000",
    28473 => x"00000000", 28474 => x"00000000", 28475 => x"00000000",
    28476 => x"00000000", 28477 => x"00000000", 28478 => x"00000000",
    28479 => x"00000000", 28480 => x"00000000", 28481 => x"00000000",
    28482 => x"00000000", 28483 => x"00000000", 28484 => x"00000000",
    28485 => x"00000000", 28486 => x"00000000", 28487 => x"00000000",
    28488 => x"00000000", 28489 => x"00000000", 28490 => x"00000000",
    28491 => x"00000000", 28492 => x"00000000", 28493 => x"00000000",
    28494 => x"00000000", 28495 => x"00000000", 28496 => x"00000000",
    28497 => x"00000000", 28498 => x"00000000", 28499 => x"00000000",
    28500 => x"00000000", 28501 => x"00000000", 28502 => x"00000000",
    28503 => x"00000000", 28504 => x"00000000", 28505 => x"00000000",
    28506 => x"00000000", 28507 => x"00000000", 28508 => x"00000000",
    28509 => x"00000000", 28510 => x"00000000", 28511 => x"00000000",
    28512 => x"00000000", 28513 => x"00000000", 28514 => x"00000000",
    28515 => x"00000000", 28516 => x"00000000", 28517 => x"00000000",
    28518 => x"00000000", 28519 => x"00000000", 28520 => x"00000000",
    28521 => x"00000000", 28522 => x"00000000", 28523 => x"00000000",
    28524 => x"00000000", 28525 => x"00000000", 28526 => x"00000000",
    28527 => x"00000000", 28528 => x"00000000", 28529 => x"00000000",
    28530 => x"00000000", 28531 => x"00000000", 28532 => x"00000000",
    28533 => x"00000000", 28534 => x"00000000", 28535 => x"00000000",
    28536 => x"00000000", 28537 => x"00000000", 28538 => x"00000000",
    28539 => x"00000000", 28540 => x"00000000", 28541 => x"00000000",
    28542 => x"00000000", 28543 => x"00000000", 28544 => x"00000000",
    28545 => x"00000000", 28546 => x"00000000", 28547 => x"00000000",
    28548 => x"00000000", 28549 => x"00000000", 28550 => x"00000000",
    28551 => x"00000000", 28552 => x"00000000", 28553 => x"00000000",
    28554 => x"00000000", 28555 => x"00000000", 28556 => x"00000000",
    28557 => x"00000000", 28558 => x"00000000", 28559 => x"00000000",
    28560 => x"00000000", 28561 => x"00000000", 28562 => x"00000000",
    28563 => x"00000000", 28564 => x"00000000", 28565 => x"00000000",
    28566 => x"00000000", 28567 => x"00000000", 28568 => x"00000000",
    28569 => x"00000000", 28570 => x"00000000", 28571 => x"00000000",
    28572 => x"00000000", 28573 => x"00000000", 28574 => x"00000000",
    28575 => x"00000000", 28576 => x"00000000", 28577 => x"00000000",
    28578 => x"00000000", 28579 => x"00000000", 28580 => x"00000000",
    28581 => x"00000000", 28582 => x"00000000", 28583 => x"00000000",
    28584 => x"00000000", 28585 => x"00000000", 28586 => x"00000000",
    28587 => x"00000000", 28588 => x"00000000", 28589 => x"00000000",
    28590 => x"00000000", 28591 => x"00000000", 28592 => x"00000000",
    28593 => x"00000000", 28594 => x"00000000", 28595 => x"00000000",
    28596 => x"00000000", 28597 => x"00000000", 28598 => x"00000000",
    28599 => x"00000000", 28600 => x"00000000", 28601 => x"00000000",
    28602 => x"00000000", 28603 => x"00000000", 28604 => x"00000000",
    28605 => x"00000000", 28606 => x"00000000", 28607 => x"00000000",
    28608 => x"00000000", 28609 => x"00000000", 28610 => x"00000000",
    28611 => x"00000000", 28612 => x"00000000", 28613 => x"00000000",
    28614 => x"00000000", 28615 => x"00000000", 28616 => x"00000000",
    28617 => x"00000000", 28618 => x"00000000", 28619 => x"00000000",
    28620 => x"00000000", 28621 => x"00000000", 28622 => x"00000000",
    28623 => x"00000000", 28624 => x"00000000", 28625 => x"00000000",
    28626 => x"00000000", 28627 => x"00000000", 28628 => x"00000000",
    28629 => x"00000000", 28630 => x"00000000", 28631 => x"00000000",
    28632 => x"00000000", 28633 => x"00000000", 28634 => x"00000000",
    28635 => x"00000000", 28636 => x"00000000", 28637 => x"00000000",
    28638 => x"00000000", 28639 => x"00000000", 28640 => x"00000000",
    28641 => x"00000000", 28642 => x"00000000", 28643 => x"00000000",
    28644 => x"00000000", 28645 => x"00000000", 28646 => x"00000000",
    28647 => x"00000000", 28648 => x"00000000", 28649 => x"00000000",
    28650 => x"00000000", 28651 => x"00000000", 28652 => x"00000000",
    28653 => x"00000000", 28654 => x"00000000", 28655 => x"00000000",
    28656 => x"00000000", 28657 => x"00000000", 28658 => x"00000000",
    28659 => x"00000000", 28660 => x"00000000", 28661 => x"00000000",
    28662 => x"00000000", 28663 => x"00000000", 28664 => x"00000000",
    28665 => x"00000000", 28666 => x"00000000", 28667 => x"00000000",
    28668 => x"00000000", 28669 => x"00000000", 28670 => x"00000000",
    28671 => x"00000000", 28672 => x"00000000", 28673 => x"00000000",
    28674 => x"00000000", 28675 => x"00000000", 28676 => x"00000000",
    28677 => x"00000000", 28678 => x"00000000", 28679 => x"00000000",
    28680 => x"00000000", 28681 => x"00000000", 28682 => x"00000000",
    28683 => x"00000000", 28684 => x"00000000", 28685 => x"00000000",
    28686 => x"00000000", 28687 => x"00000000", 28688 => x"00000000",
    28689 => x"00000000", 28690 => x"00000000", 28691 => x"00000000",
    28692 => x"00000000", 28693 => x"00000000", 28694 => x"00000000",
    28695 => x"00000000", 28696 => x"00000000", 28697 => x"00000000",
    28698 => x"00000000", 28699 => x"00000000", 28700 => x"00000000",
    28701 => x"00000000", 28702 => x"00000000", 28703 => x"00000000",
    28704 => x"00000000", 28705 => x"00000000", 28706 => x"00000000",
    28707 => x"00000000", 28708 => x"00000000", 28709 => x"00000000",
    28710 => x"00000000", 28711 => x"00000000", 28712 => x"00000000",
    28713 => x"00000000", 28714 => x"00000000", 28715 => x"00000000",
    28716 => x"00000000", 28717 => x"00000000", 28718 => x"00000000",
    28719 => x"00000000", 28720 => x"00000000", 28721 => x"00000000",
    28722 => x"00000000", 28723 => x"00000000", 28724 => x"00000000",
    28725 => x"00000000", 28726 => x"00000000", 28727 => x"00000000",
    28728 => x"00000000", 28729 => x"00000000", 28730 => x"00000000",
    28731 => x"00000000", 28732 => x"00000000", 28733 => x"00000000",
    28734 => x"00000000", 28735 => x"00000000", 28736 => x"00000000",
    28737 => x"00000000", 28738 => x"00000000", 28739 => x"00000000",
    28740 => x"00000000", 28741 => x"00000000", 28742 => x"00000000",
    28743 => x"00000000", 28744 => x"00000000", 28745 => x"00000000",
    28746 => x"00000000", 28747 => x"00000000", 28748 => x"00000000",
    28749 => x"00000000", 28750 => x"00000000", 28751 => x"00000000",
    28752 => x"00000000", 28753 => x"00000000", 28754 => x"00000000",
    28755 => x"00000000", 28756 => x"00000000", 28757 => x"00000000",
    28758 => x"00000000", 28759 => x"00000000", 28760 => x"00000000",
    28761 => x"00000000", 28762 => x"00000000", 28763 => x"00000000",
    28764 => x"00000000", 28765 => x"00000000", 28766 => x"00000000",
    28767 => x"00000000", 28768 => x"00000000", 28769 => x"00000000",
    28770 => x"00000000", 28771 => x"00000000", 28772 => x"00000000",
    28773 => x"00000000", 28774 => x"00000000", 28775 => x"00000000",
    28776 => x"00000000", 28777 => x"00000000", 28778 => x"00000000",
    28779 => x"00000000", 28780 => x"00000000", 28781 => x"00000000",
    28782 => x"00000000", 28783 => x"00000000", 28784 => x"00000000",
    28785 => x"00000000", 28786 => x"00000000", 28787 => x"00000000",
    28788 => x"00000000", 28789 => x"00000000", 28790 => x"00000000",
    28791 => x"00000000", 28792 => x"00000000", 28793 => x"00000000",
    28794 => x"00000000", 28795 => x"00000000", 28796 => x"00000000",
    28797 => x"00000000", 28798 => x"00000000", 28799 => x"00000000",
    28800 => x"00000000", 28801 => x"00000000", 28802 => x"00000000",
    28803 => x"00000000", 28804 => x"00000000", 28805 => x"00000000",
    28806 => x"00000000", 28807 => x"00000000", 28808 => x"00000000",
    28809 => x"00000000", 28810 => x"00000000", 28811 => x"00000000",
    28812 => x"00000000", 28813 => x"00000000", 28814 => x"00000000",
    28815 => x"00000000", 28816 => x"00000000", 28817 => x"00000000",
    28818 => x"00000000", 28819 => x"00000000", 28820 => x"00000000",
    28821 => x"00000000", 28822 => x"00000000", 28823 => x"00000000",
    28824 => x"00000000", 28825 => x"00000000", 28826 => x"00000000",
    28827 => x"00000000", 28828 => x"00000000", 28829 => x"00000000",
    28830 => x"00000000", 28831 => x"00000000", 28832 => x"00000000",
    28833 => x"00000000", 28834 => x"00000000", 28835 => x"00000000",
    28836 => x"00000000", 28837 => x"00000000", 28838 => x"00000000",
    28839 => x"00000000", 28840 => x"00000000", 28841 => x"00000000",
    28842 => x"00000000", 28843 => x"00000000", 28844 => x"00000000",
    28845 => x"00000000", 28846 => x"00000000", 28847 => x"00000000",
    28848 => x"00000000", 28849 => x"00000000", 28850 => x"00000000",
    28851 => x"00000000", 28852 => x"00000000", 28853 => x"00000000",
    28854 => x"00000000", 28855 => x"00000000", 28856 => x"00000000",
    28857 => x"00000000", 28858 => x"00000000", 28859 => x"00000000",
    28860 => x"00000000", 28861 => x"00000000", 28862 => x"00000000",
    28863 => x"00000000", 28864 => x"00000000", 28865 => x"00000000",
    28866 => x"00000000", 28867 => x"00000000", 28868 => x"00000000",
    28869 => x"00000000", 28870 => x"00000000", 28871 => x"00000000",
    28872 => x"00000000", 28873 => x"00000000", 28874 => x"00000000",
    28875 => x"00000000", 28876 => x"00000000", 28877 => x"00000000",
    28878 => x"00000000", 28879 => x"00000000", 28880 => x"00000000",
    28881 => x"00000000", 28882 => x"00000000", 28883 => x"00000000",
    28884 => x"00000000", 28885 => x"00000000", 28886 => x"00000000",
    28887 => x"00000000", 28888 => x"00000000", 28889 => x"00000000",
    28890 => x"00000000", 28891 => x"00000000", 28892 => x"00000000",
    28893 => x"00000000", 28894 => x"00000000", 28895 => x"00000000",
    28896 => x"00000000", 28897 => x"00000000", 28898 => x"00000000",
    28899 => x"00000000", 28900 => x"00000000", 28901 => x"00000000",
    28902 => x"00000000", 28903 => x"00000000", 28904 => x"00000000",
    28905 => x"00000000", 28906 => x"00000000", 28907 => x"00000000",
    28908 => x"00000000", 28909 => x"00000000", 28910 => x"00000000",
    28911 => x"00000000", 28912 => x"00000000", 28913 => x"00000000",
    28914 => x"00000000", 28915 => x"00000000", 28916 => x"00000000",
    28917 => x"00000000", 28918 => x"00000000", 28919 => x"00000000",
    28920 => x"00000000", 28921 => x"00000000", 28922 => x"00000000",
    28923 => x"00000000", 28924 => x"00000000", 28925 => x"00000000",
    28926 => x"00000000", 28927 => x"00000000", 28928 => x"00000000",
    28929 => x"00000000", 28930 => x"00000000", 28931 => x"00000000",
    28932 => x"00000000", 28933 => x"00000000", 28934 => x"00000000",
    28935 => x"00000000", 28936 => x"00000000", 28937 => x"00000000",
    28938 => x"00000000", 28939 => x"00000000", 28940 => x"00000000",
    28941 => x"00000000", 28942 => x"00000000", 28943 => x"00000000",
    28944 => x"00000000", 28945 => x"00000000", 28946 => x"00000000",
    28947 => x"00000000", 28948 => x"00000000", 28949 => x"00000000",
    28950 => x"00000000", 28951 => x"00000000", 28952 => x"00000000",
    28953 => x"00000000", 28954 => x"00000000", 28955 => x"00000000",
    28956 => x"00000000", 28957 => x"00000000", 28958 => x"00000000",
    28959 => x"00000000", 28960 => x"00000000", 28961 => x"00000000",
    28962 => x"00000000", 28963 => x"00000000", 28964 => x"00000000",
    28965 => x"00000000", 28966 => x"00000000", 28967 => x"00000000",
    28968 => x"00000000", 28969 => x"00000000", 28970 => x"00000000",
    28971 => x"00000000", 28972 => x"00000000", 28973 => x"00000000",
    28974 => x"00000000", 28975 => x"00000000", 28976 => x"00000000",
    28977 => x"00000000", 28978 => x"00000000", 28979 => x"00000000",
    28980 => x"00000000", 28981 => x"00000000", 28982 => x"00000000",
    28983 => x"00000000", 28984 => x"00000000", 28985 => x"00000000",
    28986 => x"00000000", 28987 => x"00000000", 28988 => x"00000000",
    28989 => x"00000000", 28990 => x"00000000", 28991 => x"00000000",
    28992 => x"00000000", 28993 => x"00000000", 28994 => x"00000000",
    28995 => x"00000000", 28996 => x"00000000", 28997 => x"00000000",
    28998 => x"00000000", 28999 => x"00000000", 29000 => x"00000000",
    29001 => x"00000000", 29002 => x"00000000", 29003 => x"00000000",
    29004 => x"00000000", 29005 => x"00000000", 29006 => x"00000000",
    29007 => x"00000000", 29008 => x"00000000", 29009 => x"00000000",
    29010 => x"00000000", 29011 => x"00000000", 29012 => x"00000000",
    29013 => x"00000000", 29014 => x"00000000", 29015 => x"00000000",
    29016 => x"00000000", 29017 => x"00000000", 29018 => x"00000000",
    29019 => x"00000000", 29020 => x"00000000", 29021 => x"00000000",
    29022 => x"00000000", 29023 => x"00000000", 29024 => x"00000000",
    29025 => x"00000000", 29026 => x"00000000", 29027 => x"00000000",
    29028 => x"00000000", 29029 => x"00000000", 29030 => x"00000000",
    29031 => x"00000000", 29032 => x"00000000", 29033 => x"00000000",
    29034 => x"00000000", 29035 => x"00000000", 29036 => x"00000000",
    29037 => x"00000000", 29038 => x"00000000", 29039 => x"00000000",
    29040 => x"00000000", 29041 => x"00000000", 29042 => x"00000000",
    29043 => x"00000000", 29044 => x"00000000", 29045 => x"00000000",
    29046 => x"00000000", 29047 => x"00000000", 29048 => x"00000000",
    29049 => x"00000000", 29050 => x"00000000", 29051 => x"00000000",
    29052 => x"00000000", 29053 => x"00000000", 29054 => x"00000000",
    29055 => x"00000000", 29056 => x"00000000", 29057 => x"00000000",
    29058 => x"00000000", 29059 => x"00000000", 29060 => x"00000000",
    29061 => x"00000000", 29062 => x"00000000", 29063 => x"00000000",
    29064 => x"00000000", 29065 => x"00000000", 29066 => x"00000000",
    29067 => x"00000000", 29068 => x"00000000", 29069 => x"00000000",
    29070 => x"00000000", 29071 => x"00000000", 29072 => x"00000000",
    29073 => x"00000000", 29074 => x"00000000", 29075 => x"00000000",
    29076 => x"00000000", 29077 => x"00000000", 29078 => x"00000000",
    29079 => x"00000000", 29080 => x"00000000", 29081 => x"00000000",
    29082 => x"00000000", 29083 => x"00000000", 29084 => x"00000000",
    29085 => x"00000000", 29086 => x"00000000", 29087 => x"00000000",
    29088 => x"00000000", 29089 => x"00000000", 29090 => x"00000000",
    29091 => x"00000000", 29092 => x"00000000", 29093 => x"00000000",
    29094 => x"00000000", 29095 => x"00000000", 29096 => x"00000000",
    29097 => x"00000000", 29098 => x"00000000", 29099 => x"00000000",
    29100 => x"00000000", 29101 => x"00000000", 29102 => x"00000000",
    29103 => x"00000000", 29104 => x"00000000", 29105 => x"00000000",
    29106 => x"00000000", 29107 => x"00000000", 29108 => x"00000000",
    29109 => x"00000000", 29110 => x"00000000", 29111 => x"00000000",
    29112 => x"00000000", 29113 => x"00000000", 29114 => x"00000000",
    29115 => x"00000000", 29116 => x"00000000", 29117 => x"00000000",
    29118 => x"00000000", 29119 => x"00000000", 29120 => x"00000000",
    29121 => x"00000000", 29122 => x"00000000", 29123 => x"00000000",
    29124 => x"00000000", 29125 => x"00000000", 29126 => x"00000000",
    29127 => x"00000000", 29128 => x"00000000", 29129 => x"00000000",
    29130 => x"00000000", 29131 => x"00000000", 29132 => x"00000000",
    29133 => x"00000000", 29134 => x"00000000", 29135 => x"00000000",
    29136 => x"00000000", 29137 => x"00000000", 29138 => x"00000000",
    29139 => x"00000000", 29140 => x"00000000", 29141 => x"00000000",
    29142 => x"00000000", 29143 => x"00000000", 29144 => x"00000000",
    29145 => x"00000000", 29146 => x"00000000", 29147 => x"00000000",
    29148 => x"00000000", 29149 => x"00000000", 29150 => x"00000000",
    29151 => x"00000000", 29152 => x"00000000", 29153 => x"00000000",
    29154 => x"00000000", 29155 => x"00000000", 29156 => x"00000000",
    29157 => x"00000000", 29158 => x"00000000", 29159 => x"00000000",
    29160 => x"00000000", 29161 => x"00000000", 29162 => x"00000000",
    29163 => x"00000000", 29164 => x"00000000", 29165 => x"00000000",
    29166 => x"00000000", 29167 => x"00000000", 29168 => x"00000000",
    29169 => x"00000000", 29170 => x"00000000", 29171 => x"00000000",
    29172 => x"00000000", 29173 => x"00000000", 29174 => x"00000000",
    29175 => x"00000000", 29176 => x"00000000", 29177 => x"00000000",
    29178 => x"00000000", 29179 => x"00000000", 29180 => x"00000000",
    29181 => x"00000000", 29182 => x"00000000", 29183 => x"00000000",
    29184 => x"00000000", 29185 => x"00000000", 29186 => x"00000000",
    29187 => x"00000000", 29188 => x"00000000", 29189 => x"00000000",
    29190 => x"00000000", 29191 => x"00000000", 29192 => x"00000000",
    29193 => x"00000000", 29194 => x"00000000", 29195 => x"00000000",
    29196 => x"00000000", 29197 => x"00000000", 29198 => x"00000000",
    29199 => x"00000000", 29200 => x"00000000", 29201 => x"00000000",
    29202 => x"00000000", 29203 => x"00000000", 29204 => x"00000000",
    29205 => x"00000000", 29206 => x"00000000", 29207 => x"00000000",
    29208 => x"00000000", 29209 => x"00000000", 29210 => x"00000000",
    29211 => x"00000000", 29212 => x"00000000", 29213 => x"00000000",
    29214 => x"00000000", 29215 => x"00000000", 29216 => x"00000000",
    29217 => x"00000000", 29218 => x"00000000", 29219 => x"00000000",
    29220 => x"00000000", 29221 => x"00000000", 29222 => x"00000000",
    29223 => x"00000000", 29224 => x"00000000", 29225 => x"00000000",
    29226 => x"00000000", 29227 => x"00000000", 29228 => x"00000000",
    29229 => x"00000000", 29230 => x"00000000", 29231 => x"00000000",
    29232 => x"00000000", 29233 => x"00000000", 29234 => x"00000000",
    29235 => x"00000000", 29236 => x"00000000", 29237 => x"00000000",
    29238 => x"00000000", 29239 => x"00000000", 29240 => x"00000000",
    29241 => x"00000000", 29242 => x"00000000", 29243 => x"00000000",
    29244 => x"00000000", 29245 => x"00000000", 29246 => x"00000000",
    29247 => x"00000000", 29248 => x"00000000", 29249 => x"00000000",
    29250 => x"00000000", 29251 => x"00000000", 29252 => x"00000000",
    29253 => x"00000000", 29254 => x"00000000", 29255 => x"00000000",
    29256 => x"00000000", 29257 => x"00000000", 29258 => x"00000000",
    29259 => x"00000000", 29260 => x"00000000", 29261 => x"00000000",
    29262 => x"00000000", 29263 => x"00000000", 29264 => x"00000000",
    29265 => x"00000000", 29266 => x"00000000", 29267 => x"00000000",
    29268 => x"00000000", 29269 => x"00000000", 29270 => x"00000000",
    29271 => x"00000000", 29272 => x"00000000", 29273 => x"00000000",
    29274 => x"00000000", 29275 => x"00000000", 29276 => x"00000000",
    29277 => x"00000000", 29278 => x"00000000", 29279 => x"00000000",
    29280 => x"00000000", 29281 => x"00000000", 29282 => x"00000000",
    29283 => x"00000000", 29284 => x"00000000", 29285 => x"00000000",
    29286 => x"00000000", 29287 => x"00000000", 29288 => x"00000000",
    29289 => x"00000000", 29290 => x"00000000", 29291 => x"00000000",
    29292 => x"00000000", 29293 => x"00000000", 29294 => x"00000000",
    29295 => x"00000000", 29296 => x"00000000", 29297 => x"00000000",
    29298 => x"00000000", 29299 => x"00000000", 29300 => x"00000000",
    29301 => x"00000000", 29302 => x"00000000", 29303 => x"00000000",
    29304 => x"00000000", 29305 => x"00000000", 29306 => x"00000000",
    29307 => x"00000000", 29308 => x"00000000", 29309 => x"00000000",
    29310 => x"00000000", 29311 => x"00000000", 29312 => x"00000000",
    29313 => x"00000000", 29314 => x"00000000", 29315 => x"00000000",
    29316 => x"00000000", 29317 => x"00000000", 29318 => x"00000000",
    29319 => x"00000000", 29320 => x"00000000", 29321 => x"00000000",
    29322 => x"00000000", 29323 => x"00000000", 29324 => x"00000000",
    29325 => x"00000000", 29326 => x"00000000", 29327 => x"00000000",
    29328 => x"00000000", 29329 => x"00000000", 29330 => x"00000000",
    29331 => x"00000000", 29332 => x"00000000", 29333 => x"00000000",
    29334 => x"00000000", 29335 => x"00000000", 29336 => x"00000000",
    29337 => x"00000000", 29338 => x"00000000", 29339 => x"00000000",
    29340 => x"00000000", 29341 => x"00000000", 29342 => x"00000000",
    29343 => x"00000000", 29344 => x"00000000", 29345 => x"00000000",
    29346 => x"00000000", 29347 => x"00000000", 29348 => x"00000000",
    29349 => x"00000000", 29350 => x"00000000", 29351 => x"00000000",
    29352 => x"00000000", 29353 => x"00000000", 29354 => x"00000000",
    29355 => x"00000000", 29356 => x"00000000", 29357 => x"00000000",
    29358 => x"00000000", 29359 => x"00000000", 29360 => x"00000000",
    29361 => x"00000000", 29362 => x"00000000", 29363 => x"00000000",
    29364 => x"00000000", 29365 => x"00000000", 29366 => x"00000000",
    29367 => x"00000000", 29368 => x"00000000", 29369 => x"00000000",
    29370 => x"00000000", 29371 => x"00000000", 29372 => x"00000000",
    29373 => x"00000000", 29374 => x"00000000", 29375 => x"00000000",
    29376 => x"00000000", 29377 => x"00000000", 29378 => x"00000000",
    29379 => x"00000000", 29380 => x"00000000", 29381 => x"00000000",
    29382 => x"00000000", 29383 => x"00000000", 29384 => x"00000000",
    29385 => x"00000000", 29386 => x"00000000", 29387 => x"00000000",
    29388 => x"00000000", 29389 => x"00000000", 29390 => x"00000000",
    29391 => x"00000000", 29392 => x"00000000", 29393 => x"00000000",
    29394 => x"00000000", 29395 => x"00000000", 29396 => x"00000000",
    29397 => x"00000000", 29398 => x"00000000", 29399 => x"00000000",
    29400 => x"00000000", 29401 => x"00000000", 29402 => x"00000000",
    29403 => x"00000000", 29404 => x"00000000", 29405 => x"00000000",
    29406 => x"00000000", 29407 => x"00000000", 29408 => x"00000000",
    29409 => x"00000000", 29410 => x"00000000", 29411 => x"00000000",
    29412 => x"00000000", 29413 => x"00000000", 29414 => x"00000000",
    29415 => x"00000000", 29416 => x"00000000", 29417 => x"00000000",
    29418 => x"00000000", 29419 => x"00000000", 29420 => x"00000000",
    29421 => x"00000000", 29422 => x"00000000", 29423 => x"00000000",
    29424 => x"00000000", 29425 => x"00000000", 29426 => x"00000000",
    29427 => x"00000000", 29428 => x"00000000", 29429 => x"00000000",
    29430 => x"00000000", 29431 => x"00000000", 29432 => x"00000000",
    29433 => x"00000000", 29434 => x"00000000", 29435 => x"00000000",
    29436 => x"00000000", 29437 => x"00000000", 29438 => x"00000000",
    29439 => x"00000000", 29440 => x"00000000", 29441 => x"00000000",
    29442 => x"00000000", 29443 => x"00000000", 29444 => x"00000000",
    29445 => x"00000000", 29446 => x"00000000", 29447 => x"00000000",
    29448 => x"00000000", 29449 => x"00000000", 29450 => x"00000000",
    29451 => x"00000000", 29452 => x"00000000", 29453 => x"00000000",
    29454 => x"00000000", 29455 => x"00000000", 29456 => x"00000000",
    29457 => x"00000000", 29458 => x"00000000", 29459 => x"00000000",
    29460 => x"00000000", 29461 => x"00000000", 29462 => x"00000000",
    29463 => x"00000000", 29464 => x"00000000", 29465 => x"00000000",
    29466 => x"00000000", 29467 => x"00000000", 29468 => x"00000000",
    29469 => x"00000000", 29470 => x"00000000", 29471 => x"00000000",
    29472 => x"00000000", 29473 => x"00000000", 29474 => x"00000000",
    29475 => x"00000000", 29476 => x"00000000", 29477 => x"00000000",
    29478 => x"00000000", 29479 => x"00000000", 29480 => x"00000000",
    29481 => x"00000000", 29482 => x"00000000", 29483 => x"00000000",
    29484 => x"00000000", 29485 => x"00000000", 29486 => x"00000000",
    29487 => x"00000000", 29488 => x"00000000", 29489 => x"00000000",
    29490 => x"00000000", 29491 => x"00000000", 29492 => x"00000000",
    29493 => x"00000000", 29494 => x"00000000", 29495 => x"00000000",
    29496 => x"00000000", 29497 => x"00000000", 29498 => x"00000000",
    29499 => x"00000000", 29500 => x"00000000", 29501 => x"00000000",
    29502 => x"00000000", 29503 => x"00000000", 29504 => x"00000000",
    29505 => x"00000000", 29506 => x"00000000", 29507 => x"00000000",
    29508 => x"00000000", 29509 => x"00000000", 29510 => x"00000000",
    29511 => x"00000000", 29512 => x"00000000", 29513 => x"00000000",
    29514 => x"00000000", 29515 => x"00000000", 29516 => x"00000000",
    29517 => x"00000000", 29518 => x"00000000", 29519 => x"00000000",
    29520 => x"00000000", 29521 => x"00000000", 29522 => x"00000000",
    29523 => x"00000000", 29524 => x"00000000", 29525 => x"00000000",
    29526 => x"00000000", 29527 => x"00000000", 29528 => x"00000000",
    29529 => x"00000000", 29530 => x"00000000", 29531 => x"00000000",
    29532 => x"00000000", 29533 => x"00000000", 29534 => x"00000000",
    29535 => x"00000000", 29536 => x"00000000", 29537 => x"00000000",
    29538 => x"00000000", 29539 => x"00000000", 29540 => x"00000000",
    29541 => x"00000000", 29542 => x"00000000", 29543 => x"00000000",
    29544 => x"00000000", 29545 => x"00000000", 29546 => x"00000000",
    29547 => x"00000000", 29548 => x"00000000", 29549 => x"00000000",
    29550 => x"00000000", 29551 => x"00000000", 29552 => x"00000000",
    29553 => x"00000000", 29554 => x"00000000", 29555 => x"00000000",
    29556 => x"00000000", 29557 => x"00000000", 29558 => x"00000000",
    29559 => x"00000000", 29560 => x"00000000", 29561 => x"00000000",
    29562 => x"00000000", 29563 => x"00000000", 29564 => x"00000000",
    29565 => x"00000000", 29566 => x"00000000", 29567 => x"00000000",
    29568 => x"00000000", 29569 => x"00000000", 29570 => x"00000000",
    29571 => x"00000000", 29572 => x"00000000", 29573 => x"00000000",
    29574 => x"00000000", 29575 => x"00000000", 29576 => x"00000000",
    29577 => x"00000000", 29578 => x"00000000", 29579 => x"00000000",
    29580 => x"00000000", 29581 => x"00000000", 29582 => x"00000000",
    29583 => x"00000000", 29584 => x"00000000", 29585 => x"00000000",
    29586 => x"00000000", 29587 => x"00000000", 29588 => x"00000000",
    29589 => x"00000000", 29590 => x"00000000", 29591 => x"00000000",
    29592 => x"00000000", 29593 => x"00000000", 29594 => x"00000000",
    29595 => x"00000000", 29596 => x"00000000", 29597 => x"00000000",
    29598 => x"00000000", 29599 => x"00000000", 29600 => x"00000000",
    29601 => x"00000000", 29602 => x"00000000", 29603 => x"00000000",
    29604 => x"00000000", 29605 => x"00000000", 29606 => x"00000000",
    29607 => x"00000000", 29608 => x"00000000", 29609 => x"00000000",
    29610 => x"00000000", 29611 => x"00000000", 29612 => x"00000000",
    29613 => x"00000000", 29614 => x"00000000", 29615 => x"00000000",
    29616 => x"00000000", 29617 => x"00000000", 29618 => x"00000000",
    29619 => x"00000000", 29620 => x"00000000", 29621 => x"00000000",
    29622 => x"00000000", 29623 => x"00000000", 29624 => x"00000000",
    29625 => x"00000000", 29626 => x"00000000", 29627 => x"00000000",
    29628 => x"00000000", 29629 => x"00000000", 29630 => x"00000000",
    29631 => x"00000000", 29632 => x"00000000", 29633 => x"00000000",
    29634 => x"00000000", 29635 => x"00000000", 29636 => x"00000000",
    29637 => x"00000000", 29638 => x"00000000", 29639 => x"00000000",
    29640 => x"00000000", 29641 => x"00000000", 29642 => x"00000000",
    29643 => x"00000000", 29644 => x"00000000", 29645 => x"00000000",
    29646 => x"00000000", 29647 => x"00000000", 29648 => x"00000000",
    29649 => x"00000000", 29650 => x"00000000", 29651 => x"00000000",
    29652 => x"00000000", 29653 => x"00000000", 29654 => x"00000000",
    29655 => x"00000000", 29656 => x"00000000", 29657 => x"00000000",
    29658 => x"00000000", 29659 => x"00000000", 29660 => x"00000000",
    29661 => x"00000000", 29662 => x"00000000", 29663 => x"00000000",
    29664 => x"00000000", 29665 => x"00000000", 29666 => x"00000000",
    29667 => x"00000000", 29668 => x"00000000", 29669 => x"00000000",
    29670 => x"00000000", 29671 => x"00000000", 29672 => x"00000000",
    29673 => x"00000000", 29674 => x"00000000", 29675 => x"00000000",
    29676 => x"00000000", 29677 => x"00000000", 29678 => x"00000000",
    29679 => x"00000000", 29680 => x"00000000", 29681 => x"00000000",
    29682 => x"00000000", 29683 => x"00000000", 29684 => x"00000000",
    29685 => x"00000000", 29686 => x"00000000", 29687 => x"00000000",
    29688 => x"00000000", 29689 => x"00000000", 29690 => x"00000000",
    29691 => x"00000000", 29692 => x"00000000", 29693 => x"00000000",
    29694 => x"00000000", 29695 => x"00000000", 29696 => x"00000000",
    29697 => x"00000000", 29698 => x"00000000", 29699 => x"00000000",
    29700 => x"00000000", 29701 => x"00000000", 29702 => x"00000000",
    29703 => x"00000000", 29704 => x"00000000", 29705 => x"00000000",
    29706 => x"00000000", 29707 => x"00000000", 29708 => x"00000000",
    29709 => x"00000000", 29710 => x"00000000", 29711 => x"00000000",
    29712 => x"00000000", 29713 => x"00000000", 29714 => x"00000000",
    29715 => x"00000000", 29716 => x"00000000", 29717 => x"00000000",
    29718 => x"00000000", 29719 => x"00000000", 29720 => x"00000000",
    29721 => x"00000000", 29722 => x"00000000", 29723 => x"00000000",
    29724 => x"00000000", 29725 => x"00000000", 29726 => x"00000000",
    29727 => x"00000000", 29728 => x"00000000", 29729 => x"00000000",
    29730 => x"00000000", 29731 => x"00000000", 29732 => x"00000000",
    29733 => x"00000000", 29734 => x"00000000", 29735 => x"00000000",
    29736 => x"00000000", 29737 => x"00000000", 29738 => x"00000000",
    29739 => x"00000000", 29740 => x"00000000", 29741 => x"00000000",
    29742 => x"00000000", 29743 => x"00000000", 29744 => x"00000000",
    29745 => x"00000000", 29746 => x"00000000", 29747 => x"00000000",
    29748 => x"00000000", 29749 => x"00000000", 29750 => x"00000000",
    29751 => x"00000000", 29752 => x"00000000", 29753 => x"00000000",
    29754 => x"00000000", 29755 => x"00000000", 29756 => x"00000000",
    29757 => x"00000000", 29758 => x"00000000", 29759 => x"00000000",
    29760 => x"00000000", 29761 => x"00000000", 29762 => x"00000000",
    29763 => x"00000000", 29764 => x"00000000", 29765 => x"00000000",
    29766 => x"00000000", 29767 => x"00000000", 29768 => x"00000000",
    29769 => x"00000000", 29770 => x"00000000", 29771 => x"00000000",
    29772 => x"00000000", 29773 => x"00000000", 29774 => x"00000000",
    29775 => x"00000000", 29776 => x"00000000", 29777 => x"00000000",
    29778 => x"00000000", 29779 => x"00000000", 29780 => x"00000000",
    29781 => x"00000000", 29782 => x"00000000", 29783 => x"00000000",
    29784 => x"00000000", 29785 => x"00000000", 29786 => x"00000000",
    29787 => x"00000000", 29788 => x"00000000", 29789 => x"00000000",
    29790 => x"00000000", 29791 => x"00000000", 29792 => x"00000000",
    29793 => x"00000000", 29794 => x"00000000", 29795 => x"00000000",
    29796 => x"00000000", 29797 => x"00000000", 29798 => x"00000000",
    29799 => x"00000000", 29800 => x"00000000", 29801 => x"00000000",
    29802 => x"00000000", 29803 => x"00000000", 29804 => x"00000000",
    29805 => x"00000000", 29806 => x"00000000", 29807 => x"00000000",
    29808 => x"00000000", 29809 => x"00000000", 29810 => x"00000000",
    29811 => x"00000000", 29812 => x"00000000", 29813 => x"00000000",
    29814 => x"00000000", 29815 => x"00000000", 29816 => x"00000000",
    29817 => x"00000000", 29818 => x"00000000", 29819 => x"00000000",
    29820 => x"00000000", 29821 => x"00000000", 29822 => x"00000000",
    29823 => x"00000000", 29824 => x"00000000", 29825 => x"00000000",
    29826 => x"00000000", 29827 => x"00000000", 29828 => x"00000000",
    29829 => x"00000000", 29830 => x"00000000", 29831 => x"00000000",
    29832 => x"00000000", 29833 => x"00000000", 29834 => x"00000000",
    29835 => x"00000000", 29836 => x"00000000", 29837 => x"00000000",
    29838 => x"00000000", 29839 => x"00000000", 29840 => x"00000000",
    29841 => x"00000000", 29842 => x"00000000", 29843 => x"00000000",
    29844 => x"00000000", 29845 => x"00000000", 29846 => x"00000000",
    29847 => x"00000000", 29848 => x"00000000", 29849 => x"00000000",
    29850 => x"00000000", 29851 => x"00000000", 29852 => x"00000000",
    29853 => x"00000000", 29854 => x"00000000", 29855 => x"00000000",
    29856 => x"00000000", 29857 => x"00000000", 29858 => x"00000000",
    29859 => x"00000000", 29860 => x"00000000", 29861 => x"00000000",
    29862 => x"00000000", 29863 => x"00000000", 29864 => x"00000000",
    29865 => x"00000000", 29866 => x"00000000", 29867 => x"00000000",
    29868 => x"00000000", 29869 => x"00000000", 29870 => x"00000000",
    29871 => x"00000000", 29872 => x"00000000", 29873 => x"00000000",
    29874 => x"00000000", 29875 => x"00000000", 29876 => x"00000000",
    29877 => x"00000000", 29878 => x"00000000", 29879 => x"00000000",
    29880 => x"00000000", 29881 => x"00000000", 29882 => x"00000000",
    29883 => x"00000000", 29884 => x"00000000", 29885 => x"00000000",
    29886 => x"00000000", 29887 => x"00000000", 29888 => x"00000000",
    29889 => x"00000000", 29890 => x"00000000", 29891 => x"00000000",
    29892 => x"00000000", 29893 => x"00000000", 29894 => x"00000000",
    29895 => x"00000000", 29896 => x"00000000", 29897 => x"00000000",
    29898 => x"00000000", 29899 => x"00000000", 29900 => x"00000000",
    29901 => x"00000000", 29902 => x"00000000", 29903 => x"00000000",
    29904 => x"00000000", 29905 => x"00000000", 29906 => x"00000000",
    29907 => x"00000000", 29908 => x"00000000", 29909 => x"00000000",
    29910 => x"00000000", 29911 => x"00000000", 29912 => x"00000000",
    29913 => x"00000000", 29914 => x"00000000", 29915 => x"00000000",
    29916 => x"00000000", 29917 => x"00000000", 29918 => x"00000000",
    29919 => x"00000000", 29920 => x"00000000", 29921 => x"00000000",
    29922 => x"00000000", 29923 => x"00000000", 29924 => x"00000000",
    29925 => x"00000000", 29926 => x"00000000", 29927 => x"00000000",
    29928 => x"00000000", 29929 => x"00000000", 29930 => x"00000000",
    29931 => x"00000000", 29932 => x"00000000", 29933 => x"00000000",
    29934 => x"00000000", 29935 => x"00000000", 29936 => x"00000000",
    29937 => x"00000000", 29938 => x"00000000", 29939 => x"00000000",
    29940 => x"00000000", 29941 => x"00000000", 29942 => x"00000000",
    29943 => x"00000000", 29944 => x"00000000", 29945 => x"00000000",
    29946 => x"00000000", 29947 => x"00000000", 29948 => x"00000000",
    29949 => x"00000000", 29950 => x"00000000", 29951 => x"00000000",
    29952 => x"00000000", 29953 => x"00000000", 29954 => x"00000000",
    29955 => x"00000000", 29956 => x"00000000", 29957 => x"00000000",
    29958 => x"00000000", 29959 => x"00000000", 29960 => x"00000000",
    29961 => x"00000000", 29962 => x"00000000", 29963 => x"00000000",
    29964 => x"00000000", 29965 => x"00000000", 29966 => x"00000000",
    29967 => x"00000000", 29968 => x"00000000", 29969 => x"00000000",
    29970 => x"00000000", 29971 => x"00000000", 29972 => x"00000000",
    29973 => x"00000000", 29974 => x"00000000", 29975 => x"00000000",
    29976 => x"00000000", 29977 => x"00000000", 29978 => x"00000000",
    29979 => x"00000000", 29980 => x"00000000", 29981 => x"00000000",
    29982 => x"00000000", 29983 => x"00000000", 29984 => x"00000000",
    29985 => x"00000000", 29986 => x"00000000", 29987 => x"00000000",
    29988 => x"00000000", 29989 => x"00000000", 29990 => x"00000000",
    29991 => x"00000000", 29992 => x"00000000", 29993 => x"00000000",
    29994 => x"00000000", 29995 => x"00000000", 29996 => x"00000000",
    29997 => x"00000000", 29998 => x"00000000", 29999 => x"00000000",
    30000 => x"00000000", 30001 => x"00000000", 30002 => x"00000000",
    30003 => x"00000000", 30004 => x"00000000", 30005 => x"00000000",
    30006 => x"00000000", 30007 => x"00000000", 30008 => x"00000000",
    30009 => x"00000000", 30010 => x"00000000", 30011 => x"00000000",
    30012 => x"00000000", 30013 => x"00000000", 30014 => x"00000000",
    30015 => x"00000000", 30016 => x"00000000", 30017 => x"00000000",
    30018 => x"00000000", 30019 => x"00000000", 30020 => x"00000000",
    30021 => x"00000000", 30022 => x"00000000", 30023 => x"00000000",
    30024 => x"00000000", 30025 => x"00000000", 30026 => x"00000000",
    30027 => x"00000000", 30028 => x"00000000", 30029 => x"00000000",
    30030 => x"00000000", 30031 => x"00000000", 30032 => x"00000000",
    30033 => x"00000000", 30034 => x"00000000", 30035 => x"00000000",
    30036 => x"00000000", 30037 => x"00000000", 30038 => x"00000000",
    30039 => x"00000000", 30040 => x"00000000", 30041 => x"00000000",
    30042 => x"00000000", 30043 => x"00000000", 30044 => x"00000000",
    30045 => x"00000000", 30046 => x"00000000", 30047 => x"00000000",
    30048 => x"00000000", 30049 => x"00000000", 30050 => x"00000000",
    30051 => x"00000000", 30052 => x"00000000", 30053 => x"00000000",
    30054 => x"00000000", 30055 => x"00000000", 30056 => x"00000000",
    30057 => x"00000000", 30058 => x"00000000", 30059 => x"00000000",
    30060 => x"00000000", 30061 => x"00000000", 30062 => x"00000000",
    30063 => x"00000000", 30064 => x"00000000", 30065 => x"00000000",
    30066 => x"00000000", 30067 => x"00000000", 30068 => x"00000000",
    30069 => x"00000000", 30070 => x"00000000", 30071 => x"00000000",
    30072 => x"00000000", 30073 => x"00000000", 30074 => x"00000000",
    30075 => x"00000000", 30076 => x"00000000", 30077 => x"00000000",
    30078 => x"00000000", 30079 => x"00000000", 30080 => x"00000000",
    30081 => x"00000000", 30082 => x"00000000", 30083 => x"00000000",
    30084 => x"00000000", 30085 => x"00000000", 30086 => x"00000000",
    30087 => x"00000000", 30088 => x"00000000", 30089 => x"00000000",
    30090 => x"00000000", 30091 => x"00000000", 30092 => x"00000000",
    30093 => x"00000000", 30094 => x"00000000", 30095 => x"00000000",
    30096 => x"00000000", 30097 => x"00000000", 30098 => x"00000000",
    30099 => x"00000000", 30100 => x"00000000", 30101 => x"00000000",
    30102 => x"00000000", 30103 => x"00000000", 30104 => x"00000000",
    30105 => x"00000000", 30106 => x"00000000", 30107 => x"00000000",
    30108 => x"00000000", 30109 => x"00000000", 30110 => x"00000000",
    30111 => x"00000000", 30112 => x"00000000", 30113 => x"00000000",
    30114 => x"00000000", 30115 => x"00000000", 30116 => x"00000000",
    30117 => x"00000000", 30118 => x"00000000", 30119 => x"00000000",
    30120 => x"00000000", 30121 => x"00000000", 30122 => x"00000000",
    30123 => x"00000000", 30124 => x"00000000", 30125 => x"00000000",
    30126 => x"00000000", 30127 => x"00000000", 30128 => x"00000000",
    30129 => x"00000000", 30130 => x"00000000", 30131 => x"00000000",
    30132 => x"00000000", 30133 => x"00000000", 30134 => x"00000000",
    30135 => x"00000000", 30136 => x"00000000", 30137 => x"00000000",
    30138 => x"00000000", 30139 => x"00000000", 30140 => x"00000000",
    30141 => x"00000000", 30142 => x"00000000", 30143 => x"00000000",
    30144 => x"00000000", 30145 => x"00000000", 30146 => x"00000000",
    30147 => x"00000000", 30148 => x"00000000", 30149 => x"00000000",
    30150 => x"00000000", 30151 => x"00000000", 30152 => x"00000000",
    30153 => x"00000000", 30154 => x"00000000", 30155 => x"00000000",
    30156 => x"00000000", 30157 => x"00000000", 30158 => x"00000000",
    30159 => x"00000000", 30160 => x"00000000", 30161 => x"00000000",
    30162 => x"00000000", 30163 => x"00000000", 30164 => x"00000000",
    30165 => x"00000000", 30166 => x"00000000", 30167 => x"00000000",
    30168 => x"00000000", 30169 => x"00000000", 30170 => x"00000000",
    30171 => x"00000000", 30172 => x"00000000", 30173 => x"00000000",
    30174 => x"00000000", 30175 => x"00000000", 30176 => x"00000000",
    30177 => x"00000000", 30178 => x"00000000", 30179 => x"00000000",
    30180 => x"00000000", 30181 => x"00000000", 30182 => x"00000000",
    30183 => x"00000000", 30184 => x"00000000", 30185 => x"00000000",
    30186 => x"00000000", 30187 => x"00000000", 30188 => x"00000000",
    30189 => x"00000000", 30190 => x"00000000", 30191 => x"00000000",
    30192 => x"00000000", 30193 => x"00000000", 30194 => x"00000000",
    30195 => x"00000000", 30196 => x"00000000", 30197 => x"00000000",
    30198 => x"00000000", 30199 => x"00000000", 30200 => x"00000000",
    30201 => x"00000000", 30202 => x"00000000", 30203 => x"00000000",
    30204 => x"00000000", 30205 => x"00000000", 30206 => x"00000000",
    30207 => x"00000000", 30208 => x"00000000", 30209 => x"00000000",
    30210 => x"00000000", 30211 => x"00000000", 30212 => x"00000000",
    30213 => x"00000000", 30214 => x"00000000", 30215 => x"00000000",
    30216 => x"00000000", 30217 => x"00000000", 30218 => x"00000000",
    30219 => x"00000000", 30220 => x"00000000", 30221 => x"00000000",
    30222 => x"00000000", 30223 => x"00000000", 30224 => x"00000000",
    30225 => x"00000000", 30226 => x"00000000", 30227 => x"00000000",
    30228 => x"00000000", 30229 => x"00000000", 30230 => x"00000000",
    30231 => x"00000000", 30232 => x"00000000", 30233 => x"00000000",
    30234 => x"00000000", 30235 => x"00000000", 30236 => x"00000000",
    30237 => x"00000000", 30238 => x"00000000", 30239 => x"00000000",
    30240 => x"00000000", 30241 => x"00000000", 30242 => x"00000000",
    30243 => x"00000000", 30244 => x"00000000", 30245 => x"00000000",
    30246 => x"00000000", 30247 => x"00000000", 30248 => x"00000000",
    30249 => x"00000000", 30250 => x"00000000", 30251 => x"00000000",
    30252 => x"00000000", 30253 => x"00000000", 30254 => x"00000000",
    30255 => x"00000000", 30256 => x"00000000", 30257 => x"00000000",
    30258 => x"00000000", 30259 => x"00000000", 30260 => x"00000000",
    30261 => x"00000000", 30262 => x"00000000", 30263 => x"00000000",
    30264 => x"00000000", 30265 => x"00000000", 30266 => x"00000000",
    30267 => x"00000000", 30268 => x"00000000", 30269 => x"00000000",
    30270 => x"00000000", 30271 => x"00000000", 30272 => x"00000000",
    30273 => x"00000000", 30274 => x"00000000", 30275 => x"00000000",
    30276 => x"00000000", 30277 => x"00000000", 30278 => x"00000000",
    30279 => x"00000000", 30280 => x"00000000", 30281 => x"00000000",
    30282 => x"00000000", 30283 => x"00000000", 30284 => x"00000000",
    30285 => x"00000000", 30286 => x"00000000", 30287 => x"00000000",
    30288 => x"00000000", 30289 => x"00000000", 30290 => x"00000000",
    30291 => x"00000000", 30292 => x"00000000", 30293 => x"00000000",
    30294 => x"00000000", 30295 => x"00000000", 30296 => x"00000000",
    30297 => x"00000000", 30298 => x"00000000", 30299 => x"00000000",
    30300 => x"00000000", 30301 => x"00000000", 30302 => x"00000000",
    30303 => x"00000000", 30304 => x"00000000", 30305 => x"00000000",
    30306 => x"00000000", 30307 => x"00000000", 30308 => x"00000000",
    30309 => x"00000000", 30310 => x"00000000", 30311 => x"00000000",
    30312 => x"00000000", 30313 => x"00000000", 30314 => x"00000000",
    30315 => x"00000000", 30316 => x"00000000", 30317 => x"00000000",
    30318 => x"00000000", 30319 => x"00000000", 30320 => x"00000000",
    30321 => x"00000000", 30322 => x"00000000", 30323 => x"00000000",
    30324 => x"00000000", 30325 => x"00000000", 30326 => x"00000000",
    30327 => x"00000000", 30328 => x"00000000", 30329 => x"00000000",
    30330 => x"00000000", 30331 => x"00000000", 30332 => x"00000000",
    30333 => x"00000000", 30334 => x"00000000", 30335 => x"00000000",
    30336 => x"00000000", 30337 => x"00000000", 30338 => x"00000000",
    30339 => x"00000000", 30340 => x"00000000", 30341 => x"00000000",
    30342 => x"00000000", 30343 => x"00000000", 30344 => x"00000000",
    30345 => x"00000000", 30346 => x"00000000", 30347 => x"00000000",
    30348 => x"00000000", 30349 => x"00000000", 30350 => x"00000000",
    30351 => x"00000000", 30352 => x"00000000", 30353 => x"00000000",
    30354 => x"00000000", 30355 => x"00000000", 30356 => x"00000000",
    30357 => x"00000000", 30358 => x"00000000", 30359 => x"00000000",
    30360 => x"00000000", 30361 => x"00000000", 30362 => x"00000000",
    30363 => x"00000000", 30364 => x"00000000", 30365 => x"00000000",
    30366 => x"00000000", 30367 => x"00000000", 30368 => x"00000000",
    30369 => x"00000000", 30370 => x"00000000", 30371 => x"00000000",
    30372 => x"00000000", 30373 => x"00000000", 30374 => x"00000000",
    30375 => x"00000000", 30376 => x"00000000", 30377 => x"00000000",
    30378 => x"00000000", 30379 => x"00000000", 30380 => x"00000000",
    30381 => x"00000000", 30382 => x"00000000", 30383 => x"00000000",
    30384 => x"00000000", 30385 => x"00000000", 30386 => x"00000000",
    30387 => x"00000000", 30388 => x"00000000", 30389 => x"00000000",
    30390 => x"00000000", 30391 => x"00000000", 30392 => x"00000000",
    30393 => x"00000000", 30394 => x"00000000", 30395 => x"00000000",
    30396 => x"00000000", 30397 => x"00000000", 30398 => x"00000000",
    30399 => x"00000000", 30400 => x"00000000", 30401 => x"00000000",
    30402 => x"00000000", 30403 => x"00000000", 30404 => x"00000000",
    30405 => x"00000000", 30406 => x"00000000", 30407 => x"00000000",
    30408 => x"00000000", 30409 => x"00000000", 30410 => x"00000000",
    30411 => x"00000000", 30412 => x"00000000", 30413 => x"00000000",
    30414 => x"00000000", 30415 => x"00000000", 30416 => x"00000000",
    30417 => x"00000000", 30418 => x"00000000", 30419 => x"00000000",
    30420 => x"00000000", 30421 => x"00000000", 30422 => x"00000000",
    30423 => x"00000000", 30424 => x"00000000", 30425 => x"00000000",
    30426 => x"00000000", 30427 => x"00000000", 30428 => x"00000000",
    30429 => x"00000000", 30430 => x"00000000", 30431 => x"00000000",
    30432 => x"00000000", 30433 => x"00000000", 30434 => x"00000000",
    30435 => x"00000000", 30436 => x"00000000", 30437 => x"00000000",
    30438 => x"00000000", 30439 => x"00000000", 30440 => x"00000000",
    30441 => x"00000000", 30442 => x"00000000", 30443 => x"00000000",
    30444 => x"00000000", 30445 => x"00000000", 30446 => x"00000000",
    30447 => x"00000000", 30448 => x"00000000", 30449 => x"00000000",
    30450 => x"00000000", 30451 => x"00000000", 30452 => x"00000000",
    30453 => x"00000000", 30454 => x"00000000", 30455 => x"00000000",
    30456 => x"00000000", 30457 => x"00000000", 30458 => x"00000000",
    30459 => x"00000000", 30460 => x"00000000", 30461 => x"00000000",
    30462 => x"00000000", 30463 => x"00000000", 30464 => x"00000000",
    30465 => x"00000000", 30466 => x"00000000", 30467 => x"00000000",
    30468 => x"00000000", 30469 => x"00000000", 30470 => x"00000000",
    30471 => x"00000000", 30472 => x"00000000", 30473 => x"00000000",
    30474 => x"00000000", 30475 => x"00000000", 30476 => x"00000000",
    30477 => x"00000000", 30478 => x"00000000", 30479 => x"00000000",
    30480 => x"00000000", 30481 => x"00000000", 30482 => x"00000000",
    30483 => x"00000000", 30484 => x"00000000", 30485 => x"00000000",
    30486 => x"00000000", 30487 => x"00000000", 30488 => x"00000000",
    30489 => x"00000000", 30490 => x"00000000", 30491 => x"00000000",
    30492 => x"00000000", 30493 => x"00000000", 30494 => x"00000000",
    30495 => x"00000000", 30496 => x"00000000", 30497 => x"00000000",
    30498 => x"00000000", 30499 => x"00000000", 30500 => x"00000000",
    30501 => x"00000000", 30502 => x"00000000", 30503 => x"00000000",
    30504 => x"00000000", 30505 => x"00000000", 30506 => x"00000000",
    30507 => x"00000000", 30508 => x"00000000", 30509 => x"00000000",
    30510 => x"00000000", 30511 => x"00000000", 30512 => x"00000000",
    30513 => x"00000000", 30514 => x"00000000", 30515 => x"00000000",
    30516 => x"00000000", 30517 => x"00000000", 30518 => x"00000000",
    30519 => x"00000000", 30520 => x"00000000", 30521 => x"00000000",
    30522 => x"00000000", 30523 => x"00000000", 30524 => x"00000000",
    30525 => x"00000000", 30526 => x"00000000", 30527 => x"00000000",
    30528 => x"00000000", 30529 => x"00000000", 30530 => x"00000000",
    30531 => x"00000000", 30532 => x"00000000", 30533 => x"00000000",
    30534 => x"00000000", 30535 => x"00000000", 30536 => x"00000000",
    30537 => x"00000000", 30538 => x"00000000", 30539 => x"00000000",
    30540 => x"00000000", 30541 => x"00000000", 30542 => x"00000000",
    30543 => x"00000000", 30544 => x"00000000", 30545 => x"00000000",
    30546 => x"00000000", 30547 => x"00000000", 30548 => x"00000000",
    30549 => x"00000000", 30550 => x"00000000", 30551 => x"00000000",
    30552 => x"00000000", 30553 => x"00000000", 30554 => x"00000000",
    30555 => x"00000000", 30556 => x"00000000", 30557 => x"00000000",
    30558 => x"00000000", 30559 => x"00000000", 30560 => x"00000000",
    30561 => x"00000000", 30562 => x"00000000", 30563 => x"00000000",
    30564 => x"00000000", 30565 => x"00000000", 30566 => x"00000000",
    30567 => x"00000000", 30568 => x"00000000", 30569 => x"00000000",
    30570 => x"00000000", 30571 => x"00000000", 30572 => x"00000000",
    30573 => x"00000000", 30574 => x"00000000", 30575 => x"00000000",
    30576 => x"00000000", 30577 => x"00000000", 30578 => x"00000000",
    30579 => x"00000000", 30580 => x"00000000", 30581 => x"00000000",
    30582 => x"00000000", 30583 => x"00000000", 30584 => x"00000000",
    30585 => x"00000000", 30586 => x"00000000", 30587 => x"00000000",
    30588 => x"00000000", 30589 => x"00000000", 30590 => x"00000000",
    30591 => x"00000000", 30592 => x"00000000", 30593 => x"00000000",
    30594 => x"00000000", 30595 => x"00000000", 30596 => x"00000000",
    30597 => x"00000000", 30598 => x"00000000", 30599 => x"00000000",
    30600 => x"00000000", 30601 => x"00000000", 30602 => x"00000000",
    30603 => x"00000000", 30604 => x"00000000", 30605 => x"00000000",
    30606 => x"00000000", 30607 => x"00000000", 30608 => x"00000000",
    30609 => x"00000000", 30610 => x"00000000", 30611 => x"00000000",
    30612 => x"00000000", 30613 => x"00000000", 30614 => x"00000000",
    30615 => x"00000000", 30616 => x"00000000", 30617 => x"00000000",
    30618 => x"00000000", 30619 => x"00000000", 30620 => x"00000000",
    30621 => x"00000000", 30622 => x"00000000", 30623 => x"00000000",
    30624 => x"00000000", 30625 => x"00000000", 30626 => x"00000000",
    30627 => x"00000000", 30628 => x"00000000", 30629 => x"00000000",
    30630 => x"00000000", 30631 => x"00000000", 30632 => x"00000000",
    30633 => x"00000000", 30634 => x"00000000", 30635 => x"00000000",
    30636 => x"00000000", 30637 => x"00000000", 30638 => x"00000000",
    30639 => x"00000000", 30640 => x"00000000", 30641 => x"00000000",
    30642 => x"00000000", 30643 => x"00000000", 30644 => x"00000000",
    30645 => x"00000000", 30646 => x"00000000", 30647 => x"00000000",
    30648 => x"00000000", 30649 => x"00000000", 30650 => x"00000000",
    30651 => x"00000000", 30652 => x"00000000", 30653 => x"00000000",
    30654 => x"00000000", 30655 => x"00000000", 30656 => x"00000000",
    30657 => x"00000000", 30658 => x"00000000", 30659 => x"00000000",
    30660 => x"00000000", 30661 => x"00000000", 30662 => x"00000000",
    30663 => x"00000000", 30664 => x"00000000", 30665 => x"00000000",
    30666 => x"00000000", 30667 => x"00000000", 30668 => x"00000000",
    30669 => x"00000000", 30670 => x"00000000", 30671 => x"00000000",
    30672 => x"00000000", 30673 => x"00000000", 30674 => x"00000000",
    30675 => x"00000000", 30676 => x"00000000", 30677 => x"00000000",
    30678 => x"00000000", 30679 => x"00000000", 30680 => x"00000000",
    30681 => x"00000000", 30682 => x"00000000", 30683 => x"00000000",
    30684 => x"00000000", 30685 => x"00000000", 30686 => x"00000000",
    30687 => x"00000000", 30688 => x"00000000", 30689 => x"00000000",
    30690 => x"00000000", 30691 => x"00000000", 30692 => x"00000000",
    30693 => x"00000000", 30694 => x"00000000", 30695 => x"00000000",
    30696 => x"00000000", 30697 => x"00000000", 30698 => x"00000000",
    30699 => x"00000000", 30700 => x"00000000", 30701 => x"00000000",
    30702 => x"00000000", 30703 => x"00000000", 30704 => x"00000000",
    30705 => x"00000000", 30706 => x"00000000", 30707 => x"00000000",
    30708 => x"00000000", 30709 => x"00000000", 30710 => x"00000000",
    30711 => x"00000000", 30712 => x"00000000", 30713 => x"00000000",
    30714 => x"00000000", 30715 => x"00000000", 30716 => x"00000000",
    30717 => x"00000000", 30718 => x"00000000", 30719 => x"00000000",
    30720 => x"00000000", 30721 => x"00000000", 30722 => x"00000000",
    30723 => x"00000000", 30724 => x"00000000", 30725 => x"00000000",
    30726 => x"00000000", 30727 => x"00000000", 30728 => x"00000000",
    30729 => x"00000000", 30730 => x"00000000", 30731 => x"00000000",
    30732 => x"00000000", 30733 => x"00000000", 30734 => x"00000000",
    30735 => x"00000000", 30736 => x"00000000", 30737 => x"00000000",
    30738 => x"00000000", 30739 => x"00000000", 30740 => x"00000000",
    30741 => x"00000000", 30742 => x"00000000", 30743 => x"00000000",
    30744 => x"00000000", 30745 => x"00000000", 30746 => x"00000000",
    30747 => x"00000000", 30748 => x"00000000", 30749 => x"00000000",
    30750 => x"00000000", 30751 => x"00000000", 30752 => x"00000000",
    30753 => x"00000000", 30754 => x"00000000", 30755 => x"00000000",
    30756 => x"00000000", 30757 => x"00000000", 30758 => x"00000000",
    30759 => x"00000000", 30760 => x"00000000", 30761 => x"00000000",
    30762 => x"00000000", 30763 => x"00000000", 30764 => x"00000000",
    30765 => x"00000000", 30766 => x"00000000", 30767 => x"00000000",
    30768 => x"00000000", 30769 => x"00000000", 30770 => x"00000000",
    30771 => x"00000000", 30772 => x"00000000", 30773 => x"00000000",
    30774 => x"00000000", 30775 => x"00000000", 30776 => x"00000000",
    30777 => x"00000000", 30778 => x"00000000", 30779 => x"00000000",
    30780 => x"00000000", 30781 => x"00000000", 30782 => x"00000000",
    30783 => x"00000000", 30784 => x"00000000", 30785 => x"00000000",
    30786 => x"00000000", 30787 => x"00000000", 30788 => x"00000000",
    30789 => x"00000000", 30790 => x"00000000", 30791 => x"00000000",
    30792 => x"00000000", 30793 => x"00000000", 30794 => x"00000000",
    30795 => x"00000000", 30796 => x"00000000", 30797 => x"00000000",
    30798 => x"00000000", 30799 => x"00000000", 30800 => x"00000000",
    30801 => x"00000000", 30802 => x"00000000", 30803 => x"00000000",
    30804 => x"00000000", 30805 => x"00000000", 30806 => x"00000000",
    30807 => x"00000000", 30808 => x"00000000", 30809 => x"00000000",
    30810 => x"00000000", 30811 => x"00000000", 30812 => x"00000000",
    30813 => x"00000000", 30814 => x"00000000", 30815 => x"00000000",
    30816 => x"00000000", 30817 => x"00000000", 30818 => x"00000000",
    30819 => x"00000000", 30820 => x"00000000", 30821 => x"00000000",
    30822 => x"00000000", 30823 => x"00000000", 30824 => x"00000000",
    30825 => x"00000000", 30826 => x"00000000", 30827 => x"00000000",
    30828 => x"00000000", 30829 => x"00000000", 30830 => x"00000000",
    30831 => x"00000000", 30832 => x"00000000", 30833 => x"00000000",
    30834 => x"00000000", 30835 => x"00000000", 30836 => x"00000000",
    30837 => x"00000000", 30838 => x"00000000", 30839 => x"00000000",
    30840 => x"00000000", 30841 => x"00000000", 30842 => x"00000000",
    30843 => x"00000000", 30844 => x"00000000", 30845 => x"00000000",
    30846 => x"00000000", 30847 => x"00000000", 30848 => x"00000000",
    30849 => x"00000000", 30850 => x"00000000", 30851 => x"00000000",
    30852 => x"00000000", 30853 => x"00000000", 30854 => x"00000000",
    30855 => x"00000000", 30856 => x"00000000", 30857 => x"00000000",
    30858 => x"00000000", 30859 => x"00000000", 30860 => x"00000000",
    30861 => x"00000000", 30862 => x"00000000", 30863 => x"00000000",
    30864 => x"00000000", 30865 => x"00000000", 30866 => x"00000000",
    30867 => x"00000000", 30868 => x"00000000", 30869 => x"00000000",
    30870 => x"00000000", 30871 => x"00000000", 30872 => x"00000000",
    30873 => x"00000000", 30874 => x"00000000", 30875 => x"00000000",
    30876 => x"00000000", 30877 => x"00000000", 30878 => x"00000000",
    30879 => x"00000000", 30880 => x"00000000", 30881 => x"00000000",
    30882 => x"00000000", 30883 => x"00000000", 30884 => x"00000000",
    30885 => x"00000000", 30886 => x"00000000", 30887 => x"00000000",
    30888 => x"00000000", 30889 => x"00000000", 30890 => x"00000000",
    30891 => x"00000000", 30892 => x"00000000", 30893 => x"00000000",
    30894 => x"00000000", 30895 => x"00000000", 30896 => x"00000000",
    30897 => x"00000000", 30898 => x"00000000", 30899 => x"00000000",
    30900 => x"00000000", 30901 => x"00000000", 30902 => x"00000000",
    30903 => x"00000000", 30904 => x"00000000", 30905 => x"00000000",
    30906 => x"00000000", 30907 => x"00000000", 30908 => x"00000000",
    30909 => x"00000000", 30910 => x"00000000", 30911 => x"00000000",
    30912 => x"00000000", 30913 => x"00000000", 30914 => x"00000000",
    30915 => x"00000000", 30916 => x"00000000", 30917 => x"00000000",
    30918 => x"00000000", 30919 => x"00000000", 30920 => x"00000000",
    30921 => x"00000000", 30922 => x"00000000", 30923 => x"00000000",
    30924 => x"00000000", 30925 => x"00000000", 30926 => x"00000000",
    30927 => x"00000000", 30928 => x"00000000", 30929 => x"00000000",
    30930 => x"00000000", 30931 => x"00000000", 30932 => x"00000000",
    30933 => x"00000000", 30934 => x"00000000", 30935 => x"00000000",
    30936 => x"00000000", 30937 => x"00000000", 30938 => x"00000000",
    30939 => x"00000000", 30940 => x"00000000", 30941 => x"00000000",
    30942 => x"00000000", 30943 => x"00000000", 30944 => x"00000000",
    30945 => x"00000000", 30946 => x"00000000", 30947 => x"00000000",
    30948 => x"00000000", 30949 => x"00000000", 30950 => x"00000000",
    30951 => x"00000000", 30952 => x"00000000", 30953 => x"00000000",
    30954 => x"00000000", 30955 => x"00000000", 30956 => x"00000000",
    30957 => x"00000000", 30958 => x"00000000", 30959 => x"00000000",
    30960 => x"00000000", 30961 => x"00000000", 30962 => x"00000000",
    30963 => x"00000000", 30964 => x"00000000", 30965 => x"00000000",
    30966 => x"00000000", 30967 => x"00000000", 30968 => x"00000000",
    30969 => x"00000000", 30970 => x"00000000", 30971 => x"00000000",
    30972 => x"00000000", 30973 => x"00000000", 30974 => x"00000000",
    30975 => x"00000000", 30976 => x"00000000", 30977 => x"00000000",
    30978 => x"00000000", 30979 => x"00000000", 30980 => x"00000000",
    30981 => x"00000000", 30982 => x"00000000", 30983 => x"00000000",
    30984 => x"00000000", 30985 => x"00000000", 30986 => x"00000000",
    30987 => x"00000000", 30988 => x"00000000", 30989 => x"00000000",
    30990 => x"00000000", 30991 => x"00000000", 30992 => x"00000000",
    30993 => x"00000000", 30994 => x"00000000", 30995 => x"00000000",
    30996 => x"00000000", 30997 => x"00000000", 30998 => x"00000000",
    30999 => x"00000000", 31000 => x"00000000", 31001 => x"00000000",
    31002 => x"00000000", 31003 => x"00000000", 31004 => x"00000000",
    31005 => x"00000000", 31006 => x"00000000", 31007 => x"00000000",
    31008 => x"00000000", 31009 => x"00000000", 31010 => x"00000000",
    31011 => x"00000000", 31012 => x"00000000", 31013 => x"00000000",
    31014 => x"00000000", 31015 => x"00000000", 31016 => x"00000000",
    31017 => x"00000000", 31018 => x"00000000", 31019 => x"00000000",
    31020 => x"00000000", 31021 => x"00000000", 31022 => x"00000000",
    31023 => x"00000000", 31024 => x"00000000", 31025 => x"00000000",
    31026 => x"00000000", 31027 => x"00000000", 31028 => x"00000000",
    31029 => x"00000000", 31030 => x"00000000", 31031 => x"00000000",
    31032 => x"00000000", 31033 => x"00000000", 31034 => x"00000000",
    31035 => x"00000000", 31036 => x"00000000", 31037 => x"00000000",
    31038 => x"00000000", 31039 => x"00000000", 31040 => x"00000000",
    31041 => x"00000000", 31042 => x"00000000", 31043 => x"00000000",
    31044 => x"00000000", 31045 => x"00000000", 31046 => x"00000000",
    31047 => x"00000000", 31048 => x"00000000", 31049 => x"00000000",
    31050 => x"00000000", 31051 => x"00000000", 31052 => x"00000000",
    31053 => x"00000000", 31054 => x"00000000", 31055 => x"00000000",
    31056 => x"00000000", 31057 => x"00000000", 31058 => x"00000000",
    31059 => x"00000000", 31060 => x"00000000", 31061 => x"00000000",
    31062 => x"00000000", 31063 => x"00000000", 31064 => x"00000000",
    31065 => x"00000000", 31066 => x"00000000", 31067 => x"00000000",
    31068 => x"00000000", 31069 => x"00000000", 31070 => x"00000000",
    31071 => x"00000000", 31072 => x"00000000", 31073 => x"00000000",
    31074 => x"00000000", 31075 => x"00000000", 31076 => x"00000000",
    31077 => x"00000000", 31078 => x"00000000", 31079 => x"00000000",
    31080 => x"00000000", 31081 => x"00000000", 31082 => x"00000000",
    31083 => x"00000000", 31084 => x"00000000", 31085 => x"00000000",
    31086 => x"00000000", 31087 => x"00000000", 31088 => x"00000000",
    31089 => x"00000000", 31090 => x"00000000", 31091 => x"00000000",
    31092 => x"00000000", 31093 => x"00000000", 31094 => x"00000000",
    31095 => x"00000000", 31096 => x"00000000", 31097 => x"00000000",
    31098 => x"00000000", 31099 => x"00000000", 31100 => x"00000000",
    31101 => x"00000000", 31102 => x"00000000", 31103 => x"00000000",
    31104 => x"00000000", 31105 => x"00000000", 31106 => x"00000000",
    31107 => x"00000000", 31108 => x"00000000", 31109 => x"00000000",
    31110 => x"00000000", 31111 => x"00000000", 31112 => x"00000000",
    31113 => x"00000000", 31114 => x"00000000", 31115 => x"00000000",
    31116 => x"00000000", 31117 => x"00000000", 31118 => x"00000000",
    31119 => x"00000000", 31120 => x"00000000", 31121 => x"00000000",
    31122 => x"00000000", 31123 => x"00000000", 31124 => x"00000000",
    31125 => x"00000000", 31126 => x"00000000", 31127 => x"00000000",
    31128 => x"00000000", 31129 => x"00000000", 31130 => x"00000000",
    31131 => x"00000000", 31132 => x"00000000", 31133 => x"00000000",
    31134 => x"00000000", 31135 => x"00000000", 31136 => x"00000000",
    31137 => x"00000000", 31138 => x"00000000", 31139 => x"00000000",
    31140 => x"00000000", 31141 => x"00000000", 31142 => x"00000000",
    31143 => x"00000000", 31144 => x"00000000", 31145 => x"00000000",
    31146 => x"00000000", 31147 => x"00000000", 31148 => x"00000000",
    31149 => x"00000000", 31150 => x"00000000", 31151 => x"00000000",
    31152 => x"00000000", 31153 => x"00000000", 31154 => x"00000000",
    31155 => x"00000000", 31156 => x"00000000", 31157 => x"00000000",
    31158 => x"00000000", 31159 => x"00000000", 31160 => x"00000000",
    31161 => x"00000000", 31162 => x"00000000", 31163 => x"00000000",
    31164 => x"00000000", 31165 => x"00000000", 31166 => x"00000000",
    31167 => x"00000000", 31168 => x"00000000", 31169 => x"00000000",
    31170 => x"00000000", 31171 => x"00000000", 31172 => x"00000000",
    31173 => x"00000000", 31174 => x"00000000", 31175 => x"00000000",
    31176 => x"00000000", 31177 => x"00000000", 31178 => x"00000000",
    31179 => x"00000000", 31180 => x"00000000", 31181 => x"00000000",
    31182 => x"00000000", 31183 => x"00000000", 31184 => x"00000000",
    31185 => x"00000000", 31186 => x"00000000", 31187 => x"00000000",
    31188 => x"00000000", 31189 => x"00000000", 31190 => x"00000000",
    31191 => x"00000000", 31192 => x"00000000", 31193 => x"00000000",
    31194 => x"00000000", 31195 => x"00000000", 31196 => x"00000000",
    31197 => x"00000000", 31198 => x"00000000", 31199 => x"00000000",
    31200 => x"00000000", 31201 => x"00000000", 31202 => x"00000000",
    31203 => x"00000000", 31204 => x"00000000", 31205 => x"00000000",
    31206 => x"00000000", 31207 => x"00000000", 31208 => x"00000000",
    31209 => x"00000000", 31210 => x"00000000", 31211 => x"00000000",
    31212 => x"00000000", 31213 => x"00000000", 31214 => x"00000000",
    31215 => x"00000000", 31216 => x"00000000", 31217 => x"00000000",
    31218 => x"00000000", 31219 => x"00000000", 31220 => x"00000000",
    31221 => x"00000000", 31222 => x"00000000", 31223 => x"00000000",
    31224 => x"00000000", 31225 => x"00000000", 31226 => x"00000000",
    31227 => x"00000000", 31228 => x"00000000", 31229 => x"00000000",
    31230 => x"00000000", 31231 => x"00000000", 31232 => x"00000000",
    31233 => x"00000000", 31234 => x"00000000", 31235 => x"00000000",
    31236 => x"00000000", 31237 => x"00000000", 31238 => x"00000000",
    31239 => x"00000000", 31240 => x"00000000", 31241 => x"00000000",
    31242 => x"00000000", 31243 => x"00000000", 31244 => x"00000000",
    31245 => x"00000000", 31246 => x"00000000", 31247 => x"00000000",
    31248 => x"00000000", 31249 => x"00000000", 31250 => x"00000000",
    31251 => x"00000000", 31252 => x"00000000", 31253 => x"00000000",
    31254 => x"00000000", 31255 => x"00000000", 31256 => x"00000000",
    31257 => x"00000000", 31258 => x"00000000", 31259 => x"00000000",
    31260 => x"00000000", 31261 => x"00000000", 31262 => x"00000000",
    31263 => x"00000000", 31264 => x"00000000", 31265 => x"00000000",
    31266 => x"00000000", 31267 => x"00000000", 31268 => x"00000000",
    31269 => x"00000000", 31270 => x"00000000", 31271 => x"00000000",
    31272 => x"00000000", 31273 => x"00000000", 31274 => x"00000000",
    31275 => x"00000000", 31276 => x"00000000", 31277 => x"00000000",
    31278 => x"00000000", 31279 => x"00000000", 31280 => x"00000000",
    31281 => x"00000000", 31282 => x"00000000", 31283 => x"00000000",
    31284 => x"00000000", 31285 => x"00000000", 31286 => x"00000000",
    31287 => x"00000000", 31288 => x"00000000", 31289 => x"00000000",
    31290 => x"00000000", 31291 => x"00000000", 31292 => x"00000000",
    31293 => x"00000000", 31294 => x"00000000", 31295 => x"00000000",
    31296 => x"00000000", 31297 => x"00000000", 31298 => x"00000000",
    31299 => x"00000000", 31300 => x"00000000", 31301 => x"00000000",
    31302 => x"00000000", 31303 => x"00000000", 31304 => x"00000000",
    31305 => x"00000000", 31306 => x"00000000", 31307 => x"00000000",
    31308 => x"00000000", 31309 => x"00000000", 31310 => x"00000000",
    31311 => x"00000000", 31312 => x"00000000", 31313 => x"00000000",
    31314 => x"00000000", 31315 => x"00000000", 31316 => x"00000000",
    31317 => x"00000000", 31318 => x"00000000", 31319 => x"00000000",
    31320 => x"00000000", 31321 => x"00000000", 31322 => x"00000000",
    31323 => x"00000000", 31324 => x"00000000", 31325 => x"00000000",
    31326 => x"00000000", 31327 => x"00000000", 31328 => x"00000000",
    31329 => x"00000000", 31330 => x"00000000", 31331 => x"00000000",
    31332 => x"00000000", 31333 => x"00000000", 31334 => x"00000000",
    31335 => x"00000000", 31336 => x"00000000", 31337 => x"00000000",
    31338 => x"00000000", 31339 => x"00000000", 31340 => x"00000000",
    31341 => x"00000000", 31342 => x"00000000", 31343 => x"00000000",
    31344 => x"00000000", 31345 => x"00000000", 31346 => x"00000000",
    31347 => x"00000000", 31348 => x"00000000", 31349 => x"00000000",
    31350 => x"00000000", 31351 => x"00000000", 31352 => x"00000000",
    31353 => x"00000000", 31354 => x"00000000", 31355 => x"00000000",
    31356 => x"00000000", 31357 => x"00000000", 31358 => x"00000000",
    31359 => x"00000000", 31360 => x"00000000", 31361 => x"00000000",
    31362 => x"00000000", 31363 => x"00000000", 31364 => x"00000000",
    31365 => x"00000000", 31366 => x"00000000", 31367 => x"00000000",
    31368 => x"00000000", 31369 => x"00000000", 31370 => x"00000000",
    31371 => x"00000000", 31372 => x"00000000", 31373 => x"00000000",
    31374 => x"00000000", 31375 => x"00000000", 31376 => x"00000000",
    31377 => x"00000000", 31378 => x"00000000", 31379 => x"00000000",
    31380 => x"00000000", 31381 => x"00000000", 31382 => x"00000000",
    31383 => x"00000000", 31384 => x"00000000", 31385 => x"00000000",
    31386 => x"00000000", 31387 => x"00000000", 31388 => x"00000000",
    31389 => x"00000000", 31390 => x"00000000", 31391 => x"00000000",
    31392 => x"00000000", 31393 => x"00000000", 31394 => x"00000000",
    31395 => x"00000000", 31396 => x"00000000", 31397 => x"00000000",
    31398 => x"00000000", 31399 => x"00000000", 31400 => x"00000000",
    31401 => x"00000000", 31402 => x"00000000", 31403 => x"00000000",
    31404 => x"00000000", 31405 => x"00000000", 31406 => x"00000000",
    31407 => x"00000000", 31408 => x"00000000", 31409 => x"00000000",
    31410 => x"00000000", 31411 => x"00000000", 31412 => x"00000000",
    31413 => x"00000000", 31414 => x"00000000", 31415 => x"00000000",
    31416 => x"00000000", 31417 => x"00000000", 31418 => x"00000000",
    31419 => x"00000000", 31420 => x"00000000", 31421 => x"00000000",
    31422 => x"00000000", 31423 => x"00000000", 31424 => x"00000000",
    31425 => x"00000000", 31426 => x"00000000", 31427 => x"00000000",
    31428 => x"00000000", 31429 => x"00000000", 31430 => x"00000000",
    31431 => x"00000000", 31432 => x"00000000", 31433 => x"00000000",
    31434 => x"00000000", 31435 => x"00000000", 31436 => x"00000000",
    31437 => x"00000000", 31438 => x"00000000", 31439 => x"00000000",
    31440 => x"00000000", 31441 => x"00000000", 31442 => x"00000000",
    31443 => x"00000000", 31444 => x"00000000", 31445 => x"00000000",
    31446 => x"00000000", 31447 => x"00000000", 31448 => x"00000000",
    31449 => x"00000000", 31450 => x"00000000", 31451 => x"00000000",
    31452 => x"00000000", 31453 => x"00000000", 31454 => x"00000000",
    31455 => x"00000000", 31456 => x"00000000", 31457 => x"00000000",
    31458 => x"00000000", 31459 => x"00000000", 31460 => x"00000000",
    31461 => x"00000000", 31462 => x"00000000", 31463 => x"00000000",
    31464 => x"00000000", 31465 => x"00000000", 31466 => x"00000000",
    31467 => x"00000000", 31468 => x"00000000", 31469 => x"00000000",
    31470 => x"00000000", 31471 => x"00000000", 31472 => x"00000000",
    31473 => x"00000000", 31474 => x"00000000", 31475 => x"00000000",
    31476 => x"00000000", 31477 => x"00000000", 31478 => x"00000000",
    31479 => x"00000000", 31480 => x"00000000", 31481 => x"00000000",
    31482 => x"00000000", 31483 => x"00000000", 31484 => x"00000000",
    31485 => x"00000000", 31486 => x"00000000", 31487 => x"00000000",
    31488 => x"00000000", 31489 => x"00000000", 31490 => x"00000000",
    31491 => x"00000000", 31492 => x"00000000", 31493 => x"00000000",
    31494 => x"00000000", 31495 => x"00000000", 31496 => x"00000000",
    31497 => x"00000000", 31498 => x"00000000", 31499 => x"00000000",
    31500 => x"00000000", 31501 => x"00000000", 31502 => x"00000000",
    31503 => x"00000000", 31504 => x"00000000", 31505 => x"00000000",
    31506 => x"00000000", 31507 => x"00000000", 31508 => x"00000000",
    31509 => x"00000000", 31510 => x"00000000", 31511 => x"00000000",
    31512 => x"00000000", 31513 => x"00000000", 31514 => x"00000000",
    31515 => x"00000000", 31516 => x"00000000", 31517 => x"00000000",
    31518 => x"00000000", 31519 => x"00000000", 31520 => x"00000000",
    31521 => x"00000000", 31522 => x"00000000", 31523 => x"00000000",
    31524 => x"00000000", 31525 => x"00000000", 31526 => x"00000000",
    31527 => x"00000000", 31528 => x"00000000", 31529 => x"00000000",
    31530 => x"00000000", 31531 => x"00000000", 31532 => x"00000000",
    31533 => x"00000000", 31534 => x"00000000", 31535 => x"00000000",
    31536 => x"00000000", 31537 => x"00000000", 31538 => x"00000000",
    31539 => x"00000000", 31540 => x"00000000", 31541 => x"00000000",
    31542 => x"00000000", 31543 => x"00000000", 31544 => x"00000000",
    31545 => x"00000000", 31546 => x"00000000", 31547 => x"00000000",
    31548 => x"00000000", 31549 => x"00000000", 31550 => x"00000000",
    31551 => x"00000000", 31552 => x"00000000", 31553 => x"00000000",
    31554 => x"00000000", 31555 => x"00000000", 31556 => x"00000000",
    31557 => x"00000000", 31558 => x"00000000", 31559 => x"00000000",
    31560 => x"00000000", 31561 => x"00000000", 31562 => x"00000000",
    31563 => x"00000000", 31564 => x"00000000", 31565 => x"00000000",
    31566 => x"00000000", 31567 => x"00000000", 31568 => x"00000000",
    31569 => x"00000000", 31570 => x"00000000", 31571 => x"00000000",
    31572 => x"00000000", 31573 => x"00000000", 31574 => x"00000000",
    31575 => x"00000000", 31576 => x"00000000", 31577 => x"00000000",
    31578 => x"00000000", 31579 => x"00000000", 31580 => x"00000000",
    31581 => x"00000000", 31582 => x"00000000", 31583 => x"00000000",
    31584 => x"00000000", 31585 => x"00000000", 31586 => x"00000000",
    31587 => x"00000000", 31588 => x"00000000", 31589 => x"00000000",
    31590 => x"00000000", 31591 => x"00000000", 31592 => x"00000000",
    31593 => x"00000000", 31594 => x"00000000", 31595 => x"00000000",
    31596 => x"00000000", 31597 => x"00000000", 31598 => x"00000000",
    31599 => x"00000000", 31600 => x"00000000", 31601 => x"00000000",
    31602 => x"00000000", 31603 => x"00000000", 31604 => x"00000000",
    31605 => x"00000000", 31606 => x"00000000", 31607 => x"00000000",
    31608 => x"00000000", 31609 => x"00000000", 31610 => x"00000000",
    31611 => x"00000000", 31612 => x"00000000", 31613 => x"00000000",
    31614 => x"00000000", 31615 => x"00000000", 31616 => x"00000000",
    31617 => x"00000000", 31618 => x"00000000", 31619 => x"00000000",
    31620 => x"00000000", 31621 => x"00000000", 31622 => x"00000000",
    31623 => x"00000000", 31624 => x"00000000", 31625 => x"00000000",
    31626 => x"00000000", 31627 => x"00000000", 31628 => x"00000000",
    31629 => x"00000000", 31630 => x"00000000", 31631 => x"00000000",
    31632 => x"00000000", 31633 => x"00000000", 31634 => x"00000000",
    31635 => x"00000000", 31636 => x"00000000", 31637 => x"00000000",
    31638 => x"00000000", 31639 => x"00000000", 31640 => x"00000000",
    31641 => x"00000000", 31642 => x"00000000", 31643 => x"00000000",
    31644 => x"00000000", 31645 => x"00000000", 31646 => x"00000000",
    31647 => x"00000000", 31648 => x"00000000", 31649 => x"00000000",
    31650 => x"00000000", 31651 => x"00000000", 31652 => x"00000000",
    31653 => x"00000000", 31654 => x"00000000", 31655 => x"00000000",
    31656 => x"00000000", 31657 => x"00000000", 31658 => x"00000000",
    31659 => x"00000000", 31660 => x"00000000", 31661 => x"00000000",
    31662 => x"00000000", 31663 => x"00000000", 31664 => x"00000000",
    31665 => x"00000000", 31666 => x"00000000", 31667 => x"00000000",
    31668 => x"00000000", 31669 => x"00000000", 31670 => x"00000000",
    31671 => x"00000000", 31672 => x"00000000", 31673 => x"00000000",
    31674 => x"00000000", 31675 => x"00000000", 31676 => x"00000000",
    31677 => x"00000000", 31678 => x"00000000", 31679 => x"00000000",
    31680 => x"00000000", 31681 => x"00000000", 31682 => x"00000000",
    31683 => x"00000000", 31684 => x"00000000", 31685 => x"00000000",
    31686 => x"00000000", 31687 => x"00000000", 31688 => x"00000000",
    31689 => x"00000000", 31690 => x"00000000", 31691 => x"00000000",
    31692 => x"00000000", 31693 => x"00000000", 31694 => x"00000000",
    31695 => x"00000000", 31696 => x"00000000", 31697 => x"00000000",
    31698 => x"00000000", 31699 => x"00000000", 31700 => x"00000000",
    31701 => x"00000000", 31702 => x"00000000", 31703 => x"00000000",
    31704 => x"00000000", 31705 => x"00000000", 31706 => x"00000000",
    31707 => x"00000000", 31708 => x"00000000", 31709 => x"00000000",
    31710 => x"00000000", 31711 => x"00000000", 31712 => x"00000000",
    31713 => x"00000000", 31714 => x"00000000", 31715 => x"00000000",
    31716 => x"00000000", 31717 => x"00000000", 31718 => x"00000000",
    31719 => x"00000000", 31720 => x"00000000", 31721 => x"00000000",
    31722 => x"00000000", 31723 => x"00000000", 31724 => x"00000000",
    31725 => x"00000000", 31726 => x"00000000", 31727 => x"00000000",
    31728 => x"00000000", 31729 => x"00000000", 31730 => x"00000000",
    31731 => x"00000000", 31732 => x"00000000", 31733 => x"00000000",
    31734 => x"00000000", 31735 => x"00000000", 31736 => x"00000000",
    31737 => x"00000000", 31738 => x"00000000", 31739 => x"00000000",
    31740 => x"00000000", 31741 => x"00000000", 31742 => x"00000000",
    31743 => x"00000000", 31744 => x"00000000", 31745 => x"00000000",
    31746 => x"00000000", 31747 => x"00000000", 31748 => x"00000000",
    31749 => x"00000000", 31750 => x"00000000", 31751 => x"00000000",
    31752 => x"00000000", 31753 => x"00000000", 31754 => x"00000000",
    31755 => x"00000000", 31756 => x"00000000", 31757 => x"00000000",
    31758 => x"00000000", 31759 => x"00000000", 31760 => x"00000000",
    31761 => x"00000000", 31762 => x"00000000", 31763 => x"00000000",
    31764 => x"00000000", 31765 => x"00000000", 31766 => x"00000000",
    31767 => x"00000000", 31768 => x"00000000", 31769 => x"00000000",
    31770 => x"00000000", 31771 => x"00000000", 31772 => x"00000000",
    31773 => x"00000000", 31774 => x"00000000", 31775 => x"00000000",
    31776 => x"00000000", 31777 => x"00000000", 31778 => x"00000000",
    31779 => x"00000000", 31780 => x"00000000", 31781 => x"00000000",
    31782 => x"00000000", 31783 => x"00000000", 31784 => x"00000000",
    31785 => x"00000000", 31786 => x"00000000", 31787 => x"00000000",
    31788 => x"00000000", 31789 => x"00000000", 31790 => x"00000000",
    31791 => x"00000000", 31792 => x"00000000", 31793 => x"00000000",
    31794 => x"00000000", 31795 => x"00000000", 31796 => x"00000000",
    31797 => x"00000000", 31798 => x"00000000", 31799 => x"00000000",
    31800 => x"00000000", 31801 => x"00000000", 31802 => x"00000000",
    31803 => x"00000000", 31804 => x"00000000", 31805 => x"00000000",
    31806 => x"00000000", 31807 => x"00000000", 31808 => x"00000000",
    31809 => x"00000000", 31810 => x"00000000", 31811 => x"00000000",
    31812 => x"00000000", 31813 => x"00000000", 31814 => x"00000000",
    31815 => x"00000000", 31816 => x"00000000", 31817 => x"00000000",
    31818 => x"00000000", 31819 => x"00000000", 31820 => x"00000000",
    31821 => x"00000000", 31822 => x"00000000", 31823 => x"00000000",
    31824 => x"00000000", 31825 => x"00000000", 31826 => x"00000000",
    31827 => x"00000000", 31828 => x"00000000", 31829 => x"00000000",
    31830 => x"00000000", 31831 => x"00000000", 31832 => x"00000000",
    31833 => x"00000000", 31834 => x"00000000", 31835 => x"00000000",
    31836 => x"00000000", 31837 => x"00000000", 31838 => x"00000000",
    31839 => x"00000000", 31840 => x"00000000", 31841 => x"00000000",
    31842 => x"00000000", 31843 => x"00000000", 31844 => x"00000000",
    31845 => x"00000000", 31846 => x"00000000", 31847 => x"00000000",
    31848 => x"00000000", 31849 => x"00000000", 31850 => x"00000000",
    31851 => x"00000000", 31852 => x"00000000", 31853 => x"00000000",
    31854 => x"00000000", 31855 => x"00000000", 31856 => x"00000000",
    31857 => x"00000000", 31858 => x"00000000", 31859 => x"00000000",
    31860 => x"00000000", 31861 => x"00000000", 31862 => x"00000000",
    31863 => x"00000000", 31864 => x"00000000", 31865 => x"00000000",
    31866 => x"00000000", 31867 => x"00000000", 31868 => x"00000000",
    31869 => x"00000000", 31870 => x"00000000", 31871 => x"00000000",
    31872 => x"00000000", 31873 => x"00000000", 31874 => x"00000000",
    31875 => x"00000000", 31876 => x"00000000", 31877 => x"00000000",
    31878 => x"00000000", 31879 => x"00000000", 31880 => x"00000000",
    31881 => x"00000000", 31882 => x"00000000", 31883 => x"00000000",
    31884 => x"00000000", 31885 => x"00000000", 31886 => x"00000000",
    31887 => x"00000000", 31888 => x"00000000", 31889 => x"00000000",
    31890 => x"00000000", 31891 => x"00000000", 31892 => x"00000000",
    31893 => x"00000000", 31894 => x"00000000", 31895 => x"00000000",
    31896 => x"00000000", 31897 => x"00000000", 31898 => x"00000000",
    31899 => x"00000000", 31900 => x"00000000", 31901 => x"00000000",
    31902 => x"00000000", 31903 => x"00000000", 31904 => x"00000000",
    31905 => x"00000000", 31906 => x"00000000", 31907 => x"00000000",
    31908 => x"00000000", 31909 => x"00000000", 31910 => x"00000000",
    31911 => x"00000000", 31912 => x"00000000", 31913 => x"00000000",
    31914 => x"00000000", 31915 => x"00000000", 31916 => x"00000000",
    31917 => x"00000000", 31918 => x"00000000", 31919 => x"00000000",
    31920 => x"00000000", 31921 => x"00000000", 31922 => x"00000000",
    31923 => x"00000000", 31924 => x"00000000", 31925 => x"00000000",
    31926 => x"00000000", 31927 => x"00000000", 31928 => x"00000000",
    31929 => x"00000000", 31930 => x"00000000", 31931 => x"00000000",
    31932 => x"00000000", 31933 => x"00000000", 31934 => x"00000000",
    31935 => x"00000000", 31936 => x"00000000", 31937 => x"00000000",
    31938 => x"00000000", 31939 => x"00000000", 31940 => x"00000000",
    31941 => x"00000000", 31942 => x"00000000", 31943 => x"00000000",
    31944 => x"00000000", 31945 => x"00000000", 31946 => x"00000000",
    31947 => x"00000000", 31948 => x"00000000", 31949 => x"00000000",
    31950 => x"00000000", 31951 => x"00000000", 31952 => x"00000000",
    31953 => x"00000000", 31954 => x"00000000", 31955 => x"00000000",
    31956 => x"00000000", 31957 => x"00000000", 31958 => x"00000000",
    31959 => x"00000000", 31960 => x"00000000", 31961 => x"00000000",
    31962 => x"00000000", 31963 => x"00000000", 31964 => x"00000000",
    31965 => x"00000000", 31966 => x"00000000", 31967 => x"00000000",
    31968 => x"00000000", 31969 => x"00000000", 31970 => x"00000000",
    31971 => x"00000000", 31972 => x"00000000", 31973 => x"00000000",
    31974 => x"00000000", 31975 => x"00000000", 31976 => x"00000000",
    31977 => x"00000000", 31978 => x"00000000", 31979 => x"00000000",
    31980 => x"00000000", 31981 => x"00000000", 31982 => x"00000000",
    31983 => x"00000000", 31984 => x"00000000", 31985 => x"00000000",
    31986 => x"00000000", 31987 => x"00000000", 31988 => x"00000000",
    31989 => x"00000000", 31990 => x"00000000", 31991 => x"00000000",
    31992 => x"00000000", 31993 => x"00000000", 31994 => x"00000000",
    31995 => x"00000000", 31996 => x"00000000", 31997 => x"00000000",
    31998 => x"00000000", 31999 => x"00000000", 32000 => x"00000000",
    32001 => x"00000000", 32002 => x"00000000", 32003 => x"00000000",
    32004 => x"00000000", 32005 => x"00000000", 32006 => x"00000000",
    32007 => x"00000000", 32008 => x"00000000", 32009 => x"00000000",
    32010 => x"00000000", 32011 => x"00000000", 32012 => x"00000000",
    32013 => x"00000000", 32014 => x"00000000", 32015 => x"00000000",
    32016 => x"00000000", 32017 => x"00000000", 32018 => x"00000000",
    32019 => x"00000000", 32020 => x"00000000", 32021 => x"00000000",
    32022 => x"00000000", 32023 => x"00000000", 32024 => x"00000000",
    32025 => x"00000000", 32026 => x"00000000", 32027 => x"00000000",
    32028 => x"00000000", 32029 => x"00000000", 32030 => x"00000000",
    32031 => x"00000000", 32032 => x"00000000", 32033 => x"00000000",
    32034 => x"00000000", 32035 => x"00000000", 32036 => x"00000000",
    32037 => x"00000000", 32038 => x"00000000", 32039 => x"00000000",
    32040 => x"00000000", 32041 => x"00000000", 32042 => x"00000000",
    32043 => x"00000000", 32044 => x"00000000", 32045 => x"00000000",
    32046 => x"00000000", 32047 => x"00000000", 32048 => x"00000000",
    32049 => x"00000000", 32050 => x"00000000", 32051 => x"00000000",
    32052 => x"00000000", 32053 => x"00000000", 32054 => x"00000000",
    32055 => x"00000000", 32056 => x"00000000", 32057 => x"00000000",
    32058 => x"00000000", 32059 => x"00000000", 32060 => x"00000000",
    32061 => x"00000000", 32062 => x"00000000", 32063 => x"00000000",
    32064 => x"00000000", 32065 => x"00000000", 32066 => x"00000000",
    32067 => x"00000000", 32068 => x"00000000", 32069 => x"00000000",
    32070 => x"00000000", 32071 => x"00000000", 32072 => x"00000000",
    32073 => x"00000000", 32074 => x"00000000", 32075 => x"00000000",
    32076 => x"00000000", 32077 => x"00000000", 32078 => x"00000000",
    32079 => x"00000000", 32080 => x"00000000", 32081 => x"00000000",
    32082 => x"00000000", 32083 => x"00000000", 32084 => x"00000000",
    32085 => x"00000000", 32086 => x"00000000", 32087 => x"00000000",
    32088 => x"00000000", 32089 => x"00000000", 32090 => x"00000000",
    32091 => x"00000000", 32092 => x"00000000", 32093 => x"00000000",
    32094 => x"00000000", 32095 => x"00000000", 32096 => x"00000000",
    32097 => x"00000000", 32098 => x"00000000", 32099 => x"00000000",
    32100 => x"00000000", 32101 => x"00000000", 32102 => x"00000000",
    32103 => x"00000000", 32104 => x"00000000", 32105 => x"00000000",
    32106 => x"00000000", 32107 => x"00000000", 32108 => x"00000000",
    32109 => x"00000000", 32110 => x"00000000", 32111 => x"00000000",
    32112 => x"00000000", 32113 => x"00000000", 32114 => x"00000000",
    32115 => x"00000000", 32116 => x"00000000", 32117 => x"00000000",
    32118 => x"00000000", 32119 => x"00000000", 32120 => x"00000000",
    32121 => x"00000000", 32122 => x"00000000", 32123 => x"00000000",
    32124 => x"00000000", 32125 => x"00000000", 32126 => x"00000000",
    32127 => x"00000000", 32128 => x"00000000", 32129 => x"00000000",
    32130 => x"00000000", 32131 => x"00000000", 32132 => x"00000000",
    32133 => x"00000000", 32134 => x"00000000", 32135 => x"00000000",
    32136 => x"00000000", 32137 => x"00000000", 32138 => x"00000000",
    32139 => x"00000000", 32140 => x"00000000", 32141 => x"00000000",
    32142 => x"00000000", 32143 => x"00000000", 32144 => x"00000000",
    32145 => x"00000000", 32146 => x"00000000", 32147 => x"00000000",
    32148 => x"00000000", 32149 => x"00000000", 32150 => x"00000000",
    32151 => x"00000000", 32152 => x"00000000", 32153 => x"00000000",
    32154 => x"00000000", 32155 => x"00000000", 32156 => x"00000000",
    32157 => x"00000000", 32158 => x"00000000", 32159 => x"00000000",
    32160 => x"00000000", 32161 => x"00000000", 32162 => x"00000000",
    32163 => x"00000000", 32164 => x"00000000", 32165 => x"00000000",
    32166 => x"00000000", 32167 => x"00000000", 32168 => x"00000000",
    32169 => x"00000000", 32170 => x"00000000", 32171 => x"00000000",
    32172 => x"00000000", 32173 => x"00000000", 32174 => x"00000000",
    32175 => x"00000000", 32176 => x"00000000", 32177 => x"00000000",
    32178 => x"00000000", 32179 => x"00000000", 32180 => x"00000000",
    32181 => x"00000000", 32182 => x"00000000", 32183 => x"00000000",
    32184 => x"00000000", 32185 => x"00000000", 32186 => x"00000000",
    32187 => x"00000000", 32188 => x"00000000", 32189 => x"00000000",
    32190 => x"00000000", 32191 => x"00000000", 32192 => x"00000000",
    32193 => x"00000000", 32194 => x"00000000", 32195 => x"00000000",
    32196 => x"00000000", 32197 => x"00000000", 32198 => x"00000000",
    32199 => x"00000000", 32200 => x"00000000", 32201 => x"00000000",
    32202 => x"00000000", 32203 => x"00000000", 32204 => x"00000000",
    32205 => x"00000000", 32206 => x"00000000", 32207 => x"00000000",
    32208 => x"00000000", 32209 => x"00000000", 32210 => x"00000000",
    32211 => x"00000000", 32212 => x"00000000", 32213 => x"00000000",
    32214 => x"00000000", 32215 => x"00000000", 32216 => x"00000000",
    32217 => x"00000000", 32218 => x"00000000", 32219 => x"00000000",
    32220 => x"00000000", 32221 => x"00000000", 32222 => x"00000000",
    32223 => x"00000000", 32224 => x"00000000", 32225 => x"00000000",
    32226 => x"00000000", 32227 => x"00000000", 32228 => x"00000000",
    32229 => x"00000000", 32230 => x"00000000", 32231 => x"00000000",
    32232 => x"00000000", 32233 => x"00000000", 32234 => x"00000000",
    32235 => x"00000000", 32236 => x"00000000", 32237 => x"00000000",
    32238 => x"00000000", 32239 => x"00000000", 32240 => x"00000000",
    32241 => x"00000000", 32242 => x"00000000", 32243 => x"00000000",
    32244 => x"00000000", 32245 => x"00000000", 32246 => x"00000000",
    32247 => x"00000000", 32248 => x"00000000", 32249 => x"00000000",
    32250 => x"00000000", 32251 => x"00000000", 32252 => x"00000000",
    32253 => x"00000000", 32254 => x"00000000", 32255 => x"00000000",
    32256 => x"00000000", 32257 => x"00000000", 32258 => x"00000000",
    32259 => x"00000000", 32260 => x"00000000", 32261 => x"00000000",
    32262 => x"00000000", 32263 => x"00000000", 32264 => x"00000000",
    32265 => x"00000000", 32266 => x"00000000", 32267 => x"00000000",
    32268 => x"00000000", 32269 => x"00000000", 32270 => x"00000000",
    32271 => x"00000000", 32272 => x"00000000", 32273 => x"00000000",
    32274 => x"00000000", 32275 => x"00000000", 32276 => x"00000000",
    32277 => x"00000000", 32278 => x"00000000", 32279 => x"00000000",
    32280 => x"00000000", 32281 => x"00000000", 32282 => x"00000000",
    32283 => x"00000000", 32284 => x"00000000", 32285 => x"00000000",
    32286 => x"00000000", 32287 => x"00000000", 32288 => x"00000000",
    32289 => x"00000000", 32290 => x"00000000", 32291 => x"00000000",
    32292 => x"00000000", 32293 => x"00000000", 32294 => x"00000000",
    32295 => x"00000000", 32296 => x"00000000", 32297 => x"00000000",
    32298 => x"00000000", 32299 => x"00000000", 32300 => x"00000000",
    32301 => x"00000000", 32302 => x"00000000", 32303 => x"00000000",
    32304 => x"00000000", 32305 => x"00000000", 32306 => x"00000000",
    32307 => x"00000000", 32308 => x"00000000", 32309 => x"00000000",
    32310 => x"00000000", 32311 => x"00000000", 32312 => x"00000000",
    32313 => x"00000000", 32314 => x"00000000", 32315 => x"00000000",
    32316 => x"00000000", 32317 => x"00000000", 32318 => x"00000000",
    32319 => x"00000000", 32320 => x"00000000", 32321 => x"00000000",
    32322 => x"00000000", 32323 => x"00000000", 32324 => x"00000000",
    32325 => x"00000000", 32326 => x"00000000", 32327 => x"00000000",
    32328 => x"00000000", 32329 => x"00000000", 32330 => x"00000000",
    32331 => x"00000000", 32332 => x"00000000", 32333 => x"00000000",
    32334 => x"00000000", 32335 => x"00000000", 32336 => x"00000000",
    32337 => x"00000000", 32338 => x"00000000", 32339 => x"00000000",
    32340 => x"00000000", 32341 => x"00000000", 32342 => x"00000000",
    32343 => x"00000000", 32344 => x"00000000", 32345 => x"00000000",
    32346 => x"00000000", 32347 => x"00000000", 32348 => x"00000000",
    32349 => x"00000000", 32350 => x"00000000", 32351 => x"00000000",
    32352 => x"00000000", 32353 => x"00000000", 32354 => x"00000000",
    32355 => x"00000000", 32356 => x"00000000", 32357 => x"00000000",
    32358 => x"00000000", 32359 => x"00000000", 32360 => x"00000000",
    32361 => x"00000000", 32362 => x"00000000", 32363 => x"00000000",
    32364 => x"00000000", 32365 => x"00000000", 32366 => x"00000000",
    32367 => x"00000000", 32368 => x"00000000", 32369 => x"00000000",
    32370 => x"00000000", 32371 => x"00000000", 32372 => x"00000000",
    32373 => x"00000000", 32374 => x"00000000", 32375 => x"00000000",
    32376 => x"00000000", 32377 => x"00000000", 32378 => x"00000000",
    32379 => x"00000000", 32380 => x"00000000", 32381 => x"00000000",
    32382 => x"00000000", 32383 => x"00000000", 32384 => x"00000000",
    32385 => x"00000000", 32386 => x"00000000", 32387 => x"00000000",
    32388 => x"00000000", 32389 => x"00000000", 32390 => x"00000000",
    32391 => x"00000000", 32392 => x"00000000", 32393 => x"00000000",
    32394 => x"00000000", 32395 => x"00000000", 32396 => x"00000000",
    32397 => x"00000000", 32398 => x"00000000", 32399 => x"00000000",
    32400 => x"00000000", 32401 => x"00000000", 32402 => x"00000000",
    32403 => x"00000000", 32404 => x"00000000", 32405 => x"00000000",
    32406 => x"00000000", 32407 => x"00000000", 32408 => x"00000000",
    32409 => x"00000000", 32410 => x"00000000", 32411 => x"00000000",
    32412 => x"00000000", 32413 => x"00000000", 32414 => x"00000000",
    32415 => x"00000000", 32416 => x"00000000", 32417 => x"00000000",
    32418 => x"00000000", 32419 => x"00000000", 32420 => x"00000000",
    32421 => x"00000000", 32422 => x"00000000", 32423 => x"00000000",
    32424 => x"00000000", 32425 => x"00000000", 32426 => x"00000000",
    32427 => x"00000000", 32428 => x"00000000", 32429 => x"00000000",
    32430 => x"00000000", 32431 => x"00000000", 32432 => x"00000000",
    32433 => x"00000000", 32434 => x"00000000", 32435 => x"00000000",
    32436 => x"00000000", 32437 => x"00000000", 32438 => x"00000000",
    32439 => x"00000000", 32440 => x"00000000", 32441 => x"00000000",
    32442 => x"00000000", 32443 => x"00000000", 32444 => x"00000000",
    32445 => x"00000000", 32446 => x"00000000", 32447 => x"00000000",
    32448 => x"00000000", 32449 => x"00000000", 32450 => x"00000000",
    32451 => x"00000000", 32452 => x"00000000", 32453 => x"00000000",
    32454 => x"00000000", 32455 => x"00000000", 32456 => x"00000000",
    32457 => x"00000000", 32458 => x"00000000", 32459 => x"00000000",
    32460 => x"00000000", 32461 => x"00000000", 32462 => x"00000000",
    32463 => x"00000000", 32464 => x"00000000", 32465 => x"00000000",
    32466 => x"00000000", 32467 => x"00000000", 32468 => x"00000000",
    32469 => x"00000000", 32470 => x"00000000", 32471 => x"00000000",
    32472 => x"00000000", 32473 => x"00000000", 32474 => x"00000000",
    32475 => x"00000000", 32476 => x"00000000", 32477 => x"00000000",
    32478 => x"00000000", 32479 => x"00000000", 32480 => x"00000000",
    32481 => x"00000000", 32482 => x"00000000", 32483 => x"00000000",
    32484 => x"00000000", 32485 => x"00000000", 32486 => x"00000000",
    32487 => x"00000000", 32488 => x"00000000", 32489 => x"00000000",
    32490 => x"00000000", 32491 => x"00000000", 32492 => x"00000000",
    32493 => x"00000000", 32494 => x"00000000", 32495 => x"00000000",
    32496 => x"00000000", 32497 => x"00000000", 32498 => x"00000000",
    32499 => x"00000000", 32500 => x"00000000", 32501 => x"00000000",
    32502 => x"00000000", 32503 => x"00000000", 32504 => x"00000000",
    32505 => x"00000000", 32506 => x"00000000", 32507 => x"00000000",
    32508 => x"00000000", 32509 => x"00000000", 32510 => x"00000000",
    32511 => x"00000000", 32512 => x"00000000", 32513 => x"00000000",
    32514 => x"00000000", 32515 => x"00000000", 32516 => x"00000000",
    32517 => x"00000000", 32518 => x"00000000", 32519 => x"00000000",
    32520 => x"00000000", 32521 => x"00000000", 32522 => x"00000000",
    32523 => x"00000000", 32524 => x"00000000", 32525 => x"00000000",
    32526 => x"00000000", 32527 => x"00000000", 32528 => x"00000000",
    32529 => x"00000000", 32530 => x"00000000", 32531 => x"00000000",
    32532 => x"00000000", 32533 => x"00000000", 32534 => x"00000000",
    32535 => x"00000000", 32536 => x"00000000", 32537 => x"00000000",
    32538 => x"00000000", 32539 => x"00000000", 32540 => x"00000000",
    32541 => x"00000000", 32542 => x"00000000", 32543 => x"00000000",
    32544 => x"00000000", 32545 => x"00000000", 32546 => x"00000000",
    32547 => x"00000000", 32548 => x"00000000", 32549 => x"00000000",
    32550 => x"00000000", 32551 => x"00000000", 32552 => x"00000000",
    32553 => x"00000000", 32554 => x"00000000", 32555 => x"00000000",
    32556 => x"00000000", 32557 => x"00000000", 32558 => x"00000000",
    32559 => x"00000000", 32560 => x"00000000", 32561 => x"00000000",
    32562 => x"00000000", 32563 => x"00000000", 32564 => x"00000000",
    32565 => x"00000000", 32566 => x"00000000", 32567 => x"00000000",
    32568 => x"00000000", 32569 => x"00000000", 32570 => x"00000000",
    32571 => x"00000000", 32572 => x"00000000", 32573 => x"00000000",
    32574 => x"00000000", 32575 => x"00000000", 32576 => x"00000000",
    32577 => x"00000000", 32578 => x"00000000", 32579 => x"00000000",
    32580 => x"00000000", 32581 => x"00000000", 32582 => x"00000000",
    32583 => x"00000000", 32584 => x"00000000", 32585 => x"00000000",
    32586 => x"00000000", 32587 => x"00000000", 32588 => x"00000000",
    32589 => x"00000000", 32590 => x"00000000", 32591 => x"00000000",
    32592 => x"00000000", 32593 => x"00000000", 32594 => x"00000000",
    32595 => x"00000000", 32596 => x"00000000", 32597 => x"00000000",
    32598 => x"00000000", 32599 => x"00000000", 32600 => x"00000000",
    32601 => x"00000000", 32602 => x"00000000", 32603 => x"00000000",
    32604 => x"00000000", 32605 => x"00000000", 32606 => x"00000000",
    32607 => x"00000000", 32608 => x"00000000", 32609 => x"00000000",
    32610 => x"00000000", 32611 => x"00000000", 32612 => x"00000000",
    32613 => x"00000000", 32614 => x"00000000", 32615 => x"00000000",
    32616 => x"00000000", 32617 => x"00000000", 32618 => x"00000000",
    32619 => x"00000000", 32620 => x"00000000", 32621 => x"00000000",
    32622 => x"00000000", 32623 => x"00000000", 32624 => x"00000000",
    32625 => x"00000000", 32626 => x"00000000", 32627 => x"00000000",
    32628 => x"00000000", 32629 => x"00000000", 32630 => x"00000000",
    32631 => x"00000000", 32632 => x"00000000", 32633 => x"00000000",
    32634 => x"00000000", 32635 => x"00000000", 32636 => x"00000000",
    32637 => x"00000000", 32638 => x"00000000", 32639 => x"00000000",
    32640 => x"00000000", 32641 => x"00000000", 32642 => x"00000000",
    32643 => x"00000000", 32644 => x"00000000", 32645 => x"00000000",
    32646 => x"00000000", 32647 => x"00000000", 32648 => x"00000000",
    32649 => x"00000000", 32650 => x"00000000", 32651 => x"00000000",
    32652 => x"00000000", 32653 => x"00000000", 32654 => x"00000000",
    32655 => x"00000000", 32656 => x"00000000", 32657 => x"00000000",
    32658 => x"00000000", 32659 => x"00000000", 32660 => x"00000000",
    32661 => x"00000000", 32662 => x"00000000", 32663 => x"00000000",
    32664 => x"00000000", 32665 => x"00000000", 32666 => x"00000000",
    32667 => x"00000000", 32668 => x"00000000", 32669 => x"00000000",
    32670 => x"00000000", 32671 => x"00000000", 32672 => x"00000000",
    32673 => x"00000000", 32674 => x"00000000", 32675 => x"00000000",
    32676 => x"00000000", 32677 => x"00000000", 32678 => x"00000000",
    32679 => x"00000000", 32680 => x"00000000", 32681 => x"00000000",
    32682 => x"00000000", 32683 => x"00000000", 32684 => x"00000000",
    32685 => x"00000000", 32686 => x"00000000", 32687 => x"00000000",
    32688 => x"00000000", 32689 => x"00000000", 32690 => x"00000000",
    32691 => x"00000000", 32692 => x"00000000", 32693 => x"00000000",
    32694 => x"00000000", 32695 => x"00000000", 32696 => x"00000000",
    32697 => x"00000000", 32698 => x"00000000", 32699 => x"00000000",
    32700 => x"00000000", 32701 => x"00000000", 32702 => x"00000000",
    32703 => x"00000000", 32704 => x"00000000", 32705 => x"00000000",
    32706 => x"00000000", 32707 => x"00000000", 32708 => x"00000000",
    32709 => x"00000000", 32710 => x"00000000", 32711 => x"00000000",
    32712 => x"00000000", 32713 => x"00000000", 32714 => x"00000000",
    32715 => x"00000000", 32716 => x"00000000", 32717 => x"00000000",
    32718 => x"00000000", 32719 => x"00000000", 32720 => x"00000000",
    32721 => x"00000000", 32722 => x"00000000", 32723 => x"00000000",
    32724 => x"00000000", 32725 => x"00000000", 32726 => x"00000000",
    32727 => x"00000000", 32728 => x"00000000", 32729 => x"00000000",
    32730 => x"00000000", 32731 => x"00000000", 32732 => x"00000000",
    32733 => x"00000000", 32734 => x"00000000", 32735 => x"00000000",
    32736 => x"00000000", 32737 => x"00000000", 32738 => x"00000000",
    32739 => x"00000000", 32740 => x"00000000", 32741 => x"00000000",
    32742 => x"00000000", 32743 => x"00000000", 32744 => x"00000000",
    32745 => x"00000000", 32746 => x"00000000", 32747 => x"00000000",
    32748 => x"00000000", 32749 => x"00000000", 32750 => x"00000000",
    32751 => x"00000000", 32752 => x"00000000", 32753 => x"00000000",
    32754 => x"00000000", 32755 => x"00000000", 32756 => x"00000000",
    32757 => x"00000000", 32758 => x"00000000", 32759 => x"00000000",
    32760 => x"00000000", 32761 => x"00000000", 32762 => x"00000000",
    32763 => x"00000000", 32764 => x"00000000", 32765 => x"00000000",
    32766 => x"00000000", 32767 => x"00000000");
end wrc_bin_pkg;

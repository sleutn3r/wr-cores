-- WRPC LM32 RAM initialization: --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.memory_loader_pkg.all;
use work.genram_pkg.all;

package wrc_bin_pkg is
  constant c_wrc_bin_init : t_ram_fast_load ( 0 to 32767 ) := (
        0 => x"98000000",     1 => x"d0000000",     2 => x"d0200000",
        3 => x"78010000",     4 => x"38210000",     5 => x"d0e10000",
        6 => x"f800003a",     7 => x"34000000",     8 => x"00000000",
        9 => x"00000000",    10 => x"00000000",    11 => x"00000000",
       12 => x"00000000",    13 => x"00000000",    14 => x"00000000",
       15 => x"00000000",    16 => x"00000000",    17 => x"00000000",
       18 => x"00000000",    19 => x"00000000",    20 => x"00000000",
       21 => x"00000000",    22 => x"00000000",    23 => x"00000000",
       24 => x"00000000",    25 => x"00000000",    26 => x"00000000",
       27 => x"00000000",    28 => x"00000000",    29 => x"00000000",
       30 => x"00000000",    31 => x"00000000",    32 => x"57525043",
       33 => x"2d2d2d2d",    34 => x"01234567",    35 => x"89abcdef",
       36 => x"00018c3c",    37 => x"00000000",    38 => x"00015e98",
       39 => x"00000000",    40 => x"00000000",    41 => x"00000000",
       42 => x"00000000",    43 => x"00000000",    44 => x"00000000",
       45 => x"00000000",    46 => x"00000000",    47 => x"00000000",
       48 => x"5b9d0000",    49 => x"f800001e",    50 => x"34010002",
       51 => x"f800459a",    52 => x"e000002e",    53 => x"34000000",
       54 => x"34000000",    55 => x"34000000",    56 => x"00000000",
       57 => x"00000000",    58 => x"00000000",    59 => x"00000000",
       60 => x"00000000",    61 => x"00000000",    62 => x"00000000",
       63 => x"00000000",    64 => x"98000000",    65 => x"781c0001",
       66 => x"3b9cfffc",    67 => x"78010001",    68 => x"38217268",
       69 => x"34020000",    70 => x"78030001",    71 => x"38638fb0",
       72 => x"c8611800",    73 => x"f8004b67",    74 => x"34010000",
       75 => x"34020000",    76 => x"34030000",    77 => x"f800010e",
       78 => x"e0000000",    79 => x"379cffc4",    80 => x"5b810004",
       81 => x"5b820008",    82 => x"5b83000c",    83 => x"5b840010",
       84 => x"5b850014",    85 => x"5b860018",    86 => x"5b87001c",
       87 => x"5b880020",    88 => x"5b890024",    89 => x"5b8a0028",
       90 => x"5b9e0034",    91 => x"5b9f0038",    92 => x"2b81003c",
       93 => x"5b810030",    94 => x"bb800800",    95 => x"3421003c",
       96 => x"5b81002c",    97 => x"c3a00000",    98 => x"2b810004",
       99 => x"2b820008",   100 => x"2b83000c",   101 => x"2b840010",
      102 => x"2b850014",   103 => x"2b860018",   104 => x"2b87001c",
      105 => x"2b880020",   106 => x"2b890024",   107 => x"2b8a0028",
      108 => x"2b9d0030",   109 => x"2b9e0034",   110 => x"2b9f0038",
      111 => x"2b9c002c",   112 => x"34000000",   113 => x"c3c00000",
      114 => x"90001000",   115 => x"3401fffe",   116 => x"a0410800",
      117 => x"d0010000",   118 => x"90201000",   119 => x"3401fffe",
      120 => x"a0410800",   121 => x"d0210000",   122 => x"c3a00000",
      123 => x"90001000",   124 => x"3401fffe",   125 => x"a0410800",
      126 => x"d0010000",   127 => x"90201000",   128 => x"38420001",
      129 => x"d0220000",   130 => x"38210001",   131 => x"d0010000",
      132 => x"c3a00000",   133 => x"379cfff0",   134 => x"5b8b0008",
      135 => x"5b9d0004",   136 => x"f8003778",   137 => x"f80040f2",
      138 => x"f80040e8",   139 => x"78010001",   140 => x"38213490",
      141 => x"f80030f2",   142 => x"34010001",   143 => x"f800369e",
      144 => x"f8003e99",   145 => x"78010001",   146 => x"38218ec0",
      147 => x"58200000",   148 => x"f8003dbf",   149 => x"f80038ad",
      150 => x"34010000",   151 => x"f800347e",   152 => x"34010000",
      153 => x"34020050",   154 => x"f8003ae0",   155 => x"3782000c",
      156 => x"34010000",   157 => x"f8003d50",   158 => x"3402ffff",
      159 => x"5c220010",   160 => x"78010001",   161 => x"382134ac",
      162 => x"f80030dd",   163 => x"34010022",   164 => x"3381000c",
      165 => x"34010033",   166 => x"3381000d",   167 => x"34010044",
      168 => x"3381000e",   169 => x"34010055",   170 => x"3381000f",
      171 => x"34010066",   172 => x"33810010",   173 => x"34010077",
      174 => x"33810011",   175 => x"4384000e",   176 => x"4385000f",
      177 => x"43860010",   178 => x"43870011",   179 => x"4383000d",
      180 => x"4382000c",   181 => x"78010001",   182 => x"382134d0",
      183 => x"f80030c8",   184 => x"378b000c",   185 => x"b9600800",
      186 => x"f8003294",   187 => x"b9600800",   188 => x"f8003894",
      189 => x"34020001",   190 => x"34010001",   191 => x"f80031e1",
      192 => x"f80034f4",   193 => x"f80039aa",   194 => x"f800029f",
      195 => x"78020001",   196 => x"38425e90",   197 => x"34010002",
      198 => x"f800384b",   199 => x"f80045c4",   200 => x"f80026fc",
      201 => x"f8002043",   202 => x"78030001",   203 => x"38635744",
      204 => x"78010001",   205 => x"28620000",   206 => x"38217268",
      207 => x"58200000",   208 => x"78010001",   209 => x"3821f800",
      210 => x"58220000",   211 => x"34010003",   212 => x"f80002eb",
      213 => x"f800029e",   214 => x"78020001",   215 => x"34010000",
      216 => x"38427270",   217 => x"f80039e1",   218 => x"2b9d0004",
      219 => x"2b8b0008",   220 => x"379c0010",   221 => x"c3a00000",
      222 => x"379cfff8",   223 => x"5b8b0008",   224 => x"5b9d0004",
      225 => x"34010000",   226 => x"f80031f0",   227 => x"b8205800",
      228 => x"78010001",   229 => x"38215e94",   230 => x"28240000",
      231 => x"7d620000",   232 => x"64830000",   233 => x"a0431800",
      234 => x"4460000d",   235 => x"78010001",   236 => x"38218f90",
      237 => x"28210000",   238 => x"34020002",   239 => x"58220004",
      240 => x"f80036aa",   241 => x"f8000282",   242 => x"78010001",
      243 => x"38218f88",   244 => x"34020001",   245 => x"58220000",
      246 => x"e0000014",   247 => x"65610000",   248 => x"7c840000",
      249 => x"a0240800",   250 => x"44230012",   251 => x"78010001",
      252 => x"38218f90",   253 => x"28210000",   254 => x"34020002",
      255 => x"58220008",   256 => x"78010001",   257 => x"38218f88",
      258 => x"58220000",   259 => x"f8000296",   260 => x"34010002",
      261 => x"34020000",   262 => x"34030001",   263 => x"f800458f",
      264 => x"34010000",   265 => x"f80039e1",   266 => x"34010001",
      267 => x"e0000008",   268 => x"fc411000",   269 => x"78010001",
      270 => x"c8021000",   271 => x"38218f88",   272 => x"20420003",
      273 => x"58220000",   274 => x"34010000",   275 => x"78020001",
      276 => x"38425e94",   277 => x"584b0000",   278 => x"2b9d0004",
      279 => x"2b8b0008",   280 => x"379c0008",   281 => x"c3a00000",
      282 => x"379cfffc",   283 => x"5b9d0004",   284 => x"f8003623",
      285 => x"78020001",   286 => x"78030001",   287 => x"38637274",
      288 => x"38427278",   289 => x"28640000",   290 => x"28450000",
      291 => x"58610000",   292 => x"340303e8",   293 => x"c8a42000",
      294 => x"b4812000",   295 => x"58440000",   296 => x"34010000",
      297 => x"50640009",   298 => x"78010000",   299 => x"382100a0",
      300 => x"3484fc18",   301 => x"58440000",   302 => x"28220000",
      303 => x"34420001",   304 => x"58220000",   305 => x"34010001",
      306 => x"2b9d0004",   307 => x"379c0004",   308 => x"c3a00000",
      309 => x"379cfffc",   310 => x"5b9d0004",   311 => x"f8003608",
      312 => x"78020001",   313 => x"38427274",   314 => x"58410000",
      315 => x"2b9d0004",   316 => x"379c0004",   317 => x"c3a00000",
      318 => x"379cfff8",   319 => x"5b8b0008",   320 => x"5b9d0004",
      321 => x"78010001",   322 => x"38217268",   323 => x"28220000",
      324 => x"34010001",   325 => x"5c41000f",   326 => x"f8001d5f",
      327 => x"b8205800",   328 => x"f8004059",   329 => x"3402001b",
      330 => x"44220005",   331 => x"78020001",   332 => x"38425e88",
      333 => x"28410000",   334 => x"5c200008",   335 => x"f8001fbd",
      336 => x"78020001",   337 => x"38427268",   338 => x"58400000",
      339 => x"e0000003",   340 => x"f8001fc2",   341 => x"b8205800",
      342 => x"b9600800",   343 => x"2b9d0004",   344 => x"2b8b0008",
      345 => x"379c0008",   346 => x"c3a00000",   347 => x"379cffe0",
      348 => x"5b8b001c",   349 => x"5b8c0018",   350 => x"5b8d0014",
      351 => x"5b8e0010",   352 => x"5b8f000c",   353 => x"5b900008",
      354 => x"5b9d0004",   355 => x"780b0001",   356 => x"780c0001",
      357 => x"f80047ec",   358 => x"396b7114",   359 => x"398c7264",
      360 => x"e0000005",   361 => x"29610008",   362 => x"44200002",
      363 => x"d8200000",   364 => x"356b001c",   365 => x"558bfffc",
      366 => x"780b0001",   367 => x"78010001",   368 => x"396b7114",
      369 => x"780f0001",   370 => x"780d0001",   371 => x"38215748",
      372 => x"39ef7264",   373 => x"39ad7270",   374 => x"282e0000",
      375 => x"b9608000",   376 => x"e0000025",   377 => x"2961000c",
      378 => x"5c200005",   379 => x"29610010",   380 => x"34210001",
      381 => x"59610010",   382 => x"e000000b",   383 => x"29620004",
      384 => x"44400003",   385 => x"28420000",   386 => x"44400007",
      387 => x"d8200000",   388 => x"29620010",   389 => x"b9606000",
      390 => x"b4411000",   391 => x"59620010",   392 => x"5c200002",
      393 => x"ba006000",   394 => x"34010000",   395 => x"37820020",
      396 => x"f800392e",   397 => x"2b820020",   398 => x"29a10000",
      399 => x"c8410800",   400 => x"4c200002",   401 => x"b42e0800",
      402 => x"29830018",   403 => x"b4230800",   404 => x"59810018",
      405 => x"51c10006",   406 => x"c82e0800",   407 => x"59810018",
      408 => x"29810014",   409 => x"34210001",   410 => x"59810014",
      411 => x"59a20000",   412 => x"356b001c",   413 => x"55ebffdc",
      414 => x"f800479a",   415 => x"ba005800",   416 => x"e3fffffd",
      417 => x"379cffbc",   418 => x"5b8b0014",   419 => x"5b8c0010",
      420 => x"5b8d000c",   421 => x"5b8e0008",   422 => x"5b9d0004",
      423 => x"5b830030",   424 => x"78030001",   425 => x"3863727c",
      426 => x"5b82002c",   427 => x"5b840034",   428 => x"5b850038",
      429 => x"5b86003c",   430 => x"5b870040",   431 => x"5b880044",
      432 => x"286d0000",   433 => x"b8205800",   434 => x"b8407000",
      435 => x"34030000",   436 => x"44200002",   437 => x"28230018",
      438 => x"b86d1800",   439 => x"0063001c",   440 => x"4460001b",
      441 => x"780c0001",   442 => x"398c727c",   443 => x"39a10001",
      444 => x"59810000",   445 => x"29610028",   446 => x"37820018",
      447 => x"28230000",   448 => x"b9600800",   449 => x"d8600000",
      450 => x"78030001",   451 => x"3863574c",   452 => x"28620000",
      453 => x"2b81001c",   454 => x"598d0000",   455 => x"296b0334",
      456 => x"f80048bc",   457 => x"780c0001",   458 => x"2b830018",
      459 => x"398c3538",   460 => x"b8202000",   461 => x"b9601000",
      462 => x"b9800800",   463 => x"f8002fb0",   464 => x"b9c00800",
      465 => x"37820030",   466 => x"f8002f8b",   467 => x"2b9d0004",
      468 => x"2b8b0014",   469 => x"2b8c0010",   470 => x"2b8d000c",
      471 => x"2b8e0008",   472 => x"379c0044",   473 => x"c3a00000",
      474 => x"379cfffc",   475 => x"5b9d0004",   476 => x"b8402800",
      477 => x"5c600005",   478 => x"78020001",   479 => x"38423554",
      480 => x"b8a01800",   481 => x"e000000c",   482 => x"34020001",
      483 => x"5c620006",   484 => x"78020001",   485 => x"38423570",
      486 => x"b8a01800",   487 => x"28240008",   488 => x"e0000005",
      489 => x"28240004",   490 => x"78020001",   491 => x"38423588",
      492 => x"b8a01800",   493 => x"fbffffb4",   494 => x"2b9d0004",
      495 => x"379c0004",   496 => x"c3a00000",   497 => x"379cffe8",
      498 => x"5b8b0018",   499 => x"5b8c0014",   500 => x"5b8d0010",
      501 => x"5b8e000c",   502 => x"5b9d0008",   503 => x"b8205800",
      504 => x"b8407000",   505 => x"b8606800",   506 => x"4460001a",
      507 => x"40480000",   508 => x"78020001",   509 => x"384264e4",
      510 => x"2108000f",   511 => x"3d030002",   512 => x"282600e4",
      513 => x"b4431000",   514 => x"28420000",   515 => x"282700e8",
      516 => x"78040001",   517 => x"5b820004",   518 => x"34030001",
      519 => x"34020005",   520 => x"388435a0",   521 => x"b9a02800",
      522 => x"f8000048",   523 => x"34010021",   524 => x"4c2d0006",
      525 => x"b9600800",   526 => x"b9c01000",   527 => x"b9a01800",
      528 => x"f8001607",   529 => x"44200003",   530 => x"340d0000",
      531 => x"340e0000",   532 => x"780c0001",   533 => x"29610000",
      534 => x"398c6374",   535 => x"e000002d",   536 => x"44410003",
      537 => x"358c000c",   538 => x"e000002a",   539 => x"59610004",
      540 => x"2961000c",   541 => x"59600008",   542 => x"44200006",
      543 => x"29820004",   544 => x"b9600800",   545 => x"34030000",
      546 => x"b9a02000",   547 => x"fbffffb7",   548 => x"29840008",
      549 => x"b9a01800",   550 => x"b9600800",   551 => x"b9c01000",
      552 => x"d8800000",   553 => x"b8201800",   554 => x"44200006",
      555 => x"29620334",   556 => x"29840004",   557 => x"78010001",
      558 => x"382135cc",   559 => x"f8002f50",   560 => x"29610004",
      561 => x"29630000",   562 => x"29820004",   563 => x"4461000a",
      564 => x"59610000",   565 => x"34010001",   566 => x"5961000c",
      567 => x"34030002",   568 => x"b9600800",   569 => x"34040000",
      570 => x"fbffffa0",   571 => x"34010000",   572 => x"e000000f",
      573 => x"b9600800",   574 => x"5960000c",   575 => x"34030001",
      576 => x"34040000",   577 => x"fbffff99",   578 => x"29610008",
      579 => x"e0000008",   580 => x"29820000",   581 => x"5c40ffd3",
      582 => x"29620334",   583 => x"78010001",   584 => x"382135e8",
      585 => x"f8002f36",   586 => x"34012710",   587 => x"2b9d0008",
      588 => x"2b8b0018",   589 => x"2b8c0014",   590 => x"2b8d0010",
      591 => x"2b8e000c",   592 => x"379c0018",   593 => x"c3a00000",
      594 => x"379cffe4",   595 => x"5b8b0008",   596 => x"5b9d0004",
      597 => x"5b84000c",   598 => x"5b850010",   599 => x"b8805800",
      600 => x"5b860014",   601 => x"78040001",   602 => x"5b870018",
      603 => x"5b88001c",   604 => x"38843608",   605 => x"34050000",
      606 => x"44200003",   607 => x"28240334",   608 => x"28250018",
      609 => x"78060001",   610 => x"38c6727c",   611 => x"28c10000",
      612 => x"3c420002",   613 => x"b8a12800",   614 => x"80a22800",
      615 => x"20a5000f",   616 => x"5465000c",   617 => x"78050001",
      618 => x"38a5580c",   619 => x"b4a22800",   620 => x"78060001",
      621 => x"28a20000",   622 => x"b8c00800",   623 => x"38213610",
      624 => x"f8002f0f",   625 => x"b9600800",   626 => x"37820010",
      627 => x"f8002eea",   628 => x"2b9d0004",   629 => x"2b8b0008",
      630 => x"379c001c",   631 => x"c3a00000",   632 => x"379cfff8",
      633 => x"5b8b0008",   634 => x"5b9d0004",   635 => x"3402001c",
      636 => x"b8201800",   637 => x"340b0000",   638 => x"3405fffc",
      639 => x"34040003",   640 => x"e0000009",   641 => x"3421ffd0",
      642 => x"202600ff",   643 => x"50860002",   644 => x"e0000008",
      645 => x"bc220800",   646 => x"34630001",   647 => x"b9615800",
      648 => x"3442fffc",   649 => x"40610000",   650 => x"44200007",
      651 => x"5c45fff6",   652 => x"78010001",   653 => x"78020001",
      654 => x"3821361c",   655 => x"384257fc",   656 => x"f8002eef",
      657 => x"b9600800",   658 => x"2b9d0004",   659 => x"2b8b0008",
      660 => x"379c0008",   661 => x"c3a00000",   662 => x"379cfffc",
      663 => x"5b9d0004",   664 => x"34030001",   665 => x"34010003",
      666 => x"34020000",   667 => x"f80043fb",   668 => x"34010000",
      669 => x"34020001",   670 => x"f800458c",   671 => x"34010000",
      672 => x"2b9d0004",   673 => x"379c0004",   674 => x"c3a00000",
      675 => x"379cfff4",   676 => x"5b8b000c",   677 => x"5b8c0008",
      678 => x"5b9d0004",   679 => x"34010000",   680 => x"b8406000",
      681 => x"f80044b7",   682 => x"45800005",   683 => x"642c0000",
      684 => x"c80c6000",   685 => x"398c0001",   686 => x"e000000f",
      687 => x"780b0001",   688 => x"396b7280",   689 => x"5c2c0004",
      690 => x"59600000",   691 => x"340cffff",   692 => x"e0000009",
      693 => x"29610000",   694 => x"340c0001",   695 => x"5c200006",
      696 => x"78020001",   697 => x"34010003",   698 => x"38425e90",
      699 => x"f8003656",   700 => x"596c0000",   701 => x"b9800800",
      702 => x"2b9d0004",   703 => x"2b8b000c",   704 => x"2b8c0008",
      705 => x"379c000c",   706 => x"c3a00000",   707 => x"34010000",
      708 => x"c3a00000",   709 => x"379cfffc",   710 => x"5b9d0004",
      711 => x"34010000",   712 => x"34020001",   713 => x"f8004561",
      714 => x"34010000",   715 => x"2b9d0004",   716 => x"379c0004",
      717 => x"c3a00000",   718 => x"379cfffc",   719 => x"5b9d0004",
      720 => x"282102c8",   721 => x"28210010",   722 => x"2823000c",
      723 => x"44430004",   724 => x"5822000c",   725 => x"b8400800",
      726 => x"f8003814",   727 => x"34010000",   728 => x"2b9d0004",
      729 => x"379c0004",   730 => x"c3a00000",   731 => x"379cfffc",
      732 => x"5b9d0004",   733 => x"f8003806",   734 => x"34020001",
      735 => x"5c200003",   736 => x"f800453a",   737 => x"7c220000",
      738 => x"b8400800",   739 => x"2b9d0004",   740 => x"379c0004",
      741 => x"c3a00000",   742 => x"379cfff8",   743 => x"5b8b0008",
      744 => x"5b9d0004",   745 => x"b8202800",   746 => x"b8220800",
      747 => x"b8402000",   748 => x"b8605800",   749 => x"44200005",
      750 => x"34010001",   751 => x"b8a01000",   752 => x"b8801800",
      753 => x"f800378b",   754 => x"45600005",   755 => x"1562001f",
      756 => x"34010002",   757 => x"b9601800",   758 => x"f8003786",
      759 => x"34010000",   760 => x"2b9d0004",   761 => x"2b8b0008",
      762 => x"379c0008",   763 => x"c3a00000",   764 => x"379cfffc",
      765 => x"5b9d0004",   766 => x"b8201000",   767 => x"3401ffff",
      768 => x"f8004471",   769 => x"34010000",   770 => x"2b9d0004",
      771 => x"379c0004",   772 => x"c3a00000",   773 => x"379cff24",
      774 => x"5b8b0014",   775 => x"5b8c0010",   776 => x"5b8d000c",
      777 => x"5b8e0008",   778 => x"5b9d0004",   779 => x"b8406000",
      780 => x"28220330",   781 => x"b8807000",   782 => x"37810018",
      783 => x"b8605800",   784 => x"b8a06800",   785 => x"f8001d54",
      786 => x"45c00005",   787 => x"78010001",   788 => x"38216d1c",
      789 => x"28210000",   790 => x"59c10000",   791 => x"45a00003",
      792 => x"2b8100cc",   793 => x"59a10000",   794 => x"2b82006c",
      795 => x"3401fffd",   796 => x"44400013",   797 => x"45800007",
      798 => x"2b820060",   799 => x"2b810058",   800 => x"b4410800",
      801 => x"2b8200a0",   802 => x"b4220800",   803 => x"59810000",
      804 => x"2b820068",   805 => x"3401fffd",   806 => x"44400009",
      807 => x"34010000",   808 => x"45600007",   809 => x"2b830064",
      810 => x"2b82005c",   811 => x"b4621000",   812 => x"2b8300a4",
      813 => x"b4431000",   814 => x"59620000",   815 => x"2b9d0004",
      816 => x"2b8b0014",   817 => x"2b8c0010",   818 => x"2b8d000c",
      819 => x"2b8e0008",   820 => x"379c00dc",   821 => x"c3a00000",
      822 => x"34010000",   823 => x"c3a00000",   824 => x"34010000",
      825 => x"c3a00000",   826 => x"379cffec",   827 => x"5b8b000c",
      828 => x"5b8c0008",   829 => x"5b9d0004",   830 => x"34040000",
      831 => x"b8406000",   832 => x"b8605800",   833 => x"37820010",
      834 => x"37830014",   835 => x"34050000",   836 => x"5b800014",
      837 => x"5b800010",   838 => x"fbffffbf",   839 => x"34010001",
      840 => x"5d810003",   841 => x"2b810010",   842 => x"e0000002",
      843 => x"2b810014",   844 => x"59610000",   845 => x"34010001",
      846 => x"2b9d0004",   847 => x"2b8b000c",   848 => x"2b8c0008",
      849 => x"379c0014",   850 => x"c3a00000",   851 => x"379cfffc",
      852 => x"5b9d0004",   853 => x"f8002fbe",   854 => x"34010000",
      855 => x"2b9d0004",   856 => x"379c0004",   857 => x"c3a00000",
      858 => x"379cfffc",   859 => x"5b9d0004",   860 => x"f8002fc2",
      861 => x"34010000",   862 => x"2b9d0004",   863 => x"379c0004",
      864 => x"c3a00000",   865 => x"379cfffc",   866 => x"5b9d0004",
      867 => x"f800349d",   868 => x"f8003e0e",   869 => x"f8003e16",
      870 => x"78010001",   871 => x"78020001",   872 => x"384236bc",
      873 => x"3821368c",   874 => x"f8002e15",   875 => x"34010000",
      876 => x"2b9d0004",   877 => x"379c0004",   878 => x"c3a00000",
      879 => x"78010001",   880 => x"38217284",   881 => x"28210000",
      882 => x"c3a00000",   883 => x"379cfff8",   884 => x"5b8b0008",
      885 => x"5b9d0004",   886 => x"78010001",   887 => x"382136d8",
      888 => x"f8002e07",   889 => x"78010001",   890 => x"78020001",
      891 => x"38426544",   892 => x"3821620c",   893 => x"780b0001",
      894 => x"f800199c",   895 => x"396b5e98",   896 => x"34030000",
      897 => x"b9600800",   898 => x"34020000",   899 => x"fbfffe6e",
      900 => x"78020001",   901 => x"38426250",   902 => x"58410000",
      903 => x"f80033b8",   904 => x"78020001",   905 => x"3842728c",
      906 => x"58410000",   907 => x"296102c8",   908 => x"28210010",
      909 => x"58200068",   910 => x"b9600800",   911 => x"f8000ad5",
      912 => x"78010001",   913 => x"38217288",   914 => x"34020001",
      915 => x"58220000",   916 => x"34010000",   917 => x"2b9d0004",
      918 => x"2b8b0008",   919 => x"379c0008",   920 => x"c3a00000",
      921 => x"379cfff4",   922 => x"5b8b000c",   923 => x"5b8c0008",
      924 => x"5b9d0004",   925 => x"780b0001",   926 => x"396b5e98",
      927 => x"296102c8",   928 => x"282c0010",   929 => x"78010001",
      930 => x"382136e4",   931 => x"f8002ddc",   932 => x"29810000",
      933 => x"34020000",   934 => x"28230034",   935 => x"b9600800",
      936 => x"d8600000",   937 => x"78010001",   938 => x"34020000",
      939 => x"340301b8",   940 => x"59800040",   941 => x"31800035",
      942 => x"38215fa8",   943 => x"f8004801",   944 => x"78010001",
      945 => x"38217288",   946 => x"58200000",   947 => x"b9600800",
      948 => x"0d60010c",   949 => x"f8000aaf",   950 => x"78010001",
      951 => x"3821620c",   952 => x"f80019ab",   953 => x"34010000",
      954 => x"2b9d0004",   955 => x"2b8b000c",   956 => x"2b8c0008",
      957 => x"379c000c",   958 => x"c3a00000",   959 => x"379cffec",
      960 => x"5b8b0014",   961 => x"5b8c0010",   962 => x"5b8d000c",
      963 => x"5b8e0008",   964 => x"5b9d0004",   965 => x"780b0001",
      966 => x"396b5e98",   967 => x"b8206000",   968 => x"296102c8",
      969 => x"282d0010",   970 => x"78010001",   971 => x"38217284",
      972 => x"58200000",   973 => x"fbffffcc",   974 => x"34010002",
      975 => x"45810016",   976 => x"34020003",   977 => x"45820026",
      978 => x"34010001",   979 => x"5d81002e",   980 => x"78010001",
      981 => x"31ac0004",   982 => x"38216544",   983 => x"340e0006",
      984 => x"316c001d",   985 => x"302e0000",   986 => x"34020000",
      987 => x"34010001",   988 => x"34030001",   989 => x"f80042b9",
      990 => x"29610020",   991 => x"2821000c",   992 => x"302e000e",
      993 => x"b9600800",   994 => x"f80012ab",   995 => x"380bea60",
      996 => x"e000001e",   997 => x"34010001",   998 => x"31a10004",
      999 => x"3161001d",  1000 => x"78010001",  1001 => x"38216544",
     1002 => x"340effbb",  1003 => x"302e0000",  1004 => x"34020000",
     1005 => x"34010002",  1006 => x"34030001",  1007 => x"f80042a7",
     1008 => x"29610020",  1009 => x"2821000c",  1010 => x"302e000e",
     1011 => x"b9600800",  1012 => x"f8001299",  1013 => x"340b0fa0",
     1014 => x"e000000c",  1015 => x"31a10004",  1016 => x"3161001d",
     1017 => x"78010001",  1018 => x"38216544",  1019 => x"3402ffff",
     1020 => x"30220000",  1021 => x"34030001",  1022 => x"34010003",
     1023 => x"34020000",  1024 => x"f8004296",  1025 => x"340b0000",
     1026 => x"f800333d",  1027 => x"78020001",  1028 => x"b8207000",
     1029 => x"b8400800",  1030 => x"382136f0",  1031 => x"f8002d78",
     1032 => x"29a20000",  1033 => x"780d0001",  1034 => x"39ad370c",
     1035 => x"28430034",  1036 => x"78020001",  1037 => x"b8400800",
     1038 => x"38215e98",  1039 => x"34020000",  1040 => x"d8600000",
     1041 => x"e000000e",  1042 => x"f8004471",  1043 => x"340103e8",
     1044 => x"f8003330",  1045 => x"f800332a",  1046 => x"c82e1000",
     1047 => x"51620006",  1048 => x"78010001",  1049 => x"382136fc",
     1050 => x"f8002d65",  1051 => x"340bff8c",  1052 => x"e0000008",
     1053 => x"b9a00800",  1054 => x"f8002d61",  1055 => x"34010000",
     1056 => x"f8004340",  1057 => x"5c200002",  1058 => x"5d61fff0",
     1059 => x"340b0000",  1060 => x"78010001",  1061 => x"38214adc",
     1062 => x"f8002d59",  1063 => x"7d620000",  1064 => x"65810001",
     1065 => x"a0410800",  1066 => x"44200005",  1067 => x"78010001",
     1068 => x"38216544",  1069 => x"34020034",  1070 => x"30220000",
     1071 => x"78010001",  1072 => x"38217284",  1073 => x"582c0000",
     1074 => x"b9600800",  1075 => x"2b9d0004",  1076 => x"2b8b0014",
     1077 => x"2b8c0010",  1078 => x"2b8d000c",  1079 => x"2b8e0008",
     1080 => x"379c0014",  1081 => x"c3a00000",  1082 => x"379cffec",
     1083 => x"5b8b0014",  1084 => x"5b8c0010",  1085 => x"5b8d000c",
     1086 => x"5b8e0008",  1087 => x"5b9d0004",  1088 => x"78010001",
     1089 => x"38217288",  1090 => x"28210000",  1091 => x"340e0000",
     1092 => x"44200024",  1093 => x"780b0001",  1094 => x"396b5e98",
     1095 => x"29610024",  1096 => x"29620038",  1097 => x"78040001",
     1098 => x"28250008",  1099 => x"3403007c",  1100 => x"b9600800",
     1101 => x"38845f7c",  1102 => x"d8a00000",  1103 => x"b8201800",
     1104 => x"4c010005",  1105 => x"29610370",  1106 => x"34210001",
     1107 => x"59610370",  1108 => x"e000000c",  1109 => x"5c20000b",
     1110 => x"780d0001",  1111 => x"f80032e8",  1112 => x"39ad728c",
     1113 => x"29a20000",  1114 => x"780c0001",  1115 => x"398c6250",
     1116 => x"c8220800",  1117 => x"29820000",  1118 => x"5441000a",
     1119 => x"e0000011",  1120 => x"78010001",  1121 => x"38215e98",
     1122 => x"28220040",  1123 => x"fbfffd8e",  1124 => x"78020001",
     1125 => x"38426250",  1126 => x"58410000",  1127 => x"340e0001",
     1128 => x"b9c00800",  1129 => x"2b9d0004",  1130 => x"2b8b0014",
     1131 => x"2b8c0010",  1132 => x"2b8d000c",  1133 => x"2b8e0008",
     1134 => x"379c0014",  1135 => x"c3a00000",  1136 => x"f80032cf",
     1137 => x"59a10000",  1138 => x"34020000",  1139 => x"b9600800",
     1140 => x"34030000",  1141 => x"fbfffd7c",  1142 => x"59810000",
     1143 => x"e3fffff0",  1144 => x"379cffe8",  1145 => x"5b9d0018",
     1146 => x"b8205000",  1147 => x"40610005",  1148 => x"40640000",
     1149 => x"40650001",  1150 => x"40660002",  1151 => x"40670003",
     1152 => x"40680004",  1153 => x"5b810004",  1154 => x"40610006",
     1155 => x"b8404800",  1156 => x"b9401000",  1157 => x"5b810008",
     1158 => x"40610007",  1159 => x"5b81000c",  1160 => x"40610008",
     1161 => x"5b810010",  1162 => x"40610009",  1163 => x"b9201800",
     1164 => x"5b810014",  1165 => x"78010001",  1166 => x"38213714",
     1167 => x"f8002cf0",  1168 => x"2b9d0018",  1169 => x"379c0018",
     1170 => x"c3a00000",  1171 => x"379cffd0",  1172 => x"5b8b0030",
     1173 => x"5b8c002c",  1174 => x"5b8d0028",  1175 => x"5b8e0024",
     1176 => x"5b8f0020",  1177 => x"5b90001c",  1178 => x"5b910018",
     1179 => x"5b920014",  1180 => x"5b930010",  1181 => x"5b94000c",
     1182 => x"5b950008",  1183 => x"5b9d0004",  1184 => x"b8603000",
     1185 => x"b8209800",  1186 => x"b8409000",  1187 => x"78010001",
     1188 => x"b880a800",  1189 => x"3821374c",  1190 => x"ba601000",
     1191 => x"ba401800",  1192 => x"b8c02000",  1193 => x"b8a0a000",
     1194 => x"78110001",  1195 => x"f8002cd4",  1196 => x"78100001",
     1197 => x"780f0001",  1198 => x"780e0001",  1199 => x"780d0001",
     1200 => x"b8205800",  1201 => x"340c0000",  1202 => x"3a313760",
     1203 => x"3a103768",  1204 => x"39ef4c00",  1205 => x"39ce4adc",
     1206 => x"39ad495c",  1207 => x"e0000017",  1208 => x"5cc00006",
     1209 => x"ba200800",  1210 => x"ba601000",  1211 => x"ba401800",
     1212 => x"f8002cc3",  1213 => x"b5615800",  1214 => x"b6ac1000",
     1215 => x"40420000",  1216 => x"ba000800",  1217 => x"358c0001",
     1218 => x"f8002cbd",  1219 => x"21820003",  1220 => x"b42b5800",
     1221 => x"b9e03000",  1222 => x"5c400005",  1223 => x"2181000f",
     1224 => x"b9c03000",  1225 => x"44220002",  1226 => x"b9a03000",
     1227 => x"b8c00800",  1228 => x"f8002cb3",  1229 => x"b5615800",
     1230 => x"2186000f",  1231 => x"4a8cffe9",  1232 => x"44c00005",
     1233 => x"78010001",  1234 => x"38214adc",  1235 => x"f8002cac",
     1236 => x"b42b5800",  1237 => x"b9600800",  1238 => x"2b9d0004",
     1239 => x"2b8b0030",  1240 => x"2b8c002c",  1241 => x"2b8d0028",
     1242 => x"2b8e0024",  1243 => x"2b8f0020",  1244 => x"2b90001c",
     1245 => x"2b910018",  1246 => x"2b920014",  1247 => x"2b930010",
     1248 => x"2b94000c",  1249 => x"2b950008",  1250 => x"379c0030",
     1251 => x"c3a00000",  1252 => x"379cffb8",  1253 => x"5b8b0048",
     1254 => x"5b8c0044",  1255 => x"5b8d0040",  1256 => x"5b8e003c",
     1257 => x"5b8f0038",  1258 => x"5b900034",  1259 => x"5b910030",
     1260 => x"5b92002c",  1261 => x"5b930028",  1262 => x"5b940024",
     1263 => x"5b950020",  1264 => x"5b96001c",  1265 => x"5b970018",
     1266 => x"5b980014",  1267 => x"5b9d0010",  1268 => x"b8608000",
     1269 => x"40430001",  1270 => x"b8206000",  1271 => x"34010002",
     1272 => x"2063000f",  1273 => x"b8406800",  1274 => x"404e0000",
     1275 => x"44610006",  1276 => x"78010001",  1277 => x"b9801000",
     1278 => x"38213770",  1279 => x"f8002c80",  1280 => x"e000013f",
     1281 => x"40450002",  1282 => x"40460003",  1283 => x"21ce000f",
     1284 => x"3ca50008",  1285 => x"78010001",  1286 => x"b8c52800",
     1287 => x"41a60004",  1288 => x"34030002",  1289 => x"b9c02000",
     1290 => x"344b0022",  1291 => x"38213790",  1292 => x"b9801000",
     1293 => x"f8002c72",  1294 => x"41a2000c",  1295 => x"41a1000d",
     1296 => x"41a4000e",  1297 => x"41a30006",  1298 => x"3c420018",
     1299 => x"3c210010",  1300 => x"41a60007",  1301 => x"41a5000f",
     1302 => x"3c840008",  1303 => x"b8220800",  1304 => x"3c630008",
     1305 => x"b8812000",  1306 => x"78010001",  1307 => x"b8c31800",
     1308 => x"b8a42000",  1309 => x"b9801000",  1310 => x"382137bc",
     1311 => x"f8002c60",  1312 => x"78020001",  1313 => x"b9800800",
     1314 => x"384237e0",  1315 => x"35a30014",  1316 => x"fbffff54",
     1317 => x"41a3001e",  1318 => x"41a4001f",  1319 => x"41a50021",
     1320 => x"3c630008",  1321 => x"78010001",  1322 => x"b8831800",
     1323 => x"41a40020",  1324 => x"382137e8",  1325 => x"b9801000",
     1326 => x"f8002c51",  1327 => x"3401000c",  1328 => x"55c100d1",
     1329 => x"78010001",  1330 => x"3dce0002",  1331 => x"3821582c",
     1332 => x"b42e0800",  1333 => x"28210000",  1334 => x"c0200000",
     1335 => x"78010001",  1336 => x"b9801000",  1337 => x"38213814",
     1338 => x"f8002c45",  1339 => x"41620002",  1340 => x"41610003",
     1341 => x"41640004",  1342 => x"3c420018",  1343 => x"3c210010",
     1344 => x"3c840008",  1345 => x"b8220800",  1346 => x"b8812000",
     1347 => x"41620006",  1348 => x"41610007",  1349 => x"41650008",
     1350 => x"3c420018",  1351 => x"3c210010",  1352 => x"3ca50008",
     1353 => x"b8220800",  1354 => x"b8a12800",  1355 => x"78030001",
     1356 => x"78010001",  1357 => x"41670005",  1358 => x"41660009",
     1359 => x"3821382c",  1360 => x"b9801000",  1361 => x"3863383c",
     1362 => x"e000001c",  1363 => x"78010001",  1364 => x"b9801000",
     1365 => x"38213848",  1366 => x"f8002c29",  1367 => x"41620002",
     1368 => x"41610003",  1369 => x"41640004",  1370 => x"3c420018",
     1371 => x"3c210010",  1372 => x"3c840008",  1373 => x"b8220800",
     1374 => x"b8812000",  1375 => x"41620006",  1376 => x"41610007",
     1377 => x"41650008",  1378 => x"3c420018",  1379 => x"3c210010",
     1380 => x"3ca50008",  1381 => x"b8220800",  1382 => x"41670005",
     1383 => x"41660009",  1384 => x"b8a12800",  1385 => x"78030001",
     1386 => x"78010001",  1387 => x"3821382c",  1388 => x"b9801000",
     1389 => x"38633864",  1390 => x"b8e42000",  1391 => x"b8c52800",
     1392 => x"f8002c0f",  1393 => x"e000008e",  1394 => x"78010001",
     1395 => x"b9801000",  1396 => x"38213874",  1397 => x"f8002c0a",
     1398 => x"41620002",  1399 => x"41610003",  1400 => x"41640004",
     1401 => x"3c420018",  1402 => x"3c210010",  1403 => x"3c840008",
     1404 => x"b8220800",  1405 => x"b8812000",  1406 => x"41620006",
     1407 => x"41610007",  1408 => x"41650008",  1409 => x"3c420018",
     1410 => x"3c210010",  1411 => x"3ca50008",  1412 => x"b8220800",
     1413 => x"b8a12800",  1414 => x"78030001",  1415 => x"78010001",
     1416 => x"41670005",  1417 => x"41660009",  1418 => x"3821382c",
     1419 => x"b9801000",  1420 => x"38633890",  1421 => x"e3ffffe1",
     1422 => x"78010001",  1423 => x"b9801000",  1424 => x"382138a0",
     1425 => x"f8002bee",  1426 => x"41620002",  1427 => x"41610003",
     1428 => x"41640004",  1429 => x"3c420018",  1430 => x"3c210010",
     1431 => x"3c840008",  1432 => x"b8220800",  1433 => x"b8812000",
     1434 => x"41620006",  1435 => x"41610007",  1436 => x"41650008",
     1437 => x"3c420018",  1438 => x"3c210010",  1439 => x"41670005",
     1440 => x"41660009",  1441 => x"3ca50008",  1442 => x"b8220800",
     1443 => x"780e0001",  1444 => x"39ce38bc",  1445 => x"b8a12800",
     1446 => x"78010001",  1447 => x"b9801000",  1448 => x"b9c01800",
     1449 => x"b8e42000",  1450 => x"b8c52800",  1451 => x"3821382c",
     1452 => x"f8002bd3",  1453 => x"3563000a",  1454 => x"b9800800",
     1455 => x"b9c01000",  1456 => x"fbfffec8",  1457 => x"340b0036",
     1458 => x"e0000080",  1459 => x"78010001",  1460 => x"b9801000",
     1461 => x"382138d0",  1462 => x"f8002bc9",  1463 => x"41620002",
     1464 => x"41610003",  1465 => x"41640004",  1466 => x"3c420018",
     1467 => x"3c210010",  1468 => x"3c840008",  1469 => x"b8220800",
     1470 => x"b8812000",  1471 => x"41620006",  1472 => x"41610007",
     1473 => x"41650008",  1474 => x"3c420018",  1475 => x"3c210010",
     1476 => x"41670005",  1477 => x"41660009",  1478 => x"3ca50008",
     1479 => x"b8220800",  1480 => x"b8a12800",  1481 => x"78030001",
     1482 => x"78010001",  1483 => x"b8e42000",  1484 => x"b8c52800",
     1485 => x"b9801000",  1486 => x"386338ec",  1487 => x"3821382c",
     1488 => x"f8002baf",  1489 => x"41660010",  1490 => x"41670011",
     1491 => x"4165000f",  1492 => x"4164000e",  1493 => x"3cc60008",
     1494 => x"78010001",  1495 => x"78030001",  1496 => x"b8e63000",
     1497 => x"b9801000",  1498 => x"38633918",  1499 => x"38213904",
     1500 => x"f8002ba3",  1501 => x"4163000d",  1502 => x"41640012",
     1503 => x"78010001",  1504 => x"b9801000",  1505 => x"3821393c",
     1506 => x"f8002b9d",  1507 => x"41610018",  1508 => x"41640013",
     1509 => x"41650014",  1510 => x"41660015",  1511 => x"41670016",
     1512 => x"41680017",  1513 => x"5b810004",  1514 => x"41610019",
     1515 => x"78030001",  1516 => x"b9801000",  1517 => x"5b810008",
     1518 => x"4161001a",  1519 => x"38633994",  1520 => x"340b0040",
     1521 => x"5b81000c",  1522 => x"78010001",  1523 => x"38213964",
     1524 => x"f8002b8b",  1525 => x"e000003d",  1526 => x"78010001",
     1527 => x"b9801000",  1528 => x"382139b4",  1529 => x"f8002b86",
     1530 => x"78020001",  1531 => x"b9800800",  1532 => x"384239d0",
     1533 => x"b9601800",  1534 => x"fbfffe7a",  1535 => x"340b002c",
     1536 => x"e0000032",  1537 => x"340b0022",  1538 => x"e0000030",
     1539 => x"55f70009",  1540 => x"78010001",  1541 => x"b9801000",
     1542 => x"ba001800",  1543 => x"b9602000",  1544 => x"b9e02800",
     1545 => x"382139ec",  1546 => x"f8002b75",  1547 => x"e0000034",
     1548 => x"b5ab7000",  1549 => x"41d60002",  1550 => x"41c10003",
     1551 => x"41c30000",  1552 => x"3ed60008",  1553 => x"41c40001",
     1554 => x"b836b000",  1555 => x"41c10008",  1556 => x"41c50004",
     1557 => x"41c60005",  1558 => x"41c70006",  1559 => x"41c80007",
     1560 => x"5b810004",  1561 => x"41c10009",  1562 => x"3c630008",
     1563 => x"36d10004",  1564 => x"5b810008",  1565 => x"b8831800",
     1566 => x"baa00800",  1567 => x"b9801000",  1568 => x"ba202000",
     1569 => x"f8002b5e",  1570 => x"4df10007",  1571 => x"ba400800",
     1572 => x"b9801000",  1573 => x"ba201800",  1574 => x"b9e02000",
     1575 => x"f8002b58",  1576 => x"e0000008",  1577 => x"b9800800",
     1578 => x"ba801000",  1579 => x"ba601800",  1580 => x"35c4000a",
     1581 => x"36c5fffa",  1582 => x"fbfffe65",  1583 => x"ba207800",
     1584 => x"b56f5800",  1585 => x"e000000b",  1586 => x"78150001",
     1587 => x"78140001",  1588 => x"78130001",  1589 => x"78120001",
     1590 => x"34180002",  1591 => x"34170009",  1592 => x"3ab53a10",
     1593 => x"3a943a7c",  1594 => x"3a733a84",  1595 => x"3a523a50",
     1596 => x"4d700003",  1597 => x"ca0b7800",  1598 => x"49f8ffc5",
     1599 => x"78020001",  1600 => x"78030001",  1601 => x"b9800800",
     1602 => x"38423a90",  1603 => x"38633a98",  1604 => x"b9a02000",
     1605 => x"ba002800",  1606 => x"fbfffe4d",  1607 => x"2b9d0010",
     1608 => x"2b8b0048",  1609 => x"2b8c0044",  1610 => x"2b8d0040",
     1611 => x"2b8e003c",  1612 => x"2b8f0038",  1613 => x"2b900034",
     1614 => x"2b910030",  1615 => x"2b92002c",  1616 => x"2b930028",
     1617 => x"2b940024",  1618 => x"2b950020",  1619 => x"2b96001c",
     1620 => x"2b970018",  1621 => x"2b980014",  1622 => x"379c0048",
     1623 => x"c3a00000",  1624 => x"379cfff0",  1625 => x"5b8b0010",
     1626 => x"5b8c000c",  1627 => x"5b8d0008",  1628 => x"5b9d0004",
     1629 => x"b8205800",  1630 => x"b8406800",  1631 => x"b8606000",
     1632 => x"4480000f",  1633 => x"2881000c",  1634 => x"78070001",
     1635 => x"28850000",  1636 => x"28860004",  1637 => x"38e75740",
     1638 => x"5c200003",  1639 => x"78070001",  1640 => x"38e73aa0",
     1641 => x"78010001",  1642 => x"38213aac",  1643 => x"b9601000",
     1644 => x"b8a01800",  1645 => x"b8a02000",  1646 => x"f8002b11",
     1647 => x"b9600800",  1648 => x"b9a01000",  1649 => x"b9801800",
     1650 => x"fbfffe72",  1651 => x"34010000",  1652 => x"2b9d0004",
     1653 => x"2b8b0010",  1654 => x"2b8c000c",  1655 => x"2b8d0008",
     1656 => x"379c0010",  1657 => x"c3a00000",  1658 => x"379cffe8",
     1659 => x"5b8b0018",  1660 => x"5b8c0014",  1661 => x"5b8d0010",
     1662 => x"5b8e000c",  1663 => x"5b8f0008",  1664 => x"5b9d0004",
     1665 => x"282d0000",  1666 => x"b8207800",  1667 => x"282e0004",
     1668 => x"b8406000",  1669 => x"340b0000",  1670 => x"34010000",
     1671 => x"34040000",  1672 => x"544d0006",  1673 => x"b9a00800",
     1674 => x"f8004447",  1675 => x"882c1000",  1676 => x"b9602000",
     1677 => x"c9a26800",  1678 => x"34030000",  1679 => x"34020001",
     1680 => x"e000000b",  1681 => x"3d850001",  1682 => x"3d6b0001",
     1683 => x"f5856000",  1684 => x"3c630001",  1685 => x"b58b5800",
     1686 => x"b8a06000",  1687 => x"3c450001",  1688 => x"f4451000",
     1689 => x"b4431800",  1690 => x"b8a01000",  1691 => x"1565001f",
     1692 => x"c8ac3000",  1693 => x"f4c53000",  1694 => x"c8ab2800",
     1695 => x"c8a62800",  1696 => x"00a5001f",  1697 => x"34060001",
     1698 => x"55ab0004",  1699 => x"5dab0002",  1700 => x"55cc0002",
     1701 => x"34060000",  1702 => x"a0a63000",  1703 => x"5cc0ffea",
     1704 => x"556d000d",  1705 => x"5d6d0002",  1706 => x"558e000b",
     1707 => x"c9cc2800",  1708 => x"f4ae7000",  1709 => x"c9ab6800",
     1710 => x"c9ae6800",  1711 => x"b8a07000",  1712 => x"b4822800",
     1713 => x"f4852000",  1714 => x"b4230800",  1715 => x"b4810800",
     1716 => x"b8a02000",  1717 => x"3c65001f",  1718 => x"00420001",
     1719 => x"00630001",  1720 => x"b8a21000",  1721 => x"b8622800",
     1722 => x"44a00006",  1723 => x"3d65001f",  1724 => x"018c0001",
     1725 => x"016b0001",  1726 => x"b8ac6000",  1727 => x"e3ffffe9",
     1728 => x"59e10000",  1729 => x"b9c00800",  1730 => x"59e40004",
     1731 => x"2b9d0004",  1732 => x"2b8b0018",  1733 => x"2b8c0014",
     1734 => x"2b8d0010",  1735 => x"2b8e000c",  1736 => x"2b8f0008",
     1737 => x"379c0018",  1738 => x"c3a00000",  1739 => x"379cfff8",
     1740 => x"5b8b0008",  1741 => x"5b9d0004",  1742 => x"b8405800",
     1743 => x"f8003070",  1744 => x"b42b0800",  1745 => x"5c200002",
     1746 => x"34010001",  1747 => x"2b9d0004",  1748 => x"2b8b0008",
     1749 => x"379c0008",  1750 => x"c3a00000",  1751 => x"379cfff8",
     1752 => x"5b8b0008",  1753 => x"5b9d0004",  1754 => x"78040001",
     1755 => x"b8405800",  1756 => x"78050001",  1757 => x"34020006",
     1758 => x"34030001",  1759 => x"38843b78",  1760 => x"38a55860",
     1761 => x"b9603000",  1762 => x"fbfffb70",  1763 => x"45600005",
     1764 => x"1562001f",  1765 => x"34010002",  1766 => x"b9601800",
     1767 => x"f8003395",  1768 => x"34010000",  1769 => x"2b9d0004",
     1770 => x"2b8b0008",  1771 => x"379c0008",  1772 => x"c3a00000",
     1773 => x"379cfff4",  1774 => x"5b8b000c",  1775 => x"5b8c0008",
     1776 => x"5b9d0004",  1777 => x"b8206000",  1778 => x"b8405800",
     1779 => x"b8603000",  1780 => x"44600008",  1781 => x"78040001",
     1782 => x"78050001",  1783 => x"34020006",  1784 => x"34030001",
     1785 => x"38843b84",  1786 => x"38a55878",  1787 => x"fbfffb57",
     1788 => x"b9800800",  1789 => x"b9601000",  1790 => x"fbffffd9",
     1791 => x"2b9d0004",  1792 => x"2b8b000c",  1793 => x"2b8c0008",
     1794 => x"379c000c",  1795 => x"c3a00000",  1796 => x"379cfff0",
     1797 => x"5b8b0010",  1798 => x"5b8c000c",  1799 => x"5b8d0008",
     1800 => x"5b9d0004",  1801 => x"b8206800",  1802 => x"44400012",
     1803 => x"284b0000",  1804 => x"284c0004",  1805 => x"34040003",
     1806 => x"1561001f",  1807 => x"b9601000",  1808 => x"b9801800",
     1809 => x"f8003389",  1810 => x"78040001",  1811 => x"78050001",
     1812 => x"b9a00800",  1813 => x"34020006",  1814 => x"34030001",
     1815 => x"38843bb0",  1816 => x"38a5588c",  1817 => x"b9603000",
     1818 => x"b9803800",  1819 => x"fbfffb37",  1820 => x"34010000",
     1821 => x"2b9d0004",  1822 => x"2b8b0010",  1823 => x"2b8c000c",
     1824 => x"2b8d0008",  1825 => x"379c0010",  1826 => x"c3a00000",
     1827 => x"379cffe8",  1828 => x"5b8b000c",  1829 => x"5b8c0008",
     1830 => x"5b9d0004",  1831 => x"b8405800",  1832 => x"b8206000",
     1833 => x"37820018",  1834 => x"37810010",  1835 => x"f800338f",
     1836 => x"78020001",  1837 => x"3842727c",  1838 => x"2b860014",
     1839 => x"2b870018",  1840 => x"28410000",  1841 => x"59660000",
     1842 => x"59670004",  1843 => x"20210001",  1844 => x"5c200009",
     1845 => x"78040001",  1846 => x"78050001",  1847 => x"b9800800",
     1848 => x"34020006",  1849 => x"34030002",  1850 => x"38843bb0",
     1851 => x"38a5589c",  1852 => x"fbfffb16",  1853 => x"34010000",
     1854 => x"2b9d0004",  1855 => x"2b8b000c",  1856 => x"2b8c0008",
     1857 => x"379c0018",  1858 => x"c3a00000",  1859 => x"379cffb0",
     1860 => x"5b8b001c",  1861 => x"5b8c0018",  1862 => x"5b8d0014",
     1863 => x"5b8e0010",  1864 => x"5b8f000c",  1865 => x"5b900008",
     1866 => x"5b9d0004",  1867 => x"28300058",  1868 => x"378c0040",
     1869 => x"b8407800",  1870 => x"b8206800",  1871 => x"78020001",
     1872 => x"340188f7",  1873 => x"b8607000",  1874 => x"0f81004c",
     1875 => x"384257f4",  1876 => x"b9800800",  1877 => x"34030006",
     1878 => x"b8805800",  1879 => x"f80043db",  1880 => x"b9801000",
     1881 => x"ba000800",  1882 => x"b9e01800",  1883 => x"b9c02000",
     1884 => x"37850020",  1885 => x"f800227f",  1886 => x"b8206000",
     1887 => x"45600011",  1888 => x"2b81003c",  1889 => x"2b870024",
     1890 => x"2b880028",  1891 => x"78040001",  1892 => x"78050001",
     1893 => x"5961000c",  1894 => x"59670000",  1895 => x"59680004",
     1896 => x"59600008",  1897 => x"b9a00800",  1898 => x"34020005",
     1899 => x"34030002",  1900 => x"38843bc0",  1901 => x"38a558ac",
     1902 => x"b9803000",  1903 => x"fbfffae3",  1904 => x"4c0c0010",
     1905 => x"78010001",  1906 => x"3821727c",  1907 => x"28220000",
     1908 => x"29a10018",  1909 => x"b8410800",  1910 => x"00210014",
     1911 => x"34020001",  1912 => x"2021000f",  1913 => x"50410007",
     1914 => x"78010001",  1915 => x"38213be0",  1916 => x"b9e01000",
     1917 => x"b9c01800",  1918 => x"b9602000",  1919 => x"fbfffed9",
     1920 => x"b9800800",  1921 => x"2b9d0004",  1922 => x"2b8b001c",
     1923 => x"2b8c0018",  1924 => x"2b8d0014",  1925 => x"2b8e0010",
     1926 => x"2b8f000c",  1927 => x"2b900008",  1928 => x"379c0050",
     1929 => x"c3a00000",  1930 => x"379cffb8",  1931 => x"5b8b0014",
     1932 => x"5b8c0010",  1933 => x"5b8d000c",  1934 => x"5b8e0008",
     1935 => x"5b9d0004",  1936 => x"b8207000",  1937 => x"28210058",
     1938 => x"b8602800",  1939 => x"b8406800",  1940 => x"b8805800",
     1941 => x"37820038",  1942 => x"b8a02000",  1943 => x"b9a01800",
     1944 => x"37850018",  1945 => x"f80021d1",  1946 => x"b8206000",
     1947 => x"4560000b",  1948 => x"2b81001c",  1949 => x"59610000",
     1950 => x"2b810020",  1951 => x"59610004",  1952 => x"2b810024",
     1953 => x"59610008",  1954 => x"2b810034",  1955 => x"5961000c",
     1956 => x"2b810030",  1957 => x"59610010",  1958 => x"4c0c0010",
     1959 => x"78040001",  1960 => x"3884727c",  1961 => x"28820000",
     1962 => x"29c10018",  1963 => x"b8410800",  1964 => x"00210014",
     1965 => x"34020001",  1966 => x"2021000f",  1967 => x"50410007",
     1968 => x"78010001",  1969 => x"38213be8",  1970 => x"b9a01000",
     1971 => x"b9801800",  1972 => x"b9602000",  1973 => x"fbfffea3",
     1974 => x"b9800800",  1975 => x"2b9d0004",  1976 => x"2b8b0014",
     1977 => x"2b8c0010",  1978 => x"2b8d000c",  1979 => x"2b8e0008",
     1980 => x"379c0048",  1981 => x"c3a00000",  1982 => x"379cfffc",
     1983 => x"5b9d0004",  1984 => x"28210058",  1985 => x"f800214f",
     1986 => x"34010000",  1987 => x"2b9d0004",  1988 => x"379c0004",
     1989 => x"c3a00000",  1990 => x"379cffd4",  1991 => x"5b8b0010",
     1992 => x"5b8c000c",  1993 => x"5b8d0008",  1994 => x"5b9d0004",
     1995 => x"b8205800",  1996 => x"28210058",  1997 => x"44200002",
     1998 => x"f8002142",  1999 => x"b9600800",  2000 => x"f8000d2a",
     2001 => x"378c0014",  2002 => x"340188f7",  2003 => x"78020001",
     2004 => x"0f810020",  2005 => x"384257f4",  2006 => x"b9800800",
     2007 => x"34030006",  2008 => x"f800435a",  2009 => x"78010001",
     2010 => x"b9801000",  2011 => x"38216340",  2012 => x"34030001",
     2013 => x"34040000",  2014 => x"f80020e9",  2015 => x"b8206000",
     2016 => x"4420000e",  2017 => x"378d0028",  2018 => x"b9a01000",
     2019 => x"f80020d3",  2020 => x"b9a01000",  2021 => x"34030006",
     2022 => x"35610060",  2023 => x"f800434b",  2024 => x"3561004c",
     2025 => x"596c0058",  2026 => x"b9a01000",  2027 => x"34030006",
     2028 => x"f8004346",  2029 => x"596c0044",  2030 => x"34010000",
     2031 => x"2b9d0004",  2032 => x"2b8b0010",  2033 => x"2b8c000c",
     2034 => x"2b8d0008",  2035 => x"379c002c",  2036 => x"c3a00000",
     2037 => x"379cfff8",  2038 => x"5b8b0008",  2039 => x"5b9d0004",
     2040 => x"78040001",  2041 => x"78050001",  2042 => x"34020002",
     2043 => x"34030002",  2044 => x"38843cd4",  2045 => x"38a5590c",
     2046 => x"b8205800",  2047 => x"fbfffa53",  2048 => x"296302c8",
     2049 => x"28610010",  2050 => x"28220064",  2051 => x"34010000",
     2052 => x"44400010",  2053 => x"34010001",  2054 => x"59610004",
     2055 => x"1061000b",  2056 => x"4062000c",  2057 => x"29640028",
     2058 => x"bc411000",  2059 => x"28830018",  2060 => x"084203e8",
     2061 => x"b9600800",  2062 => x"d8600000",  2063 => x"596102d4",
     2064 => x"296102c8",  2065 => x"28210010",  2066 => x"58200064",
     2067 => x"34010001",  2068 => x"2b9d0004",  2069 => x"2b8b0008",
     2070 => x"379c0008",  2071 => x"c3a00000",  2072 => x"379cfff4",
     2073 => x"5b8b000c",  2074 => x"5b8c0008",  2075 => x"5b9d0004",
     2076 => x"78040001",  2077 => x"78050001",  2078 => x"b8606000",
     2079 => x"34020002",  2080 => x"34030002",  2081 => x"38843cd4",
     2082 => x"38a55920",  2083 => x"b8205800",  2084 => x"fbfffa2e",
     2085 => x"29820024",  2086 => x"296102c8",  2087 => x"20430003",
     2088 => x"28210010",  2089 => x"7c640000",  2090 => x"58240038",
     2091 => x"20440008",  2092 => x"20420004",  2093 => x"7c840000",
     2094 => x"7c420000",  2095 => x"30230035",  2096 => x"58220044",
     2097 => x"58240040",  2098 => x"29610020",  2099 => x"28220010",
     2100 => x"296102c8",  2101 => x"2c210008",  2102 => x"0c41002c",
     2103 => x"2b9d0004",  2104 => x"2b8b000c",  2105 => x"2b8c0008",
     2106 => x"379c000c",  2107 => x"c3a00000",  2108 => x"379cfff8",
     2109 => x"5b8b0008",  2110 => x"5b9d0004",  2111 => x"282202c8",
     2112 => x"78040001",  2113 => x"78050001",  2114 => x"284b0010",
     2115 => x"34030002",  2116 => x"34020002",  2117 => x"38843cd4",
     2118 => x"38a55958",  2119 => x"fbfffa0b",  2120 => x"34010000",
     2121 => x"31600005",  2122 => x"2b9d0004",  2123 => x"2b8b0008",
     2124 => x"379c0008",  2125 => x"c3a00000",  2126 => x"379cfff8",
     2127 => x"5b8b0008",  2128 => x"5b9d0004",  2129 => x"78040001",
     2130 => x"78050001",  2131 => x"b8205800",  2132 => x"34020002",
     2133 => x"34010000",  2134 => x"34030002",  2135 => x"38843cd4",
     2136 => x"38a55968",  2137 => x"fbfff9f9",  2138 => x"29610024",
     2139 => x"44200006",  2140 => x"34020000",  2141 => x"34030001",
     2142 => x"34040002",  2143 => x"34060003",  2144 => x"e000001f",
     2145 => x"29610000",  2146 => x"29620040",  2147 => x"58220014",
     2148 => x"e000001d",  2149 => x"29650000",  2150 => x"08410374",
     2151 => x"b4a10800",  2152 => x"29650040",  2153 => x"58250014",
     2154 => x"28250368",  2155 => x"5ca30010",  2156 => x"4025001d",
     2157 => x"44a30004",  2158 => x"282102c8",  2159 => x"5ca40009",
     2160 => x"e0000005",  2161 => x"282102c8",  2162 => x"28210010",
     2163 => x"30230004",  2164 => x"e000000a",  2165 => x"28210010",
     2166 => x"30240004",  2167 => x"e0000007",  2168 => x"28210010",
     2169 => x"30260004",  2170 => x"e0000004",  2171 => x"282102c8",
     2172 => x"28210010",  2173 => x"30200004",  2174 => x"34420001",
     2175 => x"29610024",  2176 => x"4822ffe5",  2177 => x"34010000",
     2178 => x"2b9d0004",  2179 => x"2b8b0008",  2180 => x"379c0008",
     2181 => x"c3a00000",  2182 => x"379cfff4",  2183 => x"5b8b000c",
     2184 => x"5b8c0008",  2185 => x"5b9d0004",  2186 => x"282202c8",
     2187 => x"78040001",  2188 => x"78050001",  2189 => x"284b0010",
     2190 => x"34030002",  2191 => x"34020002",  2192 => x"38843cd4",
     2193 => x"38a55970",  2194 => x"b8206000",  2195 => x"fbfff9bf",
     2196 => x"41630004",  2197 => x"3401012c",  2198 => x"59610028",
     2199 => x"34020001",  2200 => x"34010bb8",  2201 => x"59610030",
     2202 => x"59600008",  2203 => x"31600035",  2204 => x"59600040",
     2205 => x"59620014",  2206 => x"20630003",  2207 => x"29610000",
     2208 => x"5c620004",  2209 => x"28230034",  2210 => x"b9800800",
     2211 => x"e0000004",  2212 => x"28230034",  2213 => x"34020000",
     2214 => x"b9800800",  2215 => x"d8600000",  2216 => x"34010000",
     2217 => x"2b9d0004",  2218 => x"2b8b000c",  2219 => x"2b8c0008",
     2220 => x"379c000c",  2221 => x"c3a00000",  2222 => x"379cfff0",
     2223 => x"5b8b0010",  2224 => x"5b8c000c",  2225 => x"5b8d0008",
     2226 => x"5b9d0004",  2227 => x"78040001",  2228 => x"78050001",
     2229 => x"2c2d0002",  2230 => x"b8205800",  2231 => x"b8406000",
     2232 => x"34010000",  2233 => x"34020002",  2234 => x"34030002",
     2235 => x"38843cd4",  2236 => x"38a558bc",  2237 => x"fbfff995",
     2238 => x"34010040",  2239 => x"4c2d0004",  2240 => x"b9600800",
     2241 => x"b9801000",  2242 => x"f8000466",  2243 => x"2b9d0004",
     2244 => x"2b8b0010",  2245 => x"2b8c000c",  2246 => x"2b8d0008",
     2247 => x"379c0010",  2248 => x"c3a00000",  2249 => x"379cfff8",
     2250 => x"5b8b0008",  2251 => x"5b9d0004",  2252 => x"78040001",
     2253 => x"78050001",  2254 => x"34020002",  2255 => x"34030002",
     2256 => x"38843cd4",  2257 => x"38a558d0",  2258 => x"b8205800",
     2259 => x"fbfff97f",  2260 => x"296102c8",  2261 => x"34020040",
     2262 => x"28210010",  2263 => x"40210004",  2264 => x"44200006",
     2265 => x"34030002",  2266 => x"44230004",  2267 => x"b9600800",
     2268 => x"f8000409",  2269 => x"3402004e",  2270 => x"b8400800",
     2271 => x"2b9d0004",  2272 => x"2b8b0008",  2273 => x"379c0008",
     2274 => x"c3a00000",  2275 => x"379cfff4",  2276 => x"5b8b000c",
     2277 => x"5b8c0008",  2278 => x"5b9d0004",  2279 => x"78040001",
     2280 => x"78050001",  2281 => x"34030002",  2282 => x"b8406000",
     2283 => x"38843cd4",  2284 => x"34020002",  2285 => x"38a558e4",
     2286 => x"b8205800",  2287 => x"fbfff963",  2288 => x"296102c8",
     2289 => x"34030000",  2290 => x"28210010",  2291 => x"28210008",
     2292 => x"44200007",  2293 => x"35630094",  2294 => x"59800008",
     2295 => x"b9600800",  2296 => x"b9801000",  2297 => x"f80005e9",
     2298 => x"34030001",  2299 => x"b8600800",  2300 => x"2b9d0004",
     2301 => x"2b8b000c",  2302 => x"2b8c0008",  2303 => x"379c000c",
     2304 => x"c3a00000",  2305 => x"379cfff8",  2306 => x"5b8b0008",
     2307 => x"5b9d0004",  2308 => x"78040001",  2309 => x"78050001",
     2310 => x"34020002",  2311 => x"34030002",  2312 => x"38843cd4",
     2313 => x"38a558f8",  2314 => x"b8205800",  2315 => x"fbfff947",
     2316 => x"296102c8",  2317 => x"28220010",  2318 => x"40410004",
     2319 => x"20210002",  2320 => x"4420000b",  2321 => x"40410035",
     2322 => x"20210001",  2323 => x"44200008",  2324 => x"28410008",
     2325 => x"44200003",  2326 => x"28410040",  2327 => x"5c200004",
     2328 => x"b9600800",  2329 => x"34020009",  2330 => x"f80000a1",
     2331 => x"2b9d0004",  2332 => x"2b8b0008",  2333 => x"379c0008",
     2334 => x"c3a00000",  2335 => x"379cffdc",  2336 => x"5b8b0010",
     2337 => x"5b8c000c",  2338 => x"5b8d0008",  2339 => x"5b9d0004",
     2340 => x"28220020",  2341 => x"78040001",  2342 => x"78050001",
     2343 => x"284d0010",  2344 => x"282202c8",  2345 => x"34030002",
     2346 => x"38843cd4",  2347 => x"284c0010",  2348 => x"38a55928",
     2349 => x"34020002",  2350 => x"b8205800",  2351 => x"fbfff923",
     2352 => x"29620318",  2353 => x"2963031c",  2354 => x"37810014",
     2355 => x"f80010df",  2356 => x"29810008",  2357 => x"5c200019",
     2358 => x"296200a0",  2359 => x"44410003",  2360 => x"296100b4",
     2361 => x"5c200008",  2362 => x"78040001",  2363 => x"b9600800",
     2364 => x"34020004",  2365 => x"34030001",  2366 => x"38843ce0",
     2367 => x"fbfff913",  2368 => x"e0000013",  2369 => x"b9600800",
     2370 => x"f80011d1",  2371 => x"29a20004",  2372 => x"29810000",
     2373 => x"44400005",  2374 => x"28230034",  2375 => x"34020000",
     2376 => x"b9600800",  2377 => x"e0000004",  2378 => x"28230034",
     2379 => x"34020001",  2380 => x"b9600800",  2381 => x"d8600000",
     2382 => x"29620318",  2383 => x"b9600800",  2384 => x"f80005ac",
     2385 => x"b9600800",  2386 => x"f80005d4",  2387 => x"34010000",
     2388 => x"2b9d0004",  2389 => x"2b8b0010",  2390 => x"2b8c000c",
     2391 => x"2b8d0008",  2392 => x"379c0024",  2393 => x"c3a00000",
     2394 => x"379cfff8",  2395 => x"5b8b0008",  2396 => x"5b9d0004",
     2397 => x"78040001",  2398 => x"78050001",  2399 => x"34020002",
     2400 => x"34030002",  2401 => x"38843cd4",  2402 => x"38a55938",
     2403 => x"b8205800",  2404 => x"fbfff8ee",  2405 => x"b9600800",
     2406 => x"f8000523",  2407 => x"34010000",  2408 => x"2b9d0004",
     2409 => x"2b8b0008",  2410 => x"379c0008",  2411 => x"c3a00000",
     2412 => x"379cffd8",  2413 => x"5b8b0010",  2414 => x"5b8c000c",
     2415 => x"5b8d0008",  2416 => x"5b9d0004",  2417 => x"78050001",
     2418 => x"b8806000",  2419 => x"78040001",  2420 => x"b8406800",
     2421 => x"34030002",  2422 => x"34020002",  2423 => x"38843cd4",
     2424 => x"38a55948",  2425 => x"b8205800",  2426 => x"fbfff8d8",
     2427 => x"34010001",  2428 => x"45810004",  2429 => x"3401000c",
     2430 => x"5d810036",  2431 => x"e0000022",  2432 => x"296200ec",
     2433 => x"5960031c",  2434 => x"37810024",  2435 => x"4802000c",
     2436 => x"1443001f",  2437 => x"00440010",  2438 => x"3c630010",
     2439 => x"3c420010",  2440 => x"b8641800",  2441 => x"5b820028",
     2442 => x"340203e8",  2443 => x"5b830024",  2444 => x"fbfffcee",
     2445 => x"2b810028",  2446 => x"e000000d",  2447 => x"c8021000",
     2448 => x"1443001f",  2449 => x"00440010",  2450 => x"3c630010",
     2451 => x"3c420010",  2452 => x"b8641800",  2453 => x"5b820028",
     2454 => x"340203e8",  2455 => x"5b830024",  2456 => x"fbfffce2",
     2457 => x"2b810028",  2458 => x"c8010800",  2459 => x"59610318",
     2460 => x"356200e4",  2461 => x"b9600800",  2462 => x"f8001013",
     2463 => x"340c0100",  2464 => x"e0000014",  2465 => x"296102c8",
     2466 => x"b9a01000",  2467 => x"37830014",  2468 => x"28240010",
     2469 => x"b9600800",  2470 => x"340c0100",  2471 => x"3484003c",
     2472 => x"f8000416",  2473 => x"296102c8",  2474 => x"34021000",
     2475 => x"28210010",  2476 => x"2c23003c",  2477 => x"5c620007",
     2478 => x"40210004",  2479 => x"20210001",  2480 => x"44200004",
     2481 => x"b9600800",  2482 => x"34020006",  2483 => x"f8000008",
     2484 => x"b9800800",  2485 => x"2b9d0004",  2486 => x"2b8b0010",
     2487 => x"2b8c000c",  2488 => x"2b8d0008",  2489 => x"379c0028",
     2490 => x"c3a00000",  2491 => x"282302c8",  2492 => x"34040006",
     2493 => x"28630010",  2494 => x"44440004",  2495 => x"34040009",
     2496 => x"5c440008",  2497 => x"e0000004",  2498 => x"34020001",
     2499 => x"30620005",  2500 => x"e0000007",  2501 => x"34020002",
     2502 => x"30620005",  2503 => x"e0000006",  2504 => x"40630005",
     2505 => x"34020001",  2506 => x"5c620003",  2507 => x"34020066",
     2508 => x"e0000002",  2509 => x"34020064",  2510 => x"58220004",
     2511 => x"c3a00000",  2512 => x"379cfff4",  2513 => x"5b8b000c",
     2514 => x"5b8c0008",  2515 => x"5b9d0004",  2516 => x"b8205800",
     2517 => x"282102c8",  2518 => x"78050001",  2519 => x"38a53c30",
     2520 => x"282c0010",  2521 => x"34010001",  2522 => x"41820005",
     2523 => x"5c410003",  2524 => x"78050001",  2525 => x"38a54118",
     2526 => x"78040001",  2527 => x"b9600800",  2528 => x"34020002",
     2529 => x"34030001",  2530 => x"38843d08",  2531 => x"fbfff86f",
     2532 => x"41820005",  2533 => x"34010001",  2534 => x"5c410003",
     2535 => x"34010006",  2536 => x"e0000002",  2537 => x"34010009",
     2538 => x"59610004",  2539 => x"31800005",  2540 => x"2b9d0004",
     2541 => x"2b8b000c",  2542 => x"2b8c0008",  2543 => x"379c000c",
     2544 => x"c3a00000",  2545 => x"379cfffc",  2546 => x"5b9d0004",
     2547 => x"282202c8",  2548 => x"28420010",  2549 => x"4043002c",
     2550 => x"4460000a",  2551 => x"3463ffff",  2552 => x"78040001",
     2553 => x"3043002c",  2554 => x"38843d2c",  2555 => x"34020002",
     2556 => x"34030001",  2557 => x"fbfff855",  2558 => x"34010001",
     2559 => x"e0000003",  2560 => x"fbffffd0",  2561 => x"34010000",
     2562 => x"2b9d0004",  2563 => x"379c0004",  2564 => x"c3a00000",
     2565 => x"379cffd8",  2566 => x"5b8b0018",  2567 => x"5b8c0014",
     2568 => x"5b8d0010",  2569 => x"5b8e000c",  2570 => x"5b8f0008",
     2571 => x"5b9d0004",  2572 => x"b8407000",  2573 => x"2824000c",
     2574 => x"282202c8",  2575 => x"b8205800",  2576 => x"b8607800",
     2577 => x"284d0010",  2578 => x"44800004",  2579 => x"34010003",
     2580 => x"31a1002c",  2581 => x"e000000c",  2582 => x"282202e0",
     2583 => x"44440008",  2584 => x"28220028",  2585 => x"28440018",
     2586 => x"34020000",  2587 => x"d8800000",  2588 => x"296202e0",
     2589 => x"c8220800",  2590 => x"4c20003c",  2591 => x"340c0000",
     2592 => x"e0000015",  2593 => x"29610028",  2594 => x"340203e8",
     2595 => x"28240018",  2596 => x"b9600800",  2597 => x"d8800000",
     2598 => x"596102e0",  2599 => x"296102c8",  2600 => x"29620028",
     2601 => x"4025000c",  2602 => x"1021000b",  2603 => x"28440018",
     2604 => x"bca12800",  2605 => x"b9600800",  2606 => x"08a203e8",
     2607 => x"d8800000",  2608 => x"596102d4",  2609 => x"34021000",
     2610 => x"b9600800",  2611 => x"f80003fb",  2612 => x"b8206000",
     2613 => x"45e0000e",  2614 => x"4162030d",  2615 => x"3401000c",
     2616 => x"5c41000b",  2617 => x"b9600800",  2618 => x"b9c01000",
     2619 => x"3783001c",  2620 => x"35a4003c",  2621 => x"f8000381",
     2622 => x"2da2003c",  2623 => x"34011001",  2624 => x"5c410003",
     2625 => x"34010065",  2626 => x"59610004",  2627 => x"5d800004",
     2628 => x"b9600800",  2629 => x"f8000adb",  2630 => x"e0000003",
     2631 => x"34010002",  2632 => x"59610004",  2633 => x"29620004",
     2634 => x"29610000",  2635 => x"44410002",  2636 => x"596002d4",
     2637 => x"296102c8",  2638 => x"28210010",  2639 => x"28210028",
     2640 => x"59610008",  2641 => x"b9800800",  2642 => x"2b9d0004",
     2643 => x"2b8b0018",  2644 => x"2b8c0014",  2645 => x"2b8d0010",
     2646 => x"2b8e000c",  2647 => x"2b8f0008",  2648 => x"379c0028",
     2649 => x"c3a00000",  2650 => x"b9600800",  2651 => x"34020005",
     2652 => x"f800127b",  2653 => x"b9600800",  2654 => x"596002e0",
     2655 => x"fbffff92",  2656 => x"340c0000",  2657 => x"5c20ffc0",
     2658 => x"e3ffffef",  2659 => x"379cffd8",  2660 => x"5b8b0018",
     2661 => x"5b8c0014",  2662 => x"5b8d0010",  2663 => x"5b8e000c",
     2664 => x"5b8f0008",  2665 => x"5b9d0004",  2666 => x"b8407000",
     2667 => x"2824000c",  2668 => x"282202c8",  2669 => x"b8205800",
     2670 => x"b8607800",  2671 => x"284c0010",  2672 => x"44800004",
     2673 => x"34010003",  2674 => x"3181002c",  2675 => x"e000000c",
     2676 => x"282202e0",  2677 => x"44440008",  2678 => x"28220028",
     2679 => x"28440018",  2680 => x"34020000",  2681 => x"d8800000",
     2682 => x"296202e0",  2683 => x"c8220800",  2684 => x"4c200029",
     2685 => x"340d0000",  2686 => x"e000000b",  2687 => x"34021001",
     2688 => x"b9600800",  2689 => x"f80003ad",  2690 => x"b8206800",
     2691 => x"29610028",  2692 => x"34023a98",  2693 => x"28240018",
     2694 => x"b9600800",  2695 => x"d8800000",  2696 => x"596102e0",
     2697 => x"45e0000e",  2698 => x"4162030d",  2699 => x"3401000c",
     2700 => x"5c41000b",  2701 => x"b9600800",  2702 => x"b9c01000",
     2703 => x"3783001c",  2704 => x"3584003c",  2705 => x"f800032d",
     2706 => x"2d82003c",  2707 => x"34011002",  2708 => x"5c410003",
     2709 => x"34010068",  2710 => x"59610004",  2711 => x"45a00003",
     2712 => x"34010002",  2713 => x"59610004",  2714 => x"29810028",
     2715 => x"59610008",  2716 => x"b9a00800",  2717 => x"2b9d0004",
     2718 => x"2b8b0018",  2719 => x"2b8c0014",  2720 => x"2b8d0010",
     2721 => x"2b8e000c",  2722 => x"2b8f0008",  2723 => x"379c0028",
     2724 => x"c3a00000",  2725 => x"b9600800",  2726 => x"34020005",
     2727 => x"f8001230",  2728 => x"b9600800",  2729 => x"596002e0",
     2730 => x"fbffff47",  2731 => x"340d0000",  2732 => x"5c20ffd3",
     2733 => x"e3ffffef",  2734 => x"379cfff4",  2735 => x"5b8b000c",
     2736 => x"5b8c0008",  2737 => x"5b9d0004",  2738 => x"282202c8",
     2739 => x"b8205800",  2740 => x"284c0010",  2741 => x"2822000c",
     2742 => x"44400004",  2743 => x"34010003",  2744 => x"3181002c",
     2745 => x"e000000b",  2746 => x"282302e0",  2747 => x"44620013",
     2748 => x"28220028",  2749 => x"28430018",  2750 => x"34020000",
     2751 => x"d8600000",  2752 => x"296202e0",  2753 => x"c8220800",
     2754 => x"4c200021",  2755 => x"e000000b",  2756 => x"29810000",
     2757 => x"28220000",  2758 => x"b9600800",  2759 => x"d8400000",
     2760 => x"29610028",  2761 => x"34023a98",  2762 => x"28230018",
     2763 => x"b9600800",  2764 => x"d8600000",  2765 => x"596102e0",
     2766 => x"29810000",  2767 => x"34020000",  2768 => x"28230004",
     2769 => x"b9600800",  2770 => x"d8600000",  2771 => x"34020001",
     2772 => x"5c220007",  2773 => x"34010067",  2774 => x"59610004",
     2775 => x"29810000",  2776 => x"28220008",  2777 => x"b9600800",
     2778 => x"d8400000",  2779 => x"29810028",  2780 => x"59610008",
     2781 => x"34010000",  2782 => x"2b9d0004",  2783 => x"2b8b000c",
     2784 => x"2b8c0008",  2785 => x"379c000c",  2786 => x"c3a00000",
     2787 => x"b9600800",  2788 => x"34020005",  2789 => x"f80011f2",
     2790 => x"29810000",  2791 => x"596002e0",  2792 => x"28220008",
     2793 => x"b9600800",  2794 => x"d8400000",  2795 => x"b9600800",
     2796 => x"fbffff05",  2797 => x"5c20ffd7",  2798 => x"e3ffffef",
     2799 => x"379cffd8",  2800 => x"5b8b0018",  2801 => x"5b8c0014",
     2802 => x"5b8d0010",  2803 => x"5b8e000c",  2804 => x"5b8f0008",
     2805 => x"5b9d0004",  2806 => x"b8407000",  2807 => x"2824000c",
     2808 => x"282202c8",  2809 => x"b8205800",  2810 => x"b8607800",
     2811 => x"284c0010",  2812 => x"44800004",  2813 => x"34010003",
     2814 => x"3181002c",  2815 => x"e000000c",  2816 => x"282202e0",
     2817 => x"44440008",  2818 => x"28220028",  2819 => x"28440018",
     2820 => x"34020000",  2821 => x"d8800000",  2822 => x"296202e0",
     2823 => x"c8220800",  2824 => x"4c200029",  2825 => x"340d0000",
     2826 => x"e000000b",  2827 => x"29610028",  2828 => x"29820028",
     2829 => x"28240018",  2830 => x"b9600800",  2831 => x"d8800000",
     2832 => x"596102e0",  2833 => x"34021002",  2834 => x"b9600800",
     2835 => x"f800031b",  2836 => x"b8206800",  2837 => x"45e0000e",
     2838 => x"4162030d",  2839 => x"3401000c",  2840 => x"5c41000b",
     2841 => x"b9600800",  2842 => x"b9c01000",  2843 => x"3783001c",
     2844 => x"3584003c",  2845 => x"f80002a1",  2846 => x"2d82003c",
     2847 => x"34011003",  2848 => x"5c410003",  2849 => x"3401006a",
     2850 => x"59610004",  2851 => x"45a00003",  2852 => x"34010002",
     2853 => x"59610004",  2854 => x"29810028",  2855 => x"59610008",
     2856 => x"b9a00800",  2857 => x"2b9d0004",  2858 => x"2b8b0018",
     2859 => x"2b8c0014",  2860 => x"2b8d0010",  2861 => x"2b8e000c",
     2862 => x"2b8f0008",  2863 => x"379c0028",  2864 => x"c3a00000",
     2865 => x"b9600800",  2866 => x"34020005",  2867 => x"f80011a4",
     2868 => x"b9600800",  2869 => x"596002e0",  2870 => x"fbfffebb",
     2871 => x"340d0000",  2872 => x"5c20ffd3",  2873 => x"e3ffffef",
     2874 => x"379cffec",  2875 => x"5b8b0010",  2876 => x"5b8c000c",
     2877 => x"5b8d0008",  2878 => x"5b9d0004",  2879 => x"282202c8",
     2880 => x"b8206000",  2881 => x"284b0010",  2882 => x"2822000c",
     2883 => x"44400004",  2884 => x"34010003",  2885 => x"3161002c",
     2886 => x"e000000c",  2887 => x"282302e0",  2888 => x"44620008",
     2889 => x"28220028",  2890 => x"28430018",  2891 => x"34020000",
     2892 => x"d8600000",  2893 => x"298202e0",  2894 => x"c8220800",
     2895 => x"4c2000a9",  2896 => x"340d0000",  2897 => x"e0000011",
     2898 => x"29810028",  2899 => x"29620030",  2900 => x"28230018",
     2901 => x"b9800800",  2902 => x"d8600000",  2903 => x"598102e0",
     2904 => x"34021003",  2905 => x"b9800800",  2906 => x"f80002d4",
     2907 => x"b8206800",  2908 => x"3401006c",  2909 => x"31610010",
     2910 => x"29610014",  2911 => x"44200003",  2912 => x"3401006e",
     2913 => x"31610010",  2914 => x"41660010",  2915 => x"78040001",
     2916 => x"78050001",  2917 => x"b9800800",  2918 => x"34020002",
     2919 => x"34030001",  2920 => x"38843d40",  2921 => x"38a5599c",
     2922 => x"34c6ff94",  2923 => x"fbfff6e7",  2924 => x"41620010",
     2925 => x"34010008",  2926 => x"3442ff94",  2927 => x"204200ff",
     2928 => x"5441007f",  2929 => x"78010001",  2930 => x"3c420002",
     2931 => x"38215978",  2932 => x"b4220800",  2933 => x"28210000",
     2934 => x"c0200000",  2935 => x"29610000",  2936 => x"34020000",
     2937 => x"34030000",  2938 => x"2825002c",  2939 => x"34040000",
     2940 => x"b9800800",  2941 => x"d8a00000",  2942 => x"5c200071",
     2943 => x"3401006d",  2944 => x"31610010",  2945 => x"29610000",
     2946 => x"34020001",  2947 => x"28230024",  2948 => x"b9800800",
     2949 => x"d8600000",  2950 => x"5c200069",  2951 => x"3401006e",
     2952 => x"31610010",  2953 => x"29610000",  2954 => x"34020001",
     2955 => x"37830014",  2956 => x"28240028",  2957 => x"b9800800",
     2958 => x"d8800000",  2959 => x"34020001",  2960 => x"5c22005f",
     2961 => x"2b810014",  2962 => x"78040001",  2963 => x"34020002",
     2964 => x"00250010",  2965 => x"3c210010",  2966 => x"5965001c",
     2967 => x"59610018",  2968 => x"34030001",  2969 => x"b9800800",
     2970 => x"38843d54",  2971 => x"fbfff6b7",  2972 => x"29650018",
     2973 => x"78040001",  2974 => x"b9800800",  2975 => x"34020002",
     2976 => x"34030001",  2977 => x"38843d78",  2978 => x"fbfff6b0",
     2979 => x"3401006f",  2980 => x"31610010",  2981 => x"29610000",
     2982 => x"34020001",  2983 => x"28230020",  2984 => x"b9800800",
     2985 => x"d8600000",  2986 => x"5c200045",  2987 => x"34010070",
     2988 => x"31610010",  2989 => x"29610000",  2990 => x"28220030",
     2991 => x"b9800800",  2992 => x"d8400000",  2993 => x"5c20003e",
     2994 => x"34010071",  2995 => x"31610010",  2996 => x"29610000",
     2997 => x"34020002",  2998 => x"28230024",  2999 => x"b9800800",
     3000 => x"d8600000",  3001 => x"5c200036",  3002 => x"34010072",
     3003 => x"31610010",  3004 => x"29610000",  3005 => x"34020002",
     3006 => x"37830014",  3007 => x"28240028",  3008 => x"b9800800",
     3009 => x"d8800000",  3010 => x"34020001",  3011 => x"5c22002c",
     3012 => x"2b850014",  3013 => x"78040001",  3014 => x"b9800800",
     3015 => x"34020002",  3016 => x"34030001",  3017 => x"38843d9c",
     3018 => x"fbfff688",  3019 => x"2b810014",  3020 => x"78040001",
     3021 => x"34020002",  3022 => x"00250010",  3023 => x"3c210010",
     3024 => x"59650024",  3025 => x"59610020",  3026 => x"34030001",
     3027 => x"b9800800",  3028 => x"38843db4",  3029 => x"fbfff67d",
     3030 => x"29650020",  3031 => x"78040001",  3032 => x"b9800800",
     3033 => x"34020002",  3034 => x"34030001",  3035 => x"38843dd8",
     3036 => x"fbfff676",  3037 => x"34010073",  3038 => x"31610010",
     3039 => x"29610000",  3040 => x"34020002",  3041 => x"28230020",
     3042 => x"b9800800",  3043 => x"d8600000",  3044 => x"5c20000b",
     3045 => x"34010074",  3046 => x"31610010",  3047 => x"b9800800",
     3048 => x"34021004",  3049 => x"f8000245",  3050 => x"b8206800",
     3051 => x"34010069",  3052 => x"59810004",  3053 => x"34010001",
     3054 => x"59610014",  3055 => x"29610028",  3056 => x"59810008",
     3057 => x"b9a00800",  3058 => x"2b9d0004",  3059 => x"2b8b0010",
     3060 => x"2b8c000c",  3061 => x"2b8d0008",  3062 => x"379c0014",
     3063 => x"c3a00000",  3064 => x"b9800800",  3065 => x"34020005",
     3066 => x"f80010dd",  3067 => x"b9800800",  3068 => x"598002e0",
     3069 => x"fbfffdf4",  3070 => x"340d0000",  3071 => x"5c20ff53",
     3072 => x"e3fffff1",  3073 => x"379cffdc",  3074 => x"5b8b0014",
     3075 => x"5b8c0010",  3076 => x"5b8d000c",  3077 => x"5b8e0008",
     3078 => x"5b9d0004",  3079 => x"b8406800",  3080 => x"282202c8",
     3081 => x"b8205800",  3082 => x"b8607000",  3083 => x"284c0010",
     3084 => x"2822000c",  3085 => x"44400006",  3086 => x"28220028",
     3087 => x"28440018",  3088 => x"29820028",  3089 => x"d8800000",
     3090 => x"596102e0",  3091 => x"296102e0",  3092 => x"44200009",
     3093 => x"29610028",  3094 => x"34020000",  3095 => x"28240018",
     3096 => x"b9600800",  3097 => x"d8800000",  3098 => x"296202e0",
     3099 => x"c8220800",  3100 => x"4c200023",  3101 => x"45c00018",
     3102 => x"4162030d",  3103 => x"3401000c",  3104 => x"5c410015",
     3105 => x"b9600800",  3106 => x"b9a01000",  3107 => x"37830018",
     3108 => x"3584003c",  3109 => x"f8000199",  3110 => x"2d81003c",
     3111 => x"34021003",  3112 => x"5c220006",  3113 => x"41820005",
     3114 => x"34010001",  3115 => x"5c41000a",  3116 => x"3401006a",
     3117 => x"e0000007",  3118 => x"34021005",  3119 => x"5c220006",
     3120 => x"41820005",  3121 => x"34010002",  3122 => x"5c410003",
     3123 => x"3401006b",  3124 => x"59610004",  3125 => x"29810028",
     3126 => x"59610008",  3127 => x"34010000",  3128 => x"2b9d0004",
     3129 => x"2b8b0014",  3130 => x"2b8c0010",  3131 => x"2b8d000c",
     3132 => x"2b8e0008",  3133 => x"379c0024",  3134 => x"c3a00000",
     3135 => x"b9600800",  3136 => x"34020005",  3137 => x"f8001096",
     3138 => x"b9600800",  3139 => x"596002e0",  3140 => x"fbfffd8c",
     3141 => x"e3fffff2",  3142 => x"379cffd4",  3143 => x"5b8b001c",
     3144 => x"5b8c0018",  3145 => x"5b8d0014",  3146 => x"5b8e0010",
     3147 => x"5b8f000c",  3148 => x"5b900008",  3149 => x"5b9d0004",
     3150 => x"b8407000",  3151 => x"282202c8",  3152 => x"2824000c",
     3153 => x"b8205800",  3154 => x"284c0010",  3155 => x"b8607800",
     3156 => x"2d8d0048",  3157 => x"7dad0000",  3158 => x"44800004",
     3159 => x"34010003",  3160 => x"3181002c",  3161 => x"e0000012",
     3162 => x"282202e0",  3163 => x"44440022",  3164 => x"28220028",
     3165 => x"28440018",  3166 => x"34020000",  3167 => x"d8800000",
     3168 => x"296202e0",  3169 => x"c8220800",  3170 => x"4c20003f",
     3171 => x"e000001a",  3172 => x"29810000",  3173 => x"28240030",
     3174 => x"b9600800",  3175 => x"d8800000",  3176 => x"b9600800",
     3177 => x"fbfffd88",  3178 => x"4420002d",  3179 => x"45a00008",
     3180 => x"29810000",  3181 => x"34020000",  3182 => x"34030000",
     3183 => x"2825002c",  3184 => x"34040000",  3185 => x"b9600800",
     3186 => x"d8a00000",  3187 => x"2981004c",  3188 => x"29700028",
     3189 => x"340203e8",  3190 => x"f8003e5b",  3191 => x"2a050018",
     3192 => x"b8202000",  3193 => x"b8801000",  3194 => x"b9600800",
     3195 => x"d8a00000",  3196 => x"596102e0",  3197 => x"45e00018",
     3198 => x"4162030d",  3199 => x"3401000c",  3200 => x"5c410015",
     3201 => x"b9600800",  3202 => x"b9c01000",  3203 => x"37830020",
     3204 => x"3584003c",  3205 => x"f8000139",  3206 => x"2d82003c",
     3207 => x"34011004",  3208 => x"5c41000d",  3209 => x"45a00005",
     3210 => x"29810000",  3211 => x"28220030",  3212 => x"b9600800",
     3213 => x"d8400000",  3214 => x"41820005",  3215 => x"34010001",
     3216 => x"5c410003",  3217 => x"3401006b",  3218 => x"e0000002",
     3219 => x"34010068",  3220 => x"59610004",  3221 => x"29810028",
     3222 => x"59610008",  3223 => x"34010000",  3224 => x"2b9d0004",
     3225 => x"2b8b001c",  3226 => x"2b8c0018",  3227 => x"2b8d0014",
     3228 => x"2b8e0010",  3229 => x"2b8f000c",  3230 => x"2b900008",
     3231 => x"379c002c",  3232 => x"c3a00000",  3233 => x"b9600800",
     3234 => x"34020005",  3235 => x"f8001034",  3236 => x"596002e0",
     3237 => x"45a0ffc3",  3238 => x"e3ffffbe",  3239 => x"379cfff0",
     3240 => x"5b8b0010",  3241 => x"5b8c000c",  3242 => x"5b8d0008",
     3243 => x"5b9d0004",  3244 => x"282202c8",  3245 => x"340d0001",
     3246 => x"b8206000",  3247 => x"284b0010",  3248 => x"29620000",
     3249 => x"596d0008",  3250 => x"2842000c",  3251 => x"d8400000",
     3252 => x"41610005",  3253 => x"34020000",  3254 => x"5c2d0005",
     3255 => x"34021005",  3256 => x"b9800800",  3257 => x"f8000175",
     3258 => x"b8201000",  3259 => x"34010001",  3260 => x"59610040",
     3261 => x"3401ffff",  3262 => x"5c400009",  3263 => x"41620005",
     3264 => x"34010002",  3265 => x"5c410003",  3266 => x"34010009",
     3267 => x"e0000002",  3268 => x"34010006",  3269 => x"59810004",
     3270 => x"34010000",  3271 => x"2b9d0004",  3272 => x"2b8b0010",
     3273 => x"2b8c000c",  3274 => x"2b8d0008",  3275 => x"379c0010",
     3276 => x"c3a00000",  3277 => x"00430018",  3278 => x"30220003",
     3279 => x"30230000",  3280 => x"00430010",  3281 => x"30230001",
     3282 => x"00430008",  3283 => x"30230002",  3284 => x"c3a00000",
     3285 => x"40220000",  3286 => x"40230003",  3287 => x"3c420018",
     3288 => x"b8621000",  3289 => x"40230001",  3290 => x"40210002",
     3291 => x"3c630010",  3292 => x"3c210008",  3293 => x"b8431000",
     3294 => x"b8410800",  3295 => x"c3a00000",  3296 => x"40220000",
     3297 => x"40210001",  3298 => x"3c420008",  3299 => x"b8410800",
     3300 => x"c3a00000",  3301 => x"379cfff0",  3302 => x"5b8b0010",
     3303 => x"5b8c000c",  3304 => x"5b8d0008",  3305 => x"5b9d0004",
     3306 => x"28230020",  3307 => x"282202c8",  3308 => x"b8205800",
     3309 => x"2863000c",  3310 => x"28420010",  3311 => x"282c003c",
     3312 => x"4064000e",  3313 => x"340300ba",  3314 => x"48830018",
     3315 => x"28420000",  3316 => x"28430004",  3317 => x"34020001",
     3318 => x"d8600000",  3319 => x"ec016800",  3320 => x"b9600800",
     3321 => x"f8000994",  3322 => x"29610020",  3323 => x"c80d6800",
     3324 => x"21ad002e",  3325 => x"2821000c",  3326 => x"35ad0006",
     3327 => x"4021000e",  3328 => x"45a1000a",  3329 => x"78010001",
     3330 => x"b9a01000",  3331 => x"38213dfc",  3332 => x"f800247b",
     3333 => x"29610020",  3334 => x"21ad00ff",  3335 => x"2821000c",
     3336 => x"302d000e",  3337 => x"318d0030",  3338 => x"3401004e",
     3339 => x"0d810002",  3340 => x"34010003",  3341 => x"0d810040",
     3342 => x"3401000a",  3343 => x"0d810042",  3344 => x"34010800",
     3345 => x"0d810044",  3346 => x"340130de",  3347 => x"0d810046",
     3348 => x"3401ad01",  3349 => x"0d810048",  3350 => x"34012000",
     3351 => x"0d81004a",  3352 => x"296102c8",  3353 => x"28220010",
     3354 => x"28430014",  3355 => x"40410004",  3356 => x"44600002",
     3357 => x"38210004",  3358 => x"28420008",  3359 => x"44400002",
     3360 => x"38210008",  3361 => x"0d81004c",  3362 => x"2b9d0004",
     3363 => x"2b8b0010",  3364 => x"2b8c000c",  3365 => x"2b8d0008",
     3366 => x"379c0010",  3367 => x"c3a00000",  3368 => x"379cfff4",
     3369 => x"5b8b000c",  3370 => x"5b8c0008",  3371 => x"5b9d0004",
     3372 => x"b8205800",  3373 => x"34210040",  3374 => x"b8406000",
     3375 => x"fbffffb1",  3376 => x"2d650044",  3377 => x"2d640046",
     3378 => x"78070001",  3379 => x"3ca50008",  3380 => x"00860008",
     3381 => x"38e75750",  3382 => x"b8a62800",  3383 => x"28e60000",
     3384 => x"64210003",  3385 => x"2d630048",  3386 => x"e4a62800",
     3387 => x"2d62004a",  3388 => x"a0250800",  3389 => x"44200010",
     3390 => x"3c840008",  3391 => x"00610008",  3392 => x"2084ffff",
     3393 => x"b8812000",  3394 => x"206300ff",  3395 => x"3801dead",
     3396 => x"e4812000",  3397 => x"64630001",  3398 => x"a0831800",
     3399 => x"44600006",  3400 => x"34012000",  3401 => x"5c410004",
     3402 => x"3561004c",  3403 => x"fbffff95",  3404 => x"59810024",
     3405 => x"2b9d0004",  3406 => x"2b8b000c",  3407 => x"2b8c0008",
     3408 => x"379c000c",  3409 => x"c3a00000",  3410 => x"379cfff0",
     3411 => x"5b8b0010",  3412 => x"5b8c000c",  3413 => x"5b8d0008",
     3414 => x"5b9d0004",  3415 => x"b8206000",  3416 => x"282102c8",
     3417 => x"204dffff",  3418 => x"28210010",  3419 => x"40250005",
     3420 => x"44a00003",  3421 => x"34012000",  3422 => x"5da1000a",
     3423 => x"78040001",  3424 => x"b9800800",  3425 => x"34020005",
     3426 => x"34030001",  3427 => x"38843e14",  3428 => x"b9a03000",
     3429 => x"fbfff4ed",  3430 => x"34010000",  3431 => x"e0000051",
     3432 => x"298b003c",  3433 => x"34030008",  3434 => x"41610000",
     3435 => x"202100f0",  3436 => x"3821000c",  3437 => x"31610000",
     3438 => x"34010005",  3439 => x"31610020",  3440 => x"29820020",
     3441 => x"35610022",  3442 => x"28420014",  3443 => x"f8003dbf",
     3444 => x"29810020",  3445 => x"28210014",  3446 => x"2c210008",
     3447 => x"0d6d0036",  3448 => x"00220008",  3449 => x"3161002b",
     3450 => x"34010003",  3451 => x"0d61002c",  3452 => x"34010800",
     3453 => x"0d610030",  3454 => x"340130de",  3455 => x"0d610032",
     3456 => x"3401ad01",  3457 => x"0d610034",  3458 => x"3162002a",
     3459 => x"34011003",  3460 => x"45a10005",  3461 => x"34011004",
     3462 => x"34020008",  3463 => x"5da1002d",  3464 => x"e0000017",
     3465 => x"298102c8",  3466 => x"35620038",  3467 => x"28210010",
     3468 => x"28230014",  3469 => x"44600005",  3470 => x"40210034",
     3471 => x"31610038",  3472 => x"30400001",  3473 => x"e0000007",
     3474 => x"40210034",  3475 => x"3c210008",  3476 => x"38210001",
     3477 => x"00230008",  3478 => x"31630038",  3479 => x"30410001",
     3480 => x"298102c8",  3481 => x"28220010",  3482 => x"3561003a",
     3483 => x"28420030",  3484 => x"fbffff31",  3485 => x"34020014",
     3486 => x"e0000016",  3487 => x"298102c8",  3488 => x"28220010",
     3489 => x"35610038",  3490 => x"2842001c",  3491 => x"fbffff2a",
     3492 => x"298102c8",  3493 => x"28220010",  3494 => x"3561003c",
     3495 => x"28420018",  3496 => x"fbffff25",  3497 => x"298102c8",
     3498 => x"28220010",  3499 => x"35610040",  3500 => x"28420024",
     3501 => x"fbffff20",  3502 => x"298102c8",  3503 => x"28220010",
     3504 => x"35610044",  3505 => x"28420020",  3506 => x"fbffff1b",
     3507 => x"34020018",  3508 => x"34410030",  3509 => x"31600002",
     3510 => x"31610003",  3511 => x"0d62002e",  3512 => x"2b9d0004",
     3513 => x"2b8b0010",  3514 => x"2b8c000c",  3515 => x"2b8d0008",
     3516 => x"379c0010",  3517 => x"c3a00000",  3518 => x"379cffec",
     3519 => x"5b8b0014",  3520 => x"5b8c0010",  3521 => x"5b8d000c",
     3522 => x"5b8e0008",  3523 => x"5b9d0004",  3524 => x"b8405800",
     3525 => x"b8607000",  3526 => x"34420022",  3527 => x"b8206000",
     3528 => x"b8600800",  3529 => x"34030008",  3530 => x"b8806800",
     3531 => x"f8003d67",  3532 => x"3561002a",  3533 => x"fbffff13",
     3534 => x"0dc10008",  3535 => x"3561002c",  3536 => x"fbffff10",
     3537 => x"b8202800",  3538 => x"34040003",  3539 => x"2d630030",
     3540 => x"2d620032",  3541 => x"2d610034",  3542 => x"44a40007",
     3543 => x"78040001",  3544 => x"b9800800",  3545 => x"34020005",
     3546 => x"34030001",  3547 => x"38843e48",  3548 => x"e0000022",
     3549 => x"3c650008",  3550 => x"78040001",  3551 => x"00430008",
     3552 => x"38845750",  3553 => x"b8a32800",  3554 => x"28830000",
     3555 => x"44a30007",  3556 => x"78040001",  3557 => x"b9800800",
     3558 => x"34020005",  3559 => x"34030001",  3560 => x"38843e98",
     3561 => x"e0000015",  3562 => x"3c450008",  3563 => x"00230008",
     3564 => x"20a5ffff",  3565 => x"b8a32800",  3566 => x"3802dead",
     3567 => x"44a20007",  3568 => x"78040001",  3569 => x"b9800800",
     3570 => x"34020005",  3571 => x"34030001",  3572 => x"38843ed0",
     3573 => x"e0000009",  3574 => x"202500ff",  3575 => x"34010001",
     3576 => x"44a10008",  3577 => x"78040001",  3578 => x"b9800800",
     3579 => x"34020005",  3580 => x"34030001",  3581 => x"38843f14",
     3582 => x"fbfff454",  3583 => x"e0000028",  3584 => x"2d610036",
     3585 => x"45a00002",  3586 => x"0da10000",  3587 => x"34021003",
     3588 => x"44220004",  3589 => x"34021004",  3590 => x"5c220021",
     3591 => x"e0000012",  3592 => x"298102c8",  3593 => x"356e0038",
     3594 => x"282d0010",  3595 => x"b9c00800",  3596 => x"fbfffed4",
     3597 => x"202100ff",  3598 => x"0da10048",  3599 => x"b9c00800",
     3600 => x"fbfffed0",  3601 => x"00210008",  3602 => x"31a10050",
     3603 => x"3561003a",  3604 => x"fbfffec1",  3605 => x"298202c8",
     3606 => x"28420010",  3607 => x"5841004c",  3608 => x"e000000f",
     3609 => x"298102c8",  3610 => x"282c0010",  3611 => x"35610038",
     3612 => x"fbfffeb9",  3613 => x"59810058",  3614 => x"3561003c",
     3615 => x"fbfffeb6",  3616 => x"59810054",  3617 => x"35610040",
     3618 => x"fbfffeb3",  3619 => x"59810060",  3620 => x"35610044",
     3621 => x"fbfffeb0",  3622 => x"5981005c",  3623 => x"2b9d0004",
     3624 => x"2b8b0014",  3625 => x"2b8c0010",  3626 => x"2b8d000c",
     3627 => x"2b8e0008",  3628 => x"379c0014",  3629 => x"c3a00000",
     3630 => x"379cfff4",  3631 => x"5b8b000c",  3632 => x"5b8c0008",
     3633 => x"5b9d0004",  3634 => x"2042ffff",  3635 => x"b8205800",
     3636 => x"fbffff1e",  3637 => x"b8206000",  3638 => x"29610024",
     3639 => x"29630070",  3640 => x"29620034",  3641 => x"2827000c",
     3642 => x"b5831800",  3643 => x"b9600800",  3644 => x"356400f8",
     3645 => x"34050000",  3646 => x"34060000",  3647 => x"d8e00000",
     3648 => x"78080001",  3649 => x"390864e4",  3650 => x"4c2c000b",
     3651 => x"29050030",  3652 => x"78040001",  3653 => x"b9600800",
     3654 => x"34020005",  3655 => x"34030001",  3656 => x"38843f58",
     3657 => x"3406000c",  3658 => x"fbfff408",  3659 => x"3401ffff",
     3660 => x"e000000f",  3661 => x"296600f8",  3662 => x"296700fc",
     3663 => x"29080030",  3664 => x"78040001",  3665 => x"b9600800",
     3666 => x"34020005",  3667 => x"34030001",  3668 => x"38843f78",
     3669 => x"b9802800",  3670 => x"fbfff3fc",  3671 => x"2961036c",
     3672 => x"34210001",  3673 => x"5961036c",  3674 => x"34010000",
     3675 => x"2b9d0004",  3676 => x"2b8b000c",  3677 => x"2b8c0008",
     3678 => x"379c000c",  3679 => x"c3a00000",  3680 => x"78020001",
     3681 => x"384264e0",  3682 => x"58410000",  3683 => x"c3a00000",
     3684 => x"379cffe8",  3685 => x"5b8b0018",  3686 => x"5b8c0014",
     3687 => x"5b8d0010",  3688 => x"5b8e000c",  3689 => x"5b8f0008",
     3690 => x"5b9d0004",  3691 => x"282b0014",  3692 => x"b8206800",
     3693 => x"45600014",  3694 => x"780c0001",  3695 => x"398c8f8c",
     3696 => x"29810000",  3697 => x"34020001",  3698 => x"f8001229",
     3699 => x"34020000",  3700 => x"31a0001c",  3701 => x"b9600800",
     3702 => x"34030110",  3703 => x"296f00f0",  3704 => x"296e00f4",
     3705 => x"296d00f8",  3706 => x"f8003d36",  3707 => x"29810000",
     3708 => x"596f00f0",  3709 => x"596e00f4",  3710 => x"596d00f8",
     3711 => x"34020000",  3712 => x"f800121b",  3713 => x"2b9d0004",
     3714 => x"2b8b0018",  3715 => x"2b8c0014",  3716 => x"2b8d0010",
     3717 => x"2b8e000c",  3718 => x"2b8f0008",  3719 => x"379c0018",
     3720 => x"c3a00000",  3721 => x"379cffec",  3722 => x"5b8b0014",
     3723 => x"5b8c0010",  3724 => x"5b8d000c",  3725 => x"5b8e0008",
     3726 => x"5b9d0004",  3727 => x"b8206800",  3728 => x"282102c8",
     3729 => x"780e0001",  3730 => x"39ce8f8c",  3731 => x"282c0010",
     3732 => x"29c10000",  3733 => x"34020001",  3734 => x"29ab0014",
     3735 => x"f8001204",  3736 => x"29810000",  3737 => x"34020000",
     3738 => x"34030000",  3739 => x"2826001c",  3740 => x"35640028",
     3741 => x"b9a00800",  3742 => x"3565002c",  3743 => x"d8c00000",
     3744 => x"3402ffff",  3745 => x"5c200039",  3746 => x"29810000",
     3747 => x"34020000",  3748 => x"28230034",  3749 => x"b9a00800",
     3750 => x"d8600000",  3751 => x"34030010",  3752 => x"35a20358",
     3753 => x"b9600800",  3754 => x"f8003e38",  3755 => x"29810000",
     3756 => x"596000a8",  3757 => x"28220018",  3758 => x"34010000",
     3759 => x"d8400000",  3760 => x"34010002",  3761 => x"59610014",
     3762 => x"29810058",  3763 => x"2d820054",  3764 => x"59600088",
     3765 => x"3c210010",  3766 => x"b8220800",  3767 => x"59610018",
     3768 => x"29810060",  3769 => x"2d82005c",  3770 => x"3c210010",
     3771 => x"b8220800",  3772 => x"5961001c",  3773 => x"2981001c",
     3774 => x"2d820018",  3775 => x"3c210010",  3776 => x"b8220800",
     3777 => x"59610020",  3778 => x"29810024",  3779 => x"2d820020",
     3780 => x"3c210010",  3781 => x"b8220800",  3782 => x"78020001",
     3783 => x"59610024",  3784 => x"38423f9c",  3785 => x"356100c0",
     3786 => x"f8003d78",  3787 => x"29610010",  3788 => x"34020000",
     3789 => x"596000b8",  3790 => x"38210001",  3791 => x"59610010",
     3792 => x"78010001",  3793 => x"382164e0",  3794 => x"28210000",
     3795 => x"596100bc",  3796 => x"78010001",  3797 => x"38217770",
     3798 => x"58200000",  3799 => x"29c10000",  3800 => x"f80011c3",
     3801 => x"34020000",  3802 => x"b8400800",  3803 => x"2b9d0004",
     3804 => x"2b8b0014",  3805 => x"2b8c0010",  3806 => x"2b8d000c",
     3807 => x"2b8e0008",  3808 => x"379c0014",  3809 => x"c3a00000",
     3810 => x"28460000",  3811 => x"28450004",  3812 => x"28440008",
     3813 => x"28210014",  3814 => x"28420010",  3815 => x"58260030",
     3816 => x"58220040",  3817 => x"34020001",  3818 => x"58250034",
     3819 => x"58240038",  3820 => x"5822003c",  3821 => x"28670000",
     3822 => x"28660004",  3823 => x"28650008",  3824 => x"2864000c",
     3825 => x"28630010",  3826 => x"58270044",  3827 => x"58260048",
     3828 => x"5825004c",  3829 => x"58240050",  3830 => x"58230054",
     3831 => x"78010001",  3832 => x"38217770",  3833 => x"58220000",
     3834 => x"34010000",  3835 => x"c3a00000",  3836 => x"379cfff8",
     3837 => x"5b8b0008",  3838 => x"5b9d0004",  3839 => x"282500b0",
     3840 => x"282400b4",  3841 => x"282300b8",  3842 => x"282b0014",
     3843 => x"282700a8",  3844 => x"282600ac",  3845 => x"59650060",
     3846 => x"59640064",  3847 => x"282500bc",  3848 => x"282400c0",
     3849 => x"59630068",  3850 => x"282300c4",  3851 => x"282100cc",
     3852 => x"59670058",  3853 => x"59640070",  3854 => x"5961007c",
     3855 => x"34010001",  3856 => x"59610078",  3857 => x"1441001f",
     3858 => x"59630074",  3859 => x"5966005c",  3860 => x"5965006c",
     3861 => x"34030000",  3862 => x"340403e8",  3863 => x"f8003b46",
     3864 => x"1423001f",  3865 => x"2063ffff",  3866 => x"b4621000",
     3867 => x"f4621800",  3868 => x"00420010",  3869 => x"b4610800",
     3870 => x"3c210010",  3871 => x"b8221000",  3872 => x"34010000",
     3873 => x"59620074",  3874 => x"2b9d0004",  3875 => x"2b8b0008",
     3876 => x"379c0008",  3877 => x"c3a00000",  3878 => x"379cffbc",
     3879 => x"5b8b003c",  3880 => x"5b8c0038",  3881 => x"5b8d0034",
     3882 => x"5b8e0030",  3883 => x"5b8f002c",  3884 => x"5b900028",
     3885 => x"5b910024",  3886 => x"5b920020",  3887 => x"5b93001c",
     3888 => x"5b940018",  3889 => x"5b950014",  3890 => x"5b960010",
     3891 => x"5b97000c",  3892 => x"5b980008",  3893 => x"5b9d0004",
     3894 => x"b8206000",  3895 => x"282102c8",  3896 => x"298b0014",
     3897 => x"282e0010",  3898 => x"78010001",  3899 => x"38217770",
     3900 => x"28210000",  3901 => x"44200283",  3902 => x"2963003c",
     3903 => x"44600007",  3904 => x"29610050",  3905 => x"44200005",
     3906 => x"29610064",  3907 => x"44200003",  3908 => x"29610078",
     3909 => x"5c200011",  3910 => x"78010001",  3911 => x"38217774",
     3912 => x"28220000",  3913 => x"34420001",  3914 => x"58220000",
     3915 => x"34010005",  3916 => x"4c220274",  3917 => x"29640050",
     3918 => x"29650064",  3919 => x"29660078",  3920 => x"78010001",
     3921 => x"78020001",  3922 => x"384259d8",  3923 => x"38213fbc",
     3924 => x"f800222b",  3925 => x"e000026b",  3926 => x"29c10000",
     3927 => x"28230038",  3928 => x"44600004",  3929 => x"b9600800",
     3930 => x"34020000",  3931 => x"d8600000",  3932 => x"78010001",
     3933 => x"38218f8c",  3934 => x"28210000",  3935 => x"34020001",
     3936 => x"f800113b",  3937 => x"78010001",  3938 => x"38217774",
     3939 => x"58200000",  3940 => x"296100b8",  3941 => x"356200fc",
     3942 => x"34210001",  3943 => x"596100b8",  3944 => x"29810028",
     3945 => x"28230000",  3946 => x"b9800800",  3947 => x"d8600000",
     3948 => x"78010001",  3949 => x"38217770",  3950 => x"58200000",
     3951 => x"29660030",  3952 => x"29670034",  3953 => x"29680038",
     3954 => x"2965006c",  3955 => x"29640074",  3956 => x"29610070",
     3957 => x"c8a62800",  3958 => x"c8882000",  3959 => x"c8270800",
     3960 => x"e0000002",  3961 => x"348403e8",  3962 => x"b8201800",
     3963 => x"3421ffff",  3964 => x"4804fffd",  3965 => x"b8a00800",
     3966 => x"78050001",  3967 => x"38a55748",  3968 => x"28a20000",
     3969 => x"e0000002",  3970 => x"b4621800",  3971 => x"b8205000",
     3972 => x"3421ffff",  3973 => x"4803fffd",  3974 => x"29610044",
     3975 => x"29650058",  3976 => x"29620060",  3977 => x"2969005c",
     3978 => x"c8a12800",  3979 => x"2961004c",  3980 => x"c8410800",
     3981 => x"29620048",  3982 => x"c9224800",  3983 => x"e0000002",
     3984 => x"342103e8",  3985 => x"b9201000",  3986 => x"3529ffff",
     3987 => x"4801fffd",  3988 => x"78090001",  3989 => x"39295748",
     3990 => x"292d0000",  3991 => x"e0000002",  3992 => x"b44d1000",
     3993 => x"b8a04800",  3994 => x"34a5ffff",  3995 => x"4802fffd",
     3996 => x"c8810800",  3997 => x"c9495000",  3998 => x"c8622000",
     3999 => x"e0000002",  4000 => x"342103e8",  4001 => x"b8801000",
     4002 => x"3484ffff",  4003 => x"4801fffd",  4004 => x"78040001",
     4005 => x"38845748",  4006 => x"b9401800",  4007 => x"28850000",
     4008 => x"e0000002",  4009 => x"b4451000",  4010 => x"b8602000",
     4011 => x"3463ffff",  4012 => x"4802fffd",  4013 => x"59610094",
     4014 => x"78010001",  4015 => x"3821727c",  4016 => x"59620090",
     4017 => x"28210000",  4018 => x"29820018",  4019 => x"5964008c",
     4020 => x"b8220800",  4021 => x"00210010",  4022 => x"2021000f",
     4023 => x"44200032",  4024 => x"780d0001",  4025 => x"39ad3fec",
     4026 => x"78050001",  4027 => x"b9800800",  4028 => x"34020004",
     4029 => x"34030002",  4030 => x"b9a02000",  4031 => x"38a53ffc",
     4032 => x"fbfff292",  4033 => x"29660044",  4034 => x"29670048",
     4035 => x"2968004c",  4036 => x"78050001",  4037 => x"b9800800",
     4038 => x"34020004",  4039 => x"34030002",  4040 => x"b9a02000",
     4041 => x"38a54008",  4042 => x"fbfff288",  4043 => x"29660058",
     4044 => x"2967005c",  4045 => x"29680060",  4046 => x"78050001",
     4047 => x"b9800800",  4048 => x"34020004",  4049 => x"34030002",
     4050 => x"b9a02000",  4051 => x"38a54014",  4052 => x"fbfff27e",
     4053 => x"2966006c",  4054 => x"29670070",  4055 => x"29680074",
     4056 => x"78050001",  4057 => x"b9800800",  4058 => x"34020004",
     4059 => x"34030002",  4060 => x"b9a02000",  4061 => x"38a54020",
     4062 => x"fbfff274",  4063 => x"2966008c",  4064 => x"29670090",
     4065 => x"29680094",  4066 => x"78050001",  4067 => x"b9800800",
     4068 => x"34020004",  4069 => x"34030002",  4070 => x"b9a02000",
     4071 => x"38a5402c",  4072 => x"fbfff26a",  4073 => x"2962008c",
     4074 => x"78050001",  4075 => x"38a55754",  4076 => x"28a40000",
     4077 => x"1441001f",  4078 => x"340300e8",  4079 => x"f8003a6e",
     4080 => x"b8406800",  4081 => x"29620090",  4082 => x"b8207800",
     4083 => x"34030000",  4084 => x"1441001f",  4085 => x"340403e8",
     4086 => x"f8003a67",  4087 => x"29660094",  4088 => x"b5a21800",
     4089 => x"f5a36800",  4090 => x"14c2001f",  4091 => x"b5e10800",
     4092 => x"b4663000",  4093 => x"b5a10800",  4094 => x"f4661800",
     4095 => x"b4220800",  4096 => x"29650018",  4097 => x"29620020",
     4098 => x"2964001c",  4099 => x"b4610800",  4100 => x"29630024",
     4101 => x"b4a21000",  4102 => x"b4441000",  4103 => x"b4431000",
     4104 => x"1444001f",  4105 => x"297600a0",  4106 => x"297400a4",
     4107 => x"596100a0",  4108 => x"596600a4",  4109 => x"48810004",
     4110 => x"5c810005",  4111 => x"54460002",  4112 => x"e0000003",
     4113 => x"596400a0",  4114 => x"596200a4",  4115 => x"296600a4",
     4116 => x"296100a0",  4117 => x"1477001f",  4118 => x"c8c21000",
     4119 => x"f4463000",  4120 => x"c8240800",  4121 => x"c8260800",
     4122 => x"b4652000",  4123 => x"14a6001f",  4124 => x"f4641800",
     4125 => x"b6e6b800",  4126 => x"b477b800",  4127 => x"004d0001",
     4128 => x"3c23001f",  4129 => x"00250001",  4130 => x"b86d6800",
     4131 => x"b48d6800",  4132 => x"f48d2000",  4133 => x"b6e5b800",
     4134 => x"b497b800",  4135 => x"29640028",  4136 => x"1483001f",
     4137 => x"f8003a34",  4138 => x"14350008",  4139 => x"1421001f",
     4140 => x"b5b5a800",  4141 => x"f5b56800",  4142 => x"b6e10800",
     4143 => x"b5a1b800",  4144 => x"29620030",  4145 => x"29610044",
     4146 => x"29720038",  4147 => x"29630034",  4148 => x"c8411000",
     4149 => x"2961004c",  4150 => x"ca419000",  4151 => x"29610048",
     4152 => x"c8611800",  4153 => x"e0000002",  4154 => x"365203e8",
     4155 => x"b8606800",  4156 => x"3463ffff",  4157 => x"4812fffd",
     4158 => x"78090001",  4159 => x"39295748",  4160 => x"29210000",
     4161 => x"e0000002",  4162 => x"b5a16800",  4163 => x"b8408800",
     4164 => x"3442ffff",  4165 => x"480dfffd",  4166 => x"378f0040",
     4167 => x"340203e8",  4168 => x"b9e00800",  4169 => x"5b970040",
     4170 => x"5b950044",  4171 => x"fbfff62f",  4172 => x"78030001",
     4173 => x"38635748",  4174 => x"28620000",  4175 => x"b8208000",
     4176 => x"b9e00800",  4177 => x"fbfff629",  4178 => x"2b820044",
     4179 => x"b42d6800",  4180 => x"b6509000",  4181 => x"b6221000",
     4182 => x"340103e7",  4183 => x"e0000002",  4184 => x"3652fc18",
     4185 => x"b9a08800",  4186 => x"ba408000",  4187 => x"35ad0001",
     4188 => x"4a41fffc",  4189 => x"78040001",  4190 => x"78050001",
     4191 => x"38845758",  4192 => x"38a5575c",  4193 => x"b8400800",
     4194 => x"28830000",  4195 => x"28a20000",  4196 => x"e0000002",
     4197 => x"b6228800",  4198 => x"b8207800",  4199 => x"ba206800",
     4200 => x"34210001",  4201 => x"4a23fffc",  4202 => x"2961002c",
     4203 => x"340203e8",  4204 => x"b9e0c000",  4205 => x"342103e7",
     4206 => x"f8003a16",  4207 => x"b8209800",  4208 => x"4c110008",
     4209 => x"ba200800",  4210 => x"ba601000",  4211 => x"f8003a3e",
     4212 => x"4420000a",  4213 => x"083003e8",  4214 => x"ca216800",
     4215 => x"b6128000",  4216 => x"4da00006",  4217 => x"78090001",
     4218 => x"39295748",  4219 => x"29210000",  4220 => x"35efffff",
     4221 => x"b5a16800",  4222 => x"3401ffff",  4223 => x"5de10007",
     4224 => x"4c0d0006",  4225 => x"78020001",  4226 => x"3842575c",
     4227 => x"28410000",  4228 => x"340f0000",  4229 => x"b5a16800",
     4230 => x"4da00007",  4231 => x"c8130800",  4232 => x"482d0005",
     4233 => x"5de00004",  4234 => x"b5b36800",  4235 => x"0a73fc18",
     4236 => x"b6138000",  4237 => x"78050001",  4238 => x"38a55754",
     4239 => x"28a40000",  4240 => x"1701001f",  4241 => x"bb001000",
     4242 => x"340300e8",  4243 => x"f80039ca",  4244 => x"b820c000",
     4245 => x"1621001f",  4246 => x"b8409800",  4247 => x"34030000",
     4248 => x"340403e8",  4249 => x"ba201000",  4250 => x"f80039c3",
     4251 => x"b6621800",  4252 => x"f6639800",  4253 => x"1642001f",
     4254 => x"b7010800",  4255 => x"b4729000",  4256 => x"b6610800",
     4257 => x"b4220800",  4258 => x"f4721800",  4259 => x"78020001",
     4260 => x"384264e0",  4261 => x"b4611800",  4262 => x"28410000",
     4263 => x"596300e8",  4264 => x"34020000",  4265 => x"596100bc",
     4266 => x"29c10000",  4267 => x"597200ec",  4268 => x"597700b0",
     4269 => x"28230004",  4270 => x"597500b4",  4271 => x"b9800800",
     4272 => x"d8600000",  4273 => x"34020001",  4274 => x"4422000c",
     4275 => x"78040001",  4276 => x"b9800800",  4277 => x"34020004",
     4278 => x"34030001",  4279 => x"38844038",  4280 => x"fbfff19a",
     4281 => x"29c10000",  4282 => x"34020000",  4283 => x"28230034",
     4284 => x"b9800800",  4285 => x"d8600000",  4286 => x"29c10000",
     4287 => x"28210010",  4288 => x"d8200000",  4289 => x"5c200007",
     4290 => x"29630010",  4291 => x"3402fffd",  4292 => x"a0621000",
     4293 => x"59620010",  4294 => x"5de10009",  4295 => x"e000000a",
     4296 => x"78040001",  4297 => x"b9800800",  4298 => x"34020004",
     4299 => x"34030001",  4300 => x"3884405c",  4301 => x"fbfff185",
     4302 => x"e00000e7",  4303 => x"34010002",  4304 => x"e0000003",
     4305 => x"45af0003",  4306 => x"34010001",  4307 => x"59610014",
     4308 => x"78040001",  4309 => x"b9800800",  4310 => x"34020004",
     4311 => x"b9e02800",  4312 => x"b9a03000",  4313 => x"34030002",
     4314 => x"38844068",  4315 => x"ba003800",  4316 => x"fbfff176",
     4317 => x"29620014",  4318 => x"78010001",  4319 => x"382159c0",
     4320 => x"3c420002",  4321 => x"78060001",  4322 => x"b4220800",
     4323 => x"28250000",  4324 => x"29610010",  4325 => x"38c65740",
     4326 => x"20210002",  4327 => x"44200003",  4328 => x"78060001",
     4329 => x"38c63fac",  4330 => x"78040001",  4331 => x"b9800800",
     4332 => x"34020004",  4333 => x"34030001",  4334 => x"38844088",
     4335 => x"fbfff163",  4336 => x"29620014",  4337 => x"78010001",
     4338 => x"382159c0",  4339 => x"3c420002",  4340 => x"b4221000",
     4341 => x"28420000",  4342 => x"356100c0",  4343 => x"f8003b4b",
     4344 => x"29620014",  4345 => x"34010004",  4346 => x"3442ffff",
     4347 => x"54410083",  4348 => x"78010001",  4349 => x"3c420002",
     4350 => x"382159ac",  4351 => x"b4220800",  4352 => x"28210000",
     4353 => x"c0200000",  4354 => x"29c10000",  4355 => x"b9e01000",
     4356 => x"34030000",  4357 => x"28240014",  4358 => x"15e1001f",
     4359 => x"e0000006",  4360 => x"29c10000",  4361 => x"34020000",
     4362 => x"b9a01800",  4363 => x"28240014",  4364 => x"34010000",
     4365 => x"d8800000",  4366 => x"29610010",  4367 => x"38210002",
     4368 => x"59610010",  4369 => x"e0000057",  4370 => x"296500a8",
     4371 => x"78040001",  4372 => x"b9800800",  4373 => x"34020004",
     4374 => x"34030002",  4375 => x"388440a0",  4376 => x"b9a03000",
     4377 => x"ba003800",  4378 => x"fbfff138",  4379 => x"29c20000",
     4380 => x"296100a8",  4381 => x"28420018",  4382 => x"b6010800",
     4383 => x"596100a8",  4384 => x"d8400000",  4385 => x"29610010",
     4386 => x"38210002",  4387 => x"59610010",  4388 => x"34010005",
     4389 => x"59610014",  4390 => x"e0000058",  4391 => x"78090001",
     4392 => x"39295754",  4393 => x"29240000",  4394 => x"15e1001f",
     4395 => x"b9e01000",  4396 => x"340300e8",  4397 => x"f8003930",
     4398 => x"b6027800",  4399 => x"1611001f",  4400 => x"f60f8000",
     4401 => x"b6210800",  4402 => x"b6018000",  4403 => x"15a1001f",
     4404 => x"34030000",  4405 => x"b9a01000",  4406 => x"340403e8",
     4407 => x"f8003926",  4408 => x"b5e21800",  4409 => x"f5e37800",
     4410 => x"b6010800",  4411 => x"b5e10800",  4412 => x"c8031000",
     4413 => x"48010002",  4414 => x"b8601000",  4415 => x"3401003b",
     4416 => x"4841000d",  4417 => x"29c10000",  4418 => x"34020001",
     4419 => x"28230034",  4420 => x"b9800800",  4421 => x"d8600000",
     4422 => x"296100b0",  4423 => x"59610080",  4424 => x"296100b4",
     4425 => x"59610084",  4426 => x"34010004",  4427 => x"59610014",
     4428 => x"e0000004",  4429 => x"29610088",  4430 => x"34210001",
     4431 => x"59610088",  4432 => x"29620088",  4433 => x"34010009",
     4434 => x"4c22002c",  4435 => x"59600088",  4436 => x"e0000014",
     4437 => x"296300b4",  4438 => x"29610084",  4439 => x"296400b0",
     4440 => x"29620080",  4441 => x"c8610800",  4442 => x"f4231800",
     4443 => x"596100e4",  4444 => x"78010001",  4445 => x"382164e0",
     4446 => x"c8821000",  4447 => x"28210000",  4448 => x"c8431000",
     4449 => x"596200e0",  4450 => x"4420001c",  4451 => x"1601001f",
     4452 => x"34030078",  4453 => x"98301000",  4454 => x"c8411000",
     4455 => x"4c620003",  4456 => x"34010003",  4457 => x"e3ffffbc",
     4458 => x"0021001e",  4459 => x"29c20000",  4460 => x"b4308000",
     4461 => x"296100a8",  4462 => x"16100002",  4463 => x"28420018",
     4464 => x"b6010800",  4465 => x"596100a8",  4466 => x"d8400000",
     4467 => x"296500a8",  4468 => x"78040001",  4469 => x"b9800800",
     4470 => x"34020006",  4471 => x"34030001",  4472 => x"388440bc",
     4473 => x"fbfff0d9",  4474 => x"296100b0",  4475 => x"59610080",
     4476 => x"296100b4",  4477 => x"59610084",  4478 => x"29620014",
     4479 => x"34010004",  4480 => x"44410004",  4481 => x"296100f0",
     4482 => x"34210001",  4483 => x"596100f0",  4484 => x"296400e8",
     4485 => x"296300ec",  4486 => x"1481001f",  4487 => x"98611800",
     4488 => x"c8611000",  4489 => x"98812000",  4490 => x"f4431800",
     4491 => x"c8810800",  4492 => x"c8230800",  4493 => x"48200005",
     4494 => x"5c200007",  4495 => x"340101f4",  4496 => x"54410002",
     4497 => x"e0000004",  4498 => x"296100f4",  4499 => x"34210001",
     4500 => x"596100f4",  4501 => x"296500a4",  4502 => x"296400a0",
     4503 => x"ca851800",  4504 => x"f4740800",  4505 => x"cac41000",
     4506 => x"c8411000",  4507 => x"48020007",  4508 => x"34010001",
     4509 => x"48400013",  4510 => x"5c400011",  4511 => x"340203e8",
     4512 => x"54620010",  4513 => x"e000000e",  4514 => x"c8140800",
     4515 => x"7c220000",  4516 => x"c8161800",  4517 => x"c8621800",
     4518 => x"c8251000",  4519 => x"f4410800",  4520 => x"c8641800",
     4521 => x"c8611800",  4522 => x"34010001",  4523 => x"48600005",
     4524 => x"5c600003",  4525 => x"340303e8",  4526 => x"54430002",
     4527 => x"34010000",  4528 => x"202100ff",  4529 => x"44200004",
     4530 => x"296100f8",  4531 => x"34210001",  4532 => x"596100f8",
     4533 => x"78010001",  4534 => x"38218f8c",  4535 => x"28210000",
     4536 => x"34020000",  4537 => x"f8000ee2",  4538 => x"29c10000",
     4539 => x"28230038",  4540 => x"44600004",  4541 => x"b9600800",
     4542 => x"34020001",  4543 => x"d8600000",  4544 => x"34010000",
     4545 => x"2b9d0004",  4546 => x"2b8b003c",  4547 => x"2b8c0038",
     4548 => x"2b8d0034",  4549 => x"2b8e0030",  4550 => x"2b8f002c",
     4551 => x"2b900028",  4552 => x"2b910024",  4553 => x"2b920020",
     4554 => x"2b93001c",  4555 => x"2b940018",  4556 => x"2b950014",
     4557 => x"2b960010",  4558 => x"2b97000c",  4559 => x"2b980008",
     4560 => x"379c0044",  4561 => x"c3a00000",  4562 => x"379cffe8",
     4563 => x"5b8b0018",  4564 => x"5b8c0014",  4565 => x"5b8d0010",
     4566 => x"5b8e000c",  4567 => x"5b8f0008",  4568 => x"5b9d0004",
     4569 => x"b8407800",  4570 => x"28220020",  4571 => x"b8205800",
     4572 => x"b8607000",  4573 => x"284d0008",  4574 => x"28220024",
     4575 => x"282c02c8",  4576 => x"28440000",  4577 => x"d8800000",
     4578 => x"48010058",  4579 => x"29610020",  4580 => x"34030008",
     4581 => x"2824000c",  4582 => x"4161004c",  4583 => x"30810004",
     4584 => x"4161004d",  4585 => x"30810005",  4586 => x"4161004e",
     4587 => x"30810006",  4588 => x"3401ffff",  4589 => x"30810007",
     4590 => x"3401fffe",  4591 => x"30810008",  4592 => x"4161004f",
     4593 => x"30810009",  4594 => x"41610050",  4595 => x"3081000a",
     4596 => x"41610051",  4597 => x"3081000b",  4598 => x"29610020",
     4599 => x"2824000c",  4600 => x"b9800800",  4601 => x"34820004",
     4602 => x"f8003938",  4603 => x"29610020",  4604 => x"35620374",
     4605 => x"28210000",  4606 => x"3180000a",  4607 => x"c8410800",
     4608 => x"14210002",  4609 => x"0821d775",  4610 => x"0d810008",
     4611 => x"41a10042",  4612 => x"3181000b",  4613 => x"34010014",
     4614 => x"3181000c",  4615 => x"41a10043",  4616 => x"3181000d",
     4617 => x"34010002",  4618 => x"3181000e",  4619 => x"78010001",
     4620 => x"382164ac",  4621 => x"28240000",  4622 => x"4480000f",
     4623 => x"b9600800",  4624 => x"b9e01000",  4625 => x"b9c01800",
     4626 => x"d8800000",  4627 => x"4420000a",  4628 => x"78040001",
     4629 => x"78050001",  4630 => x"b9600800",  4631 => x"34020002",
     4632 => x"34030001",  4633 => x"38844128",  4634 => x"38a559e8",
     4635 => x"fbfff037",  4636 => x"e000001e",  4637 => x"29610020",
     4638 => x"78040001",  4639 => x"34020003",  4640 => x"2825000c",
     4641 => x"34030001",  4642 => x"b9600800",  4643 => x"40a5000e",
     4644 => x"38844144",  4645 => x"fbfff02d",  4646 => x"29610020",
     4647 => x"78040001",  4648 => x"34020003",  4649 => x"2825000c",
     4650 => x"34030001",  4651 => x"b9600800",  4652 => x"40a5000f",
     4653 => x"38844158",  4654 => x"fbfff024",  4655 => x"2962003c",
     4656 => x"b9600800",  4657 => x"f8000634",  4658 => x"4162001d",
     4659 => x"34010001",  4660 => x"44410003",  4661 => x"34010004",
     4662 => x"e0000002",  4663 => x"34010006",  4664 => x"59610004",
     4665 => x"e0000003",  4666 => x"340103e8",  4667 => x"59610008",
     4668 => x"34010000",  4669 => x"2b9d0004",  4670 => x"2b8b0018",
     4671 => x"2b8c0014",  4672 => x"2b8d0010",  4673 => x"2b8e000c",
     4674 => x"2b8f0008",  4675 => x"379c0018",  4676 => x"c3a00000",
     4677 => x"379cfff4",  4678 => x"5b8b000c",  4679 => x"5b8c0008",
     4680 => x"5b9d0004",  4681 => x"2822000c",  4682 => x"b8205800",
     4683 => x"44400006",  4684 => x"28220028",  4685 => x"28430018",
     4686 => x"34020fa0",  4687 => x"d8600000",  4688 => x"596102dc",
     4689 => x"296102dc",  4690 => x"44200009",  4691 => x"29610028",
     4692 => x"34020000",  4693 => x"28230018",  4694 => x"b9600800",
     4695 => x"d8600000",  4696 => x"296202dc",  4697 => x"c8220800",
     4698 => x"4c200014",  4699 => x"296c02dc",  4700 => x"34010000",
     4701 => x"4580000a",  4702 => x"29610028",  4703 => x"34020000",
     4704 => x"28230018",  4705 => x"b9600800",  4706 => x"d8600000",
     4707 => x"c9810800",  4708 => x"a4201000",  4709 => x"1442001f",
     4710 => x"a0220800",  4711 => x"59610008",  4712 => x"34010000",
     4713 => x"2b9d0004",  4714 => x"2b8b000c",  4715 => x"2b8c0008",
     4716 => x"379c000c",  4717 => x"c3a00000",  4718 => x"b9600800",
     4719 => x"34020004",  4720 => x"f8000a67",  4721 => x"34010001",
     4722 => x"59610004",  4723 => x"e3fffff5",  4724 => x"340203e8",
     4725 => x"58220008",  4726 => x"34010000",  4727 => x"c3a00000",
     4728 => x"379cfff0",  4729 => x"5b8b0010",  4730 => x"5b8c000c",
     4731 => x"5b8d0008",  4732 => x"5b9d0004",  4733 => x"78040001",
     4734 => x"388464ac",  4735 => x"2884000c",  4736 => x"b8205800",
     4737 => x"b8406800",  4738 => x"b8606000",  4739 => x"44800003",
     4740 => x"d8800000",  4741 => x"5c20001f",  4742 => x"2961000c",
     4743 => x"4420000b",  4744 => x"296102c8",  4745 => x"29630028",
     4746 => x"4022000c",  4747 => x"1021000b",  4748 => x"28630018",
     4749 => x"bc411000",  4750 => x"b9600800",  4751 => x"084203e8",
     4752 => x"d8600000",  4753 => x"596102d4",  4754 => x"4580000f",
     4755 => x"4161030d",  4756 => x"44200008",  4757 => x"3402000b",
     4758 => x"5c22000b",  4759 => x"b9600800",  4760 => x"b9a01000",
     4761 => x"b9801800",  4762 => x"f8000352",  4763 => x"e0000005",
     4764 => x"b9600800",  4765 => x"b9a01000",  4766 => x"b9801800",
     4767 => x"f8000370",  4768 => x"5c200004",  4769 => x"b9600800",
     4770 => x"f800027e",  4771 => x"44200003",  4772 => x"34010002",
     4773 => x"59610004",  4774 => x"29620004",  4775 => x"29610000",
     4776 => x"44410002",  4777 => x"596002d4",  4778 => x"296c02d4",
     4779 => x"34010000",  4780 => x"4580000a",  4781 => x"29610028",
     4782 => x"34020000",  4783 => x"28230018",  4784 => x"b9600800",
     4785 => x"d8600000",  4786 => x"c9810800",  4787 => x"a4201000",
     4788 => x"1442001f",  4789 => x"a0220800",  4790 => x"59610008",
     4791 => x"34010000",  4792 => x"2b9d0004",  4793 => x"2b8b0010",
     4794 => x"2b8c000c",  4795 => x"2b8d0008",  4796 => x"379c0010",
     4797 => x"c3a00000",  4798 => x"34010000",  4799 => x"c3a00000",
     4800 => x"379cffec",  4801 => x"5b8b0014",  4802 => x"5b8c0010",
     4803 => x"5b8d000c",  4804 => x"5b8e0008",  4805 => x"5b9d0004",
     4806 => x"344b00b2",  4807 => x"3d6b0002",  4808 => x"b8407000",
     4809 => x"b42b5800",  4810 => x"29620004",  4811 => x"b8206000",
     4812 => x"340d0000",  4813 => x"44400008",  4814 => x"28220028",
     4815 => x"28430018",  4816 => x"34020000",  4817 => x"d8600000",
     4818 => x"29620004",  4819 => x"c8220800",  4820 => x"4c200009",
     4821 => x"b9a00800",  4822 => x"2b9d0004",  4823 => x"2b8b0014",
     4824 => x"2b8c0010",  4825 => x"2b8d000c",  4826 => x"2b8e0008",
     4827 => x"379c0014",  4828 => x"c3a00000",  4829 => x"b9800800",
     4830 => x"b9c01000",  4831 => x"f80009f8",  4832 => x"340d0001",
     4833 => x"59600004",  4834 => x"e3fffff3",  4835 => x"379cffec",
     4836 => x"5b8b0014",  4837 => x"5b8c0010",  4838 => x"5b8d000c",
     4839 => x"5b8e0008",  4840 => x"5b9d0004",  4841 => x"b8407000",
     4842 => x"2822000c",  4843 => x"b8205800",  4844 => x"b8606800",
     4845 => x"340c0000",  4846 => x"44400014",  4847 => x"282302c8",
     4848 => x"34020001",  4849 => x"1063000d",  4850 => x"f80009f4",
     4851 => x"296302c8",  4852 => x"b9600800",  4853 => x"34020003",
     4854 => x"1063000b",  4855 => x"f80009ef",  4856 => x"29630344",
     4857 => x"34020001",  4858 => x"34010000",  4859 => x"5c620002",
     4860 => x"29610340",  4861 => x"0d61007e",  4862 => x"b9600800",
     4863 => x"f80005d9",  4864 => x"b8206000",  4865 => x"48010047",
     4866 => x"b9600800",  4867 => x"34020001",  4868 => x"fbffffbc",
     4869 => x"44200010",  4870 => x"296302c8",  4871 => x"b9600800",
     4872 => x"34020001",  4873 => x"1063000d",  4874 => x"f80009dc",
     4875 => x"29630344",  4876 => x"34020001",  4877 => x"34010000",
     4878 => x"5c620002",  4879 => x"29610340",  4880 => x"0d61007e",
     4881 => x"b9600800",  4882 => x"f8000613",  4883 => x"48010046",
     4884 => x"340c0000",  4885 => x"b9600800",  4886 => x"34020003",
     4887 => x"fbffffa9",  4888 => x"44200010",  4889 => x"29630344",
     4890 => x"34020001",  4891 => x"34010000",  4892 => x"5c620002",
     4893 => x"29610340",  4894 => x"0d61007e",  4895 => x"b9600800",
     4896 => x"f80005b8",  4897 => x"48010038",  4898 => x"296302c8",
     4899 => x"b9600800",  4900 => x"34020003",  4901 => x"1063000b",
     4902 => x"340c0000",  4903 => x"f80009bf",  4904 => x"45a00020",
     4905 => x"78010001",  4906 => x"382164ac",  4907 => x"28250010",
     4908 => x"4164030d",  4909 => x"44a00007",  4910 => x"b9600800",
     4911 => x"b9c01000",  4912 => x"b9a01800",  4913 => x"d8a00000",
     4914 => x"b8202000",  4915 => x"48010042",  4916 => x"34010001",
     4917 => x"44810010",  4918 => x"3401000b",  4919 => x"44810003",
     4920 => x"5c800010",  4921 => x"e0000006",  4922 => x"b9600800",
     4923 => x"b9c01000",  4924 => x"b9a01800",  4925 => x"f80002af",
     4926 => x"e0000005",  4927 => x"b9600800",  4928 => x"b9c01000",
     4929 => x"b9a01800",  4930 => x"f80002cd",  4931 => x"b8206000",
     4932 => x"e0000004",  4933 => x"b9600800",  4934 => x"356200e4",
     4935 => x"f800066a",  4936 => x"45800006",  4937 => x"34010001",
     4938 => x"4581000f",  4939 => x"3401ffff",  4940 => x"5d81000e",
     4941 => x"e0000029",  4942 => x"29610020",  4943 => x"2821000c",
     4944 => x"4022000e",  4945 => x"340100ff",  4946 => x"44410004",
     4947 => x"4162001d",  4948 => x"34010002",  4949 => x"5c410005",
     4950 => x"34010004",  4951 => x"59610004",  4952 => x"e0000002",
     4953 => x"340c0000",  4954 => x"296e02d8",  4955 => x"340d0000",
     4956 => x"45c0000a",  4957 => x"29610028",  4958 => x"34020000",
     4959 => x"28230018",  4960 => x"b9600800",  4961 => x"d8600000",
     4962 => x"c9c16800",  4963 => x"a5a00800",  4964 => x"1421001f",
     4965 => x"a1a16800",  4966 => x"296e02d0",  4967 => x"34010000",
     4968 => x"45c0000a",  4969 => x"29610028",  4970 => x"34020000",
     4971 => x"28230018",  4972 => x"b9600800",  4973 => x"d8600000",
     4974 => x"c9c10800",  4975 => x"a4201000",  4976 => x"1442001f",
     4977 => x"a0220800",  4978 => x"4da10007",  4979 => x"b9a00800",
     4980 => x"e0000005",  4981 => x"b8206000",  4982 => x"34010002",
     4983 => x"59610004",  4984 => x"340101f4",  4985 => x"59610008",
     4986 => x"b9800800",  4987 => x"2b9d0004",  4988 => x"2b8b0014",
     4989 => x"2b8c0010",  4990 => x"2b8d000c",  4991 => x"2b8e0008",
     4992 => x"379c0014",  4993 => x"c3a00000",  4994 => x"379cfff0",
     4995 => x"5b8b000c",  4996 => x"5b8c0008",  4997 => x"5b9d0004",
     4998 => x"b8406000",  4999 => x"2822000c",  5000 => x"b8205800",
     5001 => x"4440000c",  5002 => x"282202c8",  5003 => x"28250028",
     5004 => x"4044000c",  5005 => x"1042000b",  5006 => x"bc821000",
     5007 => x"28a40018",  5008 => x"084203e8",  5009 => x"5b830010",
     5010 => x"d8800000",  5011 => x"2b830010",  5012 => x"596102d4",
     5013 => x"4460000d",  5014 => x"4161030d",  5015 => x"44200007",
     5016 => x"3402000b",  5017 => x"5c220009",  5018 => x"b9600800",
     5019 => x"b9801000",  5020 => x"f8000250",  5021 => x"e0000004",
     5022 => x"b9600800",  5023 => x"b9801000",  5024 => x"f800026f",
     5025 => x"5c200004",  5026 => x"b9600800",  5027 => x"f800017d",
     5028 => x"44200003",  5029 => x"34010002",  5030 => x"59610004",
     5031 => x"29620004",  5032 => x"29610000",  5033 => x"44410002",
     5034 => x"596002d4",  5035 => x"340103e8",  5036 => x"59610008",
     5037 => x"34010000",  5038 => x"2b9d0004",  5039 => x"2b8b000c",
     5040 => x"2b8c0008",  5041 => x"379c0010",  5042 => x"c3a00000",
     5043 => x"379cfff8",  5044 => x"5b8b0008",  5045 => x"5b9d0004",
     5046 => x"b8205800",  5047 => x"4460000d",  5048 => x"4024030d",
     5049 => x"44800007",  5050 => x"34050008",  5051 => x"44850007",
     5052 => x"3405000b",  5053 => x"5c850007",  5054 => x"f8000198",
     5055 => x"e0000004",  5056 => x"f80001b1",  5057 => x"e0000002",
     5058 => x"f80001e9",  5059 => x"5c200004",  5060 => x"b9600800",
     5061 => x"f800015b",  5062 => x"44200003",  5063 => x"34010002",
     5064 => x"59610004",  5065 => x"340103e8",  5066 => x"59610008",
     5067 => x"34010000",  5068 => x"2b9d0004",  5069 => x"2b8b0008",
     5070 => x"379c0008",  5071 => x"c3a00000",  5072 => x"379cffd4",
     5073 => x"5b8b0014",  5074 => x"5b8c0010",  5075 => x"5b8d000c",
     5076 => x"5b8e0008",  5077 => x"5b9d0004",  5078 => x"b8205800",
     5079 => x"2821000c",  5080 => x"b8407000",  5081 => x"b8606800",
     5082 => x"44200023",  5083 => x"34020000",  5084 => x"34030014",
     5085 => x"35610080",  5086 => x"f80037d2",  5087 => x"b9600800",
     5088 => x"f80006da",  5089 => x"78010001",  5090 => x"382164ac",
     5091 => x"28240014",  5092 => x"44800007",  5093 => x"b9600800",
     5094 => x"b9c01000",  5095 => x"b9a01800",  5096 => x"d8800000",
     5097 => x"b8206000",  5098 => x"5c20005f",  5099 => x"4161001c",
     5100 => x"29630028",  5101 => x"202100fd",  5102 => x"3161001c",
     5103 => x"296102c8",  5104 => x"28630018",  5105 => x"4022000c",
     5106 => x"1021000b",  5107 => x"bc411000",  5108 => x"b9600800",
     5109 => x"084203e8",  5110 => x"d8600000",  5111 => x"296302c8",
     5112 => x"596102d4",  5113 => x"34020000",  5114 => x"1063000a",
     5115 => x"b9600800",  5116 => x"f80008ea",  5117 => x"45a00049",
     5118 => x"4161030d",  5119 => x"34020008",  5120 => x"44220012",
     5121 => x"54220003",  5122 => x"5c200044",  5123 => x"e000000a",
     5124 => x"34020009",  5125 => x"44220014",  5126 => x"3402000b",
     5127 => x"5c22003f",  5128 => x"b9600800",  5129 => x"b9c01000",
     5130 => x"b9a01800",  5131 => x"f800014b",  5132 => x"e000000a",
     5133 => x"b9600800",  5134 => x"b9c01000",  5135 => x"b9a01800",
     5136 => x"f8000161",  5137 => x"e0000005",  5138 => x"b9600800",
     5139 => x"b9c01000",  5140 => x"b9a01800",  5141 => x"f8000196",
     5142 => x"b8206000",  5143 => x"5c200032",  5144 => x"e000002e",
     5145 => x"34010035",  5146 => x"340c0001",  5147 => x"4c2d002e",
     5148 => x"378c0018",  5149 => x"b9c00800",  5150 => x"b9801000",
     5151 => x"f80004a2",  5152 => x"296102c8",  5153 => x"37820024",
     5154 => x"34030008",  5155 => x"f80036ee",  5156 => x"5c20001c",
     5157 => x"2d6202f2",  5158 => x"2d61032a",  5159 => x"5c410019",
     5160 => x"296102c8",  5161 => x"2c220008",  5162 => x"2f81002c",
     5163 => x"5c410015",  5164 => x"4161001c",  5165 => x"20210001",
     5166 => x"44200012",  5167 => x"b9801000",  5168 => x"356100bc",
     5169 => x"f8000619",  5170 => x"78010001",  5171 => x"382164ac",
     5172 => x"28220018",  5173 => x"44400006",  5174 => x"b9600800",
     5175 => x"d8400000",  5176 => x"b8206000",  5177 => x"5c200010",
     5178 => x"e0000003",  5179 => x"b9600800",  5180 => x"f80006d7",
     5181 => x"4161032d",  5182 => x"316102ee",  5183 => x"e0000007",
     5184 => x"78040001",  5185 => x"b9600800",  5186 => x"34020005",
     5187 => x"34030002",  5188 => x"38844170",  5189 => x"fbffee0d",
     5190 => x"b9600800",  5191 => x"f80000d9",  5192 => x"b8206000",
     5193 => x"296102cc",  5194 => x"44200009",  5195 => x"29610028",
     5196 => x"34020000",  5197 => x"28230018",  5198 => x"b9600800",
     5199 => x"d8600000",  5200 => x"296202cc",  5201 => x"c8220800",
     5202 => x"4c200033",  5203 => x"3401ffff",  5204 => x"45810005",
     5205 => x"7d810001",  5206 => x"c8010800",  5207 => x"a1816000",
     5208 => x"e0000003",  5209 => x"34010002",  5210 => x"59610004",
     5211 => x"29620004",  5212 => x"29610000",  5213 => x"44410005",
     5214 => x"596002d4",  5215 => x"596002cc",  5216 => x"b9600800",
     5217 => x"f8000659",  5218 => x"296e02d4",  5219 => x"340d0000",
     5220 => x"45c0000a",  5221 => x"29610028",  5222 => x"34020000",
     5223 => x"28230018",  5224 => x"b9600800",  5225 => x"d8600000",
     5226 => x"c9c16800",  5227 => x"a5a00800",  5228 => x"1421001f",
     5229 => x"a1a16800",  5230 => x"296e02cc",  5231 => x"b9a00800",
     5232 => x"45c0000a",  5233 => x"29610028",  5234 => x"34020000",
     5235 => x"28230018",  5236 => x"b9600800",  5237 => x"d8600000",
     5238 => x"c9c10800",  5239 => x"a4201000",  5240 => x"1442001f",
     5241 => x"a0220800",  5242 => x"4da10002",  5243 => x"b9a00800",
     5244 => x"59610008",  5245 => x"b9800800",  5246 => x"2b9d0004",
     5247 => x"2b8b0014",  5248 => x"2b8c0010",  5249 => x"2b8d000c",
     5250 => x"2b8e0008",  5251 => x"379c002c",  5252 => x"c3a00000",
     5253 => x"b9600800",  5254 => x"34020000",  5255 => x"f8000850",
     5256 => x"b9600800",  5257 => x"596002cc",  5258 => x"f80004f6",
     5259 => x"29630100",  5260 => x"29620104",  5261 => x"296500f8",
     5262 => x"296400fc",  5263 => x"b8206000",  5264 => x"29610108",
     5265 => x"596300b0",  5266 => x"296302c8",  5267 => x"596200b4",
     5268 => x"596100b8",  5269 => x"596500a8",  5270 => x"596400ac",
     5271 => x"1063000a",  5272 => x"b9600800",  5273 => x"34020000",
     5274 => x"f800084c",  5275 => x"29620020",  5276 => x"356100a8",
     5277 => x"28430008",  5278 => x"b8201000",  5279 => x"34630018",
     5280 => x"f80005bd",  5281 => x"e3ffffb2",  5282 => x"379cfff8",
     5283 => x"5b8b0008",  5284 => x"5b9d0004",  5285 => x"282202c8",
     5286 => x"28240028",  5287 => x"b8205800",  5288 => x"4043000c",
     5289 => x"1042000b",  5290 => x"bc621000",  5291 => x"28830018",
     5292 => x"084203e8",  5293 => x"d8600000",  5294 => x"596102d4",
     5295 => x"2b9d0004",  5296 => x"2b8b0008",  5297 => x"379c0008",
     5298 => x"c3a00000",  5299 => x"379cffe4",  5300 => x"5b8b001c",
     5301 => x"5b8c0018",  5302 => x"5b8d0014",  5303 => x"5b8e0010",
     5304 => x"5b8f000c",  5305 => x"5b900008",  5306 => x"5b9d0004",
     5307 => x"340c0000",  5308 => x"b8205800",  5309 => x"b8407000",
     5310 => x"342f030c",  5311 => x"34300320",  5312 => x"e0000013",
     5313 => x"098d0058",  5314 => x"ba000800",  5315 => x"3403000a",
     5316 => x"35a20110",  5317 => x"b5621000",  5318 => x"f800364b",
     5319 => x"5c20000b",  5320 => x"b56d0800",  5321 => x"b9e01000",
     5322 => x"34030024",  5323 => x"34210144",  5324 => x"f8003666",
     5325 => x"b56d5800",  5326 => x"b9c00800",  5327 => x"3562011c",
     5328 => x"f80003be",  5329 => x"e0000020",  5330 => x"358c0001",
     5331 => x"2d63010c",  5332 => x"486cffed",  5333 => x"34010004",
     5334 => x"54610003",  5335 => x"34630001",  5336 => x"0d63010c",
     5337 => x"2d6d010c",  5338 => x"35620320",  5339 => x"3403000a",
     5340 => x"35adffff",  5341 => x"09ac0058",  5342 => x"35810110",
     5343 => x"b5610800",  5344 => x"f8003652",  5345 => x"b56c0800",
     5346 => x"34030024",  5347 => x"b9e01000",  5348 => x"34210144",
     5349 => x"f800364d",  5350 => x"b56c1000",  5351 => x"b9c00800",
     5352 => x"3442011c",  5353 => x"f80003a5",  5354 => x"78040001",
     5355 => x"b9600800",  5356 => x"34020003",  5357 => x"34030001",
     5358 => x"388441a0",  5359 => x"b9a02800",  5360 => x"fbffed62",
     5361 => x"2b9d0004",  5362 => x"2b8b001c",  5363 => x"2b8c0018",
     5364 => x"2b8d0014",  5365 => x"2b8e0010",  5366 => x"2b8f000c",
     5367 => x"2b900008",  5368 => x"379c001c",  5369 => x"c3a00000",
     5370 => x"4022001e",  5371 => x"34030001",  5372 => x"44430009",
     5373 => x"44400008",  5374 => x"34030002",  5375 => x"5c430008",
     5376 => x"34020012",  5377 => x"58220070",  5378 => x"3402000e",
     5379 => x"58220074",  5380 => x"e0000003",  5381 => x"58200070",
     5382 => x"58200074",  5383 => x"28240070",  5384 => x"2825002c",
     5385 => x"34020000",  5386 => x"b4a42800",  5387 => x"20a30003",
     5388 => x"44600003",  5389 => x"34020004",  5390 => x"c8431000",
     5391 => x"b4a22800",  5392 => x"28260030",  5393 => x"28220074",
     5394 => x"5825003c",  5395 => x"34030000",  5396 => x"b4c23000",
     5397 => x"20c70003",  5398 => x"44e00003",  5399 => x"34030004",
     5400 => x"c8671800",  5401 => x"b4c31800",  5402 => x"c8a42000",
     5403 => x"c8621000",  5404 => x"58230040",  5405 => x"58240034",
     5406 => x"58220038",  5407 => x"c3a00000",  5408 => x"379cfff4",
     5409 => x"5b8b000c",  5410 => x"5b8c0008",  5411 => x"5b9d0004",
     5412 => x"78020001",  5413 => x"384264ac",  5414 => x"28420020",
     5415 => x"b8205800",  5416 => x"44400006",  5417 => x"d8400000",
     5418 => x"b8206000",  5419 => x"34010001",  5420 => x"45810018",
     5421 => x"480c0018",  5422 => x"296102d4",  5423 => x"340c0000",
     5424 => x"44200015",  5425 => x"29610028",  5426 => x"34020000",
     5427 => x"28230018",  5428 => x"b9600800",  5429 => x"d8600000",
     5430 => x"296202d4",  5431 => x"c8220800",  5432 => x"4c200013",
     5433 => x"e000000c",  5434 => x"4162001d",  5435 => x"34010002",
     5436 => x"44410004",  5437 => x"34010006",  5438 => x"59610004",
     5439 => x"e0000006",  5440 => x"34010004",  5441 => x"59610004",
     5442 => x"b9600800",  5443 => x"fbffff5f",  5444 => x"340c0000",
     5445 => x"b9800800",  5446 => x"2b9d0004",  5447 => x"2b8b000c",
     5448 => x"2b8c0008",  5449 => x"379c000c",  5450 => x"c3a00000",
     5451 => x"b9600800",  5452 => x"34020002",  5453 => x"f800078a",
     5454 => x"29610020",  5455 => x"596002d4",  5456 => x"0d60010c",
     5457 => x"2821000c",  5458 => x"4022000e",  5459 => x"340100ff",
     5460 => x"5c41ffe6",  5461 => x"e3ffffeb",  5462 => x"379cfff4",
     5463 => x"5b8b000c",  5464 => x"5b8c0008",  5465 => x"5b9d0004",
     5466 => x"3404003f",  5467 => x"b8205800",  5468 => x"340cffff",
     5469 => x"4c83000e",  5470 => x"fbffff55",  5471 => x"b9600800",
     5472 => x"fbffff42",  5473 => x"b9600800",  5474 => x"f800015a",
     5475 => x"59610004",  5476 => x"78010001",  5477 => x"382164ac",
     5478 => x"28220024",  5479 => x"340c0000",  5480 => x"44400003",
     5481 => x"b9600800",  5482 => x"d8400000",  5483 => x"b9800800",
     5484 => x"2b9d0004",  5485 => x"2b8b000c",  5486 => x"2b8c0008",
     5487 => x"379c000c",  5488 => x"c3a00000",  5489 => x"379cffe0",
     5490 => x"5b8b0014",  5491 => x"5b8c0010",  5492 => x"5b8d000c",
     5493 => x"5b8e0008",  5494 => x"5b9d0004",  5495 => x"b8205800",
     5496 => x"3401002b",  5497 => x"b8407000",  5498 => x"340cffff",
     5499 => x"4c230028",  5500 => x"4161001c",  5501 => x"340c0000",
     5502 => x"20210001",  5503 => x"44200024",  5504 => x"296300ec",
     5505 => x"296200f0",  5506 => x"296100f4",  5507 => x"296500e4",
     5508 => x"296400e8",  5509 => x"5963009c",  5510 => x"596200a0",
     5511 => x"2963031c",  5512 => x"29620318",  5513 => x"596100a4",
     5514 => x"59650094",  5515 => x"356100d0",  5516 => x"59640098",
     5517 => x"f8000485",  5518 => x"41610313",  5519 => x"20210002",
     5520 => x"44200007",  5521 => x"4161001c",  5522 => x"38210002",
     5523 => x"3161001c",  5524 => x"2d61032a",  5525 => x"0d6102ec",
     5526 => x"e000000d",  5527 => x"378d0018",  5528 => x"b9c00800",
     5529 => x"b9a01000",  5530 => x"f80002ed",  5531 => x"4161001c",
     5532 => x"b9a01000",  5533 => x"202100fd",  5534 => x"3161001c",
     5535 => x"35610080",  5536 => x"f80004aa",  5537 => x"b9600800",
     5538 => x"f8000551",  5539 => x"b9800800",  5540 => x"2b9d0004",
     5541 => x"2b8b0014",  5542 => x"2b8c0010",  5543 => x"2b8d000c",
     5544 => x"2b8e0008",  5545 => x"379c0020",  5546 => x"c3a00000",
     5547 => x"379cffe4",  5548 => x"5b8b0010",  5549 => x"5b8c000c",
     5550 => x"5b8d0008",  5551 => x"5b9d0004",  5552 => x"b8205800",
     5553 => x"b8400800",  5554 => x"3402002b",  5555 => x"3404ffff",
     5556 => x"4c430031",  5557 => x"4162001c",  5558 => x"20430001",
     5559 => x"5c600004",  5560 => x"78010001",  5561 => x"382141c0",
     5562 => x"e0000005",  5563 => x"20420002",  5564 => x"5c400007",
     5565 => x"78010001",  5566 => x"382141fc",  5567 => x"78020001",
     5568 => x"384259f8",  5569 => x"f8001bbe",  5570 => x"e0000022",
     5571 => x"2d6402ec",  5572 => x"2d63032a",  5573 => x"44830007",
     5574 => x"78010001",  5575 => x"78020001",  5576 => x"384259f8",
     5577 => x"38214234",  5578 => x"f8001bb5",  5579 => x"e0000019",
     5580 => x"378d0014",  5581 => x"b9a01000",  5582 => x"f80002ec",
     5583 => x"4161001c",  5584 => x"356c0080",  5585 => x"b9a01000",
     5586 => x"202100fd",  5587 => x"3161001c",  5588 => x"b9800800",
     5589 => x"f8000475",  5590 => x"78030001",  5591 => x"386364ac",
     5592 => x"28640028",  5593 => x"44800009",  5594 => x"b9600800",
     5595 => x"b9801000",  5596 => x"356300d0",  5597 => x"d8800000",
     5598 => x"b8202000",  5599 => x"34010001",  5600 => x"44810004",
     5601 => x"48040004",  5602 => x"b9600800",  5603 => x"f8000510",
     5604 => x"34040000",  5605 => x"b8800800",  5606 => x"2b9d0004",
     5607 => x"2b8b0010",  5608 => x"2b8c000c",  5609 => x"2b8d0008",
     5610 => x"379c001c",  5611 => x"c3a00000",  5612 => x"379cfff0",
     5613 => x"5b8b0010",  5614 => x"5b8c000c",  5615 => x"5b8d0008",
     5616 => x"5b9d0004",  5617 => x"b8406800",  5618 => x"3402003f",
     5619 => x"b8205800",  5620 => x"340cffff",  5621 => x"4c430013",
     5622 => x"78040001",  5623 => x"34030002",  5624 => x"38844274",
     5625 => x"34020003",  5626 => x"fbffec58",  5627 => x"b9a01000",
     5628 => x"b9600800",  5629 => x"fbfffeb6",  5630 => x"b9600800",
     5631 => x"f80000bd",  5632 => x"59610004",  5633 => x"78010001",
     5634 => x"382164ac",  5635 => x"28220024",  5636 => x"340c0000",
     5637 => x"44400003",  5638 => x"b9600800",  5639 => x"d8400000",
     5640 => x"b9800800",  5641 => x"2b9d0004",  5642 => x"2b8b0010",
     5643 => x"2b8c000c",  5644 => x"2b8d0008",  5645 => x"379c0010",
     5646 => x"c3a00000",  5647 => x"34010000",  5648 => x"c3a00000",
     5649 => x"379cfffc",  5650 => x"5b9d0004",  5651 => x"34030008",
     5652 => x"f80034fd",  5653 => x"2b9d0004",  5654 => x"379c0004",
     5655 => x"c3a00000",  5656 => x"379cffe0",  5657 => x"5b8b0020",
     5658 => x"5b8c001c",  5659 => x"5b8d0018",  5660 => x"5b8e0014",
     5661 => x"5b8f0010",  5662 => x"5b90000c",  5663 => x"5b910008",
     5664 => x"5b9d0004",  5665 => x"780e0001",  5666 => x"39ce5a18",
     5667 => x"78040001",  5668 => x"b8406800",  5669 => x"b8606000",
     5670 => x"34020003",  5671 => x"34030002",  5672 => x"3884461c",
     5673 => x"b9c02800",  5674 => x"b8207800",  5675 => x"35b10021",
     5676 => x"fbffec26",  5677 => x"35900021",  5678 => x"ba200800",
     5679 => x"ba001000",  5680 => x"fbffffe1",  5681 => x"5c200033",
     5682 => x"2d81002a",  5683 => x"2dab002a",  5684 => x"c9615800",
     5685 => x"35620001",  5686 => x"34010002",  5687 => x"54410043",
     5688 => x"29e20020",  5689 => x"34030001",  5690 => x"35a10048",
     5691 => x"28420014",  5692 => x"5d63000b",  5693 => x"fbffffd4",
     5694 => x"5c20003c",  5695 => x"78040001",  5696 => x"b9e00800",
     5697 => x"34020003",  5698 => x"34030001",  5699 => x"388442a4",
     5700 => x"b9c02800",  5701 => x"3406008f",  5702 => x"e000000e",
     5703 => x"3403ffff",  5704 => x"358c0048",  5705 => x"5d63000e",
     5706 => x"b9800800",  5707 => x"fbffffc6",  5708 => x"5c20002e",
     5709 => x"78040001",  5710 => x"b9e00800",  5711 => x"34020003",
     5712 => x"34030001",  5713 => x"388442a4",  5714 => x"b9c02800",
     5715 => x"34060098",  5716 => x"fbffebfe",  5717 => x"340b0000",
     5718 => x"e0000024",  5719 => x"b9801000",  5720 => x"fbffffb9",
     5721 => x"b8205800",  5722 => x"5c200020",  5723 => x"78040001",
     5724 => x"b9e00800",  5725 => x"34020003",  5726 => x"34030001",
     5727 => x"388442b4",  5728 => x"b9c02800",  5729 => x"340600a0",
     5730 => x"fbffebf0",  5731 => x"e0000017",  5732 => x"41ab001a",
     5733 => x"4181001a",  5734 => x"5d61000e",  5735 => x"41ab001c",
     5736 => x"4181001c",  5737 => x"5d61000b",  5738 => x"41ab001d",
     5739 => x"4181001d",  5740 => x"5d610008",  5741 => x"2da2001e",
     5742 => x"2d81001e",  5743 => x"340b0000",  5744 => x"5c41000a",
     5745 => x"41ab0020",  5746 => x"41810020",  5747 => x"45610003",
     5748 => x"c9615800",  5749 => x"e0000005",  5750 => x"ba200800",
     5751 => x"ba001000",  5752 => x"fbffff99",  5753 => x"b8205800",
     5754 => x"b9600800",  5755 => x"2b9d0004",  5756 => x"2b8b0020",
     5757 => x"2b8c001c",  5758 => x"2b8d0018",  5759 => x"2b8e0014",
     5760 => x"2b8f0010",  5761 => x"2b90000c",  5762 => x"2b910008",
     5763 => x"379c0020",  5764 => x"c3a00000",  5765 => x"379cfffc",
     5766 => x"5b9d0004",  5767 => x"34020000",  5768 => x"34030014",
     5769 => x"f8003527",  5770 => x"2b9d0004",  5771 => x"379c0004",
     5772 => x"c3a00000",  5773 => x"379cfff0",  5774 => x"5b8b0010",
     5775 => x"5b8c000c",  5776 => x"5b8d0008",  5777 => x"5b9d0004",
     5778 => x"b8206800",  5779 => x"28210020",  5780 => x"282c0014",
     5781 => x"282b000c",  5782 => x"28210010",  5783 => x"0c200000",
     5784 => x"34210004",  5785 => x"fbffffec",  5786 => x"29a10020",
     5787 => x"28210010",  5788 => x"34210018",  5789 => x"fbffffe8",
     5790 => x"b9800800",  5791 => x"34020000",  5792 => x"34030020",
     5793 => x"f800350f",  5794 => x"29610004",  5795 => x"3402ffa0",
     5796 => x"59810000",  5797 => x"29610008",  5798 => x"59810004",
     5799 => x"29610004",  5800 => x"59810010",  5801 => x"29610008",
     5802 => x"59810014",  5803 => x"2d61000e",  5804 => x"0d810018",
     5805 => x"2d610010",  5806 => x"0d81001a",  5807 => x"41610012",
     5808 => x"3181001c",  5809 => x"41610013",  5810 => x"3181001d",
     5811 => x"29a10020",  5812 => x"28210018",  5813 => x"3022001c",
     5814 => x"2b9d0004",  5815 => x"2b8b0010",  5816 => x"2b8c000c",
     5817 => x"2b8d0008",  5818 => x"379c0010",  5819 => x"c3a00000",
     5820 => x"379cff8c",  5821 => x"5b8b0018",  5822 => x"5b8c0014",
     5823 => x"5b8d0010",  5824 => x"5b8e000c",  5825 => x"5b8f0008",
     5826 => x"5b9d0004",  5827 => x"2c22010c",  5828 => x"b8205800",
     5829 => x"340d0000",  5830 => x"340c0001",  5831 => x"5c400014",
     5832 => x"28230000",  5833 => x"b8406800",  5834 => x"34020006",
     5835 => x"5c620010",  5836 => x"fbffffc1",  5837 => x"29610000",
     5838 => x"e0000105",  5839 => x"09820058",  5840 => x"09a30058",
     5841 => x"b9600800",  5842 => x"34420110",  5843 => x"34630110",
     5844 => x"b5621000",  5845 => x"b5631800",  5846 => x"fbffff42",
     5847 => x"48010002",  5848 => x"e0000002",  5849 => x"b9806800",
     5850 => x"358c0001",  5851 => x"2d66010c",  5852 => x"48ccfff3",
     5853 => x"78040001",  5854 => x"b9600800",  5855 => x"34020003",
     5856 => x"34030001",  5857 => x"388442c4",  5858 => x"b9a02800",
     5859 => x"fbffeb6f",  5860 => x"1d61010e",  5861 => x"442d0022",
     5862 => x"0d6d010e",  5863 => x"296c0020",  5864 => x"340f0000",
     5865 => x"340e0001",  5866 => x"e0000015",  5867 => x"29820000",
     5868 => x"09c10374",  5869 => x"b4410800",  5870 => x"2c23010c",
     5871 => x"4460000f",  5872 => x"09e40374",  5873 => x"1c23010e",
     5874 => x"b4442000",  5875 => x"1c82010e",  5876 => x"08630058",
     5877 => x"08420058",  5878 => x"34630110",  5879 => x"b4231800",
     5880 => x"34420110",  5881 => x"b4821000",  5882 => x"fbffff1e",
     5883 => x"48010002",  5884 => x"e0000002",  5885 => x"b9c07800",
     5886 => x"35ce0001",  5887 => x"2981000c",  5888 => x"2c21000c",
     5889 => x"482effea",  5890 => x"2981001c",  5891 => x"442f0004",
     5892 => x"34010001",  5893 => x"598f001c",  5894 => x"59810020",
     5895 => x"4162001d",  5896 => x"34010002",  5897 => x"44410063",
     5898 => x"2d61010c",  5899 => x"5c200004",  5900 => x"29620000",
     5901 => x"34010004",  5902 => x"444100c5",  5903 => x"29610020",
     5904 => x"09ac0058",  5905 => x"2821000c",  5906 => x"4023000a",
     5907 => x"4022000b",  5908 => x"40290004",  5909 => x"40280005",
     5910 => x"40270006",  5911 => x"40260007",  5912 => x"40250008",
     5913 => x"40240009",  5914 => x"33830047",  5915 => x"33890041",
     5916 => x"33880042",  5917 => x"33870043",  5918 => x"33860044",
     5919 => x"33850045",  5920 => x"33840046",  5921 => x"33820048",
     5922 => x"2c22000e",  5923 => x"35830110",  5924 => x"b5631800",
     5925 => x"0f82003c",  5926 => x"2c220010",  5927 => x"0f82003e",
     5928 => x"40220012",  5929 => x"3382003a",  5930 => x"40220013",
     5931 => x"0f80004a",  5932 => x"33820040",  5933 => x"28220004",
     5934 => x"5b820068",  5935 => x"28210008",  5936 => x"37820020",
     5937 => x"5b81006c",  5938 => x"b9600800",  5939 => x"fbfffee5",
     5940 => x"4162001d",  5941 => x"34030001",  5942 => x"44430029",
     5943 => x"29620020",  5944 => x"78050001",  5945 => x"38a55a28",
     5946 => x"2844000c",  5947 => x"1086000e",  5948 => x"48060004",
     5949 => x"48010023",  5950 => x"5c200019",  5951 => x"e0000006",
     5952 => x"48010020",  5953 => x"44200004",  5954 => x"2c81000c",
     5955 => x"5c23000a",  5956 => x"e0000028",  5957 => x"78040001",
     5958 => x"b9600800",  5959 => x"34020003",  5960 => x"34030001",
     5961 => x"388442e4",  5962 => x"fbffeb08",  5963 => x"34010002",
     5964 => x"e0000087",  5965 => x"29630338",  5966 => x"2841001c",
     5967 => x"4461001d",  5968 => x"b56c1000",  5969 => x"37810041",
     5970 => x"34420131",  5971 => x"5b85001c",  5972 => x"fbfffebd",
     5973 => x"2b85001c",  5974 => x"5c20000c",  5975 => x"78040001",
     5976 => x"b9600800",  5977 => x"34020003",  5978 => x"34030001",
     5979 => x"388442f0",  5980 => x"fbffeaf6",  5981 => x"34010007",
     5982 => x"e0000075",  5983 => x"4c200003",  5984 => x"b9600800",
     5985 => x"fbffff2c",  5986 => x"78040001",  5987 => x"78050001",
     5988 => x"b9600800",  5989 => x"34020003",  5990 => x"34030001",
     5991 => x"38844300",  5992 => x"38a55a28",  5993 => x"fbffeae9",
     5994 => x"34010006",  5995 => x"e0000068",  5996 => x"09a30058",
     5997 => x"29620020",  5998 => x"b5631800",  5999 => x"2c64013a",
     6000 => x"284c0018",  6001 => x"28410014",  6002 => x"28420010",
     6003 => x"34840001",  6004 => x"0c440000",  6005 => x"34620150",
     6006 => x"28450008",  6007 => x"2844000c",  6008 => x"58250000",
     6009 => x"58240004",  6010 => x"2c420010",  6011 => x"0c220008",
     6012 => x"34620128",  6013 => x"404e0009",  6014 => x"4045000f",
     6015 => x"40440010",  6016 => x"404a000a",  6017 => x"4049000b",
     6018 => x"4048000c",  6019 => x"4047000d",  6020 => x"4046000e",
     6021 => x"302e0010",  6022 => x"30250016",  6023 => x"302a0011",
     6024 => x"30290012",  6025 => x"30280013",  6026 => x"30270014",
     6027 => x"30260015",  6028 => x"30240017",  6029 => x"28440004",
     6030 => x"346e0120",  6031 => x"58240018",  6032 => x"41c4000a",
     6033 => x"3024001c",  6034 => x"40420008",  6035 => x"3022001d",
     6036 => x"4061013c",  6037 => x"3181001c",  6038 => x"1dc50008",
     6039 => x"1d810000",  6040 => x"4425000e",  6041 => x"78040001",
     6042 => x"b9600800",  6043 => x"34020003",  6044 => x"34030001",
     6045 => x"3884430c",  6046 => x"fbffeab4",  6047 => x"2dc10008",
     6048 => x"34020000",  6049 => x"0d810000",  6050 => x"29610028",
     6051 => x"28230004",  6052 => x"b9600800",  6053 => x"d8600000",
     6054 => x"09ad0058",  6055 => x"b56d0800",  6056 => x"34210141",
     6057 => x"4022000b",  6058 => x"20420004",  6059 => x"7c420000",
     6060 => x"59820004",  6061 => x"4022000b",  6062 => x"20420002",
     6063 => x"7c420000",  6064 => x"59820008",  6065 => x"4022000b",
     6066 => x"20420001",  6067 => x"5982000c",  6068 => x"4022000b",
     6069 => x"20420010",  6070 => x"7c420000",  6071 => x"59820010",
     6072 => x"4022000b",  6073 => x"20420020",  6074 => x"7c420000",
     6075 => x"59820014",  6076 => x"4021000b",  6077 => x"20210008",
     6078 => x"7c210000",  6079 => x"59810018",  6080 => x"78010001",
     6081 => x"382164ac",  6082 => x"2824001c",  6083 => x"44800007",
     6084 => x"b56d1000",  6085 => x"b8406800",  6086 => x"b9600800",
     6087 => x"34420144",  6088 => x"35a3011c",  6089 => x"d8800000",
     6090 => x"78040001",  6091 => x"78050001",  6092 => x"b9600800",
     6093 => x"34020003",  6094 => x"34030001",  6095 => x"38844320",
     6096 => x"38a55a28",  6097 => x"fbffea81",  6098 => x"34010009",
     6099 => x"2b9d0004",  6100 => x"2b8b0018",  6101 => x"2b8c0014",
     6102 => x"2b8d0010",  6103 => x"2b8e000c",  6104 => x"2b8f0008",
     6105 => x"379c0074",  6106 => x"c3a00000",  6107 => x"379cffec",
     6108 => x"5b8b0014",  6109 => x"5b8c0010",  6110 => x"5b8d000c",
     6111 => x"5b8e0008",  6112 => x"5b9d0004",  6113 => x"b8406000",
     6114 => x"28220024",  6115 => x"b8607000",  6116 => x"28230070",
     6117 => x"2847000c",  6118 => x"28220034",  6119 => x"b8806800",
     6120 => x"b5831800",  6121 => x"342400f8",  6122 => x"b9a02800",
     6123 => x"34060000",  6124 => x"b8205800",  6125 => x"d8e00000",
     6126 => x"78070001",  6127 => x"38e764e4",  6128 => x"3dc20002",
     6129 => x"4c2c000c",  6130 => x"b4e23800",  6131 => x"28e50000",
     6132 => x"78040001",  6133 => x"b9600800",  6134 => x"34020005",
     6135 => x"34030001",  6136 => x"38843f58",  6137 => x"b9c03000",
     6138 => x"fbffea58",  6139 => x"3401ffff",  6140 => x"e0000014",
     6141 => x"b4e24000",  6142 => x"296600f8",  6143 => x"296700fc",
     6144 => x"29080000",  6145 => x"78040001",  6146 => x"b9600800",
     6147 => x"34020005",  6148 => x"34030001",  6149 => x"38843f78",
     6150 => x"b9802800",  6151 => x"fbffea4b",  6152 => x"34010001",
     6153 => x"5da10003",  6154 => x"29620104",  6155 => x"44400005",
     6156 => x"2961036c",  6157 => x"34210001",  6158 => x"5961036c",
     6159 => x"34010000",  6160 => x"2b9d0004",  6161 => x"2b8b0014",
     6162 => x"2b8c0010",  6163 => x"2b8d000c",  6164 => x"2b8e0008",
     6165 => x"379c0014",  6166 => x"c3a00000",  6167 => x"379cfff0",
     6168 => x"5b8b0010",  6169 => x"5b8c000c",  6170 => x"5b8d0008",
     6171 => x"5b9d0004",  6172 => x"b8205800",  6173 => x"40410000",
     6174 => x"b8406000",  6175 => x"34030002",  6176 => x"00210004",
     6177 => x"356d0320",  6178 => x"3161030c",  6179 => x"40410000",
     6180 => x"2021000f",  6181 => x"3161030d",  6182 => x"40410001",
     6183 => x"2021000f",  6184 => x"3161030e",  6185 => x"2c410002",
     6186 => x"0d610310",  6187 => x"40410004",  6188 => x"34420006",
     6189 => x"31610312",  6190 => x"35610313",  6191 => x"f8003303",
     6192 => x"35820008",  6193 => x"34030004",  6194 => x"3561031c",
     6195 => x"f80032ff",  6196 => x"3582000c",  6197 => x"34030004",
     6198 => x"35610318",  6199 => x"f80032fb",  6200 => x"35820014",
     6201 => x"34030008",  6202 => x"b9a00800",  6203 => x"f80032f7",
     6204 => x"2d81001c",  6205 => x"296202c8",  6206 => x"34030008",
     6207 => x"0d610328",  6208 => x"2d81001e",  6209 => x"0d61032a",
     6210 => x"41810020",  6211 => x"3161032c",  6212 => x"41810021",
     6213 => x"3161032d",  6214 => x"b9a00800",  6215 => x"f80032ca",
     6216 => x"3403ffff",  6217 => x"44200015",  6218 => x"29610020",
     6219 => x"28210014",  6220 => x"2c220008",  6221 => x"4440000a",
     6222 => x"b9a01000",  6223 => x"34030008",  6224 => x"f80032c1",
     6225 => x"5c200009",  6226 => x"29610020",  6227 => x"28210014",
     6228 => x"2c220008",  6229 => x"2d610328",  6230 => x"5c410004",
     6231 => x"4161001c",  6232 => x"38210001",  6233 => x"e0000003",
     6234 => x"4161001c",  6235 => x"202100fe",  6236 => x"3161001c",
     6237 => x"34030000",  6238 => x"b8600800",  6239 => x"2b9d0004",
     6240 => x"2b8b0010",  6241 => x"2b8c000c",  6242 => x"2b8d0008",
     6243 => x"379c0010",  6244 => x"c3a00000",  6245 => x"379cfff4",
     6246 => x"5b8b000c",  6247 => x"5b8c0008",  6248 => x"5b9d0004",
     6249 => x"30400000",  6250 => x"b8206000",  6251 => x"282102c8",
     6252 => x"b8405800",  6253 => x"34030008",  6254 => x"4021000e",
     6255 => x"30410001",  6256 => x"29810020",  6257 => x"2821000c",
     6258 => x"40210014",  6259 => x"30410004",  6260 => x"34010002",
     6261 => x"30410006",  6262 => x"34410008",  6263 => x"34020000",
     6264 => x"f8003338",  6265 => x"298202c8",  6266 => x"35610014",
     6267 => x"34030008",  6268 => x"f80032b6",  6269 => x"298102c8",
     6270 => x"2c210008",  6271 => x"0d61001c",  6272 => x"3401007f",
     6273 => x"31610021",  6274 => x"2b9d0004",  6275 => x"2b8b000c",
     6276 => x"2b8c0008",  6277 => x"379c000c",  6278 => x"c3a00000",
     6279 => x"2c230022",  6280 => x"0c430004",  6281 => x"28230024",
     6282 => x"58430000",  6283 => x"28210028",  6284 => x"58410008",
     6285 => x"c3a00000",  6286 => x"379cfff4",  6287 => x"5b8b000c",
     6288 => x"5b8c0008",  6289 => x"5b9d0004",  6290 => x"b8205800",
     6291 => x"2c210022",  6292 => x"b8406000",  6293 => x"34030008",
     6294 => x"0c410004",  6295 => x"29610024",  6296 => x"58410000",
     6297 => x"29610028",  6298 => x"58410008",  6299 => x"2d61002c",
     6300 => x"0c41000c",  6301 => x"4161002f",  6302 => x"3041000e",
     6303 => x"41610030",  6304 => x"30410010",  6305 => x"41610031",
     6306 => x"30410011",  6307 => x"2d610032",  6308 => x"0c410012",
     6309 => x"41610034",  6310 => x"30410014",  6311 => x"34410015",
     6312 => x"35620035",  6313 => x"f8003289",  6314 => x"2d61003d",
     6315 => x"0d81001e",  6316 => x"4161003f",  6317 => x"31810020",
     6318 => x"78010001",  6319 => x"382164ac",  6320 => x"28230030",
     6321 => x"44600004",  6322 => x"b9600800",  6323 => x"b9801000",
     6324 => x"d8600000",  6325 => x"2b9d0004",  6326 => x"2b8b000c",
     6327 => x"2b8c0008",  6328 => x"379c000c",  6329 => x"c3a00000",
     6330 => x"2c230022",  6331 => x"0c430004",  6332 => x"28230024",
     6333 => x"58430000",  6334 => x"28210028",  6335 => x"58410008",
     6336 => x"c3a00000",  6337 => x"379cfff4",  6338 => x"5b8b000c",
     6339 => x"5b8c0008",  6340 => x"5b9d0004",  6341 => x"b8205800",
     6342 => x"2c210022",  6343 => x"b8406000",  6344 => x"34030008",
     6345 => x"0c410004",  6346 => x"29610024",  6347 => x"58410000",
     6348 => x"29610028",  6349 => x"58410008",  6350 => x"3441000c",
     6351 => x"3562002c",  6352 => x"f8003262",  6353 => x"2d610034",
     6354 => x"0d810014",  6355 => x"2b9d0004",  6356 => x"2b8b000c",
     6357 => x"2b8c0008",  6358 => x"379c000c",  6359 => x"c3a00000",
     6360 => x"379cfff4",  6361 => x"5b8b000c",  6362 => x"5b8c0008",
     6363 => x"5b9d0004",  6364 => x"282b003c",  6365 => x"b8206000",
     6366 => x"34020000",  6367 => x"41610000",  6368 => x"3403000a",
     6369 => x"202100f0",  6370 => x"3821000b",  6371 => x"31610000",
     6372 => x"34010040",  6373 => x"0d610002",  6374 => x"2d810306",
     6375 => x"34210001",  6376 => x"2021ffff",  6377 => x"0d810306",
     6378 => x"0d61001e",  6379 => x"34010005",  6380 => x"31610020",
     6381 => x"298102c8",  6382 => x"4021000b",  6383 => x"31610021",
     6384 => x"35610022",  6385 => x"f80032bf",  6386 => x"29810020",
     6387 => x"34030008",  6388 => x"28220018",  6389 => x"28210014",
     6390 => x"2c420000",  6391 => x"0d62002c",  6392 => x"4021001c",
     6393 => x"3161002f",  6394 => x"29810020",  6395 => x"28210014",
     6396 => x"40210018",  6397 => x"31610030",  6398 => x"29810020",
     6399 => x"28210014",  6400 => x"40210019",  6401 => x"31610031",
     6402 => x"29810020",  6403 => x"28210014",  6404 => x"2c22001a",
     6405 => x"0d620032",  6406 => x"4021001d",  6407 => x"31610034",
     6408 => x"29810020",  6409 => x"28220014",  6410 => x"35610035",
     6411 => x"34420010",  6412 => x"f8003226",  6413 => x"29810020",
     6414 => x"28220010",  6415 => x"28210018",  6416 => x"2c420000",
     6417 => x"0d62003d",  6418 => x"4021001c",  6419 => x"34020040",
     6420 => x"3161003f",  6421 => x"78010001",  6422 => x"382164ac",
     6423 => x"2823002c",  6424 => x"44600004",  6425 => x"b9800800",
     6426 => x"d8600000",  6427 => x"b8201000",  6428 => x"b9800800",
     6429 => x"3403000b",  6430 => x"34040000",  6431 => x"fbfffebc",
     6432 => x"2b9d0004",  6433 => x"2b8b000c",  6434 => x"2b8c0008",
     6435 => x"379c000c",  6436 => x"c3a00000",  6437 => x"379cffc8",
     6438 => x"5b8b0018",  6439 => x"5b8c0014",  6440 => x"5b8d0010",
     6441 => x"5b8e000c",  6442 => x"5b8f0008",  6443 => x"5b9d0004",
     6444 => x"28220028",  6445 => x"378c001c",  6446 => x"b8205800",
     6447 => x"28430000",  6448 => x"b9801000",  6449 => x"378f0030",
     6450 => x"d8600000",  6451 => x"b9800800",  6452 => x"b9e01000",
     6453 => x"f8000103",  6454 => x"296c003c",  6455 => x"340efff0",
     6456 => x"340d002c",  6457 => x"41810000",  6458 => x"0d8d0002",
     6459 => x"34020000",  6460 => x"a02e0800",  6461 => x"31810000",
     6462 => x"2d6102f0",  6463 => x"34030008",  6464 => x"34210001",
     6465 => x"2021ffff",  6466 => x"0d6102f0",  6467 => x"31800020",
     6468 => x"0d81001e",  6469 => x"296102c8",  6470 => x"4021000d",
     6471 => x"31810021",  6472 => x"35810008",  6473 => x"f8003267",
     6474 => x"2f810034",  6475 => x"3402002c",  6476 => x"34030000",
     6477 => x"0d810022",  6478 => x"2b810030",  6479 => x"34040001",
     6480 => x"59810024",  6481 => x"2b810038",  6482 => x"59810028",
     6483 => x"b9600800",  6484 => x"fbfffe87",  6485 => x"5c200023",
     6486 => x"29610020",  6487 => x"356c00f8",  6488 => x"b9801000",
     6489 => x"28230008",  6490 => x"b9800800",  6491 => x"34630018",
     6492 => x"f8000101",  6493 => x"b9e01000",  6494 => x"b9800800",
     6495 => x"f80000d9",  6496 => x"2961003c",  6497 => x"34030008",
     6498 => x"34040000",  6499 => x"40220000",  6500 => x"0c2d0002",
     6501 => x"a04e7000",  6502 => x"39ce0008",  6503 => x"302e0000",
     6504 => x"2d6202f0",  6505 => x"0c22001e",  6506 => x"34020002",
     6507 => x"30220020",  6508 => x"296202c8",  6509 => x"4042000d",
     6510 => x"30220021",  6511 => x"2f820034",  6512 => x"0c220022",
     6513 => x"2b820030",  6514 => x"58220024",  6515 => x"2b820038",
     6516 => x"58220028",  6517 => x"b9600800",  6518 => x"3402002c",
     6519 => x"fbfffe64",  6520 => x"2b9d0004",  6521 => x"2b8b0018",
     6522 => x"2b8c0014",  6523 => x"2b8d0010",  6524 => x"2b8e000c",
     6525 => x"2b8f0008",  6526 => x"379c0038",  6527 => x"c3a00000",
     6528 => x"379cffd4",  6529 => x"5b8b000c",  6530 => x"5b8c0008",
     6531 => x"5b9d0004",  6532 => x"28220028",  6533 => x"378b0010",
     6534 => x"b8206000",  6535 => x"28430000",  6536 => x"b9601000",
     6537 => x"d8600000",  6538 => x"37820024",  6539 => x"b9600800",
     6540 => x"f80000ac",  6541 => x"298b003c",  6542 => x"34020000",
     6543 => x"34030008",  6544 => x"41610000",  6545 => x"202100f0",
     6546 => x"38210001",  6547 => x"31610000",  6548 => x"3401002c",
     6549 => x"0d610002",  6550 => x"2d8102f2",  6551 => x"34210001",
     6552 => x"2021ffff",  6553 => x"0d8102f2",  6554 => x"0d61001e",
     6555 => x"34010001",  6556 => x"31610020",  6557 => x"3401007f",
     6558 => x"31610021",  6559 => x"35610008",  6560 => x"f8003210",
     6561 => x"2f810028",  6562 => x"3402002c",  6563 => x"34030001",
     6564 => x"0d610022",  6565 => x"2b810024",  6566 => x"34040001",
     6567 => x"59610024",  6568 => x"2b81002c",  6569 => x"59610028",
     6570 => x"b9800800",  6571 => x"fbfffe30",  6572 => x"2b9d0004",
     6573 => x"2b8b000c",  6574 => x"2b8c0008",  6575 => x"379c002c",
     6576 => x"c3a00000",  6577 => x"379cffe8",  6578 => x"5b8b000c",
     6579 => x"5b8c0008",  6580 => x"5b9d0004",  6581 => x"b8206000",
     6582 => x"b8400800",  6583 => x"37820010",  6584 => x"f8000080",
     6585 => x"298b003c",  6586 => x"34020000",  6587 => x"34030008",
     6588 => x"41610000",  6589 => x"202100f0",  6590 => x"38210009",
     6591 => x"31610000",  6592 => x"34010036",  6593 => x"0d610002",
     6594 => x"41810312",  6595 => x"31610004",  6596 => x"35610008",
     6597 => x"f80031eb",  6598 => x"2981031c",  6599 => x"35820320",
     6600 => x"34030008",  6601 => x"59610008",  6602 => x"29810318",
     6603 => x"5961000c",  6604 => x"2d81032a",  6605 => x"0d61001e",
     6606 => x"34010003",  6607 => x"31610020",  6608 => x"298102c8",
     6609 => x"4021000a",  6610 => x"31610021",  6611 => x"2f810014",
     6612 => x"0d610022",  6613 => x"2b810010",  6614 => x"59610024",
     6615 => x"2b810018",  6616 => x"59610028",  6617 => x"3561002c",
     6618 => x"f8003158",  6619 => x"2d810328",  6620 => x"34020036",
     6621 => x"34030009",  6622 => x"0d610034",  6623 => x"34040000",
     6624 => x"b9800800",  6625 => x"fbfffdfa",  6626 => x"2b9d0004",
     6627 => x"2b8b000c",  6628 => x"2b8c0008",  6629 => x"379c0018",
     6630 => x"c3a00000",  6631 => x"379cfff0",  6632 => x"5b8b0010",
     6633 => x"5b8c000c",  6634 => x"5b8d0008",  6635 => x"5b9d0004",
     6636 => x"78030001",  6637 => x"282d0004",  6638 => x"38635748",
     6639 => x"28620000",  6640 => x"b8205800",  6641 => x"b9a00800",
     6642 => x"f8003092",  6643 => x"78030001",  6644 => x"296c0000",
     6645 => x"38635748",  6646 => x"28620000",  6647 => x"b42c6000",
     6648 => x"596c0000",  6649 => x"b9a00800",  6650 => x"f80030b7",
     6651 => x"59610004",  6652 => x"4c0c0007",  6653 => x"4c20000f",
     6654 => x"358cffff",  6655 => x"78030001",  6656 => x"596c0000",
     6657 => x"38635748",  6658 => x"e0000007",  6659 => x"45800009",
     6660 => x"4c010008",  6661 => x"358c0001",  6662 => x"78030001",
     6663 => x"596c0000",  6664 => x"3863575c",  6665 => x"28620000",
     6666 => x"b4220800",  6667 => x"59610004",  6668 => x"2b9d0004",
     6669 => x"2b8b0010",  6670 => x"2b8c000c",  6671 => x"2b8d0008",
     6672 => x"379c0010",  6673 => x"c3a00000",  6674 => x"379cffe8",
     6675 => x"5b8b0008",  6676 => x"5b9d0004",  6677 => x"5b82000c",
     6678 => x"5b830010",  6679 => x"5b830014",  6680 => x"5b820018",
     6681 => x"b8205800",  6682 => x"4c600006",  6683 => x"78010001",
     6684 => x"78020001",  6685 => x"382143a0",  6686 => x"38425a3c",
     6687 => x"f8001760",  6688 => x"2b810018",  6689 => x"38028000",
     6690 => x"2b830014",  6691 => x"b4221000",  6692 => x"f4220800",
     6693 => x"00420010",  6694 => x"b4230800",  6695 => x"3c230010",
     6696 => x"00210010",  6697 => x"b8431000",  6698 => x"78030001",
     6699 => x"38635748",  6700 => x"5b820018",  6701 => x"28620000",
     6702 => x"5b810014",  6703 => x"37810014",  6704 => x"fbffec4a",
     6705 => x"59610004",  6706 => x"2b810018",  6707 => x"59610000",
     6708 => x"2b9d0004",  6709 => x"2b8b0008",  6710 => x"379c0018",
     6711 => x"c3a00000",  6712 => x"379cfffc",  6713 => x"5b9d0004",
     6714 => x"28230000",  6715 => x"48030003",  6716 => x"28210004",
     6717 => x"4c200006",  6718 => x"78010001",  6719 => x"382143cc",
     6720 => x"f800173f",  6721 => x"3401ffff",  6722 => x"e0000005",
     6723 => x"58410008",  6724 => x"58430000",  6725 => x"0c400004",
     6726 => x"34010000",  6727 => x"2b9d0004",  6728 => x"379c0004",
     6729 => x"c3a00000",  6730 => x"379cfffc",  6731 => x"5b9d0004",
     6732 => x"78050001",  6733 => x"38a55760",  6734 => x"28430000",
     6735 => x"28a40000",  6736 => x"54640006",  6737 => x"28420008",
     6738 => x"58230000",  6739 => x"58220004",  6740 => x"34010000",
     6741 => x"e0000005",  6742 => x"78010001",  6743 => x"38214408",
     6744 => x"f8001727",  6745 => x"3401ffff",  6746 => x"2b9d0004",
     6747 => x"379c0004",  6748 => x"c3a00000",  6749 => x"379cfffc",
     6750 => x"5b9d0004",  6751 => x"28660000",  6752 => x"28450000",
     6753 => x"28630004",  6754 => x"28420004",  6755 => x"b4c52800",
     6756 => x"58250000",  6757 => x"b4621000",  6758 => x"58220004",
     6759 => x"fbffff80",  6760 => x"2b9d0004",  6761 => x"379c0004",
     6762 => x"c3a00000",  6763 => x"379cfffc",  6764 => x"5b9d0004",
     6765 => x"28460000",  6766 => x"28650000",  6767 => x"c8c52800",
     6768 => x"58250000",  6769 => x"28450004",  6770 => x"28620004",
     6771 => x"c8a21000",  6772 => x"58220004",  6773 => x"fbffff72",
     6774 => x"2b9d0004",  6775 => x"379c0004",  6776 => x"c3a00000",
     6777 => x"379cfffc",  6778 => x"5b9d0004",  6779 => x"78040001",
     6780 => x"38845764",  6781 => x"28230000",  6782 => x"28820000",
     6783 => x"a0621000",  6784 => x"4c400005",  6785 => x"3442ffff",
     6786 => x"3404fffe",  6787 => x"b8441000",  6788 => x"34420001",
     6789 => x"78050001",  6790 => x"38a55748",  6791 => x"28a40000",
     6792 => x"88441000",  6793 => x"28240004",  6794 => x"b4441000",
     6795 => x"0064001f",  6796 => x"b4831800",  6797 => x"14630001",
     6798 => x"58230000",  6799 => x"0043001f",  6800 => x"b4621000",
     6801 => x"14420001",  6802 => x"58220004",  6803 => x"fbffff54",
     6804 => x"2b9d0004",  6805 => x"379c0004",  6806 => x"c3a00000",
     6807 => x"379cfff8",  6808 => x"5b8b0008",  6809 => x"5b9d0004",
     6810 => x"28250000",  6811 => x"78030001",  6812 => x"b8201000",
     6813 => x"38634458",  6814 => x"4805000a",  6815 => x"78030001",
     6816 => x"38634c00",  6817 => x"5ca00007",  6818 => x"28210004",
     6819 => x"78030001",  6820 => x"38634458",  6821 => x"48a10003",
     6822 => x"78030001",  6823 => x"38634c00",  6824 => x"28410004",
     6825 => x"14a4001f",  6826 => x"780b0001",  6827 => x"1426001f",
     6828 => x"98853800",  6829 => x"396b7778",  6830 => x"98c12800",
     6831 => x"78020001",  6832 => x"b9600800",  6833 => x"3842445c",
     6834 => x"c8e42000",  6835 => x"c8a62800",  6836 => x"f80016bd",
     6837 => x"b9600800",  6838 => x"2b9d0004",  6839 => x"2b8b0008",
     6840 => x"379c0008",  6841 => x"c3a00000",  6842 => x"379cfff8",
     6843 => x"5b8b0008",  6844 => x"5b9d0004",  6845 => x"28220020",
     6846 => x"28240028",  6847 => x"b8205800",  6848 => x"28430004",
     6849 => x"58600038",  6850 => x"28430014",  6851 => x"0c20010c",
     6852 => x"0c600008",  6853 => x"28830014",  6854 => x"44600013",
     6855 => x"d8600000",  6856 => x"3402ffff",  6857 => x"5c220008",
     6858 => x"78040001",  6859 => x"b9600800",  6860 => x"34020004",
     6861 => x"34030001",  6862 => x"38844468",  6863 => x"fbffe783",
     6864 => x"34010000",  6865 => x"29620020",  6866 => x"c8010800",
     6867 => x"3c21000a",  6868 => x"28420004",  6869 => x"1423001f",
     6870 => x"5841002c",  6871 => x"58430028",  6872 => x"e000000d",
     6873 => x"28420008",  6874 => x"28420038",  6875 => x"20420001",
     6876 => x"5c430005",  6877 => x"28840008",  6878 => x"34020000",
     6879 => x"34030000",  6880 => x"d8800000",  6881 => x"29610020",
     6882 => x"28210004",  6883 => x"58200028",  6884 => x"5820002c",
     6885 => x"29610020",  6886 => x"78040001",  6887 => x"34020004",
     6888 => x"28260004",  6889 => x"34030001",  6890 => x"b9600800",
     6891 => x"28c50028",  6892 => x"28c6002c",  6893 => x"38844484",
     6894 => x"fbffe764",  6895 => x"2b9d0004",  6896 => x"2b8b0008",
     6897 => x"379c0008",  6898 => x"c3a00000",  6899 => x"379cfff0",
     6900 => x"5b8b0010",  6901 => x"5b8c000c",  6902 => x"5b8d0008",
     6903 => x"5b9d0004",  6904 => x"b8205800",  6905 => x"28210020",
     6906 => x"35620094",  6907 => x"35630080",  6908 => x"282d0004",
     6909 => x"356c00d0",  6910 => x"b9a00800",  6911 => x"fbffff6c",
     6912 => x"b9a01000",  6913 => x"b9801800",  6914 => x"b9a00800",
     6915 => x"fbffff68",  6916 => x"b9800800",  6917 => x"fbffff92",
     6918 => x"78040001",  6919 => x"b8202800",  6920 => x"34020004",
     6921 => x"b9600800",  6922 => x"34030003",  6923 => x"388444a4",
     6924 => x"fbffe746",  6925 => x"2b9d0004",  6926 => x"2b8b0010",
     6927 => x"2b8c000c",  6928 => x"2b8d0008",  6929 => x"379c0010",
     6930 => x"c3a00000",  6931 => x"379cffb8",  6932 => x"5b8b0024",
     6933 => x"5b8c0020",  6934 => x"5b8d001c",  6935 => x"5b8e0018",
     6936 => x"5b8f0014",  6937 => x"5b900010",  6938 => x"5b91000c",
     6939 => x"5b920008",  6940 => x"5b9d0004",  6941 => x"28220020",
     6942 => x"b8205800",  6943 => x"284d0004",  6944 => x"284c0010",
     6945 => x"28220080",  6946 => x"5c400008",  6947 => x"28230084",
     6948 => x"5c620006",  6949 => x"78040001",  6950 => x"34020004",
     6951 => x"34030002",  6952 => x"388444bc",  6953 => x"e000006e",
     6954 => x"35af0014",  6955 => x"357000bc",  6956 => x"357100a8",
     6957 => x"b9e00800",  6958 => x"ba001000",  6959 => x"ba201800",
     6960 => x"fbffff3b",  6961 => x"357200d0",  6962 => x"b9e01000",
     6963 => x"ba401800",  6964 => x"b9e00800",  6965 => x"fbffff36",
     6966 => x"ba400800",  6967 => x"fbffff60",  6968 => x"78040001",
     6969 => x"b8202800",  6970 => x"34020004",  6971 => x"34030003",
     6972 => x"388444dc",  6973 => x"b9600800",  6974 => x"fbffe714",
     6975 => x"35610080",  6976 => x"fbffff57",  6977 => x"78040001",
     6978 => x"b8202800",  6979 => x"34020004",  6980 => x"34030002",
     6981 => x"388444f4",  6982 => x"b9600800",  6983 => x"fbffe70b",
     6984 => x"35610094",  6985 => x"fbffff4e",  6986 => x"78040001",
     6987 => x"b8202800",  6988 => x"34020004",  6989 => x"34030002",
     6990 => x"388444fc",  6991 => x"b9600800",  6992 => x"fbffe702",
     6993 => x"ba200800",  6994 => x"fbffff45",  6995 => x"78040001",
     6996 => x"b8202800",  6997 => x"34020004",  6998 => x"34030002",
     6999 => x"38844504",  7000 => x"b9600800",  7001 => x"fbffe6f9",
     7002 => x"ba000800",  7003 => x"fbffff3c",  7004 => x"78040001",
     7005 => x"b8202800",  7006 => x"34020004",  7007 => x"34030002",
     7008 => x"3884450c",  7009 => x"b9600800",  7010 => x"fbffe6f0",
     7011 => x"b9a00800",  7012 => x"fbffff33",  7013 => x"78040001",
     7014 => x"b8202800",  7015 => x"34020004",  7016 => x"34030001",
     7017 => x"38844514",  7018 => x"b9600800",  7019 => x"fbffe6e7",
     7020 => x"b9e00800",  7021 => x"fbffff2a",  7022 => x"78040001",
     7023 => x"b8202800",  7024 => x"3884452c",  7025 => x"b9600800",
     7026 => x"34020004",  7027 => x"34030001",  7028 => x"fbffe6de",
     7029 => x"29610020",  7030 => x"358e0018",  7031 => x"28220004",
     7032 => x"b9c00800",  7033 => x"34430014",  7034 => x"fbfffee3",
     7035 => x"b9c00800",  7036 => x"fbfffefd",  7037 => x"b9c00800",
     7038 => x"fbffff19",  7039 => x"78040001",  7040 => x"b8202800",
     7041 => x"34020004",  7042 => x"b9600800",  7043 => x"34030001",
     7044 => x"38844544",  7045 => x"fbffe6cd",  7046 => x"29610020",
     7047 => x"28220010",  7048 => x"28260004",  7049 => x"28420018",
     7050 => x"5c400142",  7051 => x"28210008",  7052 => x"28270030",
     7053 => x"44e2013c",  7054 => x"28c20000",  7055 => x"5c400003",
     7056 => x"28c30014",  7057 => x"44620008",  7058 => x"78040001",
     7059 => x"b9600800",  7060 => x"34020004",  7061 => x"34030001",
     7062 => x"38844558",  7063 => x"fbffe6bb",  7064 => x"e0000134",
     7065 => x"28c50004",  7066 => x"48a70003",  7067 => x"28c20018",
     7068 => x"4ce2012d",  7069 => x"28c60018",  7070 => x"78040001",
     7071 => x"b9600800",  7072 => x"34020004",  7073 => x"34030001",
     7074 => x"38844584",  7075 => x"fbffe6af",  7076 => x"e0000128",
     7077 => x"2982001c",  7078 => x"59a20034",  7079 => x"1c220040",
     7080 => x"29a10034",  7081 => x"3444ffff",  7082 => x"1423001f",
     7083 => x"98612800",  7084 => x"c8a32800",  7085 => x"3403001f",
     7086 => x"c8621800",  7087 => x"94a33800",  7088 => x"34820001",
     7089 => x"34630001",  7090 => x"3484ffff",  7091 => x"5ce0fffc",
     7092 => x"34030001",  7093 => x"bc621000",  7094 => x"4c460002",
     7095 => x"59a20038",  7096 => x"29a30038",  7097 => x"4c620003",
     7098 => x"34630001",  7099 => x"59a30038",  7100 => x"2982001c",
     7101 => x"4c400002",  7102 => x"5981001c",  7103 => x"2982001c",
     7104 => x"4c400002",  7105 => x"5980001c",  7106 => x"2985001c",
     7107 => x"08210003",  7108 => x"4c25000d",  7109 => x"78040001",
     7110 => x"b9600800",  7111 => x"34020004",  7112 => x"34030001",
     7113 => x"388445c8",  7114 => x"fbffe688",  7115 => x"29a10034",
     7116 => x"29a20038",  7117 => x"3c210001",  7118 => x"34420001",
     7119 => x"b4410800",  7120 => x"5981001c",  7121 => x"29af0038",
     7122 => x"29a20034",  7123 => x"35900004",  7124 => x"35e1ffff",
     7125 => x"88220800",  7126 => x"2982001c",  7127 => x"b4220800",
     7128 => x"b9e01000",  7129 => x"f8002eab",  7130 => x"59a10034",
     7131 => x"78040001",  7132 => x"b8203000",  7133 => x"b9e02800",
     7134 => x"388445e0",  7135 => x"5981001c",  7136 => x"34020004",
     7137 => x"b9600800",  7138 => x"34030001",  7139 => x"fbffe66f",
     7140 => x"b9a01000",  7141 => x"b9c01800",  7142 => x"ba000800",
     7143 => x"fbfffe84",  7144 => x"ba000800",  7145 => x"fbfffeae",
     7146 => x"78040001",  7147 => x"b8202800",  7148 => x"34020004",
     7149 => x"b9600800",  7150 => x"34030001",  7151 => x"38844604",
     7152 => x"fbffe662",  7153 => x"296f0020",  7154 => x"29e10008",
     7155 => x"2825002c",  7156 => x"44a00011",  7157 => x"29820004",
     7158 => x"44400007",  7159 => x"78040001",  7160 => x"b9600800",
     7161 => x"34020004",  7162 => x"34030001",  7163 => x"38844620",
     7164 => x"e3ffff9b",  7165 => x"29820008",  7166 => x"4ca20007",
     7167 => x"78040001",  7168 => x"b9600800",  7169 => x"34020004",
     7170 => x"34030001",  7171 => x"38844650",  7172 => x"e00000c3",
     7173 => x"29820004",  7174 => x"44400031",  7175 => x"28220038",
     7176 => x"20410001",  7177 => x"5c2000c3",  7178 => x"20420002",
     7179 => x"5c410019",  7180 => x"296300c4",  7181 => x"296200c8",
     7182 => x"296100cc",  7183 => x"5b830030",  7184 => x"29e30010",
     7185 => x"296500bc",  7186 => x"296400c0",  7187 => x"378c0028",
     7188 => x"5b820034",  7189 => x"5b810038",  7190 => x"b9801000",
     7191 => x"b9800800",  7192 => x"34630018",  7193 => x"5b850028",
     7194 => x"5b84002c",  7195 => x"fbfffe42",  7196 => x"29610028",
     7197 => x"b9801000",  7198 => x"28230004",  7199 => x"b9600800",
     7200 => x"d8600000",  7201 => x"b9600800",  7202 => x"fbfffe98",
     7203 => x"e00000a9",  7204 => x"29820008",  7205 => x"78030001",
     7206 => x"38635768",  7207 => x"28610000",  7208 => x"ec021000",
     7209 => x"78050001",  7210 => x"c8021000",  7211 => x"38a5576c",
     7212 => x"a0411000",  7213 => x"28a10000",  7214 => x"b4411000",
     7215 => x"29610028",  7216 => x"c8021000",  7217 => x"28230010",
     7218 => x"5c600002",  7219 => x"2823000c",  7220 => x"b9600800",
     7221 => x"d8600000",  7222 => x"e0000096",  7223 => x"29830008",
     7224 => x"29ed0004",  7225 => x"78050001",  7226 => x"1462001f",
     7227 => x"29b0002c",  7228 => x"00640016",  7229 => x"3c63000a",
     7230 => x"29ae0028",  7231 => x"3c42000a",  7232 => x"b4708000",
     7233 => x"b8821000",  7234 => x"f4701800",  7235 => x"b44e1000",
     7236 => x"b4627000",  7237 => x"1c22003e",  7238 => x"38a5576c",
     7239 => x"28a40000",  7240 => x"1441001f",  7241 => x"34030000",
     7242 => x"59ae0028",  7243 => x"59b0002c",  7244 => x"f8002e11",
     7245 => x"00430016",  7246 => x"3c21000a",  7247 => x"3c42000a",
     7248 => x"b8610800",  7249 => x"49c1000b",  7250 => x"5dc10002",
     7251 => x"56020009",  7252 => x"c8021000",  7253 => x"7c430000",
     7254 => x"c8010800",  7255 => x"c8230800",  7256 => x"482e0004",
     7257 => x"5c2e0005",  7258 => x"54500002",  7259 => x"e0000003",
     7260 => x"59a10028",  7261 => x"59a2002c",  7262 => x"29a10028",
     7263 => x"29a2002c",  7264 => x"48200003",  7265 => x"5c200004",
     7266 => x"44410003",  7267 => x"340d0000",  7268 => x"e0000002",
     7269 => x"340dffff",  7270 => x"5b810044",  7271 => x"5b820048",
     7272 => x"45a00007",  7273 => x"c8021000",  7274 => x"7c430000",
     7275 => x"c8010800",  7276 => x"c8230800",  7277 => x"5b810044",
     7278 => x"5b820048",  7279 => x"29e20008",  7280 => x"37810044",
     7281 => x"1c42003e",  7282 => x"fbffea08",  7283 => x"45a00009",
     7284 => x"2b810048",  7285 => x"2b820044",  7286 => x"c8010800",
     7287 => x"7c230000",  7288 => x"c8021000",  7289 => x"c8431000",
     7290 => x"5b820044",  7291 => x"5b810048",  7292 => x"29820008",
     7293 => x"1441001f",  7294 => x"00430016",  7295 => x"3c21000a",
     7296 => x"ec026000",  7297 => x"3c42000a",  7298 => x"b8610800",
     7299 => x"c80c6000",  7300 => x"5b81003c",  7301 => x"5b820040",
     7302 => x"45800007",  7303 => x"c8021000",  7304 => x"7c430000",
     7305 => x"c8010800",  7306 => x"c8230800",  7307 => x"5b81003c",
     7308 => x"5b820040",  7309 => x"29610020",  7310 => x"28220008",
     7311 => x"3781003c",  7312 => x"1c42003c",  7313 => x"fbffe9e9",
     7314 => x"45800009",  7315 => x"2b810040",  7316 => x"2b82003c",
     7317 => x"c8010800",  7318 => x"7c230000",  7319 => x"c8021000",
     7320 => x"c8431000",  7321 => x"5b82003c",  7322 => x"5b810040",
     7323 => x"2b830048",  7324 => x"2b820040",  7325 => x"2b81003c",
     7326 => x"2b840044",  7327 => x"b4621000",  7328 => x"f4621800",
     7329 => x"b4810800",  7330 => x"b4610800",  7331 => x"48200003",
     7332 => x"5c200006",  7333 => x"44410005",  7334 => x"3c210016",
     7335 => x"0042000a",  7336 => x"b8221000",  7337 => x"e0000009",
     7338 => x"c8021000",  7339 => x"7c430000",  7340 => x"c8010800",
     7341 => x"c8230800",  7342 => x"3c210016",  7343 => x"0042000a",
     7344 => x"b8221000",  7345 => x"c8021000",  7346 => x"29610020",
     7347 => x"28210008",  7348 => x"28250038",  7349 => x"20a50001",
     7350 => x"5ca00008",  7351 => x"29640028",  7352 => x"c8021000",
     7353 => x"28830010",  7354 => x"5c650002",  7355 => x"2883000c",
     7356 => x"b9600800",  7357 => x"d8600000",  7358 => x"29610020",
     7359 => x"78040001",  7360 => x"34020004",  7361 => x"28210004",
     7362 => x"34030002",  7363 => x"3884468c",  7364 => x"2825002c",
     7365 => x"b9600800",  7366 => x"14a5000a",  7367 => x"fbffe58b",
     7368 => x"e0000004",  7369 => x"29a60038",  7370 => x"4c06fedb",
     7371 => x"e3fffedc",  7372 => x"2b9d0004",  7373 => x"2b8b0024",
     7374 => x"2b8c0020",  7375 => x"2b8d001c",  7376 => x"2b8e0018",
     7377 => x"2b8f0014",  7378 => x"2b900010",  7379 => x"2b91000c",
     7380 => x"2b920008",  7381 => x"379c0048",  7382 => x"c3a00000",
     7383 => x"379cfffc",  7384 => x"5b9d0004",  7385 => x"78030001",
     7386 => x"3c420002",  7387 => x"38636524",  7388 => x"b4622800",
     7389 => x"28a50000",  7390 => x"78040001",  7391 => x"34020006",
     7392 => x"34030001",  7393 => x"388446a4",  7394 => x"fbffe570",
     7395 => x"2b9d0004",  7396 => x"379c0004",  7397 => x"c3a00000",
     7398 => x"379cfff0",  7399 => x"5b8b0010",  7400 => x"5b8c000c",
     7401 => x"5b8d0008",  7402 => x"5b9d0004",  7403 => x"b8205800",
     7404 => x"78010001",  7405 => x"38217790",  7406 => x"b8406800",
     7407 => x"28220000",  7408 => x"5c400005",  7409 => x"29620020",
     7410 => x"2844000c",  7411 => x"28820008",  7412 => x"58220000",
     7413 => x"78040001",  7414 => x"78010001",  7415 => x"38847790",
     7416 => x"38215770",  7417 => x"28260000",  7418 => x"28850000",
     7419 => x"340c0190",  7420 => x"bd836000",  7421 => x"88a62800",
     7422 => x"b9801000",  7423 => x"34a53039",  7424 => x"00a10010",
     7425 => x"88a62800",  7426 => x"202107ff",  7427 => x"34a53039",
     7428 => x"58850000",  7429 => x"00a50010",  7430 => x"3c24000a",
     7431 => x"20a103ff",  7432 => x"b8240800",  7433 => x"f8002dd8",
     7434 => x"3d820001",  7435 => x"b4221000",  7436 => x"29610028",
     7437 => x"28230018",  7438 => x"b9600800",  7439 => x"d8600000",
     7440 => x"35a200b2",  7441 => x"3c420002",  7442 => x"b5625800",
     7443 => x"59610004",  7444 => x"2b9d0004",  7445 => x"2b8b0010",
     7446 => x"2b8c000c",  7447 => x"2b8d0008",  7448 => x"379c0010",
     7449 => x"c3a00000",  7450 => x"379cfff0",  7451 => x"5b8b0010",
     7452 => x"5b8c000c",  7453 => x"5b8d0008",  7454 => x"5b9d0004",
     7455 => x"282b000c",  7456 => x"b8206000",  7457 => x"34010001",
     7458 => x"59610000",  7459 => x"29810024",  7460 => x"48200002",
     7461 => x"34010001",  7462 => x"0d61000c",  7463 => x"29810008",
     7464 => x"5c200002",  7465 => x"59820008",  7466 => x"298d0008",
     7467 => x"3561000e",  7468 => x"34030004",  7469 => x"b9a01000",
     7470 => x"f8002e04",  7471 => x"2d62000c",  7472 => x"34010001",
     7473 => x"5c410004",  7474 => x"29810000",  7475 => x"4021001d",
     7476 => x"64210002",  7477 => x"59610018",  7478 => x"41a10044",
     7479 => x"2d67000c",  7480 => x"34060002",  7481 => x"31610012",
     7482 => x"41a10045",  7483 => x"34050001",  7484 => x"3404ffff",
     7485 => x"31610013",  7486 => x"41a10046",  7487 => x"31610014",
     7488 => x"34010000",  7489 => x"e000000c",  7490 => x"08220374",
     7491 => x"29880000",  7492 => x"b5021000",  7493 => x"44600004",
     7494 => x"4043001d",  7495 => x"44660002",  7496 => x"59600018",
     7497 => x"58410338",  7498 => x"58450000",  7499 => x"0c44010e",
     7500 => x"34210001",  7501 => x"29630018",  7502 => x"48e1fff4",
     7503 => x"44600006",  7504 => x"78010001",  7505 => x"38214734",
     7506 => x"f800142d",  7507 => x"3401ffff",  7508 => x"3161000e",
     7509 => x"78010001",  7510 => x"382164ac",  7511 => x"28230004",
     7512 => x"34010000",  7513 => x"44600004",  7514 => x"b9800800",
     7515 => x"b9a01000",  7516 => x"d8600000",  7517 => x"2b9d0004",
     7518 => x"2b8b0010",  7519 => x"2b8c000c",  7520 => x"2b8d0008",
     7521 => x"379c0010",  7522 => x"c3a00000",  7523 => x"379cfffc",
     7524 => x"5b9d0004",  7525 => x"78020001",  7526 => x"384264ac",
     7527 => x"28430008",  7528 => x"34020000",  7529 => x"44600003",
     7530 => x"d8600000",  7531 => x"b8201000",  7532 => x"b8400800",
     7533 => x"2b9d0004",  7534 => x"379c0004",  7535 => x"c3a00000",
     7536 => x"78010001",  7537 => x"38216590",  7538 => x"28220000",
     7539 => x"78010001",  7540 => x"38216374",  7541 => x"e0000004",
     7542 => x"28440000",  7543 => x"44640004",  7544 => x"3421000c",
     7545 => x"28230000",  7546 => x"5c60fffc",  7547 => x"28210004",
     7548 => x"c3a00000",  7549 => x"379cfff4",  7550 => x"5b9d0004",
     7551 => x"5b810008",  7552 => x"5b82000c",  7553 => x"b8401800",
     7554 => x"5c20000b",  7555 => x"78020001",  7556 => x"38425758",
     7557 => x"28410000",  7558 => x"54610007",  7559 => x"78010001",
     7560 => x"78020001",  7561 => x"38424758",  7562 => x"38217798",
     7563 => x"f80013e6",  7564 => x"e000000d",  7565 => x"78030001",
     7566 => x"38635748",  7567 => x"28620000",  7568 => x"37810008",
     7569 => x"fbffe8e9",  7570 => x"2b83000c",  7571 => x"b8202000",
     7572 => x"78020001",  7573 => x"78010001",  7574 => x"38217798",
     7575 => x"3842475c",  7576 => x"f80013d9",  7577 => x"78010001",
     7578 => x"38217798",  7579 => x"2b9d0004",  7580 => x"379c000c",
     7581 => x"c3a00000",  7582 => x"379cff18",  7583 => x"5b8b000c",
     7584 => x"5b8c0008",  7585 => x"5b9d0004",  7586 => x"78010001",
     7587 => x"38216590",  7588 => x"28210000",  7589 => x"282b0014",
     7590 => x"78010001",  7591 => x"38218f7c",  7592 => x"28220000",
     7593 => x"34010000",  7594 => x"444000ce",  7595 => x"780c0001",
     7596 => x"398c7794",  7597 => x"29810000",  7598 => x"5c200008",
     7599 => x"f8001990",  7600 => x"78020001",  7601 => x"38425e88",
     7602 => x"28420000",  7603 => x"a4401000",  7604 => x"b4410800",
     7605 => x"59810000",  7606 => x"78010001",  7607 => x"38218c1c",
     7608 => x"28210000",  7609 => x"296200b8",  7610 => x"5c220007",
     7611 => x"78010001",  7612 => x"38217284",  7613 => x"28230000",
     7614 => x"34020003",  7615 => x"34010000",  7616 => x"446200b8",
     7617 => x"f800197e",  7618 => x"78030001",  7619 => x"78020001",
     7620 => x"38635e88",  7621 => x"38427794",  7622 => x"28630000",
     7623 => x"28420000",  7624 => x"b4621000",  7625 => x"c8220800",
     7626 => x"4c200007",  7627 => x"78010001",  7628 => x"38217284",
     7629 => x"28230000",  7630 => x"34020003",  7631 => x"34010000",
     7632 => x"5c6200a8",  7633 => x"f800196e",  7634 => x"78020001",
     7635 => x"38427794",  7636 => x"58410000",  7637 => x"296200b8",
     7638 => x"78010001",  7639 => x"38218c1c",  7640 => x"58220000",
     7641 => x"378100d8",  7642 => x"378200e0",  7643 => x"f8001cdf",
     7644 => x"34020000",  7645 => x"37810010",  7646 => x"f8000287",
     7647 => x"378100e8",  7648 => x"378200e4",  7649 => x"f8001945",
     7650 => x"2b8300e4",  7651 => x"2b8400e8",  7652 => x"2b82003c",
     7653 => x"78010001",  7654 => x"38214764",  7655 => x"f8001398",
     7656 => x"2b820044",  7657 => x"78010001",  7658 => x"38214778",
     7659 => x"7c420000",  7660 => x"f8001393",  7661 => x"fbffff83",
     7662 => x"b8201000",  7663 => x"78010001",  7664 => x"38214784",
     7665 => x"f800138e",  7666 => x"78010001",  7667 => x"38217284",
     7668 => x"28220000",  7669 => x"34010003",  7670 => x"5c41000a",
     7671 => x"29620010",  7672 => x"78010001",  7673 => x"3821478c",
     7674 => x"20420001",  7675 => x"f8001384",  7676 => x"78010001",
     7677 => x"38214794",  7678 => x"356200c0",  7679 => x"f8001380",
     7680 => x"34010000",  7681 => x"f8002a4f",  7682 => x"b8201000",
     7683 => x"78010001",  7684 => x"382147a0",  7685 => x"f800137a",
     7686 => x"2b8200dc",  7687 => x"2b8300e0",  7688 => x"78010001",
     7689 => x"382147a8",  7690 => x"f8001375",  7691 => x"78010001",
     7692 => x"38217284",  7693 => x"28220000",  7694 => x"34010003",
     7695 => x"5c41004b",  7696 => x"296200a4",  7697 => x"296100a0",
     7698 => x"fbffff6b",  7699 => x"b8201000",  7700 => x"78010001",
     7701 => x"382147b8",  7702 => x"f8001369",  7703 => x"296200b4",
     7704 => x"296100b0",  7705 => x"fbffff64",  7706 => x"b8201000",
     7707 => x"78010001",  7708 => x"382147c0",  7709 => x"f8001362",
     7710 => x"29620018",  7711 => x"2963001c",  7712 => x"78010001",
     7713 => x"382147c8",  7714 => x"f800135d",  7715 => x"29620020",
     7716 => x"29630024",  7717 => x"78010001",  7718 => x"382147dc",
     7719 => x"f8001358",  7720 => x"296200b4",  7721 => x"296300a4",
     7722 => x"78010001",  7723 => x"3c420001",  7724 => x"382147f0",
     7725 => x"c8621000",  7726 => x"f8001351",  7727 => x"29620018",
     7728 => x"296100a4",  7729 => x"296300a0",  7730 => x"1444001f",
     7731 => x"c8221000",  7732 => x"f4410800",  7733 => x"c8641800",
     7734 => x"c8611800",  7735 => x"2961001c",  7736 => x"1424001f",
     7737 => x"c8410800",  7738 => x"f4221000",  7739 => x"c8641800",
     7740 => x"c8621000",  7741 => x"29630020",  7742 => x"1464001f",
     7743 => x"c8231800",  7744 => x"f4610800",  7745 => x"c8441000",
     7746 => x"c8410800",  7747 => x"29620024",  7748 => x"1444001f",
     7749 => x"c8621000",  7750 => x"f4431800",  7751 => x"c8240800",
     7752 => x"c8230800",  7753 => x"fbffff34",  7754 => x"b8201000",
     7755 => x"78010001",  7756 => x"382147fc",  7757 => x"f8001332",
     7758 => x"296200ec",  7759 => x"78010001",  7760 => x"38214808",
     7761 => x"f800132e",  7762 => x"296200a8",  7763 => x"78010001",
     7764 => x"38214810",  7765 => x"f800132a",  7766 => x"296200b8",
     7767 => x"78010001",  7768 => x"3821481c",  7769 => x"f8001326",
     7770 => x"3401ffff",  7771 => x"f8002a00",  7772 => x"b8206000",
     7773 => x"34010000",  7774 => x"f80029fd",  7775 => x"b8205800",
     7776 => x"34010001",  7777 => x"f80029fa",  7778 => x"78050001",
     7779 => x"b8202000",  7780 => x"b8a00800",  7781 => x"b9801000",
     7782 => x"b9601800",  7783 => x"38214828",  7784 => x"f8001317",
     7785 => x"78010001",  7786 => x"3821483c",  7787 => x"f8001b4a",
     7788 => x"2023ffff",  7789 => x"08632710",  7790 => x"b8201000",
     7791 => x"14420010",  7792 => x"14630010",  7793 => x"78010001",
     7794 => x"38214840",  7795 => x"f800130c",  7796 => x"78010001",
     7797 => x"38214adc",  7798 => x"f8001309",  7799 => x"34010001",
     7800 => x"2b9d0004",  7801 => x"2b8b000c",  7802 => x"2b8c0008",
     7803 => x"379c00e8",  7804 => x"c3a00000",  7805 => x"379cfff4",
     7806 => x"5b8b000c",  7807 => x"5b8c0008",  7808 => x"5b9d0004",
     7809 => x"780b0001",  7810 => x"396b6590",  7811 => x"29610000",
     7812 => x"78020001",  7813 => x"38424850",  7814 => x"282c0014",
     7815 => x"34010004",  7816 => x"f80008c8",  7817 => x"fbfffee7",
     7818 => x"78020001",  7819 => x"b8201800",  7820 => x"38424860",
     7821 => x"34010007",  7822 => x"f80008c2",  7823 => x"29810010",
     7824 => x"44200005",  7825 => x"29610000",  7826 => x"28220000",
     7827 => x"34010009",  7828 => x"44410007",  7829 => x"78020001",
     7830 => x"34010001",  7831 => x"38424864",  7832 => x"f80008b8",
     7833 => x"34010000",  7834 => x"e0000006",  7835 => x"78020001",
     7836 => x"34010004",  7837 => x"3842487c",  7838 => x"f80008b2",
     7839 => x"34010001",  7840 => x"2b9d0004",  7841 => x"2b8b000c",
     7842 => x"2b8c0008",  7843 => x"379c000c",  7844 => x"c3a00000",
     7845 => x"379cfef0",  7846 => x"5b8b0018",  7847 => x"5b8c0014",
     7848 => x"5b8d0010",  7849 => x"5b8e000c",  7850 => x"5b8f0008",
     7851 => x"5b9d0004",  7852 => x"78010001",  7853 => x"38216590",
     7854 => x"28210000",  7855 => x"780c0001",  7856 => x"398c77b4",
     7857 => x"282b0014",  7858 => x"29810000",  7859 => x"5c200008",
     7860 => x"f800188b",  7861 => x"78020001",  7862 => x"38425e88",
     7863 => x"28420000",  7864 => x"a4401000",  7865 => x"b4410800",
     7866 => x"59810000",  7867 => x"f8001884",  7868 => x"78030001",
     7869 => x"78020001",  7870 => x"38635e88",  7871 => x"384277b4",
     7872 => x"28630000",  7873 => x"28420000",  7874 => x"b4621000",
     7875 => x"c8220800",  7876 => x"4c200007",  7877 => x"78010001",
     7878 => x"382177b0",  7879 => x"28210000",  7880 => x"296200b8",
     7881 => x"340d0000",  7882 => x"44220192",  7883 => x"f8001874",
     7884 => x"78020001",  7885 => x"384277b4",  7886 => x"58410000",
     7887 => x"296200b8",  7888 => x"78010001",  7889 => x"382177b0",
     7890 => x"58220000",  7891 => x"f80008c3",  7892 => x"78040001",
     7893 => x"34010001",  7894 => x"34020001",  7895 => x"34030004",
     7896 => x"38844898",  7897 => x"f8000896",  7898 => x"78040001",
     7899 => x"388448b8",  7900 => x"34030087",  7901 => x"34010002",
     7902 => x"34020001",  7903 => x"f8000890",  7904 => x"378100fc",
     7905 => x"37820108",  7906 => x"f8001bd8",  7907 => x"78020001",
     7908 => x"34010004",  7909 => x"384248c4",  7910 => x"f800086a",
     7911 => x"2b820100",  7912 => x"2b8100fc",  7913 => x"34030000",
     7914 => x"f80007b5",  7915 => x"78020001",  7916 => x"b8201800",
     7917 => x"38424860",  7918 => x"34010007",  7919 => x"f8000861",
     7920 => x"34020000",  7921 => x"37810020",  7922 => x"f8000173",
     7923 => x"78040001",  7924 => x"34010004",  7925 => x"34020001",
     7926 => x"34030004",  7927 => x"388448e4",  7928 => x"f8000877",
     7929 => x"78040001",  7930 => x"78050001",  7931 => x"34010006",
     7932 => x"34020001",  7933 => x"34030007",  7934 => x"388448f4",
     7935 => x"38a548fc",  7936 => x"f800086f",  7937 => x"2b81004c",
     7938 => x"44200005",  7939 => x"78020001",  7940 => x"34010002",
     7941 => x"38424904",  7942 => x"e0000004",  7943 => x"78020001",
     7944 => x"34010001",  7945 => x"38424910",  7946 => x"f8000846",
     7947 => x"2b81004c",  7948 => x"4420014c",  7949 => x"37810110",
     7950 => x"3782010c",  7951 => x"f8001817",  7952 => x"2b83010c",
     7953 => x"2b840110",  7954 => x"78020001",  7955 => x"34010087",
     7956 => x"3842491c",  7957 => x"780c0001",  7958 => x"f800083a",
     7959 => x"398c6590",  7960 => x"29810000",  7961 => x"282102c8",
     7962 => x"28210010",  7963 => x"282e0008",  7964 => x"5dc00039",
     7965 => x"78020001",  7966 => x"34010001",  7967 => x"38424938",
     7968 => x"f8000830",  7969 => x"fbffff5c",  7970 => x"340d0001",
     7971 => x"442e0139",  7972 => x"78020001",  7973 => x"34010087",
     7974 => x"38424940",  7975 => x"f8000829",  7976 => x"29810000",
     7977 => x"28210020",  7978 => x"28240010",  7979 => x"28830004",
     7980 => x"4460000b",  7981 => x"78020001",  7982 => x"38424960",
     7983 => x"28840008",  7984 => x"4c030003",  7985 => x"34010007",
     7986 => x"e0000003",  7987 => x"34010007",  7988 => x"c8042000",
     7989 => x"f800081b",  7990 => x"e0000126",  7991 => x"28830008",
     7992 => x"780b0001",  7993 => x"396b496c",  7994 => x"b9601000",
     7995 => x"34010007",  7996 => x"f8000814",  7997 => x"78020001",
     7998 => x"34010087",  7999 => x"38424974",  8000 => x"f8000810",
     8001 => x"29810000",  8002 => x"b9601000",  8003 => x"28210020",
     8004 => x"28230010",  8005 => x"34010007",  8006 => x"2863001c",
     8007 => x"f8000809",  8008 => x"78020001",  8009 => x"34010087",
     8010 => x"38424994",  8011 => x"f8000805",  8012 => x"29810000",
     8013 => x"b9601000",  8014 => x"28210020",  8015 => x"28240004",
     8016 => x"34010007",  8017 => x"28830028",  8018 => x"2884002c",
     8019 => x"f80007fd",  8020 => x"e0000108",  8021 => x"78010001",
     8022 => x"38217284",  8023 => x"28210000",  8024 => x"34020001",
     8025 => x"4841000e",  8026 => x"34020002",  8027 => x"4c410004",
     8028 => x"34020003",  8029 => x"5c22000a",  8030 => x"e0000005",
     8031 => x"78020001",  8032 => x"34010007",  8033 => x"384249b4",
     8034 => x"e0000008",  8035 => x"78020001",  8036 => x"34010007",
     8037 => x"384249c0",  8038 => x"e0000004",  8039 => x"78020001",
     8040 => x"34010001",  8041 => x"384249cc",  8042 => x"f80007e6",
     8043 => x"2b810054",  8044 => x"44200005",  8045 => x"78020001",
     8046 => x"34010002",  8047 => x"384249dc",  8048 => x"e0000004",
     8049 => x"78020001",  8050 => x"34010001",  8051 => x"384249e8",
     8052 => x"f80007dc",  8053 => x"2b810070",  8054 => x"44200007",
     8055 => x"2b810074",  8056 => x"44200005",  8057 => x"78020001",
     8058 => x"34010002",  8059 => x"384249f4",  8060 => x"e0000004",
     8061 => x"78020001",  8062 => x"34010001",  8063 => x"38424a04",
     8064 => x"f80007d0",  8065 => x"78020001",  8066 => x"38424a14",
     8067 => x"34010007",  8068 => x"f80007cc",  8069 => x"378c0104",
     8070 => x"b9800800",  8071 => x"f8000b58",  8072 => x"378300e8",
     8073 => x"b8600800",  8074 => x"b9801000",  8075 => x"5b83001c",
     8076 => x"f800067c",  8077 => x"78010001",  8078 => x"38217a80",
     8079 => x"28210000",  8080 => x"34020001",  8081 => x"2b83001c",
     8082 => x"4422000a",  8083 => x"44200004",  8084 => x"34020002",
     8085 => x"5c22000f",  8086 => x"e000000a",  8087 => x"78020001",
     8088 => x"34010001",  8089 => x"38424a1c",  8090 => x"f80007b6",
     8091 => x"e0000009",  8092 => x"78020001",  8093 => x"34010002",
     8094 => x"38424a2c",  8095 => x"e0000004",  8096 => x"78020001",
     8097 => x"34010002",  8098 => x"38424a3c",  8099 => x"f80007ad",
     8100 => x"fbfffed9",  8101 => x"340d0001",  8102 => x"442000b6",
     8103 => x"78020001",  8104 => x"34010087",  8105 => x"38424a54",
     8106 => x"f80007a6",  8107 => x"78020001",  8108 => x"34010007",
     8109 => x"3842461c",  8110 => x"356300c0",  8111 => x"f80007a1",
     8112 => x"78020001",  8113 => x"34010087",  8114 => x"38424a70",
     8115 => x"f800079d",  8116 => x"296100bc",  8117 => x"44200005",
     8118 => x"78020001",  8119 => x"34010002",  8120 => x"38424a8c",
     8121 => x"e0000004",  8122 => x"78020001",  8123 => x"34010001",
     8124 => x"38424a90",  8125 => x"f8000793",  8126 => x"78020001",
     8127 => x"34010087",  8128 => x"38424a98",  8129 => x"f800078f",
     8130 => x"34010000",  8131 => x"f800288d",  8132 => x"b8206000",
     8133 => x"20210001",  8134 => x"44200005",  8135 => x"78020001",
     8136 => x"34010002",  8137 => x"38424ab4",  8138 => x"f8000786",
     8139 => x"218c0002",  8140 => x"45800005",  8141 => x"78020001",
     8142 => x"34010002",  8143 => x"38424abc",  8144 => x"f8000780",
     8145 => x"78010001",  8146 => x"38214adc",  8147 => x"f80011ac",
     8148 => x"78020001",  8149 => x"34010004",  8150 => x"38424ac8",
     8151 => x"f8000779",  8152 => x"78020001",  8153 => x"34010087",
     8154 => x"38424ae0",  8155 => x"f8000775",  8156 => x"296200a4",
     8157 => x"296100a0",  8158 => x"780d0001",  8159 => x"39ad4afc",
     8160 => x"fbfffd9d",  8161 => x"b8201800",  8162 => x"b9a01000",
     8163 => x"34010007",  8164 => x"f800076c",  8165 => x"78020001",
     8166 => x"34010087",  8167 => x"38424b04",  8168 => x"f8000768",
     8169 => x"296200b4",  8170 => x"296100b0",  8171 => x"780c0001",
     8172 => x"398c4b3c",  8173 => x"fbfffd90",  8174 => x"b8201800",
     8175 => x"b9a01000",  8176 => x"34010007",  8177 => x"f800075f",
     8178 => x"78020001",  8179 => x"34010087",  8180 => x"38424b20",
     8181 => x"f800075b",  8182 => x"29630018",  8183 => x"2964001c",
     8184 => x"b9801000",  8185 => x"34010007",  8186 => x"f8000756",
     8187 => x"78020001",  8188 => x"34010087",  8189 => x"38424b54",
     8190 => x"f8000752",  8191 => x"29640024",  8192 => x"29630020",
     8193 => x"b9801000",  8194 => x"34010007",  8195 => x"f800074d",
     8196 => x"296e00b4",  8197 => x"296100a4",  8198 => x"78020001",
     8199 => x"3dce0001",  8200 => x"38424b70",  8201 => x"c82e7000",
     8202 => x"780c0001",  8203 => x"34010087",  8204 => x"f8000744",
     8205 => x"398c4b8c",  8206 => x"b9c01800",  8207 => x"34010007",
     8208 => x"b9801000",  8209 => x"f800073f",  8210 => x"29610018",
     8211 => x"296200a4",  8212 => x"296f00a0",  8213 => x"1423001f",
     8214 => x"c8410800",  8215 => x"f4221000",  8216 => x"c9e37800",
     8217 => x"c9e27800",  8218 => x"2962001c",  8219 => x"296e0024",
     8220 => x"1443001f",  8221 => x"c8221000",  8222 => x"f4410800",
     8223 => x"c9e37800",  8224 => x"c9e17800",  8225 => x"29610020",
     8226 => x"1423001f",  8227 => x"c8410800",  8228 => x"f4221000",
     8229 => x"c9e37800",  8230 => x"15c3001f",  8231 => x"c82e7000",
     8232 => x"c9e27800",  8233 => x"f5c10800",  8234 => x"c9e37800",
     8235 => x"78020001",  8236 => x"c9e17800",  8237 => x"38424b94",
     8238 => x"34010087",  8239 => x"f8000721",  8240 => x"b9c01000",
     8241 => x"b9e00800",  8242 => x"fbfffd4b",  8243 => x"b8201800",
     8244 => x"b9a01000",  8245 => x"34010007",  8246 => x"f800071a",
     8247 => x"78020001",  8248 => x"34010087",  8249 => x"38424bb0",
     8250 => x"f8000716",  8251 => x"296300ec",  8252 => x"34010007",
     8253 => x"b9801000",  8254 => x"f8000712",  8255 => x"78020001",
     8256 => x"34010087",  8257 => x"38424bcc",  8258 => x"f800070e",
     8259 => x"296300a8",  8260 => x"34010007",  8261 => x"b9801000",
     8262 => x"f800070a",  8263 => x"78020001",  8264 => x"34010087",
     8265 => x"38424be8",  8266 => x"f8000706",  8267 => x"296300e4",
     8268 => x"34010007",  8269 => x"b9801000",  8270 => x"f8000702",
     8271 => x"78020001",  8272 => x"34010087",  8273 => x"38424c04",
     8274 => x"f80006fe",  8275 => x"296300b8",  8276 => x"78020001",
     8277 => x"34010007",  8278 => x"38424c20",  8279 => x"f80006f9",
     8280 => x"78010001",  8281 => x"38214c28",  8282 => x"f8001125",
     8283 => x"340d0001",  8284 => x"b9a00800",  8285 => x"2b9d0004",
     8286 => x"2b8b0018",  8287 => x"2b8c0014",  8288 => x"2b8d0010",
     8289 => x"2b8e000c",  8290 => x"2b8f0008",  8291 => x"379c0110",
     8292 => x"c3a00000",  8293 => x"379cfff4",  8294 => x"5b8b0008",
     8295 => x"5b9d0004",  8296 => x"b8205800",  8297 => x"fbffe306",
     8298 => x"34020003",  8299 => x"5c220003",  8300 => x"34010002",
     8301 => x"e0000002",  8302 => x"34010001",  8303 => x"59610028",
     8304 => x"3562004c",  8305 => x"35610048",  8306 => x"f8001288",
     8307 => x"34010000",  8308 => x"59600040",  8309 => x"59600044",
     8310 => x"59600088",  8311 => x"5960008c",  8312 => x"3782000c",
     8313 => x"34030000",  8314 => x"f800274b",  8315 => x"44200006",
     8316 => x"2b81000c",  8317 => x"596100a0",  8318 => x"34010001",
     8319 => x"596100a4",  8320 => x"e0000003",  8321 => x"596000a0",
     8322 => x"596000a4",  8323 => x"34010000",  8324 => x"f800124e",
     8325 => x"5961002c",  8326 => x"34010001",  8327 => x"59610054",
     8328 => x"59610050",  8329 => x"34010000",  8330 => x"f80026d6",
     8331 => x"59610034",  8332 => x"34011f40",  8333 => x"596100b4",
     8334 => x"78010001",  8335 => x"38215e90",  8336 => x"28210000",
     8337 => x"596100b8",  8338 => x"596100bc",  8339 => x"35610014",
     8340 => x"f80011f3",  8341 => x"34010000",  8342 => x"5960001c",
     8343 => x"2b9d0004",  8344 => x"2b8b0008",  8345 => x"379c000c",
     8346 => x"c3a00000",  8347 => x"c3a00000",  8348 => x"379cfffc",
     8349 => x"5b9d0004",  8350 => x"b8201000",  8351 => x"78010001",
     8352 => x"38214c3c",  8353 => x"f80010de",  8354 => x"2b9d0004",
     8355 => x"379c0004",  8356 => x"c3a00000",  8357 => x"379cffcc",
     8358 => x"5b8b0010",  8359 => x"5b8c000c",  8360 => x"5b8d0008",
     8361 => x"5b9d0004",  8362 => x"378b0014",  8363 => x"34020000",
     8364 => x"34030024",  8365 => x"b9600800",  8366 => x"f8002b02",
     8367 => x"78030001",  8368 => x"b9600800",  8369 => x"34040000",
     8370 => x"34020000",  8371 => x"386377b8",  8372 => x"34080020",
     8373 => x"34070008",  8374 => x"e0000004",  8375 => x"34840001",
     8376 => x"34210004",  8377 => x"44870017",  8378 => x"b4432800",
     8379 => x"e0000004",  8380 => x"30a00000",  8381 => x"34420001",
     8382 => x"34a50001",  8383 => x"40a60000",  8384 => x"44c8fffc",
     8385 => x"44c0000d",  8386 => x"b4432800",  8387 => x"58250000",
     8388 => x"e0000002",  8389 => x"34420001",  8390 => x"b4432800",
     8391 => x"40a50000",  8392 => x"7ca90000",  8393 => x"7ca60020",
     8394 => x"a1263000",  8395 => x"5cc0fffa",  8396 => x"5ca6ffeb",
     8397 => x"e0000003",  8398 => x"340c0000",  8399 => x"448c0021",
     8400 => x"2b810014",  8401 => x"340c0000",  8402 => x"40220000",
     8403 => x"34010023",  8404 => x"4441001c",  8405 => x"780b0001",
     8406 => x"780c0001",  8407 => x"396b7058",  8408 => x"398c7108",
     8409 => x"e0000011",  8410 => x"29610000",  8411 => x"f8002b16",
     8412 => x"b8206800",  8413 => x"5c20000c",  8414 => x"29620004",
     8415 => x"37810018",  8416 => x"d8400000",  8417 => x"b8206000",
     8418 => x"4c2d000e",  8419 => x"29620000",  8420 => x"78010001",
     8421 => x"b9801800",  8422 => x"38214c44",  8423 => x"f8001098",
     8424 => x"e0000008",  8425 => x"356b0008",  8426 => x"2b820014",
     8427 => x"558bffef",  8428 => x"78010001",  8429 => x"38214c5c",
     8430 => x"f8001091",  8431 => x"340cffea",  8432 => x"b9800800",
     8433 => x"2b9d0004",  8434 => x"2b8b0010",  8435 => x"2b8c000c",
     8436 => x"2b8d0008",  8437 => x"379c0034",  8438 => x"c3a00000",
     8439 => x"379cfff8",  8440 => x"5b8b0008",  8441 => x"5b9d0004",
     8442 => x"780b0001",  8443 => x"396b780c",  8444 => x"29650000",
     8445 => x"78020001",  8446 => x"34240001",  8447 => x"b8201800",
     8448 => x"384277b8",  8449 => x"b4220800",  8450 => x"c8a31800",
     8451 => x"b4821000",  8452 => x"f8002a67",  8453 => x"29610000",
     8454 => x"3421ffff",  8455 => x"59610000",  8456 => x"2b9d0004",
     8457 => x"2b8b0008",  8458 => x"379c0008",  8459 => x"c3a00000",
     8460 => x"78010001",  8461 => x"38217814",  8462 => x"58200000",
     8463 => x"78010001",  8464 => x"3821780c",  8465 => x"58200000",
     8466 => x"78010001",  8467 => x"38217810",  8468 => x"58200000",
     8469 => x"c3a00000",  8470 => x"379cfff4",  8471 => x"5b8b000c",
     8472 => x"5b8c0008",  8473 => x"5b9d0004",  8474 => x"780b0001",
     8475 => x"396b7810",  8476 => x"29610000",  8477 => x"340c0001",
     8478 => x"442c0010",  8479 => x"34020002",  8480 => x"4422009d",
     8481 => x"34020000",  8482 => x"5c2000a5",  8483 => x"78010001",
     8484 => x"38214c78",  8485 => x"f800105a",  8486 => x"78010001",
     8487 => x"38217814",  8488 => x"58200000",  8489 => x"78010001",
     8490 => x"3821780c",  8491 => x"58200000",  8492 => x"596c0000",
     8493 => x"e000008e",  8494 => x"f8002073",  8495 => x"34020000",
     8496 => x"48010097",  8497 => x"3402001b",  8498 => x"44220008",
     8499 => x"78020001",  8500 => x"38427818",  8501 => x"28430000",
     8502 => x"6424005b",  8503 => x"00650010",  8504 => x"a0a42000",
     8505 => x"44800006",  8506 => x"78010001",  8507 => x"38217818",
     8508 => x"78020001",  8509 => x"58220000",  8510 => x"e0000003",
     8511 => x"b8230800",  8512 => x"58410000",  8513 => x"78010001",
     8514 => x"38217818",  8515 => x"282b0000",  8516 => x"34020001",
     8517 => x"216100ff",  8518 => x"44200081",  8519 => x"3401007e",
     8520 => x"4561002e",  8521 => x"49610006",  8522 => x"34010009",
     8523 => x"4561006d",  8524 => x"3401000d",  8525 => x"5d610042",
     8526 => x"e0000020",  8527 => x"78020001",  8528 => x"38425774",
     8529 => x"28410000",  8530 => x"45610010",  8531 => x"78020001",
     8532 => x"38425778",  8533 => x"28410000",  8534 => x"45610004",
     8535 => x"3401007f",  8536 => x"5d610037",  8537 => x"e0000027",
     8538 => x"78010001",  8539 => x"38217814",  8540 => x"28220000",
     8541 => x"4c02005b",  8542 => x"3442ffff",  8543 => x"58220000",
     8544 => x"34010044",  8545 => x"e000000b",  8546 => x"78010001",
     8547 => x"78020001",  8548 => x"38217814",  8549 => x"3842780c",
     8550 => x"28230000",  8551 => x"28420000",  8552 => x"4c620050",
     8553 => x"34630001",  8554 => x"58230000",  8555 => x"34010043",
     8556 => x"fbffff30",  8557 => x"e000004b",  8558 => x"78010001",
     8559 => x"38214adc",  8560 => x"f800100f",  8561 => x"78010001",
     8562 => x"38217810",  8563 => x"34020002",  8564 => x"58220000",
     8565 => x"e0000043",  8566 => x"78010001",  8567 => x"78020001",
     8568 => x"38217814",  8569 => x"3842780c",  8570 => x"28210000",
     8571 => x"28420000",  8572 => x"4422003c",  8573 => x"fbffff7a",
     8574 => x"34010050",  8575 => x"e3ffffed",  8576 => x"780b0001",
     8577 => x"396b7814",  8578 => x"29610000",  8579 => x"4c010035",
     8580 => x"34010044",  8581 => x"fbffff17",  8582 => x"34010050",
     8583 => x"fbffff15",  8584 => x"29610000",  8585 => x"3421ffff",
     8586 => x"fbffff6d",  8587 => x"29610000",  8588 => x"3421ffff",
     8589 => x"59610000",  8590 => x"e000002a",  8591 => x"78010001",
     8592 => x"a1610800",  8593 => x"5c200027",  8594 => x"78010001",
     8595 => x"3821780c",  8596 => x"28240000",  8597 => x"3401004f",
     8598 => x"48810022",  8599 => x"78010001",  8600 => x"38217814",
     8601 => x"28230000",  8602 => x"44640008",  8603 => x"78020001",
     8604 => x"34610001",  8605 => x"384277b8",  8606 => x"b4220800",
     8607 => x"b4621000",  8608 => x"c8831800",  8609 => x"f80029ca",
     8610 => x"78010001",  8611 => x"38217814",  8612 => x"28230000",
     8613 => x"78020001",  8614 => x"384277b8",  8615 => x"b4431000",
     8616 => x"304b0000",  8617 => x"34620001",  8618 => x"58220000",
     8619 => x"78010001",  8620 => x"3821780c",  8621 => x"28220000",
     8622 => x"34420001",  8623 => x"58220000",  8624 => x"34010040",
     8625 => x"fbfffeeb",  8626 => x"78020001",  8627 => x"38427818",
     8628 => x"28420000",  8629 => x"78010001",  8630 => x"38214c80",
     8631 => x"f8000fc8",  8632 => x"78010001",  8633 => x"38217818",
     8634 => x"58200000",  8635 => x"34020001",  8636 => x"e000000b",
     8637 => x"78020001",  8638 => x"3842780c",  8639 => x"28420000",
     8640 => x"78010001",  8641 => x"382177b8",  8642 => x"b4220800",
     8643 => x"30200000",  8644 => x"fbfffee1",  8645 => x"59600000",
     8646 => x"e3fffff5",  8647 => x"b8400800",  8648 => x"2b9d0004",
     8649 => x"2b8b000c",  8650 => x"2b8c0008",  8651 => x"379c000c",
     8652 => x"c3a00000",  8653 => x"34030000",  8654 => x"34070009",
     8655 => x"34050005",  8656 => x"e0000014",  8657 => x"3486ffd0",
     8658 => x"20c800ff",  8659 => x"55070004",  8660 => x"3c630004",
     8661 => x"b4c31800",  8662 => x"e000000d",  8663 => x"3486ffbf",
     8664 => x"20c600ff",  8665 => x"54c50004",  8666 => x"3c630004",
     8667 => x"3484ffc9",  8668 => x"e0000006",  8669 => x"3486ff9f",
     8670 => x"20c600ff",  8671 => x"54c50007",  8672 => x"3c630004",
     8673 => x"3484ffa9",  8674 => x"b4831800",  8675 => x"34210001",
     8676 => x"40240000",  8677 => x"5c80ffec",  8678 => x"58430000",
     8679 => x"c3a00000",  8680 => x"34030000",  8681 => x"34050009",
     8682 => x"e0000007",  8683 => x"3484ffd0",  8684 => x"208600ff",
     8685 => x"54c50006",  8686 => x"0863000a",  8687 => x"34210001",
     8688 => x"b4831800",  8689 => x"40240000",  8690 => x"5c80fff9",
     8691 => x"58430000",  8692 => x"c3a00000",  8693 => x"379cffec",
     8694 => x"5b8b0014",  8695 => x"5b8c0010",  8696 => x"5b8d000c",
     8697 => x"5b8e0008",  8698 => x"5b9d0004",  8699 => x"78010001",
     8700 => x"38218bec",  8701 => x"40210000",  8702 => x"4420001b",
     8703 => x"780b0001",  8704 => x"780e0001",  8705 => x"780d0001",
     8706 => x"340c0000",  8707 => x"396b77b8",  8708 => x"39ce780c",
     8709 => x"39ad4c9c",  8710 => x"b9600800",  8711 => x"34020050",
     8712 => x"b9801800",  8713 => x"f8001b89",  8714 => x"59c10000",
     8715 => x"48200006",  8716 => x"5d80000d",  8717 => x"78010001",
     8718 => x"38214c84",  8719 => x"f8000f70",  8720 => x"e0000009",
     8721 => x"b5610800",  8722 => x"3020ffff",  8723 => x"b9601000",
     8724 => x"b9a00800",  8725 => x"f8000f6a",  8726 => x"fbfffe8f",
     8727 => x"340c0001",  8728 => x"e3ffffee",  8729 => x"2b9d0004",
     8730 => x"2b8b0014",  8731 => x"2b8c0010",  8732 => x"2b8d000c",
     8733 => x"2b8e0008",  8734 => x"379c0014",  8735 => x"c3a00000",
     8736 => x"379cfff8",  8737 => x"5b8b0008",  8738 => x"5b9d0004",
     8739 => x"78010001",  8740 => x"38218f90",  8741 => x"28210000",
     8742 => x"78030001",  8743 => x"38635e78",  8744 => x"28620000",
     8745 => x"282b000c",  8746 => x"78030001",  8747 => x"78010001",
     8748 => x"38634cc4",  8749 => x"38214cac",  8750 => x"f8000f51",
     8751 => x"78050001",  8752 => x"78030001",  8753 => x"78040001",
     8754 => x"38a55e7c",  8755 => x"38635e80",  8756 => x"38845e84",
     8757 => x"28a20000",  8758 => x"28630000",  8759 => x"28840000",
     8760 => x"78010001",  8761 => x"38214ce4",  8762 => x"f8000f45",
     8763 => x"216b000f",  8764 => x"356b0001",  8765 => x"78010001",
     8766 => x"34020080",  8767 => x"3d6b0004",  8768 => x"38214cf8",
     8769 => x"34030800",  8770 => x"f8000f3d",  8771 => x"3561ff80",
     8772 => x"3402000f",  8773 => x"50410006",  8774 => x"78010001",
     8775 => x"38214d20",  8776 => x"b9601000",  8777 => x"35630010",
     8778 => x"f8000f35",  8779 => x"34010000",  8780 => x"2b9d0004",
     8781 => x"2b8b0008",  8782 => x"379c0008",  8783 => x"c3a00000",
     8784 => x"379cfff8",  8785 => x"5b8b0008",  8786 => x"5b9d0004",
     8787 => x"b8205800",  8788 => x"28210000",  8789 => x"78020001",
     8790 => x"38424d50",  8791 => x"f800299a",  8792 => x"5c200003",
     8793 => x"fbffe11a",  8794 => x"e0000008",  8795 => x"29610000",
     8796 => x"78020001",  8797 => x"38424d58",  8798 => x"f8002993",
     8799 => x"3402ffea",  8800 => x"5c200003",  8801 => x"fbffe138",
     8802 => x"b8201000",  8803 => x"b8400800",  8804 => x"2b9d0004",
     8805 => x"2b8b0008",  8806 => x"379c0008",  8807 => x"c3a00000",
     8808 => x"379cfff8",  8809 => x"5b8b0008",  8810 => x"5b9d0004",
     8811 => x"b8205800",  8812 => x"28210000",  8813 => x"78020001",
     8814 => x"38424d60",  8815 => x"f8002982",  8816 => x"34020001",
     8817 => x"44200018",  8818 => x"29610000",  8819 => x"78020001",
     8820 => x"38424118",  8821 => x"f800297c",  8822 => x"34020002",
     8823 => x"44200012",  8824 => x"29610000",  8825 => x"78020001",
     8826 => x"38423c30",  8827 => x"f8002976",  8828 => x"34020003",
     8829 => x"4420000c",  8830 => x"fbffe0f1",  8831 => x"3c210002",
     8832 => x"78020001",  8833 => x"38425a54",  8834 => x"b4411000",
     8835 => x"28420000",  8836 => x"78010001",  8837 => x"3821461c",
     8838 => x"f8000ef9",  8839 => x"34010000",  8840 => x"e0000003",
     8841 => x"b8400800",  8842 => x"fbffe135",  8843 => x"2b9d0004",
     8844 => x"2b8b0008",  8845 => x"379c0008",  8846 => x"c3a00000",
     8847 => x"379cfff0",  8848 => x"5b8b0010",  8849 => x"5b8c000c",
     8850 => x"5b8d0008",  8851 => x"5b9d0004",  8852 => x"78010001",
     8853 => x"38214d78",  8854 => x"780b0001",  8855 => x"780d0001",
     8856 => x"780c0001",  8857 => x"f8000ee6",  8858 => x"396b7058",
     8859 => x"39ad7108",  8860 => x"398c4d90",  8861 => x"e0000005",
     8862 => x"29620000",  8863 => x"b9800800",  8864 => x"356b0008",
     8865 => x"f8000ede",  8866 => x"55abfffc",  8867 => x"34010000",
     8868 => x"2b9d0004",  8869 => x"2b8b0010",  8870 => x"2b8c000c",
     8871 => x"2b8d0008",  8872 => x"379c0010",  8873 => x"c3a00000",
     8874 => x"379cffec",  8875 => x"5b8b0010",  8876 => x"5b8c000c",
     8877 => x"5b8d0008",  8878 => x"5b9d0004",  8879 => x"340b0000",
     8880 => x"b8406800",  8881 => x"340c0006",  8882 => x"37820014",
     8883 => x"fbffff1a",  8884 => x"2b830014",  8885 => x"b5ab1000",
     8886 => x"356b0001",  8887 => x"30430000",  8888 => x"40220000",
     8889 => x"6442003a",  8890 => x"b4220800",  8891 => x"5d6cfff7",
     8892 => x"2b9d0004",  8893 => x"2b8b0010",  8894 => x"2b8c000c",
     8895 => x"2b8d0008",  8896 => x"379c0014",  8897 => x"c3a00000",
     8898 => x"379cfff8",  8899 => x"5b8b0008",  8900 => x"5b9d0004",
     8901 => x"b8404000",  8902 => x"41030000",  8903 => x"41040001",
     8904 => x"41050002",  8905 => x"41060003",  8906 => x"41070004",
     8907 => x"41080005",  8908 => x"78020001",  8909 => x"38424da0",
     8910 => x"b8205800",  8911 => x"f8000ea2",  8912 => x"b9600800",
     8913 => x"2b9d0004",  8914 => x"2b8b0008",  8915 => x"379c0008",
     8916 => x"c3a00000",  8917 => x"379cffd0",  8918 => x"5b8b0008",
     8919 => x"5b9d0004",  8920 => x"b8205800",  8921 => x"28210000",
     8922 => x"44200005",  8923 => x"78020001",  8924 => x"38424dc0",
     8925 => x"f8002914",  8926 => x"5c200004",  8927 => x"3781002c",
     8928 => x"f8000fa7",  8929 => x"e000002b",  8930 => x"29610000",
     8931 => x"78020001",  8932 => x"38424dc4",  8933 => x"f800290c",
     8934 => x"5c200008",  8935 => x"378b002c",  8936 => x"b9600800",
     8937 => x"f8000f9e",  8938 => x"b9601000",  8939 => x"34010000",
     8940 => x"f8001b01",  8941 => x"e000001f",  8942 => x"29610000",
     8943 => x"78020001",  8944 => x"38424dcc",  8945 => x"f8002900",
     8946 => x"5c20000b",  8947 => x"29630004",  8948 => x"44610009",
     8949 => x"378b002c",  8950 => x"b8600800",  8951 => x"b9601000",
     8952 => x"fbffffb2",  8953 => x"b9600800",  8954 => x"f8000f79",
     8955 => x"f8001074",  8956 => x"e0000010",  8957 => x"29610000",
     8958 => x"78020001",  8959 => x"38424dd0",  8960 => x"f80028f1",
     8961 => x"b8201800",  8962 => x"3402ffea",  8963 => x"5c200011",
     8964 => x"29610004",  8965 => x"4423000f",  8966 => x"378b002c",
     8967 => x"b9601000",  8968 => x"fbffffa2",  8969 => x"34010000",
     8970 => x"b9601000",  8971 => x"f8001ad9",  8972 => x"3782002c",
     8973 => x"3781000c",  8974 => x"fbffffb4",  8975 => x"b8201000",
     8976 => x"78010001",  8977 => x"38214dd8",  8978 => x"f8000e6d",
     8979 => x"34020000",  8980 => x"b8400800",  8981 => x"2b9d0004",
     8982 => x"2b8b0008",  8983 => x"379c0030",  8984 => x"c3a00000",
     8985 => x"379cffe8",  8986 => x"5b8b0018",  8987 => x"5b8c0014",
     8988 => x"5b8d0010",  8989 => x"5b8e000c",  8990 => x"5b8f0008",
     8991 => x"5b9d0004",  8992 => x"28210000",  8993 => x"44200010",
     8994 => x"78020001",  8995 => x"38424df0",  8996 => x"f80028cd",
     8997 => x"5c20000c",  8998 => x"78010001",  8999 => x"78020001",
     9000 => x"38217114",  9001 => x"38427264",  9002 => x"e0000005",
     9003 => x"58200018",  9004 => x"58200014",  9005 => x"58200010",
     9006 => x"3421001c",  9007 => x"5441fffc",  9008 => x"e0000018",
     9009 => x"78010001",  9010 => x"38214df8",  9011 => x"780b0001",
     9012 => x"780d0001",  9013 => x"780c0001",  9014 => x"f8000e49",
     9015 => x"396b7114",  9016 => x"39ad7264",  9017 => x"398c4e20",
     9018 => x"e000000d",  9019 => x"29610018",  9020 => x"340203e8",
     9021 => x"296f0010",  9022 => x"f8002793",  9023 => x"296e0014",
     9024 => x"29650000",  9025 => x"b8202000",  9026 => x"b9e01000",
     9027 => x"b9800800",  9028 => x"b9c01800",  9029 => x"f8000e3a",
     9030 => x"356b001c",  9031 => x"55abfff4",  9032 => x"34010000",
     9033 => x"2b9d0004",  9034 => x"2b8b0018",  9035 => x"2b8c0014",
     9036 => x"2b8d0010",  9037 => x"2b8e000c",  9038 => x"2b8f0008",
     9039 => x"379c0018",  9040 => x"c3a00000",  9041 => x"379cfff8",
     9042 => x"5b9d0004",  9043 => x"b8201000",  9044 => x"28210000",
     9045 => x"4420000d",  9046 => x"28420004",  9047 => x"5c40000b",
     9048 => x"37820008",  9049 => x"fbfffe8f",  9050 => x"2b820008",
     9051 => x"78010001",  9052 => x"38215e88",  9053 => x"084203e8",
     9054 => x"58220000",  9055 => x"78010001",  9056 => x"38214adc",
     9057 => x"e0000003",  9058 => x"78010001",  9059 => x"38214e40",
     9060 => x"f8000e1b",  9061 => x"34010000",  9062 => x"2b9d0004",
     9063 => x"379c0008",  9064 => x"c3a00000",  9065 => x"379cfff8",
     9066 => x"5b8b0008",  9067 => x"5b9d0004",  9068 => x"b8205800",
     9069 => x"28210000",  9070 => x"5c200011",  9071 => x"78010001",
     9072 => x"38218f7c",  9073 => x"28220000",  9074 => x"340b0000",
     9075 => x"64420000",  9076 => x"58220000",  9077 => x"78010001",
     9078 => x"38218c1c",  9079 => x"28230000",  9080 => x"3463ffff",
     9081 => x"58230000",  9082 => x"5c4b002b",  9083 => x"78010001",
     9084 => x"38214e64",  9085 => x"f8000e02",  9086 => x"e0000027",
     9087 => x"78020001",  9088 => x"38424e78",  9089 => x"f8002870",
     9090 => x"5c200007",  9091 => x"f8000f6d",  9092 => x"b8201000",
     9093 => x"78010001",  9094 => x"382154ac",  9095 => x"f8000df8",
     9096 => x"e000001c",  9097 => x"29610000",  9098 => x"78020001",
     9099 => x"38423cd0",  9100 => x"f8002865",  9101 => x"5c20000b",
     9102 => x"78010001",  9103 => x"38218f7c",  9104 => x"34020001",
     9105 => x"58220000",  9106 => x"78010001",  9107 => x"38218c1c",
     9108 => x"28220000",  9109 => x"3442ffff",  9110 => x"58220000",
     9111 => x"e000000d",  9112 => x"29610000",  9113 => x"78020001",
     9114 => x"38424e7c",  9115 => x"f8002856",  9116 => x"340bffea",
     9117 => x"5c200008",  9118 => x"78010001",  9119 => x"38218f7c",
     9120 => x"58200000",  9121 => x"78010001",  9122 => x"38214e64",
     9123 => x"f8000ddc",  9124 => x"340b0000",  9125 => x"b9600800",
     9126 => x"2b9d0004",  9127 => x"2b8b0008",  9128 => x"379c0008",
     9129 => x"c3a00000",  9130 => x"379cffb8",  9131 => x"5b8b0028",
     9132 => x"5b8c0024",  9133 => x"5b8d0020",  9134 => x"5b8e001c",
     9135 => x"5b8f0018",  9136 => x"5b900014",  9137 => x"5b910010",
     9138 => x"5b92000c",  9139 => x"5b930008",  9140 => x"5b9d0004",
     9141 => x"b8205800",  9142 => x"28210000",  9143 => x"442000c8",
     9144 => x"78020001",  9145 => x"38424e9c",  9146 => x"f8002837",
     9147 => x"5c200008",  9148 => x"f80017df",  9149 => x"3403ffff",
     9150 => x"34020000",  9151 => x"5c2300c4",  9152 => x"78010001",
     9153 => x"38214ea4",  9154 => x"e000003c",  9155 => x"29610010",
     9156 => x"44200045",  9157 => x"29610000",  9158 => x"78020001",
     9159 => x"38424eb8",  9160 => x"f8002829",  9161 => x"5c200040",
     9162 => x"29610004",  9163 => x"34020010",  9164 => x"356c0004",
     9165 => x"f8002948",  9166 => x"3c210018",  9167 => x"34030000",
     9168 => x"14210018",  9169 => x"3784002c",  9170 => x"e0000007",
     9171 => x"29820000",  9172 => x"b4832800",  9173 => x"b4431000",
     9174 => x"40420000",  9175 => x"34630001",  9176 => x"30a20000",
     9177 => x"b0601000",  9178 => x"4822fff9",  9179 => x"b4820800",
     9180 => x"34030020",  9181 => x"3404000f",  9182 => x"e0000005",
     9183 => x"34420001",  9184 => x"30230000",  9185 => x"b0401000",
     9186 => x"34210001",  9187 => x"4c82fffc",  9188 => x"29610008",
     9189 => x"f80003b9",  9190 => x"5b810040",  9191 => x"2961000c",
     9192 => x"f80003b6",  9193 => x"5b810044",  9194 => x"29610010",
     9195 => x"f80003b3",  9196 => x"5b81003c",  9197 => x"34020001",
     9198 => x"3781002c",  9199 => x"34030000",  9200 => x"f80017c4",
     9201 => x"3c220018",  9202 => x"3401fffe",  9203 => x"14420018",
     9204 => x"5c410006",  9205 => x"78010001",  9206 => x"38214ebc",
     9207 => x"f8000d88",  9208 => x"3402ffe4",  9209 => x"e000008a",
     9210 => x"3401ffff",  9211 => x"5c410006",  9212 => x"78010001",
     9213 => x"38214ecc",  9214 => x"f8000d81",  9215 => x"3402fffb",
     9216 => x"e0000083",  9217 => x"4c400004",  9218 => x"78010001",
     9219 => x"38214ed8",  9220 => x"e0000023",  9221 => x"78010001",
     9222 => x"38214ef4",  9223 => x"f8000d78",  9224 => x"e0000075",
     9225 => x"29610000",  9226 => x"78020001",  9227 => x"38424f04",
     9228 => x"f80027e5",  9229 => x"5c200030",  9230 => x"78100001",
     9231 => x"780f0001",  9232 => x"780e0001",  9233 => x"340c0000",
     9234 => x"34110000",  9235 => x"3792002c",  9236 => x"3a104f20",
     9237 => x"3793003c",  9238 => x"39ef4c80",  9239 => x"39ce4f28",
     9240 => x"ba400800",  9241 => x"34020000",  9242 => x"b9801800",
     9243 => x"f8001799",  9244 => x"3c2b0018",  9245 => x"156b0018",
     9246 => x"5d600005",  9247 => x"78010001",  9248 => x"38214f0c",
     9249 => x"f8000d5e",  9250 => x"e000005b",  9251 => x"4d600007",
     9252 => x"78010001",  9253 => x"38214ed8",  9254 => x"b9601000",
     9255 => x"f8000d58",  9256 => x"3402fff2",  9257 => x"e000005a",
     9258 => x"358c0001",  9259 => x"ba000800",  9260 => x"b9801000",
     9261 => x"f8000d52",  9262 => x"ba406800",  9263 => x"41a20000",
     9264 => x"b9e00800",  9265 => x"35ad0001",  9266 => x"f8000d4d",
     9267 => x"5db3fffc",  9268 => x"2b820040",  9269 => x"2b830044",
     9270 => x"2b84003c",  9271 => x"36310001",  9272 => x"b9c00800",
     9273 => x"b2208800",  9274 => x"f8000d45",  9275 => x"4971ffdd",
     9276 => x"e0000041",  9277 => x"29610000",  9278 => x"78020001",
     9279 => x"38424f48",  9280 => x"f80027b1",  9281 => x"5c200032",
     9282 => x"f8001358",  9283 => x"3c2c0018",  9284 => x"3401ffed",
     9285 => x"158c0018",  9286 => x"5d810006",  9287 => x"78010001",
     9288 => x"38214f50",  9289 => x"f8000d36",  9290 => x"3402ffed",
     9291 => x"e0000038",  9292 => x"780b0001",  9293 => x"396b8c24",
     9294 => x"780d0001",  9295 => x"3401fffb",  9296 => x"356e0010",
     9297 => x"39ad4c80",  9298 => x"5d810004",  9299 => x"78010001",
     9300 => x"38214f5c",  9301 => x"e3ffffa9",  9302 => x"41620000",
     9303 => x"b9a00800",  9304 => x"356b0001",  9305 => x"f8000d26",
     9306 => x"5d6efffc",  9307 => x"78010001",  9308 => x"38214adc",
     9309 => x"f8000d22",  9310 => x"3401fffa",  9311 => x"5d810006",
     9312 => x"78010001",  9313 => x"38214f6c",  9314 => x"f8000d1d",
     9315 => x"3402fffa",  9316 => x"e000001f",  9317 => x"78020001",
     9318 => x"78030001",  9319 => x"78040001",  9320 => x"38428bb8",
     9321 => x"38638bbc",  9322 => x"38846d1c",  9323 => x"28420000",
     9324 => x"28630000",  9325 => x"28840000",  9326 => x"78010001",
     9327 => x"38214f84",  9328 => x"f8000d0f",  9329 => x"b9801000",
     9330 => x"e0000011",  9331 => x"29610004",  9332 => x"4420000b",
     9333 => x"29610000",  9334 => x"78020001",  9335 => x"38424fac",
     9336 => x"f8002779",  9337 => x"5c200006",  9338 => x"29610004",
     9339 => x"f8000323",  9340 => x"f8000ec1",  9341 => x"34020000",
     9342 => x"e0000005",  9343 => x"78010001",  9344 => x"38214e88",
     9345 => x"f8000cfe",  9346 => x"3402ffea",  9347 => x"b8400800",
     9348 => x"2b9d0004",  9349 => x"2b8b0028",  9350 => x"2b8c0024",
     9351 => x"2b8d0020",  9352 => x"2b8e001c",  9353 => x"2b8f0018",
     9354 => x"2b900014",  9355 => x"2b910010",  9356 => x"2b92000c",
     9357 => x"2b930008",  9358 => x"379c0048",  9359 => x"c3a00000",
     9360 => x"379cffe8",  9361 => x"5b8b0010",  9362 => x"5b8c000c",
     9363 => x"5b8d0008",  9364 => x"5b9d0004",  9365 => x"b8205800",
     9366 => x"28210000",  9367 => x"78020001",  9368 => x"38424fb4",
     9369 => x"f8002758",  9370 => x"5c200011",  9371 => x"2963000c",
     9372 => x"3402ffea",  9373 => x"44610086",  9374 => x"29610004",
     9375 => x"f80002ff",  9376 => x"b8206800",  9377 => x"29610008",
     9378 => x"f80002fc",  9379 => x"b8206000",  9380 => x"2961000c",
     9381 => x"f80002f9",  9382 => x"b8201800",  9383 => x"b9801000",
     9384 => x"b9a00800",  9385 => x"f80021ed",  9386 => x"e0000078",
     9387 => x"29610000",  9388 => x"78020001",  9389 => x"38424fbc",
     9390 => x"f8002743",  9391 => x"b8201800",  9392 => x"5c200007",
     9393 => x"29610004",  9394 => x"3402ffea",  9395 => x"44230070",
     9396 => x"f80002ea",  9397 => x"f80022ab",  9398 => x"e0000060",
     9399 => x"29610000",  9400 => x"78020001",  9401 => x"38424e80",
     9402 => x"f8002737",  9403 => x"5c200003",  9404 => x"f800233e",
     9405 => x"e0000065",  9406 => x"29610000",  9407 => x"78020001",
     9408 => x"38424fc0",  9409 => x"f8002730",  9410 => x"5c20000d",
     9411 => x"29630008",  9412 => x"3402ffea",  9413 => x"4461005e",
     9414 => x"29610004",  9415 => x"f80002d7",  9416 => x"b8206000",
     9417 => x"29610008",  9418 => x"f80002d4",  9419 => x"b8201000",
     9420 => x"b9800800",  9421 => x"f80022a4",  9422 => x"e0000054",
     9423 => x"29610000",  9424 => x"78020001",  9425 => x"38424fc4",
     9426 => x"f800271f",  9427 => x"b8201800",  9428 => x"5c20000e",
     9429 => x"29610004",  9430 => x"3402ffea",  9431 => x"4423004c",
     9432 => x"f80002c6",  9433 => x"37820018",  9434 => x"37830014",
     9435 => x"f80022be",  9436 => x"2b820018",  9437 => x"2b830014",
     9438 => x"78010001",  9439 => x"38214fc8",  9440 => x"f8000c9f",
     9441 => x"e0000041",  9442 => x"29610000",  9443 => x"78020001",
     9444 => x"38424d50",  9445 => x"f800270c",  9446 => x"b8201800",
     9447 => x"5c200007",  9448 => x"29610004",  9449 => x"3402ffea",
     9450 => x"44230039",  9451 => x"f80002b3",  9452 => x"f8002256",
     9453 => x"e0000035",  9454 => x"29610000",  9455 => x"78020001",
     9456 => x"38424d58",  9457 => x"f8002700",  9458 => x"b8201800",
     9459 => x"5c200007",  9460 => x"29610004",  9461 => x"3402ffea",
     9462 => x"4423002d",  9463 => x"f80002a7",  9464 => x"f800225b",
     9465 => x"e0000029",  9466 => x"29610000",  9467 => x"78020001",
     9468 => x"38424fd0",  9469 => x"f80026f4",  9470 => x"5c20000d",
     9471 => x"29630008",  9472 => x"3402ffea",  9473 => x"44610022",
     9474 => x"29610004",  9475 => x"f800029b",  9476 => x"b8206000",
     9477 => x"29610008",  9478 => x"f8000298",  9479 => x"b8201000",
     9480 => x"b9800800",  9481 => x"f8002361",  9482 => x"e0000018",
     9483 => x"29610000",  9484 => x"78020001",  9485 => x"38424fd8",
     9486 => x"f80026e3",  9487 => x"b8201800",  9488 => x"5c20000b",
     9489 => x"29610004",  9490 => x"3402ffea",  9491 => x"44230010",
     9492 => x"f800028a",  9493 => x"f8002346",  9494 => x"b8201000",
     9495 => x"78010001",  9496 => x"38214c58",  9497 => x"f8000c66",
     9498 => x"e0000008",  9499 => x"29610000",  9500 => x"78020001",
     9501 => x"38424fe0",  9502 => x"f80026d3",  9503 => x"3402ffea",
     9504 => x"5c200003",  9505 => x"f80023f8",  9506 => x"34020000",
     9507 => x"b8400800",  9508 => x"2b9d0004",  9509 => x"2b8b0010",
     9510 => x"2b8c000c",  9511 => x"2b8d0008",  9512 => x"379c0018",
     9513 => x"c3a00000",  9514 => x"379cfff0",  9515 => x"5b8b000c",
     9516 => x"5b8c0008",  9517 => x"5b9d0004",  9518 => x"b8205800",
     9519 => x"28210000",  9520 => x"4420000b",  9521 => x"78020001",
     9522 => x"38424ff0",  9523 => x"f80026be",  9524 => x"b8206000",
     9525 => x"5c200006",  9526 => x"37810010",  9527 => x"f80013ae",
     9528 => x"340bffff",  9529 => x"49810021",  9530 => x"e000001c",
     9531 => x"29610000",  9532 => x"340b0000",  9533 => x"5c20001d",
     9534 => x"37810010",  9535 => x"34020000",  9536 => x"f800174d",
     9537 => x"4d61000a",  9538 => x"2b820010",  9539 => x"78010001",
     9540 => x"38214ff8",  9541 => x"f8000c3a",  9542 => x"2b820010",
     9543 => x"78010001",  9544 => x"38215e90",  9545 => x"58220000",
     9546 => x"e0000010",  9547 => x"78010001",  9548 => x"38215020",
     9549 => x"f8000c32",  9550 => x"37810010",  9551 => x"f8001396",
     9552 => x"340bffff",  9553 => x"48010009",  9554 => x"2b820010",
     9555 => x"78010001",  9556 => x"38215e90",  9557 => x"58220000",
     9558 => x"37810010",  9559 => x"34020001",  9560 => x"f8001735",
     9561 => x"b8205800",  9562 => x"b9600800",  9563 => x"2b9d0004",
     9564 => x"2b8b000c",  9565 => x"2b8c0008",  9566 => x"379c0010",
     9567 => x"c3a00000",  9568 => x"379cffe8",  9569 => x"5b8b000c",
     9570 => x"5b8c0008",  9571 => x"5b9d0004",  9572 => x"b8205800",
     9573 => x"37820018",  9574 => x"37810010",  9575 => x"f8001553",
     9576 => x"29610008",  9577 => x"44200014",  9578 => x"29610000",
     9579 => x"78020001",  9580 => x"38424dcc",  9581 => x"f8002684",
     9582 => x"5c20000f",  9583 => x"fbffde00",  9584 => x"34030003",
     9585 => x"3402fff0",  9586 => x"44230040",  9587 => x"29610004",
     9588 => x"f800022a",  9589 => x"b8206000",  9590 => x"29610008",
     9591 => x"f8000227",  9592 => x"b8201800",  9593 => x"b9801000",
     9594 => x"1581001f",  9595 => x"34040003",  9596 => x"e0000020",
     9597 => x"29610000",  9598 => x"4420000f",  9599 => x"78020001",
     9600 => x"38425054",  9601 => x"f8002670",  9602 => x"5c20000b",
     9603 => x"fbffddec",  9604 => x"34020003",  9605 => x"44220023",
     9606 => x"29610004",  9607 => x"f8000217",  9608 => x"b8201000",
     9609 => x"34030000",  9610 => x"1421001f",  9611 => x"34040001",
     9612 => x"e0000010",  9613 => x"29610000",  9614 => x"44200010",
     9615 => x"78020001",  9616 => x"3842505c",  9617 => x"f8002660",
     9618 => x"5c20000c",  9619 => x"fbffdddc",  9620 => x"34020003",
     9621 => x"44220013",  9622 => x"29610004",  9623 => x"f8000207",
     9624 => x"b8201800",  9625 => x"34020000",  9626 => x"34010000",
     9627 => x"34040002",  9628 => x"f80014fe",  9629 => x"e0000014",
     9630 => x"29610000",  9631 => x"44200009",  9632 => x"78020001",
     9633 => x"38425064",  9634 => x"f800264f",  9635 => x"5c200005",
     9636 => x"78010001",  9637 => x"38214fc8",  9638 => x"2b820014",
     9639 => x"e0000008",  9640 => x"2b820014",  9641 => x"2b810010",
     9642 => x"34030000",  9643 => x"f80000f4",  9644 => x"b8201000",
     9645 => x"78010001",  9646 => x"38215068",  9647 => x"2b830018",
     9648 => x"f8000bcf",  9649 => x"34020000",  9650 => x"b8400800",
     9651 => x"2b9d0004",  9652 => x"2b8b000c",  9653 => x"2b8c0008",
     9654 => x"379c0018",  9655 => x"c3a00000",  9656 => x"78010001",
     9657 => x"38217268",  9658 => x"34020001",  9659 => x"58220000",
     9660 => x"34010000",  9661 => x"c3a00000",  9662 => x"379cfffc",
     9663 => x"5b9d0004",  9664 => x"f800120e",  9665 => x"34010000",
     9666 => x"2b9d0004",  9667 => x"379c0004",  9668 => x"c3a00000",
     9669 => x"379cfff8",  9670 => x"5b8b0008",  9671 => x"5b9d0004",
     9672 => x"b8205800",  9673 => x"28210000",  9674 => x"4420000c",
     9675 => x"78020001",  9676 => x"38425098",  9677 => x"f8002624",
     9678 => x"5c200008",  9679 => x"34010001",  9680 => x"fbffe890",
     9681 => x"78010001",  9682 => x"38215e8c",  9683 => x"34020001",
     9684 => x"58220000",  9685 => x"e000000b",  9686 => x"29610000",
     9687 => x"44200009",  9688 => x"78020001",  9689 => x"384250a0",
     9690 => x"f8002617",  9691 => x"5c200005",  9692 => x"fbffe884",
     9693 => x"78010001",  9694 => x"38215e8c",  9695 => x"58200000",
     9696 => x"78010001",  9697 => x"38215e8c",  9698 => x"28210000",
     9699 => x"78020001",  9700 => x"38425094",  9701 => x"44200003",
     9702 => x"78020001",  9703 => x"38425090",  9704 => x"78010001",
     9705 => x"382150a8",  9706 => x"f8000b95",  9707 => x"34010000",
     9708 => x"2b9d0004",  9709 => x"2b8b0008",  9710 => x"379c0008",
     9711 => x"c3a00000",  9712 => x"379cffec",  9713 => x"5b8b0010",
     9714 => x"5b8c000c",  9715 => x"5b8d0008",  9716 => x"5b9d0004",
     9717 => x"340b0000",  9718 => x"b8406800",  9719 => x"340c0004",
     9720 => x"37820014",  9721 => x"fbfffbef",  9722 => x"2b830014",
     9723 => x"b5ab1000",  9724 => x"356b0001",  9725 => x"30430000",
     9726 => x"40220000",  9727 => x"6442002e",  9728 => x"b4220800",
     9729 => x"5d6cfff7",  9730 => x"2b9d0004",  9731 => x"2b8b0010",
     9732 => x"2b8c000c",  9733 => x"2b8d0008",  9734 => x"379c0014",
     9735 => x"c3a00000",  9736 => x"379cfff8",  9737 => x"5b8b0008",
     9738 => x"5b9d0004",  9739 => x"b8403000",  9740 => x"40c30000",
     9741 => x"40c40001",  9742 => x"40c50002",  9743 => x"40c60003",
     9744 => x"78020001",  9745 => x"384250c4",  9746 => x"b8205800",
     9747 => x"f8000b5e",  9748 => x"b9600800",  9749 => x"2b9d0004",
     9750 => x"2b8b0008",  9751 => x"379c0008",  9752 => x"c3a00000",
     9753 => x"379cffe0",  9754 => x"5b8b0008",  9755 => x"5b9d0004",
     9756 => x"b8205800",  9757 => x"28210000",  9758 => x"44200005",
     9759 => x"78020001",  9760 => x"38424dc0",  9761 => x"f80025d0",
     9762 => x"5c200004",  9763 => x"37810020",  9764 => x"f80004bb",
     9765 => x"e0000012",  9766 => x"29610000",  9767 => x"78020001",
     9768 => x"38424dcc",  9769 => x"f80025c8",  9770 => x"b8201800",
     9771 => x"3402ffea",  9772 => x"5c200024",  9773 => x"29610004",
     9774 => x"44230022",  9775 => x"78020001",  9776 => x"38427a80",
     9777 => x"34030002",  9778 => x"58430000",  9779 => x"37820020",
     9780 => x"fbffffbc",  9781 => x"37810020",  9782 => x"f80004b2",
     9783 => x"378b000c",  9784 => x"37820020",  9785 => x"b9600800",
     9786 => x"fbffffce",  9787 => x"78010001",  9788 => x"38217a80",
     9789 => x"28210000",  9790 => x"34020001",  9791 => x"44220009",
     9792 => x"44200004",  9793 => x"34020002",  9794 => x"5c22000d",
     9795 => x"e0000008",  9796 => x"78010001",  9797 => x"382150d0",
     9798 => x"f8000b39",  9799 => x"e0000008",  9800 => x"78010001",
     9801 => x"382150ec",  9802 => x"e0000003",  9803 => x"78010001",
     9804 => x"3821510c",  9805 => x"b9601000",  9806 => x"f8000b31",
     9807 => x"34020000",  9808 => x"b8400800",  9809 => x"2b9d0004",
     9810 => x"2b8b0008",  9811 => x"379c0020",  9812 => x"c3a00000",
     9813 => x"379cfffc",  9814 => x"5b9d0004",  9815 => x"28210000",
     9816 => x"44200005",  9817 => x"fbffdc1f",  9818 => x"78020001",
     9819 => x"3842727c",  9820 => x"58410000",  9821 => x"78020001",
     9822 => x"3842727c",  9823 => x"28420000",  9824 => x"78010001",
     9825 => x"38215134",  9826 => x"f8000b1d",  9827 => x"34010000",
     9828 => x"2b9d0004",  9829 => x"379c0004",  9830 => x"c3a00000",
     9831 => x"379cfff4",  9832 => x"5b8b000c",  9833 => x"5b8c0008",
     9834 => x"5b9d0004",  9835 => x"b8205800",  9836 => x"28210000",
     9837 => x"4420000b",  9838 => x"78020001",  9839 => x"38424e9c",
     9840 => x"f8002581",  9841 => x"b8206000",  9842 => x"5c200006",
     9843 => x"f800164f",  9844 => x"4c2c0025",  9845 => x"78010001",
     9846 => x"38215154",  9847 => x"e000000e",  9848 => x"29610004",
     9849 => x"44200011",  9850 => x"29610000",  9851 => x"78020001",
     9852 => x"38424eb8",  9853 => x"f8002574",  9854 => x"b8206000",
     9855 => x"5c20000b",  9856 => x"b9600800",  9857 => x"f8001656",
     9858 => x"4c2c0005",  9859 => x"78010001",  9860 => x"38215174",
     9861 => x"f8000afa",  9862 => x"e0000013",  9863 => x"78010001",
     9864 => x"38215190",  9865 => x"e3fffffc",  9866 => x"29610000",
     9867 => x"44200007",  9868 => x"78020001",  9869 => x"38424f04",
     9870 => x"f8002563",  9871 => x"5c200003",  9872 => x"f80016c1",
     9873 => x"e0000008",  9874 => x"29610000",  9875 => x"44200006",
     9876 => x"78020001",  9877 => x"38425198",  9878 => x"f800255b",
     9879 => x"5c200002",  9880 => x"fbfffb5d",  9881 => x"34010000",
     9882 => x"2b9d0004",  9883 => x"2b8b000c",  9884 => x"2b8c0008",
     9885 => x"379c000c",  9886 => x"c3a00000",  9887 => x"379cffd0",
     9888 => x"5b8b0030",  9889 => x"5b8c002c",  9890 => x"5b8d0028",
     9891 => x"5b8e0024",  9892 => x"5b8f0020",  9893 => x"5b90001c",
     9894 => x"5b910018",  9895 => x"5b920014",  9896 => x"5b930010",
     9897 => x"5b94000c",  9898 => x"5b9d0008",  9899 => x"b8609000",
     9900 => x"78030001",  9901 => x"3863577c",  9902 => x"b8406000",
     9903 => x"b8400800",  9904 => x"28620000",  9905 => x"f8002430",
     9906 => x"78030001",  9907 => x"3863577c",  9908 => x"28620000",
     9909 => x"b8205800",  9910 => x"b9800800",  9911 => x"f800241a",
     9912 => x"b820a000",  9913 => x"3402003c",  9914 => x"b9600800",
     9915 => x"f8002426",  9916 => x"34020e10",  9917 => x"b8207800",
     9918 => x"b9600800",  9919 => x"f8002422",  9920 => x"3402003c",
     9921 => x"f8002410",  9922 => x"b8208000",  9923 => x"34020e10",
     9924 => x"b9600800",  9925 => x"f800240c",  9926 => x"b8208800",
     9927 => x"ba807000",  9928 => x"340b07b2",  9929 => x"e000000f",
     9930 => x"3402016d",  9931 => x"5d80000b",  9932 => x"34020064",
     9933 => x"b9600800",  9934 => x"f80023e3",  9935 => x"3402016e",
     9936 => x"5c2c0006",  9937 => x"34020190",  9938 => x"b9600800",
     9939 => x"f80023de",  9940 => x"64220000",  9941 => x"3442016d",
     9942 => x"c9c27000",  9943 => x"356b0001",  9944 => x"216c0003",
     9945 => x"3402016d",  9946 => x"5d80000b",  9947 => x"34020064",
     9948 => x"b9600800",  9949 => x"f80023d4",  9950 => x"3402016e",
     9951 => x"5c2c0006",  9952 => x"34020190",  9953 => x"b9600800",
     9954 => x"f80023cf",  9955 => x"64220000",  9956 => x"3442016d",
     9957 => x"51c2ffe5",  9958 => x"34020064",  9959 => x"b9600800",
     9960 => x"f80023c9",  9961 => x"34020190",  9962 => x"b8209800",
     9963 => x"b9600800",  9964 => x"f80023c5",  9965 => x"78020001",
     9966 => x"340d0000",  9967 => x"64250000",  9968 => x"38425a64",
     9969 => x"e000000d",  9970 => x"34040000",  9971 => x"5d800004",
     9972 => x"34040001",  9973 => x"5e6c0002",  9974 => x"b8a02000",
     9975 => x"0884000c",  9976 => x"b48d2000",  9977 => x"3c840002",
     9978 => x"35ad0001",  9979 => x"b4442000",  9980 => x"28810000",
     9981 => x"c9c17000",  9982 => x"34040000",  9983 => x"5d800004",
     9984 => x"34040001",  9985 => x"5e6c0002",  9986 => x"b8a02000",
     9987 => x"0884000c",  9988 => x"b48d2000",  9989 => x"3c840002",
     9990 => x"b4442000",  9991 => x"28810000",  9992 => x"51c1ffea",
     9993 => x"34010001",  9994 => x"35ce0001",  9995 => x"4641001d",
     9996 => x"780c0001",  9997 => x"34010002",  9998 => x"398c781c",
     9999 => x"46410028", 10000 => x"36810004", 10001 => x"34020007",
    10002 => x"f80023cf", 10003 => x"3c210002", 10004 => x"78130001",
    10005 => x"78020001", 10006 => x"3dad0002", 10007 => x"38425ae0",
    10008 => x"3a735ac4", 10009 => x"b6619800", 10010 => x"b44d6800",
    10011 => x"78120001", 10012 => x"2a630000", 10013 => x"29a40000",
    10014 => x"3a5251a0", 10015 => x"b9800800", 10016 => x"ba401000",
    10017 => x"b9c02800", 10018 => x"b9603000", 10019 => x"ba203800",
    10020 => x"ba004000", 10021 => x"5b8f0004", 10022 => x"f8000a4b",
    10023 => x"e000001a", 10024 => x"78010001", 10025 => x"3dad0002",
    10026 => x"38215ae0", 10027 => x"b42d6800", 10028 => x"29a30000",
    10029 => x"78010001", 10030 => x"78020001", 10031 => x"384251c0",
    10032 => x"b9c02000", 10033 => x"ba202800", 10034 => x"ba003000",
    10035 => x"b9e03800", 10036 => x"3821781c", 10037 => x"f8000a3c",
    10038 => x"e000000b", 10039 => x"78020001", 10040 => x"b9800800",
    10041 => x"384251d8", 10042 => x"b9601800", 10043 => x"35a40001",
    10044 => x"b9c02800", 10045 => x"ba203000", 10046 => x"ba003800",
    10047 => x"b9e04000", 10048 => x"f8000a31", 10049 => x"78010001",
    10050 => x"3821781c", 10051 => x"2b9d0008", 10052 => x"2b8b0030",
    10053 => x"2b8c002c", 10054 => x"2b8d0028", 10055 => x"2b8e0024",
    10056 => x"2b8f0020", 10057 => x"2b90001c", 10058 => x"2b910018",
    10059 => x"2b920014", 10060 => x"2b930010", 10061 => x"2b94000c",
    10062 => x"379c0030", 10063 => x"c3a00000", 10064 => x"379cffdc",
    10065 => x"5b8b0008", 10066 => x"5b9d0004", 10067 => x"5b840014",
    10068 => x"20240080", 10069 => x"64840000", 10070 => x"5b830010",
    10071 => x"78030001", 10072 => x"b8204800", 10073 => x"b8600800",
    10074 => x"34030002", 10075 => x"5b82000c", 10076 => x"b8405800",
    10077 => x"382151f8", 10078 => x"c8641000", 10079 => x"2123007f",
    10080 => x"5b850018", 10081 => x"5b86001c", 10082 => x"5b870020",
    10083 => x"5b880024", 10084 => x"f8000a1b", 10085 => x"37820010",
    10086 => x"b9600800", 10087 => x"f80009f6", 10088 => x"78010001",
    10089 => x"38215204", 10090 => x"f8000a15", 10091 => x"2b9d0004",
    10092 => x"2b8b0008", 10093 => x"379c0024", 10094 => x"c3a00000",
    10095 => x"379cffe0", 10096 => x"5b8b000c", 10097 => x"5b8c0008",
    10098 => x"5b9d0004", 10099 => x"b8404800", 10100 => x"78020001",
    10101 => x"b8205000", 10102 => x"b8400800", 10103 => x"b8605800",
    10104 => x"b9401000", 10105 => x"b9201800", 10106 => x"38215208",
    10107 => x"b8806000", 10108 => x"5b840010", 10109 => x"5b850014",
    10110 => x"5b860018", 10111 => x"5b87001c", 10112 => x"5b880020",
    10113 => x"f80009fe", 10114 => x"21620080", 10115 => x"78030001",
    10116 => x"64420000", 10117 => x"b8600800", 10118 => x"34030002",
    10119 => x"c8621000", 10120 => x"382151f8", 10121 => x"2163007f",
    10122 => x"f80009f5", 10123 => x"37820014", 10124 => x"b9800800",
    10125 => x"f80009d0", 10126 => x"78010001", 10127 => x"38215204",
    10128 => x"f80009ef", 10129 => x"2b9d0004", 10130 => x"2b8b000c",
    10131 => x"2b8c0008", 10132 => x"379c0020", 10133 => x"c3a00000",
    10134 => x"379cfffc", 10135 => x"5b9d0004", 10136 => x"78010001",
    10137 => x"38215214", 10138 => x"f80009e5", 10139 => x"2b9d0004",
    10140 => x"379c0004", 10141 => x"c3a00000", 10142 => x"40240000",
    10143 => x"3402002d", 10144 => x"34030001", 10145 => x"5c820003",
    10146 => x"34210001", 10147 => x"3403ffff", 10148 => x"34020000",
    10149 => x"34050009", 10150 => x"e0000004", 10151 => x"0842000a",
    10152 => x"34210001", 10153 => x"b4821000", 10154 => x"40240000",
    10155 => x"3484ffd0", 10156 => x"208600ff", 10157 => x"50a6fffa",
    10158 => x"88430800", 10159 => x"c3a00000", 10160 => x"379cfff4",
    10161 => x"5b8b000c", 10162 => x"5b8c0008", 10163 => x"5b9d0004",
    10164 => x"b8206000", 10165 => x"f8000f8a", 10166 => x"342b0001",
    10167 => x"f8000f88", 10168 => x"5c2bffff", 10169 => x"b9800800",
    10170 => x"e0000002", 10171 => x"3421ffff", 10172 => x"4820ffff",
    10173 => x"f8000f82", 10174 => x"c82b0800", 10175 => x"2b9d0004",
    10176 => x"2b8b000c", 10177 => x"2b8c0008", 10178 => x"379c000c",
    10179 => x"c3a00000", 10180 => x"379cfff0", 10181 => x"5b8b0010",
    10182 => x"5b8c000c", 10183 => x"5b8d0008", 10184 => x"5b9d0004",
    10185 => x"340b0400", 10186 => x"340c0400", 10187 => x"e0000003",
    10188 => x"b58b6000", 10189 => x"3d6b0001", 10190 => x"b9800800",
    10191 => x"fbffffe1", 10192 => x"4420fffc", 10193 => x"158c0001",
    10194 => x"156b0002", 10195 => x"e0000009", 10196 => x"b56c6800",
    10197 => x"b9a00800", 10198 => x"fbffffda", 10199 => x"5c200002",
    10200 => x"b9a06000", 10201 => x"0161001f", 10202 => x"b42b5800",
    10203 => x"156b0001", 10204 => x"5d60fff8", 10205 => x"78010001",
    10206 => x"3821785c", 10207 => x"582c0000", 10208 => x"78010001",
    10209 => x"b9801000", 10210 => x"3821526c", 10211 => x"f800099c",
    10212 => x"2b9d0004", 10213 => x"2b8b0010", 10214 => x"2b8c000c",
    10215 => x"2b8d0008", 10216 => x"379c0010", 10217 => x"c3a00000",
    10218 => x"379cfffc", 10219 => x"5b9d0004", 10220 => x"78020001",
    10221 => x"3842785c", 10222 => x"28430000", 10223 => x"34042710",
    10224 => x"0865000a", 10225 => x"e0000004", 10226 => x"3442ffff",
    10227 => x"4840ffff", 10228 => x"3421d8f0", 10229 => x"50810003",
    10230 => x"b8a01000", 10231 => x"e3fffffc", 10232 => x"88230800",
    10233 => x"340203e8", 10234 => x"f80022d7", 10235 => x"e0000002",
    10236 => x"3421ffff", 10237 => x"4820ffff", 10238 => x"34010000",
    10239 => x"2b9d0004", 10240 => x"379c0004", 10241 => x"c3a00000",
    10242 => x"b8202800", 10243 => x"5c800002", 10244 => x"b8602000",
    10245 => x"b8803000", 10246 => x"50640002", 10247 => x"b8603000",
    10248 => x"b4260800", 10249 => x"e000000e", 10250 => x"2c460002",
    10251 => x"2847000c", 10252 => x"b4e63800", 10253 => x"40e60000",
    10254 => x"30a60000", 10255 => x"2c470002", 10256 => x"2c460006",
    10257 => x"34a50001", 10258 => x"34e70001", 10259 => x"20e7ffff",
    10260 => x"0c470002", 10261 => x"5cc70002", 10262 => x"0c400002",
    10263 => x"5ca1fff3", 10264 => x"5083000b", 10265 => x"2c410002",
    10266 => x"b4610800", 10267 => x"c8242000", 10268 => x"0c440002",
    10269 => x"2c410006", 10270 => x"e0000003", 10271 => x"c8812000",
    10272 => x"0c440002", 10273 => x"2c440002", 10274 => x"5481fffd",
    10275 => x"b8600800", 10276 => x"c3a00000", 10277 => x"b4432800",
    10278 => x"e000000d", 10279 => x"2c240000", 10280 => x"2826000c",
    10281 => x"40470000", 10282 => x"34420001", 10283 => x"b4c43000",
    10284 => x"30c70000", 10285 => x"34840001", 10286 => x"2c260006",
    10287 => x"2084ffff", 10288 => x"0c240000", 10289 => x"5cc40002",
    10290 => x"0c200000", 10291 => x"5c45fff4", 10292 => x"b8600800",
    10293 => x"c3a00000", 10294 => x"379cffc8", 10295 => x"5b8b001c",
    10296 => x"5b8c0018", 10297 => x"5b8d0014", 10298 => x"5b8e0010",
    10299 => x"5b8f000c", 10300 => x"5b900008", 10301 => x"5b9d0004",
    10302 => x"780b0001", 10303 => x"780c0001", 10304 => x"396b7a70",
    10305 => x"398c7890", 10306 => x"b9600800", 10307 => x"b9801000",
    10308 => x"340301e0", 10309 => x"37840020", 10310 => x"f8000d94",
    10311 => x"b8206800", 10312 => x"340f0000", 10313 => x"4c010061",
    10314 => x"2d62000c", 10315 => x"0f800038", 10316 => x"38018100",
    10317 => x"5c41000e", 10318 => x"b9801000", 10319 => x"34030002",
    10320 => x"37810038", 10321 => x"f80022e1", 10322 => x"78010001",
    10323 => x"78020001", 10324 => x"38217a7c", 10325 => x"38427892",
    10326 => x"34030002", 10327 => x"780c0001", 10328 => x"f80022da",
    10329 => x"35adfffc", 10330 => x"398c7894", 10331 => x"78010001",
    10332 => x"2f820038", 10333 => x"3821726c", 10334 => x"28210000",
    10335 => x"20420fff", 10336 => x"340f0000", 10337 => x"5c410049",
    10338 => x"41820000", 10339 => x"34010045", 10340 => x"34030000",
    10341 => x"5c410008", 10342 => x"41820009", 10343 => x"34010011",
    10344 => x"5c410005", 10345 => x"41830016", 10346 => x"41810017",
    10347 => x"3c630008", 10348 => x"b8611800", 10349 => x"78010001",
    10350 => x"78020001", 10351 => x"38217a70", 10352 => x"38427860",
    10353 => x"2c27000c", 10354 => x"34460030", 10355 => x"34040000",
    10356 => x"340b0000", 10357 => x"e000000c", 10358 => x"28410000",
    10359 => x"44200009", 10360 => x"2c25000c", 10361 => x"5ca70007",
    10362 => x"2c25000e", 10363 => x"5c600003", 10364 => x"44a30038",
    10365 => x"e0000003", 10366 => x"5ca30002", 10367 => x"b8202000",
    10368 => x"34420004", 10369 => x"5c46fff5", 10370 => x"44800002",
    10371 => x"b8805800", 10372 => x"340f0001", 10373 => x"45600025",
    10374 => x"2d700028", 10375 => x"35a10028", 10376 => x"48300022",
    10377 => x"356e0024", 10378 => x"3782003a", 10379 => x"34030002",
    10380 => x"b9c00800", 10381 => x"0f8d003a", 10382 => x"fbffff97",
    10383 => x"ca016800", 10384 => x"21adffff", 10385 => x"0d6d0028",
    10386 => x"37820020", 10387 => x"34030018", 10388 => x"b9c00800",
    10389 => x"fbffff90", 10390 => x"c9a16800", 10391 => x"21adffff",
    10392 => x"78020001", 10393 => x"0d6d0028", 10394 => x"38427a70",
    10395 => x"3403000e", 10396 => x"b9c00800", 10397 => x"fbffff88",
    10398 => x"c9a16800", 10399 => x"2f83003a", 10400 => x"21adffff",
    10401 => x"0d6d0028", 10402 => x"b9c00800", 10403 => x"b9801000",
    10404 => x"fbffff81", 10405 => x"c9a10800", 10406 => x"0d610028",
    10407 => x"2d61002c", 10408 => x"34210001", 10409 => x"0d61002c",
    10410 => x"b9e00800", 10411 => x"2b9d0004", 10412 => x"2b8b001c",
    10413 => x"2b8c0018", 10414 => x"2b8d0014", 10415 => x"2b8e0010",
    10416 => x"2b8f000c", 10417 => x"2b900008", 10418 => x"379c0038",
    10419 => x"c3a00000", 10420 => x"b8205800", 10421 => x"e3ffffcb",
    10422 => x"379cfffc", 10423 => x"5b9d0004", 10424 => x"b8400800",
    10425 => x"f80009ce", 10426 => x"34010000", 10427 => x"2b9d0004",
    10428 => x"379c0004", 10429 => x"c3a00000", 10430 => x"78020001",
    10431 => x"38427860", 10432 => x"34430030", 10433 => x"e0000004",
    10434 => x"28440000", 10435 => x"34420004", 10436 => x"5881001c",
    10437 => x"5c43fffd", 10438 => x"c3a00000", 10439 => x"379cff24",
    10440 => x"5b8b0014", 10441 => x"5b8c0010", 10442 => x"5b8d000c",
    10443 => x"5b8e0008", 10444 => x"5b9d0004", 10445 => x"78050001",
    10446 => x"b8205800", 10447 => x"b8406000", 10448 => x"b8607000",
    10449 => x"b8806800", 10450 => x"38a57860", 10451 => x"34010000",
    10452 => x"3402000c", 10453 => x"28a30000", 10454 => x"34a50004",
    10455 => x"5c600009", 10456 => x"3c220002", 10457 => x"78050001",
    10458 => x"38a57860", 10459 => x"b4a22800", 10460 => x"58ab0000",
    10461 => x"3402000c", 10462 => x"5c22000a", 10463 => x"e0000003",
    10464 => x"34210001", 10465 => x"5c22fff4", 10466 => x"78010001",
    10467 => x"78020001", 10468 => x"38425b10", 10469 => x"38215284",
    10470 => x"f8000899", 10471 => x"e0000020", 10472 => x"78020001",
    10473 => x"37810018", 10474 => x"384252a0", 10475 => x"fbfff77a",
    10476 => x"4801001b", 10477 => x"b9600800", 10478 => x"34020000",
    10479 => x"34030012", 10480 => x"f80022c0", 10481 => x"45800005",
    10482 => x"b9600800", 10483 => x"b9801000", 10484 => x"34030012",
    10485 => x"f800223d", 10486 => x"0d60000e", 10487 => x"5dc00004",
    10488 => x"34010800", 10489 => x"0d61000c", 10490 => x"0d6d000e",
    10491 => x"35610012", 10492 => x"f800098b", 10493 => x"2b8100d0",
    10494 => x"0d600026", 10495 => x"0d600024", 10496 => x"5961001c",
    10497 => x"2b8100b8", 10498 => x"0d60002c", 10499 => x"59610020",
    10500 => x"2d61002a", 10501 => x"0d610028", 10502 => x"e0000002",
    10503 => x"340b0000", 10504 => x"b9600800", 10505 => x"2b9d0004",
    10506 => x"2b8b0014", 10507 => x"2b8c0010", 10508 => x"2b8d000c",
    10509 => x"2b8e0008", 10510 => x"379c00dc", 10511 => x"c3a00000",
    10512 => x"78020001", 10513 => x"38427860", 10514 => x"34430030",
    10515 => x"e0000005", 10516 => x"28440000", 10517 => x"5c810002",
    10518 => x"58400000", 10519 => x"34420004", 10520 => x"5c43fffc",
    10521 => x"34010000", 10522 => x"c3a00000", 10523 => x"379cffe8",
    10524 => x"5b8b0018", 10525 => x"5b8c0014", 10526 => x"5b8d0010",
    10527 => x"5b8e000c", 10528 => x"5b8f0008", 10529 => x"5b9d0004",
    10530 => x"b8205800", 10531 => x"59620010", 10532 => x"b8407000",
    10533 => x"b8807800", 10534 => x"b8a06000", 10535 => x"282d0008",
    10536 => x"44600005", 10537 => x"b8a00800", 10538 => x"3402fc18",
    10539 => x"f8002159", 10540 => x"b42d6800", 10541 => x"c9cf2000",
    10542 => x"b8801800", 10543 => x"4c800002", 10544 => x"b48c1800",
    10545 => x"0181001f", 10546 => x"b42c0800", 10547 => x"14210001",
    10548 => x"b4242000", 10549 => x"4c800002", 10550 => x"b48c2000",
    10551 => x"49840002", 10552 => x"c88c2000", 10553 => x"09820003",
    10554 => x"1445001f", 10555 => x"00a5001e", 10556 => x"b4a21000",
    10557 => x"14420002", 10558 => x"48620006", 10559 => x"1582001f",
    10560 => x"0042001e", 10561 => x"b44c1000", 10562 => x"14420002",
    10563 => x"4c62000d", 10564 => x"b4812000", 10565 => x"596d0008",
    10566 => x"5964000c", 10567 => x"4984000a", 10568 => x"c88c2000",
    10569 => x"5964000c", 10570 => x"b9800800", 10571 => x"340203e8",
    10572 => x"f8002138", 10573 => x"b5a10800", 10574 => x"59610008",
    10575 => x"e0000002", 10576 => x"5963000c", 10577 => x"78030001",
    10578 => x"38635758", 10579 => x"29610008", 10580 => x"28620000",
    10581 => x"4c41000d", 10582 => x"78030001", 10583 => x"3863575c",
    10584 => x"28620000", 10585 => x"29630000", 10586 => x"b4220800",
    10587 => x"29620004", 10588 => x"59610008", 10589 => x"34410001",
    10590 => x"f4411000", 10591 => x"59610004", 10592 => x"b4431000",
    10593 => x"59620000", 10594 => x"2b9d0004", 10595 => x"2b8b0018",
    10596 => x"2b8c0014", 10597 => x"2b8d0010", 10598 => x"2b8e000c",
    10599 => x"2b8f0008", 10600 => x"379c0018", 10601 => x"c3a00000",
    10602 => x"379cffb4", 10603 => x"5b8b0024", 10604 => x"5b8c0020",
    10605 => x"5b8d001c", 10606 => x"5b8e0018", 10607 => x"5b8f0014",
    10608 => x"5b900010", 10609 => x"5b91000c", 10610 => x"5b920008",
    10611 => x"5b9d0004", 10612 => x"b8406800", 10613 => x"2c22002c",
    10614 => x"b8a05800", 10615 => x"b8206000", 10616 => x"b8609000",
    10617 => x"b8807800", 10618 => x"34050000", 10619 => x"44400055",
    10620 => x"342e0024", 10621 => x"2c310028", 10622 => x"3442ffff",
    10623 => x"0c22002c", 10624 => x"34030002", 10625 => x"b9c01000",
    10626 => x"34040000", 10627 => x"3781004e", 10628 => x"fbfffe7e",
    10629 => x"b6218800", 10630 => x"2231ffff", 10631 => x"0d910028",
    10632 => x"b9c01000", 10633 => x"34030018", 10634 => x"34040000",
    10635 => x"37810028", 10636 => x"fbfffe76", 10637 => x"b6218800",
    10638 => x"2231ffff", 10639 => x"37900040", 10640 => x"0d910028",
    10641 => x"b9c01000", 10642 => x"3403000e", 10643 => x"34040000",
    10644 => x"ba000800", 10645 => x"fbfffe6d", 10646 => x"b6218800",
    10647 => x"2f83004e", 10648 => x"2231ffff", 10649 => x"b9c01000",
    10650 => x"b9e02000", 10651 => x"0d910028", 10652 => x"ba400800",
    10653 => x"fbfffe65", 10654 => x"b6210800", 10655 => x"0d810028",
    10656 => x"2f81004c", 10657 => x"78030001", 10658 => x"3863726c",
    10659 => x"0da1000c", 10660 => x"28610000", 10661 => x"37820046",
    10662 => x"34030006", 10663 => x"0da10010", 10664 => x"b9a00800",
    10665 => x"f8002189", 10666 => x"35a10006", 10667 => x"ba001000",
    10668 => x"34030006", 10669 => x"f8002185", 10670 => x"4560001e",
    10671 => x"2b810038", 10672 => x"59610014", 10673 => x"2b81002c",
    10674 => x"59610018", 10675 => x"34010000", 10676 => x"f8001e66",
    10677 => x"b8206800", 10678 => x"35620010", 10679 => x"34030000",
    10680 => x"34010000", 10681 => x"f8001e0c", 10682 => x"2b810030",
    10683 => x"43820028", 10684 => x"2b83002c", 10685 => x"59610000",
    10686 => x"2b810034", 10687 => x"2984001c", 10688 => x"5960000c",
    10689 => x"59610004", 10690 => x"2b810038", 10691 => x"34051f40",
    10692 => x"59610008", 10693 => x"21a100ff", 10694 => x"64210000",
    10695 => x"a0220800", 10696 => x"29620010", 10697 => x"5961001c",
    10698 => x"b9600800", 10699 => x"fbffff50", 10700 => x"2f81004e",
    10701 => x"b9e02800", 10702 => x"502f0002", 10703 => x"b8202800",
    10704 => x"b8a00800", 10705 => x"2b9d0004", 10706 => x"2b8b0024",
    10707 => x"2b8c0020", 10708 => x"2b8d001c", 10709 => x"2b8e0018",
    10710 => x"2b8f0014", 10711 => x"2b900010", 10712 => x"2b91000c",
    10713 => x"2b920008", 10714 => x"379c004c", 10715 => x"c3a00000",
    10716 => x"379cffc0", 10717 => x"5b8b0014", 10718 => x"5b8c0010",
    10719 => x"5b8d000c", 10720 => x"5b8e0008", 10721 => x"5b9d0004",
    10722 => x"b8206000", 10723 => x"b8607000", 10724 => x"37810030",
    10725 => x"34030006", 10726 => x"b8a05800", 10727 => x"b8806800",
    10728 => x"f800214a", 10729 => x"37810036", 10730 => x"35820012",
    10731 => x"34030006", 10732 => x"f8002146", 10733 => x"78010001",
    10734 => x"3821726c", 10735 => x"28250000", 10736 => x"2d81000c",
    10737 => x"44a00009", 10738 => x"34028100", 10739 => x"0f82003c",
    10740 => x"2d820018", 10741 => x"0f810040", 10742 => x"3c42000d",
    10743 => x"b8452800", 10744 => x"0f85003e", 10745 => x"e0000002",
    10746 => x"0f81003c", 10747 => x"37810030", 10748 => x"b9c01000",
    10749 => x"b9a01800", 10750 => x"37840018", 10751 => x"f8000c86",
    10752 => x"4560000a", 10753 => x"2b820020", 10754 => x"5960000c",
    10755 => x"59620000", 10756 => x"2b820024", 10757 => x"59620004",
    10758 => x"2b820028", 10759 => x"59620008", 10760 => x"43820018",
    10761 => x"5962001c", 10762 => x"2b9d0004", 10763 => x"2b8b0014",
    10764 => x"2b8c0010", 10765 => x"2b8d000c", 10766 => x"2b8e0008",
    10767 => x"379c0040", 10768 => x"c3a00000", 10769 => x"c3a00000",
    10770 => x"379cffe4", 10771 => x"5b8b0008", 10772 => x"5b9d0004",
    10773 => x"78010001", 10774 => x"34020000", 10775 => x"34030000",
    10776 => x"34040044", 10777 => x"38216594", 10778 => x"fbfffead",
    10779 => x"78020001", 10780 => x"38427a84", 10781 => x"58410000",
    10782 => x"78010001", 10783 => x"34040025", 10784 => x"34020000",
    10785 => x"34030000", 10786 => x"382165c8", 10787 => x"fbfffea4",
    10788 => x"78020001", 10789 => x"378b000c", 10790 => x"38427a94",
    10791 => x"58410000", 10792 => x"34030012", 10793 => x"b9600800",
    10794 => x"34020000", 10795 => x"f8002185", 10796 => x"34010800",
    10797 => x"0f810018", 10798 => x"78010001", 10799 => x"b9601000",
    10800 => x"34030001", 10801 => x"34040000", 10802 => x"382165fc",
    10803 => x"fbfffe94", 10804 => x"78020001", 10805 => x"38427a90",
    10806 => x"58410000", 10807 => x"fbffffda", 10808 => x"2b9d0004",
    10809 => x"2b8b0008", 10810 => x"379c001c", 10811 => x"c3a00000",
    10812 => x"34010000", 10813 => x"c3a00000", 10814 => x"379cfe34",
    10815 => x"5b8b001c", 10816 => x"5b8c0018", 10817 => x"5b8d0014",
    10818 => x"5b8e0010", 10819 => x"5b8f000c", 10820 => x"5b900008",
    10821 => x"5b9d0004", 10822 => x"78010001", 10823 => x"38218f88",
    10824 => x"28220000", 10825 => x"34010001", 10826 => x"5c410006",
    10827 => x"78010001", 10828 => x"38217a80", 10829 => x"28230000",
    10830 => x"5c620002", 10831 => x"58200000", 10832 => x"78020001",
    10833 => x"38427a84", 10834 => x"28410000", 10835 => x"378b0020",
    10836 => x"378201b0", 10837 => x"34040190", 10838 => x"b9601800",
    10839 => x"34050000", 10840 => x"fbffff12", 10841 => x"78040001",
    10842 => x"38847a80", 10843 => x"b8201000", 10844 => x"28810000",
    10845 => x"340c0000", 10846 => x"5c200023", 10847 => x"4c220003",
    10848 => x"b9600800", 10849 => x"f800027a", 10850 => x"f8000cdd",
    10851 => x"78020001", 10852 => x"38427a88", 10853 => x"28430000",
    10854 => x"5c600003", 10855 => x"58410000", 10856 => x"e0000006",
    10857 => x"346303e8", 10858 => x"c8230800", 10859 => x"340c0000",
    10860 => x"48010015", 10861 => x"58430000", 10862 => x"78010001",
    10863 => x"38217a8c", 10864 => x"28230000", 10865 => x"378c01b0",
    10866 => x"378b0020", 10867 => x"34630001", 10868 => x"58230000",
    10869 => x"b9601000", 10870 => x"b9800800", 10871 => x"f8000200",
    10872 => x"78050001", 10873 => x"38a57a84", 10874 => x"b8202000",
    10875 => x"28a10000", 10876 => x"b9801000", 10877 => x"b9601800",
    10878 => x"34050000", 10879 => x"fbffff5d", 10880 => x"340c0001",
    10881 => x"780b0001", 10882 => x"396b7a90", 10883 => x"29610000",
    10884 => x"378e01b0", 10885 => x"378d0020", 10886 => x"34040080",
    10887 => x"b9c01000", 10888 => x"b9a01800", 10889 => x"34050000",
    10890 => x"fbfffee0", 10891 => x"b8202000", 10892 => x"340f0000",
    10893 => x"4c010010", 10894 => x"78030001", 10895 => x"38637a80",
    10896 => x"28610000", 10897 => x"4420000c", 10898 => x"b8801000",
    10899 => x"b9a00800", 10900 => x"f8000108", 10901 => x"b8202000",
    10902 => x"340f0001", 10903 => x"4c010006", 10904 => x"29610000",
    10905 => x"b9c01000", 10906 => x"b9a01800", 10907 => x"34050000",
    10908 => x"fbffff40", 10909 => x"780b0001", 10910 => x"396b7a94",
    10911 => x"29610000", 10912 => x"379001b0", 10913 => x"378d0020",
    10914 => x"ba001000", 10915 => x"b9a01800", 10916 => x"34040020",
    10917 => x"34050000", 10918 => x"fbfffec4", 10919 => x"340e0000",
    10920 => x"4c010019", 10921 => x"378101c4", 10922 => x"34020000",
    10923 => x"f800100f", 10924 => x"78020001", 10925 => x"38425780",
    10926 => x"28410000", 10927 => x"2b8201c8", 10928 => x"34030004",
    10929 => x"340e0001", 10930 => x"b4410800", 10931 => x"5b8101cc",
    10932 => x"378201cc", 10933 => x"3781003c", 10934 => x"f800207c",
    10935 => x"b9a00800", 10936 => x"34020020", 10937 => x"34030000",
    10938 => x"f8000143", 10939 => x"29610000", 10940 => x"ba001000",
    10941 => x"b9a01800", 10942 => x"34040020", 10943 => x"34050000",
    10944 => x"fbffff1c", 10945 => x"fbffff7b", 10946 => x"b5ec6000",
    10947 => x"b5810800", 10948 => x"b42e7000", 10949 => x"7dc10000",
    10950 => x"2b9d0004", 10951 => x"2b8b001c", 10952 => x"2b8c0018",
    10953 => x"2b8d0014", 10954 => x"2b8e0010", 10955 => x"2b8f000c",
    10956 => x"2b900008", 10957 => x"379c01cc", 10958 => x"c3a00000",
    10959 => x"34030000", 10960 => x"34040000", 10961 => x"e0000005",
    10962 => x"2c250000", 10963 => x"34840001", 10964 => x"34210002",
    10965 => x"b4651800", 10966 => x"4844fffc", 10967 => x"00610010",
    10968 => x"2063ffff", 10969 => x"b4611800", 10970 => x"00610010",
    10971 => x"b4231800", 10972 => x"a4600800", 10973 => x"2021ffff",
    10974 => x"c3a00000", 10975 => x"379cfffc", 10976 => x"5b9d0004",
    10977 => x"78020001", 10978 => x"38427a98", 10979 => x"34030004",
    10980 => x"f800204e", 10981 => x"2b9d0004", 10982 => x"379c0004",
    10983 => x"c3a00000", 10984 => x"379cfff0", 10985 => x"5b8b0010",
    10986 => x"5b8c000c", 10987 => x"5b8d0008", 10988 => x"5b9d0004",
    10989 => x"78030001", 10990 => x"780b0001", 10991 => x"396b7a98",
    10992 => x"b8206000", 10993 => x"38638fa0", 10994 => x"286d0000",
    10995 => x"b9600800", 10996 => x"b9801000", 10997 => x"34030004",
    10998 => x"f800203c", 10999 => x"41620000", 11000 => x"41610001",
    11001 => x"3c420018", 11002 => x"3c210010", 11003 => x"b8411000",
    11004 => x"41610003", 11005 => x"b8411000", 11006 => x"41610002",
    11007 => x"3c210008", 11008 => x"b8415800", 11009 => x"29a10018",
    11010 => x"b9800800", 11011 => x"f8000e61", 11012 => x"5d600004",
    11013 => x"78010001", 11014 => x"38217a80", 11015 => x"58200000",
    11016 => x"78010001", 11017 => x"38217a8c", 11018 => x"58200000",
    11019 => x"2b9d0004", 11020 => x"2b8b0010", 11021 => x"2b8c000c",
    11022 => x"2b8d0008", 11023 => x"379c0010", 11024 => x"c3a00000",
    11025 => x"379cfffc", 11026 => x"5b9d0004", 11027 => x"b8201000",
    11028 => x"3401ffff", 11029 => x"44400006", 11030 => x"34410010",
    11031 => x"78020001", 11032 => x"38427a98", 11033 => x"34030004",
    11034 => x"f8001ff7", 11035 => x"2b9d0004", 11036 => x"379c0004",
    11037 => x"c3a00000", 11038 => x"379cff34", 11039 => x"5b8b0028",
    11040 => x"5b8c0024", 11041 => x"5b8d0020", 11042 => x"5b8e001c",
    11043 => x"5b8f0018", 11044 => x"5b900014", 11045 => x"5b910010",
    11046 => x"5b92000c", 11047 => x"5b930008", 11048 => x"5b9d0004",
    11049 => x"78010001", 11050 => x"38217a80", 11051 => x"28210000",
    11052 => x"340b0000", 11053 => x"44200047", 11054 => x"780c0001",
    11055 => x"398c7d7c", 11056 => x"29810000", 11057 => x"378f00ac",
    11058 => x"378e002c", 11059 => x"b9e01000", 11060 => x"b9c01800",
    11061 => x"34040080", 11062 => x"34050000", 11063 => x"fbfffe33",
    11064 => x"4c01003c", 11065 => x"3402001b", 11066 => x"340b0001",
    11067 => x"4c410039", 11068 => x"378d00c8", 11069 => x"b9a00800",
    11070 => x"fbffffa1", 11071 => x"43810032", 11072 => x"5c200034",
    11073 => x"43810033", 11074 => x"5c2b0032", 11075 => x"37900044",
    11076 => x"ba000800", 11077 => x"b9a01000", 11078 => x"34030004",
    11079 => x"f8001fca", 11080 => x"5c20002c", 11081 => x"379100c0",
    11082 => x"37930034", 11083 => x"ba601000", 11084 => x"34030006",
    11085 => x"ba200800", 11086 => x"f8001fe4", 11087 => x"3792003a",
    11088 => x"ba401000", 11089 => x"34030004", 11090 => x"378100cc",
    11091 => x"f8001fdf", 11092 => x"34010008", 11093 => x"3381002e",
    11094 => x"34010006", 11095 => x"33810030", 11096 => x"34010004",
    11097 => x"33810031", 11098 => x"34010002", 11099 => x"33810033",
    11100 => x"ba600800", 11101 => x"3380002c", 11102 => x"338b002d",
    11103 => x"3380002f", 11104 => x"33800032", 11105 => x"f8000726",
    11106 => x"b9a01000", 11107 => x"34030004", 11108 => x"ba400800",
    11109 => x"f8001fcd", 11110 => x"ba201000", 11111 => x"34030006",
    11112 => x"3781003e", 11113 => x"f8001fc9", 11114 => x"378200cc",
    11115 => x"34030004", 11116 => x"ba000800", 11117 => x"f8001fc5",
    11118 => x"29810000", 11119 => x"b9e01000", 11120 => x"b9c01800",
    11121 => x"3404001c", 11122 => x"34050000", 11123 => x"fbfffe69",
    11124 => x"b9600800", 11125 => x"2b9d0004", 11126 => x"2b8b0028",
    11127 => x"2b8c0024", 11128 => x"2b8d0020", 11129 => x"2b8e001c",
    11130 => x"2b8f0018", 11131 => x"2b900014", 11132 => x"2b910010",
    11133 => x"2b92000c", 11134 => x"2b930008", 11135 => x"379c00cc",
    11136 => x"c3a00000", 11137 => x"379cffe4", 11138 => x"5b8b0008",
    11139 => x"5b9d0004", 11140 => x"378b000c", 11141 => x"b9600800",
    11142 => x"34020000", 11143 => x"34030012", 11144 => x"f8002028",
    11145 => x"b9600800", 11146 => x"340200ff", 11147 => x"34030006",
    11148 => x"f8002024", 11149 => x"34010806", 11150 => x"0f810018",
    11151 => x"78010001", 11152 => x"b9601000", 11153 => x"34030001",
    11154 => x"34040000", 11155 => x"38216630", 11156 => x"fbfffd33",
    11157 => x"78020001", 11158 => x"38427d7c", 11159 => x"58410000",
    11160 => x"2b9d0004", 11161 => x"2b8b0008", 11162 => x"379c001c",
    11163 => x"c3a00000", 11164 => x"379cffe0", 11165 => x"5b8b0018",
    11166 => x"5b8c0014", 11167 => x"5b8d0010", 11168 => x"5b8e000c",
    11169 => x"5b8f0008", 11170 => x"5b9d0004", 11171 => x"378d001c",
    11172 => x"b8205800", 11173 => x"b9a00800", 11174 => x"fbffff39",
    11175 => x"41620000", 11176 => x"34010045", 11177 => x"340c0000",
    11178 => x"5c41004a", 11179 => x"356e0010", 11180 => x"b9a01000",
    11181 => x"b9c00800", 11182 => x"34030004", 11183 => x"f8001f62",
    11184 => x"b8201000", 11185 => x"5c200043", 11186 => x"41640009",
    11187 => x"34030001", 11188 => x"416d0002", 11189 => x"41610003",
    11190 => x"b8406000", 11191 => x"5c83003d", 11192 => x"41630014",
    11193 => x"34020008", 11194 => x"5c62003a", 11195 => x"3dad0008",
    11196 => x"b9a16800", 11197 => x"35adffe8", 11198 => x"34010040",
    11199 => x"4c2d0002", 11200 => x"340d0040", 11201 => x"356f000c",
    11202 => x"b9e01000", 11203 => x"34030004", 11204 => x"37810020",
    11205 => x"f8001f6d", 11206 => x"35ac0018", 11207 => x"34010045",
    11208 => x"31610000", 11209 => x"15810008", 11210 => x"3782001c",
    11211 => x"31610002", 11212 => x"3401003f", 11213 => x"31610008",
    11214 => x"34010001", 11215 => x"31610009", 11216 => x"34030004",
    11217 => x"31600001", 11218 => x"316c0003", 11219 => x"31600004",
    11220 => x"31600005", 11221 => x"31600006", 11222 => x"31600007",
    11223 => x"3160000a", 11224 => x"3160000b", 11225 => x"b9e00800",
    11226 => x"f8001f58", 11227 => x"34030004", 11228 => x"37820020",
    11229 => x"b9c00800", 11230 => x"f8001f54", 11231 => x"35ad0005",
    11232 => x"01a1001f", 11233 => x"31600014", 11234 => x"b42d6800",
    11235 => x"15a20001", 11236 => x"31600015", 11237 => x"31600016",
    11238 => x"31600017", 11239 => x"35610014", 11240 => x"fbfffee7",
    11241 => x"2021ffff", 11242 => x"00220008", 11243 => x"31610017",
    11244 => x"31620016", 11245 => x"b9600800", 11246 => x"3402000a",
    11247 => x"fbfffee0", 11248 => x"2021ffff", 11249 => x"00220008",
    11250 => x"3161000b", 11251 => x"3162000a", 11252 => x"b9800800",
    11253 => x"2b9d0004", 11254 => x"2b8b0018", 11255 => x"2b8c0014",
    11256 => x"2b8d0010", 11257 => x"2b8e000c", 11258 => x"2b8f0008",
    11259 => x"379c0020", 11260 => x"c3a00000", 11261 => x"379cffcc",
    11262 => x"5b8b0028", 11263 => x"5b8c0024", 11264 => x"5b8d0020",
    11265 => x"5b8e001c", 11266 => x"5b8f0018", 11267 => x"5b900014",
    11268 => x"5b910010", 11269 => x"5b92000c", 11270 => x"5b930008",
    11271 => x"5b9d0004", 11272 => x"b8205800", 11273 => x"b8406800",
    11274 => x"b8606000", 11275 => x"5c600012", 11276 => x"3562000c",
    11277 => x"34030004", 11278 => x"37810030", 11279 => x"f8001f23",
    11280 => x"378c002c", 11281 => x"35620010", 11282 => x"34030004",
    11283 => x"b9800800", 11284 => x"f8001f1e", 11285 => x"35620014",
    11286 => x"34030002", 11287 => x"37810036", 11288 => x"f8001f1a",
    11289 => x"37810034", 11290 => x"35620016", 11291 => x"34030002",
    11292 => x"f8001f16", 11293 => x"35700008", 11294 => x"b9801000",
    11295 => x"34030004", 11296 => x"ba000800", 11297 => x"f8001f11",
    11298 => x"35b1ffec", 11299 => x"356f000c", 11300 => x"358e0004",
    11301 => x"b9c01000", 11302 => x"34030004", 11303 => x"16320008",
    11304 => x"b9e00800", 11305 => x"f8001f09", 11306 => x"34010011",
    11307 => x"225200ff", 11308 => x"223100ff", 11309 => x"31610011",
    11310 => x"35820008", 11311 => x"34030002", 11312 => x"31600010",
    11313 => x"31720012", 11314 => x"31710013", 11315 => x"35610014",
    11316 => x"f8001efe", 11317 => x"34030002", 11318 => x"3582000a",
    11319 => x"35610016", 11320 => x"f8001efa", 11321 => x"b56d0800",
    11322 => x"31720018", 11323 => x"31710019", 11324 => x"3160001a",
    11325 => x"3160001b", 11326 => x"35a2fff9", 11327 => x"30200000",
    11328 => x"0041001f", 11329 => x"35730010", 11330 => x"b4221000",
    11331 => x"14420001", 11332 => x"ba000800", 11333 => x"fbfffe8a",
    11334 => x"2023ffff", 11335 => x"5c600002", 11336 => x"3803ffff",
    11337 => x"00610008", 11338 => x"3163001b", 11339 => x"3161001a",
    11340 => x"34010045", 11341 => x"31610000", 11342 => x"15a10008",
    11343 => x"b9801000", 11344 => x"31610002", 11345 => x"3401003f",
    11346 => x"31610008", 11347 => x"34010011", 11348 => x"31610009",
    11349 => x"31600001", 11350 => x"316d0003", 11351 => x"31600004",
    11352 => x"31600005", 11353 => x"31600006", 11354 => x"31600007",
    11355 => x"3160000a", 11356 => x"3160000b", 11357 => x"b9e00800",
    11358 => x"34030004", 11359 => x"f8001ed3", 11360 => x"b9c01000",
    11361 => x"34030004", 11362 => x"ba600800", 11363 => x"f8001ecf",
    11364 => x"b9600800", 11365 => x"3402000a", 11366 => x"fbfffe69",
    11367 => x"2021ffff", 11368 => x"00220008", 11369 => x"3161000b",
    11370 => x"3162000a", 11371 => x"2b9d0004", 11372 => x"2b8b0028",
    11373 => x"2b8c0024", 11374 => x"2b8d0020", 11375 => x"2b8e001c",
    11376 => x"2b8f0018", 11377 => x"2b900014", 11378 => x"2b910010",
    11379 => x"2b92000c", 11380 => x"2b930008", 11381 => x"379c0034",
    11382 => x"c3a00000", 11383 => x"379cffe4", 11384 => x"5b8b0010",
    11385 => x"5b8c000c", 11386 => x"5b8d0008", 11387 => x"5b9d0004",
    11388 => x"b8405800", 11389 => x"b8206800", 11390 => x"34020001",
    11391 => x"34010006", 11392 => x"3162001c", 11393 => x"3162001d",
    11394 => x"3161001e", 11395 => x"3160001f", 11396 => x"35610020",
    11397 => x"b8606000", 11398 => x"f8000601", 11399 => x"41620024",
    11400 => x"41610020", 11401 => x"34030002", 11402 => x"98410800",
    11403 => x"31610020", 11404 => x"41620025", 11405 => x"41610021",
    11406 => x"316c0025", 11407 => x"98410800", 11408 => x"31610021",
    11409 => x"41610022", 11410 => x"15820008", 11411 => x"98410800",
    11412 => x"31610022", 11413 => x"41610023", 11414 => x"31620024",
    11415 => x"34020000", 11416 => x"982c0800", 11417 => x"31610023",
    11418 => x"35610026", 11419 => x"f8001f15", 11420 => x"35610028",
    11421 => x"34020000", 11422 => x"34030004", 11423 => x"f8001f11",
    11424 => x"3561002c", 11425 => x"34020000", 11426 => x"34030004",
    11427 => x"f8001f0d", 11428 => x"35610030", 11429 => x"34020000",
    11430 => x"34030004", 11431 => x"f8001f09", 11432 => x"35610034",
    11433 => x"34020000", 11434 => x"34030004", 11435 => x"f8001f05",
    11436 => x"356c0038", 11437 => x"34020000", 11438 => x"34030010",
    11439 => x"b9800800", 11440 => x"f8001f00", 11441 => x"b9800800",
    11442 => x"f80005d5", 11443 => x"35610048", 11444 => x"34020000",
    11445 => x"34030040", 11446 => x"f8001efa", 11447 => x"35610088",
    11448 => x"34020000", 11449 => x"34030080", 11450 => x"f8001ef6",
    11451 => x"35610108", 11452 => x"34020000", 11453 => x"34030040",
    11454 => x"f8001ef2", 11455 => x"378c0014", 11456 => x"b9800800",
    11457 => x"34020000", 11458 => x"34030004", 11459 => x"f8001eed",
    11460 => x"37810018", 11461 => x"340200ff", 11462 => x"34030004",
    11463 => x"f8001ee9", 11464 => x"34010044", 11465 => x"0f81001c",
    11466 => x"34010043", 11467 => x"0f81001e", 11468 => x"b9801800",
    11469 => x"b9600800", 11470 => x"34020148", 11471 => x"fbffff2e",
    11472 => x"b9a00800", 11473 => x"340200ff", 11474 => x"34030006",
    11475 => x"f8001edd", 11476 => x"34010148", 11477 => x"2b9d0004",
    11478 => x"2b8b0010", 11479 => x"2b8c000c", 11480 => x"2b8d0008",
    11481 => x"379c001c", 11482 => x"c3a00000", 11483 => x"379cffe0",
    11484 => x"5b8b0014", 11485 => x"5b8c0010", 11486 => x"5b8d000c",
    11487 => x"5b8e0008", 11488 => x"5b9d0004", 11489 => x"378d0018",
    11490 => x"b8205800", 11491 => x"b9a00800", 11492 => x"b8407000",
    11493 => x"f80005a2", 11494 => x"34010148", 11495 => x"340c0000",
    11496 => x"5dc1001b", 11497 => x"41610014", 11498 => x"5c200019",
    11499 => x"41620015", 11500 => x"34010043", 11501 => x"5c410016",
    11502 => x"35610038", 11503 => x"b9a01000", 11504 => x"34030006",
    11505 => x"f8001e20", 11506 => x"5c200011", 11507 => x"78010001",
    11508 => x"34020001", 11509 => x"38217a80", 11510 => x"58220000",
    11511 => x"3561002c", 11512 => x"fbfffdf0", 11513 => x"37810020",
    11514 => x"fbfffde5", 11515 => x"43820020", 11516 => x"43830021",
    11517 => x"43840022", 11518 => x"43850023", 11519 => x"78010001",
    11520 => x"382152b8", 11521 => x"f800047e", 11522 => x"340c0001",
    11523 => x"b9800800", 11524 => x"2b9d0004", 11525 => x"2b8b0014",
    11526 => x"2b8c0010", 11527 => x"2b8d000c", 11528 => x"2b8e0008",
    11529 => x"379c0020", 11530 => x"c3a00000", 11531 => x"379cfffc",
    11532 => x"5b8b0004", 11533 => x"78040001", 11534 => x"38845b48",
    11535 => x"3442ffff", 11536 => x"348a001c", 11537 => x"34030000",
    11538 => x"340900fd", 11539 => x"340800f9", 11540 => x"340700ff",
    11541 => x"3406ffa2", 11542 => x"e0000011", 11543 => x"40850000",
    11544 => x"5ca90004", 11545 => x"b4232800", 11546 => x"30a60000",
    11547 => x"e000000a", 11548 => x"5ca80005", 11549 => x"b4232800",
    11550 => x"40a50000", 11551 => x"b4651800", 11552 => x"e0000005",
    11553 => x"5ca70004", 11554 => x"b4232800", 11555 => x"c8435800",
    11556 => x"30ab0000", 11557 => x"34630001", 11558 => x"34840001",
    11559 => x"5c8afff0", 11560 => x"2b8b0004", 11561 => x"379c0004",
    11562 => x"c3a00000", 11563 => x"379cfff8", 11564 => x"5b8b0008",
    11565 => x"5b9d0004", 11566 => x"40230006", 11567 => x"34040020",
    11568 => x"4c830002", 11569 => x"34030020", 11570 => x"206b00ff",
    11571 => x"b42b1800", 11572 => x"3404ffa2", 11573 => x"30640007",
    11574 => x"4063000a", 11575 => x"34040004", 11576 => x"4c830002",
    11577 => x"34030004", 11578 => x"b5635800", 11579 => x"216b00ff",
    11580 => x"b42b1800", 11581 => x"3062000d", 11582 => x"34020001",
    11583 => x"30620010", 11584 => x"40620016", 11585 => x"34030028",
    11586 => x"4c620002", 11587 => x"34020028", 11588 => x"b5621000",
    11589 => x"204200ff", 11590 => x"b4221800", 11591 => x"34420019",
    11592 => x"34040005", 11593 => x"204b00ff", 11594 => x"30640017",
    11595 => x"30600018", 11596 => x"b9601000", 11597 => x"fbffffbe",
    11598 => x"b9600800", 11599 => x"2b9d0004", 11600 => x"2b8b0008",
    11601 => x"379c0008", 11602 => x"c3a00000", 11603 => x"379cfefc",
    11604 => x"5b8b0028", 11605 => x"5b8c0024", 11606 => x"5b8d0020",
    11607 => x"5b8e001c", 11608 => x"5b8f0018", 11609 => x"5b900014",
    11610 => x"5b910010", 11611 => x"5b92000c", 11612 => x"5b930008",
    11613 => x"5b9d0004", 11614 => x"78010001", 11615 => x"38217e00",
    11616 => x"28210000", 11617 => x"378b002c", 11618 => x"378200f4",
    11619 => x"b9601800", 11620 => x"340400c8", 11621 => x"34050000",
    11622 => x"fbfffc04", 11623 => x"34020038", 11624 => x"340c0000",
    11625 => x"504100a6", 11626 => x"b9600800", 11627 => x"fbfffda6",
    11628 => x"5c2000a3", 11629 => x"78010001", 11630 => x"78020001",
    11631 => x"38218f84", 11632 => x"38425b48", 11633 => x"78030001",
    11634 => x"40250000", 11635 => x"344e001c", 11636 => x"b9600800",
    11637 => x"34040000", 11638 => x"340d0006", 11639 => x"38635b2c",
    11640 => x"340b00a0", 11641 => x"340a00a1", 11642 => x"340900a3",
    11643 => x"34080001", 11644 => x"e0000028", 11645 => x"40460000",
    11646 => x"34c70007", 11647 => x"20e700ff", 11648 => x"54ed0014",
    11649 => x"3ce70002", 11650 => x"b4673800", 11651 => x"28e60000",
    11652 => x"c0c00000", 11653 => x"b4813000", 11654 => x"40c6001c",
    11655 => x"b4862000", 11656 => x"e000001a", 11657 => x"b4812800",
    11658 => x"40a5001c", 11659 => x"51050017", 11660 => x"e000000b",
    11661 => x"b4813000", 11662 => x"40c6001c", 11663 => x"44cb000e",
    11664 => x"44ca000f", 11665 => x"44c90010", 11666 => x"5d800010",
    11667 => x"e0000004", 11668 => x"b4813800", 11669 => x"40e7001c",
    11670 => x"44e6000c", 11671 => x"78010001", 11672 => x"38218f84",
    11673 => x"30250000", 11674 => x"34020005", 11675 => x"37810048",
    11676 => x"e000005b", 11677 => x"340c0002", 11678 => x"e0000004",
    11679 => x"340c0004", 11680 => x"e0000002", 11681 => x"340c0001",
    11682 => x"34840001", 11683 => x"34420001", 11684 => x"5c4effd9",
    11685 => x"78010001", 11686 => x"38218f84", 11687 => x"30250000",
    11688 => x"37810048", 11689 => x"b4246800", 11690 => x"780b0001",
    11691 => x"34840001", 11692 => x"b4247800", 11693 => x"396b6684",
    11694 => x"21930003", 11695 => x"21900004", 11696 => x"39920008",
    11697 => x"e000003f", 11698 => x"41b10000", 11699 => x"46600002",
    11700 => x"5431003b", 11701 => x"222200ff", 11702 => x"50220002",
    11703 => x"b8208800", 11704 => x"29610000", 11705 => x"223100ff",
    11706 => x"b9e01000", 11707 => x"ba201800", 11708 => x"f8001d55",
    11709 => x"3c250018", 11710 => x"b9807000", 11711 => x"14a50018",
    11712 => x"4600000a", 11713 => x"48a00007", 11714 => x"4163000c",
    11715 => x"41a10000", 11716 => x"64a20000", 11717 => x"f0610800",
    11718 => x"a0410800", 11719 => x"44200003", 11720 => x"4171000c",
    11721 => x"ba407000", 11722 => x"4163000c", 11723 => x"64a10000",
    11724 => x"e4711000", 11725 => x"a0411000", 11726 => x"5c400003",
    11727 => x"21c10008", 11728 => x"4422001e", 11729 => x"5e000003",
    11730 => x"21c10008", 11731 => x"44300004", 11732 => x"29620000",
    11733 => x"b9e00800", 11734 => x"f8001d5c", 11735 => x"29650004",
    11736 => x"29630008", 11737 => x"b9a00800", 11738 => x"ba201000",
    11739 => x"b9c02000", 11740 => x"d8a00000", 11741 => x"4c01000c",
    11742 => x"5e000003", 11743 => x"21ce0008", 11744 => x"45d00005",
    11745 => x"41a30000", 11746 => x"4162000c", 11747 => x"b4621000",
    11748 => x"31a20000", 11749 => x"4164000c", 11750 => x"b5e47800",
    11751 => x"b5e17800", 11752 => x"e000000a", 11753 => x"44200006",
    11754 => x"c8011000", 11755 => x"204200ff", 11756 => x"37810048",
    11757 => x"e000000a", 11758 => x"48a10007", 11759 => x"356b0010",
    11760 => x"4161000c", 11761 => x"5c20ffc1", 11762 => x"45600003",
    11763 => x"4161000c", 11764 => x"5c200006", 11765 => x"37810048",
    11766 => x"34020002", 11767 => x"fbffff34", 11768 => x"b8205800",
    11769 => x"e0000007", 11770 => x"37810048", 11771 => x"c9e15800",
    11772 => x"b9601000", 11773 => x"fbffff0e", 11774 => x"340c0000",
    11775 => x"480b0010", 11776 => x"378c002c", 11777 => x"356b001c",
    11778 => x"b9800800", 11779 => x"b9601000", 11780 => x"34030000",
    11781 => x"fbfffdf8", 11782 => x"78050001", 11783 => x"38a57e00",
    11784 => x"28a10000", 11785 => x"b9801800", 11786 => x"378200f4",
    11787 => x"b9602000", 11788 => x"34050000", 11789 => x"fbfffbcf",
    11790 => x"340c0001", 11791 => x"b9800800", 11792 => x"2b9d0004",
    11793 => x"2b8b0028", 11794 => x"2b8c0024", 11795 => x"2b8d0020",
    11796 => x"2b8e001c", 11797 => x"2b8f0018", 11798 => x"2b900014",
    11799 => x"2b910010", 11800 => x"2b92000c", 11801 => x"2b930008",
    11802 => x"379c0104", 11803 => x"c3a00000", 11804 => x"379cffec",
    11805 => x"5b8b0010", 11806 => x"5b8c000c", 11807 => x"5b8d0008",
    11808 => x"5b9d0004", 11809 => x"b8403000", 11810 => x"40c50011",
    11811 => x"40220000", 11812 => x"b8606000", 11813 => x"402b0001",
    11814 => x"3404fffd", 11815 => x"5ca2001e", 11816 => x"34220002",
    11817 => x"34010004", 11818 => x"44a10013", 11819 => x"34010042",
    11820 => x"44a10004", 11821 => x"34010002", 11822 => x"34040000",
    11823 => x"5ca10016", 11824 => x"340d0004", 11825 => x"3404fffd",
    11826 => x"556d0013", 11827 => x"37810014", 11828 => x"b9601800",
    11829 => x"5b800014", 11830 => x"f8001cfc", 11831 => x"2b810014",
    11832 => x"c9ab6800", 11833 => x"3dad0003", 11834 => x"802d6800",
    11835 => x"598d0000", 11836 => x"e0000008", 11837 => x"40c10013",
    11838 => x"55610007", 11839 => x"b8600800", 11840 => x"b58b6000",
    11841 => x"b9601800", 11842 => x"f8001cf0", 11843 => x"31800000",
    11844 => x"35640002", 11845 => x"b8800800", 11846 => x"2b9d0004",
    11847 => x"2b8b0010", 11848 => x"2b8c000c", 11849 => x"2b8d0008",
    11850 => x"379c0014", 11851 => x"c3a00000", 11852 => x"379cfffc",
    11853 => x"5b9d0004", 11854 => x"40430012", 11855 => x"2844000c",
    11856 => x"b4831800", 11857 => x"fbffffcb", 11858 => x"2b9d0004",
    11859 => x"379c0004", 11860 => x"c3a00000", 11861 => x"379cffcc",
    11862 => x"5b8b0020", 11863 => x"5b8c001c", 11864 => x"5b8d0018",
    11865 => x"5b8e0014", 11866 => x"5b8f0010", 11867 => x"5b90000c",
    11868 => x"5b910008", 11869 => x"5b9d0004", 11870 => x"402e0000",
    11871 => x"204200ff", 11872 => x"208400ff", 11873 => x"344c0001",
    11874 => x"c9c27000", 11875 => x"20820001", 11876 => x"b8207800",
    11877 => x"b42c6000", 11878 => x"3401fffc", 11879 => x"5c400068",
    11880 => x"208d0004", 11881 => x"7dad0000", 11882 => x"20900008",
    11883 => x"7e100000", 11884 => x"b8605800", 11885 => x"21b100ff",
    11886 => x"e0000023", 11887 => x"b9c01800", 11888 => x"4c2e0002",
    11889 => x"b8201800", 11890 => x"29610000", 11891 => x"b9801000",
    11892 => x"206300ff", 11893 => x"f8001c9c", 11894 => x"5e00000a",
    11895 => x"b0200800", 11896 => x"64220000", 11897 => x"a0511800",
    11898 => x"44700003", 11899 => x"41630010", 11900 => x"4c6e0004",
    11901 => x"68210000", 11902 => x"a2210800", 11903 => x"4420000b",
    11904 => x"29620000", 11905 => x"41630010", 11906 => x"b9800800",
    11907 => x"340e0000", 11908 => x"f8001cae", 11909 => x"41610010",
    11910 => x"34020001", 11911 => x"b5810800", 11912 => x"30220000",
    11913 => x"e000000d", 11914 => x"44410006", 11915 => x"41610010",
    11916 => x"34210001", 11917 => x"45c10006", 11918 => x"45a00002",
    11919 => x"49c10006", 11920 => x"356b0014", 11921 => x"41610010",
    11922 => x"5c20ffdd", 11923 => x"b9a07000", 11924 => x"e0000002",
    11925 => x"340e0001", 11926 => x"41620010", 11927 => x"34010000",
    11928 => x"44400037", 11929 => x"41610011", 11930 => x"33820034",
    11931 => x"5b8c0024", 11932 => x"33810035", 11933 => x"2961000c",
    11934 => x"5b810030", 11935 => x"45c00004", 11936 => x"41810001",
    11937 => x"34210001", 11938 => x"31810001", 11939 => x"41610010",
    11940 => x"29630004", 11941 => x"37910024", 11942 => x"34210001",
    11943 => x"b5810800", 11944 => x"ba201000", 11945 => x"d8600000",
    11946 => x"64230000", 11947 => x"a06e7000", 11948 => x"45c00019",
    11949 => x"356b0014", 11950 => x"41630010", 11951 => x"34010000",
    11952 => x"4460001f", 11953 => x"29620000", 11954 => x"b9800800",
    11955 => x"f8001c7f", 11956 => x"41610010", 11957 => x"34020001",
    11958 => x"b5810800", 11959 => x"30220000", 11960 => x"41620011",
    11961 => x"41610010", 11962 => x"29630004", 11963 => x"33820035",
    11964 => x"2962000c", 11965 => x"33810034", 11966 => x"34210001",
    11967 => x"5b820030", 11968 => x"b5810800", 11969 => x"ba201000",
    11970 => x"d8600000", 11971 => x"5c200003", 11972 => x"e000000b",
    11973 => x"5c6e0009", 11974 => x"48010009", 11975 => x"41620010",
    11976 => x"ba0d6800", 11977 => x"34420001", 11978 => x"b4220800",
    11979 => x"45a00004", 11980 => x"31e20000", 11981 => x"e0000002",
    11982 => x"34010000", 11983 => x"2b9d0004", 11984 => x"2b8b0020",
    11985 => x"2b8c001c", 11986 => x"2b8d0018", 11987 => x"2b8e0014",
    11988 => x"2b8f0010", 11989 => x"2b90000c", 11990 => x"2b910008",
    11991 => x"379c0034", 11992 => x"c3a00000", 11993 => x"379cffd0",
    11994 => x"5b8b0030", 11995 => x"5b8c002c", 11996 => x"5b8d0028",
    11997 => x"5b8e0024", 11998 => x"5b8f0020", 11999 => x"5b90001c",
    12000 => x"5b910018", 12001 => x"5b920014", 12002 => x"5b930010",
    12003 => x"5b94000c", 12004 => x"5b950008", 12005 => x"5b9d0004",
    12006 => x"208400ff", 12007 => x"40310000", 12008 => x"204200ff",
    12009 => x"008d0003", 12010 => x"344e0001", 12011 => x"208f0004",
    12012 => x"b8208000", 12013 => x"ca228800", 12014 => x"b42e7000",
    12015 => x"21ad0001", 12016 => x"b8605800", 12017 => x"340c0000",
    12018 => x"20950003", 12019 => x"20940001", 12020 => x"7df30000",
    12021 => x"e0000034", 12022 => x"b8a09000", 12023 => x"5da00005",
    12024 => x"ba209000", 12025 => x"4cb10002", 12026 => x"b8a09000",
    12027 => x"225200ff", 12028 => x"46a00002", 12029 => x"5e25002b",
    12030 => x"5da0000c", 12031 => x"29610000", 12032 => x"b9c01000",
    12033 => x"ba401800", 12034 => x"f8001c0f", 12035 => x"3c2c0018",
    12036 => x"158c0018", 12037 => x"5d8d0006", 12038 => x"45ec0009",
    12039 => x"41610010", 12040 => x"5c320007", 12041 => x"e000001f",
    12042 => x"45800005", 12043 => x"69810000", 12044 => x"a0331000",
    12045 => x"5c400002", 12046 => x"45a20019", 12047 => x"45e00007",
    12048 => x"29620000", 12049 => x"41630010", 12050 => x"b9c00800",
    12051 => x"f8001c1f", 12052 => x"41610010", 12053 => x"32010000",
    12054 => x"46800008", 12055 => x"29630008", 12056 => x"44600014",
    12057 => x"41610010", 12058 => x"b9601000", 12059 => x"b5c10800",
    12060 => x"d8600000", 12061 => x"48010012", 12062 => x"41610010",
    12063 => x"29630004", 12064 => x"b9601000", 12065 => x"b5c10800",
    12066 => x"d8600000", 12067 => x"44200005", 12068 => x"41620010",
    12069 => x"b4220800", 12070 => x"e0000009", 12071 => x"5c2d0007",
    12072 => x"356b0014", 12073 => x"41650010", 12074 => x"5ca0ffcc",
    12075 => x"e0000003", 12076 => x"3401fffc", 12077 => x"e0000002",
    12078 => x"34010000", 12079 => x"2b9d0004", 12080 => x"2b8b0030",
    12081 => x"2b8c002c", 12082 => x"2b8d0028", 12083 => x"2b8e0024",
    12084 => x"2b8f0020", 12085 => x"2b90001c", 12086 => x"2b910018",
    12087 => x"2b920014", 12088 => x"2b930010", 12089 => x"2b94000c",
    12090 => x"2b950008", 12091 => x"379c0030", 12092 => x"c3a00000",
    12093 => x"379cffe4", 12094 => x"5b8b0010", 12095 => x"5b8c000c",
    12096 => x"5b8d0008", 12097 => x"5b9d0004", 12098 => x"b8206000",
    12099 => x"342d0002", 12100 => x"30220000", 12101 => x"34010043",
    12102 => x"b8605800", 12103 => x"54410008", 12104 => x"34010041",
    12105 => x"50410009", 12106 => x"34010002", 12107 => x"44410007",
    12108 => x"34010004", 12109 => x"5c410029", 12110 => x"e000001c",
    12111 => x"34010046", 12112 => x"5c410026", 12113 => x"e0000009",
    12114 => x"29610000", 12115 => x"3782001c", 12116 => x"34030004",
    12117 => x"5b81001c", 12118 => x"b9a00800", 12119 => x"f8001bdb",
    12120 => x"34010004", 12121 => x"e000000f", 12122 => x"78010001",
    12123 => x"38218f84", 12124 => x"40210000", 12125 => x"34020000",
    12126 => x"44200019", 12127 => x"28610000", 12128 => x"37820014",
    12129 => x"5b810014", 12130 => x"28610004", 12131 => x"34030008",
    12132 => x"5b810018", 12133 => x"b9a00800", 12134 => x"f8001bcc",
    12135 => x"34010008", 12136 => x"31810001", 12137 => x"e000000a",
    12138 => x"b8600800", 12139 => x"3402001f", 12140 => x"f8001da9",
    12141 => x"202300ff", 12142 => x"31830001", 12143 => x"b9a00800",
    12144 => x"b9601000", 12145 => x"34630001", 12146 => x"f8001bc0",
    12147 => x"41820001", 12148 => x"34420002", 12149 => x"e0000002",
    12150 => x"34020000", 12151 => x"b8400800", 12152 => x"2b9d0004",
    12153 => x"2b8b0010", 12154 => x"2b8c000c", 12155 => x"2b8d0008",
    12156 => x"379c001c", 12157 => x"c3a00000", 12158 => x"379cff98",
    12159 => x"5b8b0034", 12160 => x"5b8c0030", 12161 => x"5b8d002c",
    12162 => x"5b8e0028", 12163 => x"5b8f0024", 12164 => x"5b900020",
    12165 => x"5b91001c", 12166 => x"5b920018", 12167 => x"5b930014",
    12168 => x"5b940010", 12169 => x"5b95000c", 12170 => x"5b960008",
    12171 => x"5b9d0004", 12172 => x"b8208000", 12173 => x"28410000",
    12174 => x"b8407000", 12175 => x"340d0000", 12176 => x"40360001",
    12177 => x"402c0000", 12178 => x"340b0001", 12179 => x"378f0038",
    12180 => x"3415ffff", 12181 => x"34140002", 12182 => x"34130003",
    12183 => x"34120004", 12184 => x"34110005", 12185 => x"21a300ff",
    12186 => x"b9e00800", 12187 => x"34020000", 12188 => x"f8000c18",
    12189 => x"b8201800", 12190 => x"4420001c", 12191 => x"4435001b",
    12192 => x"5ecb000d", 12193 => x"5d940009", 12194 => x"378b0058",
    12195 => x"34030010", 12196 => x"b9600800", 12197 => x"b9e01000",
    12198 => x"f8001b8c", 12199 => x"b9601800", 12200 => x"33800068",
    12201 => x"e000000d", 12202 => x"45930007", 12203 => x"45920008",
    12204 => x"45910009", 12205 => x"356b0001", 12206 => x"35ad0001",
    12207 => x"4c6bffea", 12208 => x"e000000a", 12209 => x"3783004c",
    12210 => x"e0000004", 12211 => x"37830050", 12212 => x"e0000002",
    12213 => x"37830048", 12214 => x"41c20011", 12215 => x"ba000800",
    12216 => x"fbffff85", 12217 => x"e0000002", 12218 => x"34010000",
    12219 => x"2b9d0004", 12220 => x"2b8b0034", 12221 => x"2b8c0030",
    12222 => x"2b8d002c", 12223 => x"2b8e0028", 12224 => x"2b8f0024",
    12225 => x"2b900020", 12226 => x"2b91001c", 12227 => x"2b920018",
    12228 => x"2b930014", 12229 => x"2b940010", 12230 => x"2b95000c",
    12231 => x"2b960008", 12232 => x"379c0068", 12233 => x"c3a00000",
    12234 => x"379cffe8", 12235 => x"5b8b0010", 12236 => x"5b8c000c",
    12237 => x"5b8d0008", 12238 => x"5b9d0004", 12239 => x"b8405800",
    12240 => x"2842000c", 12241 => x"34030001", 12242 => x"b8206800",
    12243 => x"44430019", 12244 => x"34030002", 12245 => x"5c43002e",
    12246 => x"78020001", 12247 => x"38427e04", 12248 => x"28430000",
    12249 => x"286400b4", 12250 => x"286500b0", 12251 => x"c8042000",
    12252 => x"7c820000", 12253 => x"c8052800", 12254 => x"c8a22800",
    12255 => x"3c820001", 12256 => x"3ca50001", 12257 => x"f4822000",
    12258 => x"b4852000", 12259 => x"286500a0", 12260 => x"286300a4",
    12261 => x"b4852000", 12262 => x"b4431800", 12263 => x"f4431000",
    12264 => x"5b830018", 12265 => x"b4441000", 12266 => x"5b820014",
    12267 => x"e0000014", 12268 => x"78020001", 12269 => x"38427e04",
    12270 => x"284c0000", 12271 => x"78050001", 12272 => x"38a55748",
    12273 => x"298200fc", 12274 => x"28a40000", 12275 => x"34030000",
    12276 => x"1441001f", 12277 => x"f8001a68", 12278 => x"29830100",
    12279 => x"1464001f", 12280 => x"b4431800", 12281 => x"f4431000",
    12282 => x"b4242000", 12283 => x"b4442000", 12284 => x"5b840014",
    12285 => x"5b830018", 12286 => x"b9a00800", 12287 => x"41620011",
    12288 => x"37830014", 12289 => x"fbffff3c", 12290 => x"e0000002",
    12291 => x"3401ffff", 12292 => x"2b9d0004", 12293 => x"2b8b0010",
    12294 => x"2b8c000c", 12295 => x"2b8d0008", 12296 => x"379c0018",
    12297 => x"c3a00000", 12298 => x"379cfff8", 12299 => x"5b9d0004",
    12300 => x"2843000c", 12301 => x"40450011", 12302 => x"40420012",
    12303 => x"28630000", 12304 => x"b4621000", 12305 => x"28440000",
    12306 => x"28430004", 12307 => x"4880000e", 12308 => x"5c800005",
    12309 => x"78060001", 12310 => x"38c65760", 12311 => x"28c20000",
    12312 => x"54620009", 12313 => x"3402ffff", 12314 => x"4844000b",
    12315 => x"5c82000b", 12316 => x"78040001", 12317 => x"38845764",
    12318 => x"28820000", 12319 => x"54430006", 12320 => x"e0000006",
    12321 => x"78060001", 12322 => x"38c65784", 12323 => x"28c30000",
    12324 => x"e0000002", 12325 => x"78038000", 12326 => x"5b830008",
    12327 => x"b8a01000", 12328 => x"37830008", 12329 => x"fbffff14",
    12330 => x"2b9d0004", 12331 => x"379c0008", 12332 => x"c3a00000",
    12333 => x"379cfffc", 12334 => x"5b9d0004", 12335 => x"2844000c",
    12336 => x"40430012", 12337 => x"40420011", 12338 => x"28840000",
    12339 => x"b4831800", 12340 => x"fbffff09", 12341 => x"2b9d0004",
    12342 => x"379c0004", 12343 => x"c3a00000", 12344 => x"379cfffc",
    12345 => x"5b9d0004", 12346 => x"2844000c", 12347 => x"40430012",
    12348 => x"40420011", 12349 => x"b4831800", 12350 => x"fbfffeff",
    12351 => x"2b9d0004", 12352 => x"379c0004", 12353 => x"c3a00000",
    12354 => x"379cfff0", 12355 => x"5b8b000c", 12356 => x"5b8c0008",
    12357 => x"5b9d0004", 12358 => x"b8405800", 12359 => x"2842000c",
    12360 => x"b8206000", 12361 => x"34010001", 12362 => x"5c41000a",
    12363 => x"34010000", 12364 => x"f8000286", 12365 => x"34220001",
    12366 => x"5b820010", 12367 => x"41620011", 12368 => x"b9800800",
    12369 => x"37830010", 12370 => x"fbfffeeb", 12371 => x"e0000002",
    12372 => x"3401ffff", 12373 => x"2b9d0004", 12374 => x"2b8b000c",
    12375 => x"2b8c0008", 12376 => x"379c0010", 12377 => x"c3a00000",
    12378 => x"379cfff4", 12379 => x"5b8b000c", 12380 => x"5b8c0008",
    12381 => x"5b9d0004", 12382 => x"284b000c", 12383 => x"b9601800",
    12384 => x"fbfffdbc", 12385 => x"b8206000", 12386 => x"4c01000a",
    12387 => x"29620000", 12388 => x"34010001", 12389 => x"5c410005",
    12390 => x"fbffd333", 12391 => x"fbffd30c", 12392 => x"34010064",
    12393 => x"e0000002", 12394 => x"340100c8", 12395 => x"59610000",
    12396 => x"b9800800", 12397 => x"2b9d0004", 12398 => x"2b8b000c",
    12399 => x"2b8c0008", 12400 => x"379c000c", 12401 => x"c3a00000",
    12402 => x"379cfff0", 12403 => x"5b8b0010", 12404 => x"5b8c000c",
    12405 => x"5b8d0008", 12406 => x"5b9d0004", 12407 => x"284b000c",
    12408 => x"b9601800", 12409 => x"fbfffda3", 12410 => x"b8206800",
    12411 => x"4c010050", 12412 => x"29620000", 12413 => x"34010002",
    12414 => x"4441001e", 12415 => x"48410004", 12416 => x"34010001",
    12417 => x"5c410048", 12418 => x"e0000020", 12419 => x"34010003",
    12420 => x"44410004", 12421 => x"34010032", 12422 => x"5c410043",
    12423 => x"e000003d", 12424 => x"78020001", 12425 => x"38427e08",
    12426 => x"28410014", 12427 => x"78030001", 12428 => x"38638bb8",
    12429 => x"58610000", 12430 => x"28410018", 12431 => x"78030001",
    12432 => x"38638bbc", 12433 => x"58610000", 12434 => x"28410010",
    12435 => x"78030001", 12436 => x"38636d1c", 12437 => x"58610000",
    12438 => x"78010001", 12439 => x"382152e0", 12440 => x"f80000e7",
    12441 => x"fbffd300", 12442 => x"fbffd2d9", 12443 => x"e000002c",
    12444 => x"78010001", 12445 => x"78020001", 12446 => x"38217e08",
    12447 => x"38428c24", 12448 => x"34030010", 12449 => x"f8001a91",
    12450 => x"780c0001", 12451 => x"398c7e08", 12452 => x"41810000",
    12453 => x"5c200003", 12454 => x"340100cb", 12455 => x"e0000023",
    12456 => x"34020010", 12457 => x"b9800800", 12458 => x"f8001c6b",
    12459 => x"b8201000", 12460 => x"3403000f", 12461 => x"34010020",
    12462 => x"e0000004", 12463 => x"b44c2000", 12464 => x"30810000",
    12465 => x"34420001", 12466 => x"4c62fffd", 12467 => x"34020001",
    12468 => x"b9800800", 12469 => x"34030000", 12470 => x"f8000afe",
    12471 => x"b8201000", 12472 => x"3401fffe", 12473 => x"5c410003",
    12474 => x"340100ca", 12475 => x"e000000f", 12476 => x"3401ffff",
    12477 => x"5c410003", 12478 => x"340100c9", 12479 => x"e000000b",
    12480 => x"f80006da", 12481 => x"44200006", 12482 => x"34010065",
    12483 => x"e0000007", 12484 => x"f8000ad7", 12485 => x"3402ffff",
    12486 => x"44220003", 12487 => x"34010064", 12488 => x"e0000002",
    12489 => x"340100c8", 12490 => x"59610000", 12491 => x"b9a00800",
    12492 => x"2b9d0004", 12493 => x"2b8b0010", 12494 => x"2b8c000c",
    12495 => x"2b8d0008", 12496 => x"379c0010", 12497 => x"c3a00000",
    12498 => x"379cffc8", 12499 => x"5b8b0024", 12500 => x"5b8c0020",
    12501 => x"5b8d001c", 12502 => x"5b8e0018", 12503 => x"5b8f0014",
    12504 => x"5b900010", 12505 => x"5b91000c", 12506 => x"5b920008",
    12507 => x"5b9d0004", 12508 => x"b8207800", 12509 => x"28410000",
    12510 => x"b8406800", 12511 => x"340c0001", 12512 => x"40320001",
    12513 => x"402e0000", 12514 => x"34010000", 12515 => x"f80008f2",
    12516 => x"b8202000", 12517 => x"34110002", 12518 => x"34100003",
    12519 => x"e0000025", 12520 => x"5e4c0020", 12521 => x"288b0004",
    12522 => x"5dd10007", 12523 => x"28830000", 12524 => x"78020001",
    12525 => x"37810028", 12526 => x"38424860", 12527 => x"f8000082",
    12528 => x"e000001f", 12529 => x"5dd00017", 12530 => x"78018000",
    12531 => x"5d610006", 12532 => x"78020001", 12533 => x"37810028",
    12534 => x"3842530c", 12535 => x"f800007a", 12536 => x"e0000017",
    12537 => x"4d600006", 12538 => x"78020001", 12539 => x"37810028",
    12540 => x"38424458", 12541 => x"c80b5800", 12542 => x"f8000073",
    12543 => x"2164ffff", 12544 => x"08842710", 12545 => x"78020001",
    12546 => x"15630010", 12547 => x"00840010", 12548 => x"37810028",
    12549 => x"38425314", 12550 => x"f800006b", 12551 => x"e0000008",
    12552 => x"b8800800", 12553 => x"f80008cc", 12554 => x"b8202000",
    12555 => x"358c0001", 12556 => x"5c80ffdc", 12557 => x"34010000",
    12558 => x"e0000005", 12559 => x"41a20011", 12560 => x"b9e00800",
    12561 => x"37830028", 12562 => x"fbfffe2b", 12563 => x"2b9d0004",
    12564 => x"2b8b0024", 12565 => x"2b8c0020", 12566 => x"2b8d001c",
    12567 => x"2b8e0018", 12568 => x"2b8f0014", 12569 => x"2b900010",
    12570 => x"2b91000c", 12571 => x"2b920008", 12572 => x"379c0038",
    12573 => x"c3a00000", 12574 => x"379cffe4", 12575 => x"5b8b0010",
    12576 => x"5b8c000c", 12577 => x"5b8d0008", 12578 => x"5b9d0004",
    12579 => x"284d000c", 12580 => x"b8206000", 12581 => x"b8405800",
    12582 => x"21a10002", 12583 => x"44200009", 12584 => x"f8000617",
    12585 => x"3402000a", 12586 => x"f80019a7", 12587 => x"5b81001c",
    12588 => x"41620011", 12589 => x"b9800800", 12590 => x"3783001c",
    12591 => x"e0000013", 12592 => x"21a20004", 12593 => x"44410004",
    12594 => x"37810014", 12595 => x"34020000", 12596 => x"f8000986",
    12597 => x"21ad0001", 12598 => x"45a00009", 12599 => x"2b820018",
    12600 => x"2b810014", 12601 => x"34030002", 12602 => x"fbfff565",
    12603 => x"b8201800", 12604 => x"41620011", 12605 => x"b9800800",
    12606 => x"e0000004", 12607 => x"41620011", 12608 => x"b9800800",
    12609 => x"37830014", 12610 => x"fbfffdfb", 12611 => x"2b9d0004",
    12612 => x"2b8b0010", 12613 => x"2b8c000c", 12614 => x"2b8d0008",
    12615 => x"379c001c", 12616 => x"c3a00000", 12617 => x"379cfffc",
    12618 => x"5b9d0004", 12619 => x"78010001", 12620 => x"34020000",
    12621 => x"34030000", 12622 => x"340400a1", 12623 => x"38216714",
    12624 => x"fbfff777", 12625 => x"78020001", 12626 => x"38427e00",
    12627 => x"58410000", 12628 => x"78010001", 12629 => x"38215e98",
    12630 => x"28210014", 12631 => x"78020001", 12632 => x"38427e04",
    12633 => x"58410000", 12634 => x"2b9d0004", 12635 => x"379c0004",
    12636 => x"c3a00000", 12637 => x"379cfff4", 12638 => x"5b8b000c",
    12639 => x"5b8c0008", 12640 => x"5b9d0004", 12641 => x"780b0001",
    12642 => x"b8202000", 12643 => x"396b7f30", 12644 => x"b8401800",
    12645 => x"b9600800", 12646 => x"b8801000", 12647 => x"f8000027",
    12648 => x"b8206000", 12649 => x"b9600800", 12650 => x"f8001025",
    12651 => x"b9800800", 12652 => x"2b9d0004", 12653 => x"2b8b000c",
    12654 => x"2b8c0008", 12655 => x"379c000c", 12656 => x"c3a00000",
    12657 => x"379cffe0", 12658 => x"5b9d0004", 12659 => x"5b83000c",
    12660 => x"3783000c", 12661 => x"5b820008", 12662 => x"5b840010",
    12663 => x"5b850014", 12664 => x"5b860018", 12665 => x"5b87001c",
    12666 => x"5b880020", 12667 => x"f8000013", 12668 => x"2b9d0004",
    12669 => x"379c0020", 12670 => x"c3a00000", 12671 => x"379cffdc",
    12672 => x"5b9d0004", 12673 => x"5b82000c", 12674 => x"3782000c",
    12675 => x"5b810008", 12676 => x"5b830010", 12677 => x"5b840014",
    12678 => x"5b850018", 12679 => x"5b86001c", 12680 => x"5b870020",
    12681 => x"5b880024", 12682 => x"fbffffd3", 12683 => x"2b9d0004",
    12684 => x"379c0024", 12685 => x"c3a00000", 12686 => x"379cff94",
    12687 => x"5b8b0044", 12688 => x"5b8c0040", 12689 => x"5b8d003c",
    12690 => x"5b8e0038", 12691 => x"5b8f0034", 12692 => x"5b900030",
    12693 => x"5b91002c", 12694 => x"5b920028", 12695 => x"5b930024",
    12696 => x"5b940020", 12697 => x"5b95001c", 12698 => x"5b960018",
    12699 => x"5b970014", 12700 => x"5b980010", 12701 => x"5b99000c",
    12702 => x"5b9b0008", 12703 => x"5b9d0004", 12704 => x"78160001",
    12705 => x"b820c800", 12706 => x"b840a000", 12707 => x"b8209800",
    12708 => x"34180025", 12709 => x"34090069", 12710 => x"34080070",
    12711 => x"34070058", 12712 => x"34060063", 12713 => x"34050064",
    12714 => x"341b002a", 12715 => x"340a0030", 12716 => x"34170010",
    12717 => x"37950060", 12718 => x"3ad6533c", 12719 => x"e0000093",
    12720 => x"34110001", 12721 => x"34100020", 12722 => x"340e000a",
    12723 => x"44380004", 12724 => x"32610000", 12725 => x"e0000038",
    12726 => x"34100030", 12727 => x"36940001", 12728 => x"42810000",
    12729 => x"4429003c", 12730 => x"5429000d", 12731 => x"44270037",
    12732 => x"54270008", 12733 => x"443b0018", 12734 => x"543b0004",
    12735 => x"44200085", 12736 => x"5c380017", 12737 => x"e000002b",
    12738 => x"5c2a0015", 12739 => x"e3fffff3", 12740 => x"44260019",
    12741 => x"5c250012", 12742 => x"e000002f", 12743 => x"4428002b",
    12744 => x"54280006", 12745 => x"3402006e", 12746 => x"44220077",
    12747 => x"3404006f", 12748 => x"5c24000b", 12749 => x"e0000022",
    12750 => x"34020075", 12751 => x"44220026", 12752 => x"34040078",
    12753 => x"44240021", 12754 => x"34020073", 12755 => x"5c220004",
    12756 => x"e000000e", 12757 => x"286e0000", 12758 => x"34630004",
    12759 => x"3422ffcf", 12760 => x"204200ff", 12761 => x"34040008",
    12762 => x"5444ffdd", 12763 => x"3431ffd0", 12764 => x"e3ffffdb",
    12765 => x"28610000", 12766 => x"34630004", 12767 => x"32610000",
    12768 => x"36730001", 12769 => x"e0000060", 12770 => x"b8600800",
    12771 => x"28210000", 12772 => x"34630004", 12773 => x"e0000004",
    12774 => x"32620000", 12775 => x"34210001", 12776 => x"36730001",
    12777 => x"40220000", 12778 => x"5c40fffc", 12779 => x"e0000056",
    12780 => x"32780000", 12781 => x"36730001", 12782 => x"e0000053",
    12783 => x"3401000a", 12784 => x"45c10004", 12785 => x"e0000004",
    12786 => x"340e0010", 12787 => x"e0000002", 12788 => x"340e0008",
    12789 => x"286d0000", 12790 => x"34720004", 12791 => x"65c3000a",
    12792 => x"01a4001f", 12793 => x"340f0000", 12794 => x"a0831800",
    12795 => x"44600003", 12796 => x"c80d6800", 12797 => x"340f0001",
    12798 => x"340c0010", 12799 => x"e0000019", 12800 => x"b9a00800",
    12801 => x"b9c01000", 12802 => x"5b85004c", 12803 => x"5b860050",
    12804 => x"5b870054", 12805 => x"5b880058", 12806 => x"5b89005c",
    12807 => x"5b8a0048", 12808 => x"f80018d9", 12809 => x"b6c11800",
    12810 => x"40630000", 12811 => x"358cffff", 12812 => x"b6ac5800",
    12813 => x"b9a00800", 12814 => x"31630000", 12815 => x"b9c01000",
    12816 => x"f80018c1", 12817 => x"2b8a0048", 12818 => x"2b89005c",
    12819 => x"2b880058", 12820 => x"2b870054", 12821 => x"2b860050",
    12822 => x"2b85004c", 12823 => x"b8206800", 12824 => x"7d840000",
    12825 => x"7da30000", 12826 => x"a0831800", 12827 => x"5c60ffe5",
    12828 => x"5d970004", 12829 => x"34020030", 12830 => x"3382006f",
    12831 => x"340c000f", 12832 => x"66020020", 12833 => x"a1e21000",
    12834 => x"4440000b", 12835 => x"358cffff", 12836 => x"b6ac1000",
    12837 => x"3403002d", 12838 => x"30430000", 12839 => x"340f0000",
    12840 => x"e0000005", 12841 => x"358cffff", 12842 => x"b6ac1000",
    12843 => x"30500000", 12844 => x"e0000003", 12845 => x"caf10800",
    12846 => x"b42f0800", 12847 => x"4981fffa", 12848 => x"45e00005",
    12849 => x"358cffff", 12850 => x"b6ac0800", 12851 => x"3402002d",
    12852 => x"30220000", 12853 => x"caec1800", 12854 => x"ba600800",
    12855 => x"3404000f", 12856 => x"e0000006", 12857 => x"b6ac1000",
    12858 => x"40420000", 12859 => x"358c0001", 12860 => x"30220000",
    12861 => x"34210001", 12862 => x"4c8cfffb", 12863 => x"b6639800",
    12864 => x"ba401800", 12865 => x"36940001", 12866 => x"42810000",
    12867 => x"5c20ff6d", 12868 => x"ca790800", 12869 => x"32600000",
    12870 => x"2b9d0004", 12871 => x"2b8b0044", 12872 => x"2b8c0040",
    12873 => x"2b8d003c", 12874 => x"2b8e0038", 12875 => x"2b8f0034",
    12876 => x"2b900030", 12877 => x"2b91002c", 12878 => x"2b920028",
    12879 => x"2b930024", 12880 => x"2b940020", 12881 => x"2b95001c",
    12882 => x"2b960018", 12883 => x"2b970014", 12884 => x"2b980010",
    12885 => x"2b99000c", 12886 => x"2b9b0008", 12887 => x"379c006c",
    12888 => x"c3a00000", 12889 => x"78020001", 12890 => x"14210002",
    12891 => x"38428f94", 12892 => x"28420000", 12893 => x"202100ff",
    12894 => x"3c210010", 12895 => x"5841002c", 12896 => x"28410030",
    12897 => x"4c20ffff", 12898 => x"28410030", 12899 => x"2021ffff",
    12900 => x"c3a00000", 12901 => x"14210002", 12902 => x"78030001",
    12903 => x"38638f94", 12904 => x"202100ff", 12905 => x"28630000",
    12906 => x"2042ffff", 12907 => x"78048000", 12908 => x"3c210010",
    12909 => x"b8441000", 12910 => x"b8411000", 12911 => x"5862002c",
    12912 => x"28610030", 12913 => x"4c20ffff", 12914 => x"c3a00000",
    12915 => x"40240002", 12916 => x"40230003", 12917 => x"78020001",
    12918 => x"3c840018", 12919 => x"3c630010", 12920 => x"38428f94",
    12921 => x"b8831800", 12922 => x"40240005", 12923 => x"28420000",
    12924 => x"b8641800", 12925 => x"40240004", 12926 => x"3c840008",
    12927 => x"b8641800", 12928 => x"58430028", 12929 => x"40230001",
    12930 => x"40210000", 12931 => x"3c210008", 12932 => x"b8610800",
    12933 => x"58410024", 12934 => x"c3a00000", 12935 => x"78020001",
    12936 => x"38428f94", 12937 => x"28430000", 12938 => x"28630028",
    12939 => x"30230005", 12940 => x"28430000", 12941 => x"28630028",
    12942 => x"00630008", 12943 => x"30230004", 12944 => x"28430000",
    12945 => x"28630028", 12946 => x"00630010", 12947 => x"30230003",
    12948 => x"28430000", 12949 => x"28630028", 12950 => x"00630018",
    12951 => x"30230002", 12952 => x"28430000", 12953 => x"28630024",
    12954 => x"30230001", 12955 => x"28420000", 12956 => x"28420024",
    12957 => x"00420008", 12958 => x"30220000", 12959 => x"c3a00000",
    12960 => x"379cfff4", 12961 => x"5b8b000c", 12962 => x"5b8c0008",
    12963 => x"5b9d0004", 12964 => x"780b0001", 12965 => x"b8406000",
    12966 => x"396b8f94", 12967 => x"5c200004", 12968 => x"29610000",
    12969 => x"58200000", 12970 => x"e0000022", 12971 => x"29610000",
    12972 => x"58200000", 12973 => x"28220034", 12974 => x"78010001",
    12975 => x"38215350", 12976 => x"fbfffecf", 12977 => x"f80000be",
    12978 => x"29610000", 12979 => x"340200e0", 12980 => x"58220000",
    12981 => x"78010001", 12982 => x"38217fb0", 12983 => x"34020800",
    12984 => x"582c0000", 12985 => x"34010000", 12986 => x"fbffffab",
    12987 => x"340100c8", 12988 => x"f8000488", 12989 => x"34010000",
    12990 => x"38028000", 12991 => x"fbffffa6", 12992 => x"34010000",
    12993 => x"34020000", 12994 => x"fbffffa3", 12995 => x"34010010",
    12996 => x"34020000", 12997 => x"fbffffa0", 12998 => x"7d820000",
    12999 => x"34010000", 13000 => x"c8021000", 13001 => x"20421200",
    13002 => x"34420140", 13003 => x"fbffff9a", 13004 => x"34010000",
    13005 => x"2b9d0004", 13006 => x"2b8b000c", 13007 => x"2b8c0008",
    13008 => x"379c000c", 13009 => x"c3a00000", 13010 => x"379cfff0",
    13011 => x"5b8b000c", 13012 => x"5b8c0008", 13013 => x"5b9d0004",
    13014 => x"78020001", 13015 => x"38427fb0", 13016 => x"284b0000",
    13017 => x"b8206000", 13018 => x"34010004", 13019 => x"fbffff7e",
    13020 => x"7d6b0000", 13021 => x"0f810012", 13022 => x"34010004",
    13023 => x"c80b5800", 13024 => x"fbffff79", 13025 => x"216b0020",
    13026 => x"0f810012", 13027 => x"356b0004", 13028 => x"45800004",
    13029 => x"34010014", 13030 => x"fbffff73", 13031 => x"0d810000",
    13032 => x"2f810012", 13033 => x"a1610800", 13034 => x"e42b0800",
    13035 => x"2b9d0004", 13036 => x"2b8b000c", 13037 => x"2b8c0008",
    13038 => x"379c0010", 13039 => x"c3a00000", 13040 => x"379cfffc",
    13041 => x"5b9d0004", 13042 => x"34010040", 13043 => x"fbffff66",
    13044 => x"00210004", 13045 => x"2021001f", 13046 => x"08210320",
    13047 => x"2b9d0004", 13048 => x"379c0004", 13049 => x"c3a00000",
    13050 => x"379cfff4", 13051 => x"5b8b000c", 13052 => x"5b8c0008",
    13053 => x"5b9d0004", 13054 => x"78030001", 13055 => x"38638bb8",
    13056 => x"b8405800", 13057 => x"28620000", 13058 => x"58220000",
    13059 => x"78010001", 13060 => x"38218bbc", 13061 => x"282c0000",
    13062 => x"34010040", 13063 => x"fbffff52", 13064 => x"00210004",
    13065 => x"2021001f", 13066 => x"08210320", 13067 => x"b42c0800",
    13068 => x"59610000", 13069 => x"34010000", 13070 => x"2b9d0004",
    13071 => x"2b8b000c", 13072 => x"2b8c0008", 13073 => x"379c000c",
    13074 => x"c3a00000", 13075 => x"379cfffc", 13076 => x"5b9d0004",
    13077 => x"34010040", 13078 => x"fbffff43", 13079 => x"38220001",
    13080 => x"34010040", 13081 => x"fbffff4c", 13082 => x"34010000",
    13083 => x"2b9d0004", 13084 => x"379c0004", 13085 => x"c3a00000",
    13086 => x"379cfffc", 13087 => x"5b9d0004", 13088 => x"34010040",
    13089 => x"fbffff38", 13090 => x"3402fffe", 13091 => x"a0221000",
    13092 => x"34010040", 13093 => x"fbffff40", 13094 => x"34010000",
    13095 => x"2b9d0004", 13096 => x"379c0004", 13097 => x"c3a00000",
    13098 => x"379cfff8", 13099 => x"5b8b0008", 13100 => x"5b9d0004",
    13101 => x"780b0001", 13102 => x"396b8f94", 13103 => x"29610000",
    13104 => x"28220004", 13105 => x"38420010", 13106 => x"58220004",
    13107 => x"34010001", 13108 => x"f8000410", 13109 => x"29610000",
    13110 => x"28210004", 13111 => x"20210020", 13112 => x"7c210000",
    13113 => x"2b9d0004", 13114 => x"2b8b0008", 13115 => x"379c0008",
    13116 => x"c3a00000", 13117 => x"379cfff8", 13118 => x"5b8b0008",
    13119 => x"5b9d0004", 13120 => x"b8205800", 13121 => x"34010044",
    13122 => x"fbffff17", 13123 => x"38220020", 13124 => x"45600003",
    13125 => x"3402ffdf", 13126 => x"a0221000", 13127 => x"34010044",
    13128 => x"fbffff1d", 13129 => x"34010000", 13130 => x"2b9d0004",
    13131 => x"2b8b0008", 13132 => x"379c0008", 13133 => x"c3a00000",
    13134 => x"379cfff8", 13135 => x"5b8b0008", 13136 => x"5b9d0004",
    13137 => x"78020001", 13138 => x"38428c18", 13139 => x"28420000",
    13140 => x"780b0001", 13141 => x"396b8f94", 13142 => x"59620000",
    13143 => x"fbffff1c", 13144 => x"34010001", 13145 => x"fbffffe4",
    13146 => x"78020001", 13147 => x"38425788", 13148 => x"28410000",
    13149 => x"78040001", 13150 => x"3884578c", 13151 => x"58200000",
    13152 => x"29610000", 13153 => x"28830000", 13154 => x"34020003",
    13155 => x"58200000", 13156 => x"5822000c", 13157 => x"58230008",
    13158 => x"78030001", 13159 => x"38635790", 13160 => x"58220004",
    13161 => x"28620000", 13162 => x"5822003c", 13163 => x"2b9d0004",
    13164 => x"2b8b0008", 13165 => x"379c0008", 13166 => x"c3a00000",
    13167 => x"379cffec", 13168 => x"5b8b000c", 13169 => x"5b8c0008",
    13170 => x"5b9d0004", 13171 => x"78010001", 13172 => x"3821726c",
    13173 => x"28220000", 13174 => x"78010001", 13175 => x"38216cfc",
    13176 => x"44400003", 13177 => x"78010001", 13178 => x"38216d04",
    13179 => x"282b0000", 13180 => x"5d600004", 13181 => x"78010001",
    13182 => x"38215358", 13183 => x"e0000036", 13184 => x"78030001",
    13185 => x"38635794", 13186 => x"282c0004", 13187 => x"29620000",
    13188 => x"28610000", 13189 => x"44410011", 13190 => x"b9600800",
    13191 => x"780400ff", 13192 => x"e000000d", 13193 => x"28230000",
    13194 => x"3c660018", 13195 => x"00650018", 13196 => x"b8c52800",
    13197 => x"a0643000", 13198 => x"00c60008", 13199 => x"2063ff00",
    13200 => x"3c630008", 13201 => x"b8a62800", 13202 => x"b8a31800",
    13203 => x"58230000", 13204 => x"34210004", 13205 => x"5581fff4",
    13206 => x"78040001", 13207 => x"38845794", 13208 => x"29630000",
    13209 => x"28810000", 13210 => x"44610005", 13211 => x"78010001",
    13212 => x"38215370", 13213 => x"fbfffde2", 13214 => x"e000008c",
    13215 => x"78010001", 13216 => x"38217fb4", 13217 => x"28220000",
    13218 => x"356b0004", 13219 => x"5c400016", 13220 => x"29630008",
    13221 => x"34021234", 13222 => x"0063000d", 13223 => x"2063ffff",
    13224 => x"5c62000b", 13225 => x"29630010", 13226 => x"34025678",
    13227 => x"0063000d", 13228 => x"2063ffff", 13229 => x"5c620006",
    13230 => x"29630018", 13231 => x"34424444", 13232 => x"0063000d",
    13233 => x"2063ffff", 13234 => x"44620005", 13235 => x"78010001",
    13236 => x"38215398", 13237 => x"fbfffdca", 13238 => x"e0000074",
    13239 => x"34020001", 13240 => x"58220000", 13241 => x"37810010",
    13242 => x"fbfffecd", 13243 => x"78050001", 13244 => x"38a55798",
    13245 => x"28a20000", 13246 => x"29640008", 13247 => x"29630010",
    13248 => x"29610018", 13249 => x"a0822000", 13250 => x"a0621800",
    13251 => x"a0220800", 13252 => x"59640008", 13253 => x"59630010",
    13254 => x"59610018", 13255 => x"43850010", 13256 => x"43860011",
    13257 => x"3ca50008", 13258 => x"b8a62800", 13259 => x"3ca5000d",
    13260 => x"3806cafe", 13261 => x"b8852000", 13262 => x"59640008",
    13263 => x"43840012", 13264 => x"43850013", 13265 => x"3c840008",
    13266 => x"b8852000", 13267 => x"3c84000d", 13268 => x"34050001",
    13269 => x"b8641800", 13270 => x"59630010", 13271 => x"43830014",
    13272 => x"43840015", 13273 => x"3c630008", 13274 => x"b8641800",
    13275 => x"3c63000d", 13276 => x"b8230800", 13277 => x"78030001",
    13278 => x"3863579c", 13279 => x"59610018", 13280 => x"28640000",
    13281 => x"b9600800", 13282 => x"e000000b", 13283 => x"28230000",
    13284 => x"0067000d", 13285 => x"20e7ffff", 13286 => x"5ce60006",
    13287 => x"20670007", 13288 => x"5ce50004", 13289 => x"a0621800",
    13290 => x"b8641800", 13291 => x"58230000", 13292 => x"34210008",
    13293 => x"5581fff6", 13294 => x"78040001", 13295 => x"38845798",
    13296 => x"78030001", 13297 => x"b9600800", 13298 => x"34020000",
    13299 => x"34070aaa", 13300 => x"34060007", 13301 => x"28850000",
    13302 => x"3863726c", 13303 => x"e0000010", 13304 => x"28240000",
    13305 => x"0088000d", 13306 => x"2108ffff", 13307 => x"5d07000b",
    13308 => x"00880007", 13309 => x"2108001f", 13310 => x"5d060008",
    13311 => x"a0852000", 13312 => x"58240000", 13313 => x"28620000",
    13314 => x"3c42000d", 13315 => x"b8442000", 13316 => x"58240000",
    13317 => x"b8201000", 13318 => x"34210008", 13319 => x"5581fff1",
    13320 => x"78010001", 13321 => x"38218f94", 13322 => x"28210000",
    13323 => x"34030000", 13324 => x"58200014", 13325 => x"e000000f",
    13326 => x"29640000", 13327 => x"29660004", 13328 => x"356b0008",
    13329 => x"20850fff", 13330 => x"3cc60014", 13331 => x"0084000c",
    13332 => x"58250018", 13333 => x"b8c42000", 13334 => x"3c840008",
    13335 => x"2066003f", 13336 => x"38840040", 13337 => x"b8862000",
    13338 => x"58240014", 13339 => x"34630001", 13340 => x"558bfff2",
    13341 => x"4440000b", 13342 => x"78050001", 13343 => x"38a55798",
    13344 => x"28440000", 13345 => x"28a30000", 13346 => x"78050001",
    13347 => x"38a557a0", 13348 => x"a0831800", 13349 => x"28a40000",
    13350 => x"b8641800", 13351 => x"58430000", 13352 => x"34020080",
    13353 => x"58220014", 13354 => x"2b9d0004", 13355 => x"2b8b000c",
    13356 => x"2b8c0008", 13357 => x"379c0014", 13358 => x"c3a00000",
    13359 => x"78030001", 13360 => x"38638f90", 13361 => x"44400004",
    13362 => x"28620000", 13363 => x"58410004", 13364 => x"c3a00000",
    13365 => x"28620000", 13366 => x"58410008", 13367 => x"c3a00000",
    13368 => x"78030001", 13369 => x"38638f90", 13370 => x"44400004",
    13371 => x"28620000", 13372 => x"58410004", 13373 => x"c3a00000",
    13374 => x"28620000", 13375 => x"58410008", 13376 => x"c3a00000",
    13377 => x"3401012c", 13378 => x"34000000", 13379 => x"3421ffff",
    13380 => x"5c20fffe", 13381 => x"c3a00000", 13382 => x"379cfff8",
    13383 => x"5b8b0008", 13384 => x"5b9d0004", 13385 => x"202100ff",
    13386 => x"3c2b0003", 13387 => x"78020001", 13388 => x"38426d0c",
    13389 => x"b44b5800", 13390 => x"29610004", 13391 => x"34020000",
    13392 => x"fbffffdf", 13393 => x"fbfffff0", 13394 => x"29610000",
    13395 => x"34020000", 13396 => x"fbffffdb", 13397 => x"fbffffec",
    13398 => x"2b9d0004", 13399 => x"2b8b0008", 13400 => x"379c0008",
    13401 => x"c3a00000", 13402 => x"379cfff8", 13403 => x"5b8b0008",
    13404 => x"5b9d0004", 13405 => x"202100ff", 13406 => x"3c2b0003",
    13407 => x"78020001", 13408 => x"38426d0c", 13409 => x"b44b5800",
    13410 => x"29610004", 13411 => x"34020001", 13412 => x"fbffffcb",
    13413 => x"fbffffdc", 13414 => x"29610000", 13415 => x"34020001",
    13416 => x"fbffffc7", 13417 => x"fbffffd8", 13418 => x"29610004",
    13419 => x"34020000", 13420 => x"fbffffc3", 13421 => x"fbffffd4",
    13422 => x"29610000", 13423 => x"34020000", 13424 => x"fbffffbf",
    13425 => x"fbffffd0", 13426 => x"2b9d0004", 13427 => x"2b8b0008",
    13428 => x"379c0008", 13429 => x"c3a00000", 13430 => x"379cfff8",
    13431 => x"5b8b0008", 13432 => x"5b9d0004", 13433 => x"202100ff",
    13434 => x"3c2b0003", 13435 => x"78020001", 13436 => x"38426d0c",
    13437 => x"b44b5800", 13438 => x"29610004", 13439 => x"34020000",
    13440 => x"fbffffaf", 13441 => x"fbffffc0", 13442 => x"29610000",
    13443 => x"34020001", 13444 => x"fbffffab", 13445 => x"fbffffbc",
    13446 => x"29610004", 13447 => x"34020001", 13448 => x"fbffffa7",
    13449 => x"fbffffb8", 13450 => x"2b9d0004", 13451 => x"2b8b0008",
    13452 => x"379c0008", 13453 => x"c3a00000", 13454 => x"379cffec",
    13455 => x"5b8b0014", 13456 => x"5b8c0010", 13457 => x"5b8d000c",
    13458 => x"5b8e0008", 13459 => x"5b9d0004", 13460 => x"202100ff",
    13461 => x"78030001", 13462 => x"3c2b0003", 13463 => x"38636d0c",
    13464 => x"204e00ff", 13465 => x"340d0008", 13466 => x"b46b5800",
    13467 => x"29610004", 13468 => x"21c20080", 13469 => x"35adffff",
    13470 => x"fbffff91", 13471 => x"fbffffa2", 13472 => x"29610000",
    13473 => x"34020001", 13474 => x"3dce0001", 13475 => x"fbffff8c",
    13476 => x"fbffff9d", 13477 => x"29610000", 13478 => x"34020000",
    13479 => x"21ad00ff", 13480 => x"fbffff87", 13481 => x"356c0004",
    13482 => x"fbffff97", 13483 => x"21ce00ff", 13484 => x"5da0ffef",
    13485 => x"29810000", 13486 => x"34020001", 13487 => x"fbffff80",
    13488 => x"fbffff91", 13489 => x"29610000", 13490 => x"34020001",
    13491 => x"fbffff7c", 13492 => x"fbffff8d", 13493 => x"78010001",
    13494 => x"38218f90", 13495 => x"28210000", 13496 => x"298d0000",
    13497 => x"34020000", 13498 => x"28210004", 13499 => x"a02d6800",
    13500 => x"29610000", 13501 => x"fbffff72", 13502 => x"fbffff83",
    13503 => x"29810000", 13504 => x"34020000", 13505 => x"fbffff6e",
    13506 => x"fbffff7f", 13507 => x"7da10000", 13508 => x"2b9d0004",
    13509 => x"2b8b0014", 13510 => x"2b8c0010", 13511 => x"2b8d000c",
    13512 => x"2b8e0008", 13513 => x"379c0014", 13514 => x"c3a00000",
    13515 => x"379cffe0", 13516 => x"5b8b0020", 13517 => x"5b8c001c",
    13518 => x"5b8d0018", 13519 => x"5b8e0014", 13520 => x"5b8f0010",
    13521 => x"5b90000c", 13522 => x"5b910008", 13523 => x"5b9d0004",
    13524 => x"202100ff", 13525 => x"3c2b0003", 13526 => x"78040001",
    13527 => x"38846d0c", 13528 => x"b48b5800", 13529 => x"29610004",
    13530 => x"b8407800", 13531 => x"34020001", 13532 => x"207000ff",
    13533 => x"fbffff52", 13534 => x"fbffff63", 13535 => x"29610000",
    13536 => x"34020000", 13537 => x"780d0001", 13538 => x"fbffff4d",
    13539 => x"340c0000", 13540 => x"fbffff5d", 13541 => x"340e0000",
    13542 => x"39ad8f90", 13543 => x"34110008", 13544 => x"29610000",
    13545 => x"34020001", 13546 => x"3d8c0001", 13547 => x"fbffff44",
    13548 => x"fbffff55", 13549 => x"29a10000", 13550 => x"29620004",
    13551 => x"218c00ff", 13552 => x"28210004", 13553 => x"a0220800",
    13554 => x"44200002", 13555 => x"398c0001", 13556 => x"29610000",
    13557 => x"34020000", 13558 => x"35ce0001", 13559 => x"fbffff38",
    13560 => x"fbffff49", 13561 => x"5dd1ffef", 13562 => x"46000004",
    13563 => x"29610004", 13564 => x"34020001", 13565 => x"e0000003",
    13566 => x"29610004", 13567 => x"34020000", 13568 => x"fbffff2f",
    13569 => x"fbffff40", 13570 => x"29610000", 13571 => x"34020001",
    13572 => x"fbffff2b", 13573 => x"fbffff3c", 13574 => x"29610000",
    13575 => x"34020000", 13576 => x"fbffff27", 13577 => x"fbffff38",
    13578 => x"31ec0000", 13579 => x"2b9d0004", 13580 => x"2b8b0020",
    13581 => x"2b8c001c", 13582 => x"2b8d0018", 13583 => x"2b8e0014",
    13584 => x"2b8f0010", 13585 => x"2b90000c", 13586 => x"2b910008",
    13587 => x"379c0020", 13588 => x"c3a00000", 13589 => x"379cfff8",
    13590 => x"5b8b0008", 13591 => x"5b9d0004", 13592 => x"202100ff",
    13593 => x"3c2b0003", 13594 => x"78020001", 13595 => x"38426d0c",
    13596 => x"b44b5800", 13597 => x"29610000", 13598 => x"34020001",
    13599 => x"fbffff10", 13600 => x"fbffff21", 13601 => x"29610004",
    13602 => x"34020001", 13603 => x"fbffff0c", 13604 => x"fbffff1d",
    13605 => x"2b9d0004", 13606 => x"2b8b0008", 13607 => x"379c0008",
    13608 => x"c3a00000", 13609 => x"379cfff4", 13610 => x"5b8b000c",
    13611 => x"5b8c0008", 13612 => x"5b9d0004", 13613 => x"202b00ff",
    13614 => x"b9600800", 13615 => x"204c00ff", 13616 => x"fbffff16",
    13617 => x"3d820001", 13618 => x"b9600800", 13619 => x"204200fe",
    13620 => x"fbffff5a", 13621 => x"b8206000", 13622 => x"b9600800",
    13623 => x"fbffff3f", 13624 => x"65810000", 13625 => x"2b9d0004",
    13626 => x"2b8b000c", 13627 => x"2b8c0008", 13628 => x"379c000c",
    13629 => x"c3a00000", 13630 => x"379cffe8", 13631 => x"5b8b0018",
    13632 => x"5b8c0014", 13633 => x"5b8d0010", 13634 => x"5b8e000c",
    13635 => x"5b8f0008", 13636 => x"5b9d0004", 13637 => x"780b0001",
    13638 => x"396b8f4c", 13639 => x"296d000c", 13640 => x"296f0004",
    13641 => x"b8206000", 13642 => x"3dad0002", 13643 => x"c84f0800",
    13644 => x"b9a01000", 13645 => x"b8607000", 13646 => x"f8001593",
    13647 => x"b42f1000", 13648 => x"b5af6800", 13649 => x"b44e0800",
    13650 => x"542d0006", 13651 => x"b9800800", 13652 => x"b9c01800",
    13653 => x"f80015dd", 13654 => x"b8206000", 13655 => x"e0000009",
    13656 => x"c9a26800", 13657 => x"b9a01800", 13658 => x"b9800800",
    13659 => x"f80015d7", 13660 => x"29620004", 13661 => x"b58d0800",
    13662 => x"c9cd1800", 13663 => x"f80015d3", 13664 => x"b9800800",
    13665 => x"2b9d0004", 13666 => x"2b8b0018", 13667 => x"2b8c0014",
    13668 => x"2b8d0010", 13669 => x"2b8e000c", 13670 => x"2b8f0008",
    13671 => x"379c0018", 13672 => x"c3a00000", 13673 => x"379cffe8",
    13674 => x"5b8b0018", 13675 => x"5b8c0014", 13676 => x"5b8d0010",
    13677 => x"5b8e000c", 13678 => x"5b8f0008", 13679 => x"5b9d0004",
    13680 => x"780b0001", 13681 => x"396b8f4c", 13682 => x"296f000c",
    13683 => x"296e0004", 13684 => x"b8406800", 13685 => x"3def0002",
    13686 => x"c82e0800", 13687 => x"b9e01000", 13688 => x"f8001569",
    13689 => x"b42e6000", 13690 => x"b58d0800", 13691 => x"b5ee7000",
    13692 => x"542e0006", 13693 => x"b9800800", 13694 => x"34020000",
    13695 => x"b9a01800", 13696 => x"f8001630", 13697 => x"e000000b",
    13698 => x"c9cc7000", 13699 => x"34020000", 13700 => x"b9c01800",
    13701 => x"b9800800", 13702 => x"f800162a", 13703 => x"29610004",
    13704 => x"34020000", 13705 => x"c9ae1800", 13706 => x"f8001626",
    13707 => x"b9800800", 13708 => x"2b9d0004", 13709 => x"2b8b0018",
    13710 => x"2b8c0014", 13711 => x"2b8d0010", 13712 => x"2b8e000c",
    13713 => x"2b8f0008", 13714 => x"379c0018", 13715 => x"c3a00000",
    13716 => x"379cfff4", 13717 => x"5b8b000c", 13718 => x"5b8c0008",
    13719 => x"5b9d0004", 13720 => x"780c0001", 13721 => x"398c8fa4",
    13722 => x"29810000", 13723 => x"780b0001", 13724 => x"396b8f4c",
    13725 => x"58200000", 13726 => x"34020200", 13727 => x"78010001",
    13728 => x"382183b8", 13729 => x"5962000c", 13730 => x"34020800",
    13731 => x"59610004", 13732 => x"59610000", 13733 => x"fbffffc4",
    13734 => x"29620004", 13735 => x"29810000", 13736 => x"58220008",
    13737 => x"2962000c", 13738 => x"5822000c", 13739 => x"34020002",
    13740 => x"5822004c", 13741 => x"34020400", 13742 => x"58220000",
    13743 => x"2b9d0004", 13744 => x"2b8b000c", 13745 => x"2b8c0008",
    13746 => x"379c000c", 13747 => x"c3a00000", 13748 => x"379cfff4",
    13749 => x"5b8b000c", 13750 => x"5b8c0008", 13751 => x"5b9d0004",
    13752 => x"780b0001", 13753 => x"396b8fa4", 13754 => x"29630000",
    13755 => x"340c0002", 13756 => x"78010001", 13757 => x"586c0040",
    13758 => x"78020001", 13759 => x"586c004c", 13760 => x"38218f4c",
    13761 => x"384283b8", 13762 => x"58220004", 13763 => x"00420002",
    13764 => x"34040800", 13765 => x"5824000c", 13766 => x"344401ff",
    13767 => x"3c840010", 13768 => x"2042ffff", 13769 => x"b8821000",
    13770 => x"58620020", 13771 => x"78020001", 13772 => x"38427fb8",
    13773 => x"58220014", 13774 => x"34020100", 13775 => x"5822001c",
    13776 => x"58200020", 13777 => x"58200024", 13778 => x"fbffffc2",
    13779 => x"29610000", 13780 => x"582c0044", 13781 => x"2b9d0004",
    13782 => x"2b8b000c", 13783 => x"2b8c0008", 13784 => x"379c000c",
    13785 => x"c3a00000", 13786 => x"379cffc8", 13787 => x"5b8b0024",
    13788 => x"5b8c0020", 13789 => x"5b8d001c", 13790 => x"5b8e0018",
    13791 => x"5b8f0014", 13792 => x"5b900010", 13793 => x"5b91000c",
    13794 => x"5b920008", 13795 => x"5b9d0004", 13796 => x"b8805800",
    13797 => x"78040001", 13798 => x"38848fa4", 13799 => x"b8608000",
    13800 => x"28830000", 13801 => x"b8209000", 13802 => x"b8408800",
    13803 => x"2861004c", 13804 => x"340d0000", 13805 => x"20210002",
    13806 => x"4420008b", 13807 => x"780e0001", 13808 => x"39ce8f4c",
    13809 => x"29c20000", 13810 => x"28440000", 13811 => x"4804000a",
    13812 => x"28610000", 13813 => x"20210200", 13814 => x"5c200005",
    13815 => x"78010001", 13816 => x"382153c0", 13817 => x"b8801800",
    13818 => x"fbfffb85", 13819 => x"fbffff99", 13820 => x"e000007d",
    13821 => x"20810001", 13822 => x"208c0ffe", 13823 => x"c9816000",
    13824 => x"358f0003", 13825 => x"01ef0002", 13826 => x"78034000",
    13827 => x"a0831800", 13828 => x"35ef0001", 13829 => x"340dffff",
    13830 => x"5c600054", 13831 => x"7d610000", 13832 => x"0084001d",
    13833 => x"a0812000", 13834 => x"4483003e", 13835 => x"b44c1000",
    13836 => x"34030004", 13837 => x"37810034", 13838 => x"fbffff30",
    13839 => x"29c30000", 13840 => x"358dfffa", 13841 => x"358cfffe",
    13842 => x"b46c1000", 13843 => x"3781003a", 13844 => x"34030002",
    13845 => x"fbffff29", 13846 => x"78010001", 13847 => x"382157a4",
    13848 => x"282c0000", 13849 => x"37820030", 13850 => x"37810028",
    13851 => x"2b8e0034", 13852 => x"f800049e", 13853 => x"78020001",
    13854 => x"384257a8", 13855 => x"28410000", 13856 => x"a1cc6000",
    13857 => x"01ce001c", 13858 => x"502c000e", 13859 => x"78030001",
    13860 => x"386357ac", 13861 => x"2b820030", 13862 => x"28610000",
    13863 => x"54410009", 13864 => x"2b82002c", 13865 => x"2b810028",
    13866 => x"3444ffff", 13867 => x"f4441000", 13868 => x"3421ffff",
    13869 => x"b4410800", 13870 => x"5b810028", 13871 => x"5b84002c",
    13872 => x"78020001", 13873 => x"38425784", 13874 => x"28410000",
    13875 => x"2b82002c", 13876 => x"2183000f", 13877 => x"c86e1800",
    13878 => x"a0410800", 13879 => x"5961000c", 13880 => x"6461fff1",
    13881 => x"64630001", 13882 => x"59600008", 13883 => x"b8231800",
    13884 => x"44600004", 13885 => x"34010001", 13886 => x"59610004",
    13887 => x"e0000002", 13888 => x"59600004", 13889 => x"2f81003a",
    13890 => x"3d8c0003", 13891 => x"20210800", 13892 => x"64210000",
    13893 => x"596c0010", 13894 => x"31610000", 13895 => x"b9a06000",
    13896 => x"358dfff2", 13897 => x"520d0002", 13898 => x"ba006800",
    13899 => x"780b0001", 13900 => x"396b8f4c", 13901 => x"29610024",
    13902 => x"29620000", 13903 => x"3403000e", 13904 => x"34210001",
    13905 => x"59610024", 13906 => x"34420004", 13907 => x"ba400800",
    13908 => x"fbfffeea", 13909 => x"29630000", 13910 => x"ba200800",
    13911 => x"34620012", 13912 => x"b9a01800", 13913 => x"fbfffee5",
    13914 => x"780b0001", 13915 => x"396b8f4c", 13916 => x"3dee0002",
    13917 => x"29610000", 13918 => x"b9c01000", 13919 => x"fbffff0a",
    13920 => x"78030001", 13921 => x"38638fa4", 13922 => x"286c0000",
    13923 => x"29610000", 13924 => x"598f0010", 13925 => x"2962000c",
    13926 => x"296f0004", 13927 => x"3c420002", 13928 => x"c82f0800",
    13929 => x"b42e0800", 13930 => x"f8001477", 13931 => x"b42f0800",
    13932 => x"59610000", 13933 => x"29820010", 13934 => x"28210000",
    13935 => x"4801000a", 13936 => x"29810000", 13937 => x"20210200",
    13938 => x"44200002", 13939 => x"fbffff21", 13940 => x"78010001",
    13941 => x"38218fa4", 13942 => x"28210000", 13943 => x"34020002",
    13944 => x"5822004c", 13945 => x"b9a00800", 13946 => x"2b9d0004",
    13947 => x"2b8b0024", 13948 => x"2b8c0020", 13949 => x"2b8d001c",
    13950 => x"2b8e0018", 13951 => x"2b8f0014", 13952 => x"2b900010",
    13953 => x"2b91000c", 13954 => x"2b920008", 13955 => x"379c0038",
    13956 => x"c3a00000", 13957 => x"379cffd4", 13958 => x"5b8b0020",
    13959 => x"5b8c001c", 13960 => x"5b8d0018", 13961 => x"5b8e0014",
    13962 => x"5b8f0010", 13963 => x"5b90000c", 13964 => x"5b910008",
    13965 => x"5b9d0004", 13966 => x"780b0001", 13967 => x"78050001",
    13968 => x"396b8f4c", 13969 => x"38a58fa4", 13970 => x"b8208000",
    13971 => x"34010100", 13972 => x"5961001c", 13973 => x"59610018",
    13974 => x"b8806000", 13975 => x"28a10000", 13976 => x"78040001",
    13977 => x"38847fb8", 13978 => x"2e0e000c", 13979 => x"59640014",
    13980 => x"59640010", 13981 => x"58240004", 13982 => x"38018100",
    13983 => x"fdc17000", 13984 => x"3401fffc", 13985 => x"c80e7000",
    13986 => x"a1c17000", 13987 => x"35ce0012", 13988 => x"b5c36800",
    13989 => x"b8800800", 13990 => x"b8408800", 13991 => x"b8607800",
    13992 => x"34020000", 13993 => x"35a30004", 13994 => x"f8001506",
    13995 => x"29610010", 13996 => x"b9c01800", 13997 => x"ba001000",
    13998 => x"34210004", 13999 => x"f8001483", 14000 => x"29610010",
    14001 => x"35ce0004", 14002 => x"ba201000", 14003 => x"b42e0800",
    14004 => x"b9e01800", 14005 => x"f800147d", 14006 => x"3401003b",
    14007 => x"502d0002", 14008 => x"e0000002", 14009 => x"340d003c",
    14010 => x"35a30001", 14011 => x"7d810000", 14012 => x"00630001",
    14013 => x"3c21001e", 14014 => x"78048000", 14015 => x"b8642000",
    14016 => x"b8812000", 14017 => x"78010001", 14018 => x"38218f4c",
    14019 => x"28220010", 14020 => x"3c630002", 14021 => x"78010001",
    14022 => x"58440000", 14023 => x"38218fa4", 14024 => x"b4431000",
    14025 => x"58400000", 14026 => x"28220000", 14027 => x"340b0000",
    14028 => x"b8207800", 14029 => x"28430000", 14030 => x"341003e8",
    14031 => x"38630001", 14032 => x"58430000", 14033 => x"29e10000",
    14034 => x"282e0000", 14035 => x"21c10002", 14036 => x"5c200009",
    14037 => x"34010001", 14038 => x"356b0001", 14039 => x"f800006d",
    14040 => x"5d70fff9", 14041 => x"78010001", 14042 => x"382153e0",
    14043 => x"b9c01000", 14044 => x"fbfffaa3", 14045 => x"4580003e",
    14046 => x"780b0001", 14047 => x"340e0000", 14048 => x"396b8fa4",
    14049 => x"340f0064", 14050 => x"29610000", 14051 => x"28220000",
    14052 => x"20420800", 14053 => x"5c40000a", 14054 => x"34010001",
    14055 => x"35ce0001", 14056 => x"f800005c", 14057 => x"5dcffff9",
    14058 => x"78010001", 14059 => x"38215410", 14060 => x"fbfffa93",
    14061 => x"340e0000", 14062 => x"e0000003", 14063 => x"282e0014",
    14064 => x"21ce0001", 14065 => x"78010001", 14066 => x"38218fa4",
    14067 => x"28210000", 14068 => x"78020001", 14069 => x"384257a4",
    14070 => x"282b0018", 14071 => x"28210014", 14072 => x"28410000",
    14073 => x"3782002c", 14074 => x"a1615800", 14075 => x"37810024",
    14076 => x"f80003be", 14077 => x"78030001", 14078 => x"386357a8",
    14079 => x"28610000", 14080 => x"502b000e", 14081 => x"78030001",
    14082 => x"386357ac", 14083 => x"2b82002c", 14084 => x"28610000",
    14085 => x"54410009", 14086 => x"2b830028", 14087 => x"2b820024",
    14088 => x"3461ffff", 14089 => x"f4611800", 14090 => x"3442ffff",
    14091 => x"b4621000", 14092 => x"5b820024", 14093 => x"5b810028",
    14094 => x"2b810024", 14095 => x"318e0000", 14096 => x"3d6b0003",
    14097 => x"59810008", 14098 => x"2b810028", 14099 => x"59800004",
    14100 => x"598b0010", 14101 => x"5981000c", 14102 => x"78010001",
    14103 => x"38218f4c", 14104 => x"28220020", 14105 => x"34420001",
    14106 => x"58220020", 14107 => x"b9a00800", 14108 => x"2b9d0004",
    14109 => x"2b8b0020", 14110 => x"2b8c001c", 14111 => x"2b8d0018",
    14112 => x"2b8e0014", 14113 => x"2b8f0010", 14114 => x"2b90000c",
    14115 => x"2b910008", 14116 => x"379c002c", 14117 => x"c3a00000",
    14118 => x"78030001", 14119 => x"38638f4c", 14120 => x"28640020",
    14121 => x"58240000", 14122 => x"28610024", 14123 => x"58410000",
    14124 => x"c3a00000", 14125 => x"78020001", 14126 => x"38428fa8",
    14127 => x"28420000", 14128 => x"78030001", 14129 => x"38638f90",
    14130 => x"58620000", 14131 => x"44200005", 14132 => x"28430010",
    14133 => x"78018000", 14134 => x"b8610800", 14135 => x"e0000006",
    14136 => x"78040001", 14137 => x"38845784", 14138 => x"28430010",
    14139 => x"28810000", 14140 => x"a0610800", 14141 => x"58410010",
    14142 => x"c3a00000", 14143 => x"78010001", 14144 => x"38218f90",
    14145 => x"28210000", 14146 => x"28210014", 14147 => x"c3a00000",
    14148 => x"78020001", 14149 => x"38428f90", 14150 => x"28420000",
    14151 => x"28430014", 14152 => x"b4230800", 14153 => x"28430014",
    14154 => x"c8611800", 14155 => x"4803fffe", 14156 => x"c3a00000",
    14157 => x"78010001", 14158 => x"38218f90", 14159 => x"28210000",
    14160 => x"28210004", 14161 => x"20210080", 14162 => x"64210000",
    14163 => x"c3a00000", 14164 => x"379cffe0", 14165 => x"5b8b001c",
    14166 => x"5b8c0018", 14167 => x"5b8d0014", 14168 => x"5b8e0010",
    14169 => x"5b8f000c", 14170 => x"5b900008", 14171 => x"5b9d0004",
    14172 => x"b8208000", 14173 => x"34010001", 14174 => x"fbfffdb7",
    14175 => x"34010001", 14176 => x"fbfffce6", 14177 => x"340200a0",
    14178 => x"34010001", 14179 => x"fbfffd2b", 14180 => x"34020000",
    14181 => x"34010001", 14182 => x"fbfffd28", 14183 => x"34010001",
    14184 => x"fbfffcf2", 14185 => x"340200a1", 14186 => x"34010001",
    14187 => x"fbfffd23", 14188 => x"378d0023", 14189 => x"b9a01000",
    14190 => x"34030001", 14191 => x"34010001", 14192 => x"fbfffd5b",
    14193 => x"34010001", 14194 => x"fbfffd04", 14195 => x"34010001",
    14196 => x"438c0023", 14197 => x"fbfffcd1", 14198 => x"34010001",
    14199 => x"340200a1", 14200 => x"fbfffd16", 14201 => x"340bffd9",
    14202 => x"340f000f", 14203 => x"340e0017", 14204 => x"34030000",
    14205 => x"34010001", 14206 => x"b9a01000", 14207 => x"fbfffd4c",
    14208 => x"43830023", 14209 => x"b5836000", 14210 => x"218c00ff",
    14211 => x"556f0003", 14212 => x"b60b0800", 14213 => x"30230000",
    14214 => x"356b0001", 14215 => x"5d6efff5", 14216 => x"37820023",
    14217 => x"34030001", 14218 => x"34010001", 14219 => x"fbfffd40",
    14220 => x"34010001", 14221 => x"fbfffce9", 14222 => x"43810023",
    14223 => x"fc2c6000", 14224 => x"c80c0800", 14225 => x"2b9d0004",
    14226 => x"2b8b001c", 14227 => x"2b8c0018", 14228 => x"2b8d0014",
    14229 => x"2b8e0010", 14230 => x"2b8f000c", 14231 => x"2b900008",
    14232 => x"379c0020", 14233 => x"c3a00000", 14234 => x"379cffd0",
    14235 => x"5b8b0010", 14236 => x"5b8c000c", 14237 => x"5b8d0008",
    14238 => x"5b9d0004", 14239 => x"780b0001", 14240 => x"396b8c24",
    14241 => x"31600000", 14242 => x"fbffffab", 14243 => x"3403ffed",
    14244 => x"44200023", 14245 => x"b9600800", 14246 => x"fbffffae",
    14247 => x"b8206000", 14248 => x"3403fffb", 14249 => x"5c20001e",
    14250 => x"378d0014", 14251 => x"b9601000", 14252 => x"34030010",
    14253 => x"b9a00800", 14254 => x"f8001534", 14255 => x"b9a00800",
    14256 => x"f80004a2", 14257 => x"78020001", 14258 => x"38428bc0",
    14259 => x"5c2c0005", 14260 => x"34010001", 14261 => x"58410000",
    14262 => x"3403fffa", 14263 => x"e0000010", 14264 => x"2b830028",
    14265 => x"78010001", 14266 => x"38218bb8", 14267 => x"58230000",
    14268 => x"2b83002c", 14269 => x"78010001", 14270 => x"38218bbc",
    14271 => x"58230000", 14272 => x"2b830024", 14273 => x"78010001",
    14274 => x"38216d1c", 14275 => x"58230000", 14276 => x"34010002",
    14277 => x"58410000", 14278 => x"34030000", 14279 => x"b8600800",
    14280 => x"2b9d0004", 14281 => x"2b8b0010", 14282 => x"2b8c000c",
    14283 => x"2b8d0008", 14284 => x"379c0030", 14285 => x"c3a00000",
    14286 => x"379cffe0", 14287 => x"5b9b0008", 14288 => x"341b0020",
    14289 => x"b77cd800", 14290 => x"5b8b0020", 14291 => x"5b8c001c",
    14292 => x"5b8d0018", 14293 => x"5b8e0014", 14294 => x"5b8f0010",
    14295 => x"5b90000c", 14296 => x"5b9d0004", 14297 => x"780b0001",
    14298 => x"780c0001", 14299 => x"bb807800", 14300 => x"34020001",
    14301 => x"396b6df8", 14302 => x"398c5440", 14303 => x"e0000012",
    14304 => x"bb808000", 14305 => x"379cffe4", 14306 => x"378e000b",
    14307 => x"01ce0003", 14308 => x"35a2002c", 14309 => x"3dce0003",
    14310 => x"34030014", 14311 => x"b9c00800", 14312 => x"f800134a",
    14313 => x"31c00013", 14314 => x"29a20020", 14315 => x"29630074",
    14316 => x"b9800800", 14317 => x"b9c02000", 14318 => x"fbfff991",
    14319 => x"34020000", 14320 => x"ba00e000", 14321 => x"b9600800",
    14322 => x"f80011a9", 14323 => x"b8206800", 14324 => x"5c20ffec",
    14325 => x"b9e0e000", 14326 => x"2b9d0004", 14327 => x"2b8b0020",
    14328 => x"2b8c001c", 14329 => x"2b8d0018", 14330 => x"2b8e0014",
    14331 => x"2b8f0010", 14332 => x"2b90000c", 14333 => x"2b9b0008",
    14334 => x"379c0020", 14335 => x"c3a00000", 14336 => x"379cffec",
    14337 => x"5b8b0014", 14338 => x"5b8c0010", 14339 => x"5b8d000c",
    14340 => x"5b8e0008", 14341 => x"5b9d0004", 14342 => x"780b0001",
    14343 => x"396b8bc4", 14344 => x"29610000", 14345 => x"5c200007",
    14346 => x"78010001", 14347 => x"38216df8", 14348 => x"f800116d",
    14349 => x"29610000", 14350 => x"34210001", 14351 => x"59610000",
    14352 => x"780b0001", 14353 => x"396b6d20", 14354 => x"780c0001",
    14355 => x"356d00d8", 14356 => x"398c6df8", 14357 => x"e0000009",
    14358 => x"29620008", 14359 => x"2963000c", 14360 => x"29640010",
    14361 => x"296e0000", 14362 => x"b9800800", 14363 => x"f8001232",
    14364 => x"59c10000", 14365 => x"356b0018", 14366 => x"5d6dfff8",
    14367 => x"2b9d0004", 14368 => x"2b8b0014", 14369 => x"2b8c0010",
    14370 => x"2b8d000c", 14371 => x"2b8e0008", 14372 => x"379c0014",
    14373 => x"c3a00000", 14374 => x"379cfff4", 14375 => x"5b8b000c",
    14376 => x"5b8c0008", 14377 => x"5b9d0004", 14378 => x"34020000",
    14379 => x"b8206000", 14380 => x"f8000461", 14381 => x"b8205800",
    14382 => x"4c200005", 14383 => x"78010001", 14384 => x"38215468",
    14385 => x"b9601000", 14386 => x"e0000004", 14387 => x"29820000",
    14388 => x"78010001", 14389 => x"38215494", 14390 => x"fbfff949",
    14391 => x"b9600800", 14392 => x"2b9d0004", 14393 => x"2b8b000c",
    14394 => x"2b8c0008", 14395 => x"379c000c", 14396 => x"c3a00000",
    14397 => x"379cfffc", 14398 => x"5b9d0004", 14399 => x"78010001",
    14400 => x"38218bc8", 14401 => x"58200000", 14402 => x"78020001",
    14403 => x"78010001", 14404 => x"38218bdc", 14405 => x"38428bcc",
    14406 => x"3403ffff", 14407 => x"58230000", 14408 => x"58430000",
    14409 => x"58200008", 14410 => x"58400008", 14411 => x"58400004",
    14412 => x"58200004", 14413 => x"5840000c", 14414 => x"5820000c",
    14415 => x"34020000", 14416 => x"34010000", 14417 => x"f8000f20",
    14418 => x"2b9d0004", 14419 => x"379c0004", 14420 => x"c3a00000",
    14421 => x"379cfff4", 14422 => x"5b8b000c", 14423 => x"5b8c0008",
    14424 => x"5b9d0004", 14425 => x"b8206000", 14426 => x"34010000",
    14427 => x"f8000fbf", 14428 => x"b8205800", 14429 => x"34020000",
    14430 => x"5c200081", 14431 => x"fbfffacb", 14432 => x"78030001",
    14433 => x"38638bcc", 14434 => x"28650008", 14435 => x"78020001",
    14436 => x"38428bc8", 14437 => x"b8202000", 14438 => x"28420000",
    14439 => x"44ab0004", 14440 => x"34010001", 14441 => x"5ca1001d",
    14442 => x"e0000010", 14443 => x"34010001", 14444 => x"44810005",
    14445 => x"28610004", 14446 => x"34210001", 14447 => x"58610004",
    14448 => x"e0000002", 14449 => x"58600004", 14450 => x"78030001",
    14451 => x"38638bcc", 14452 => x"28650004", 14453 => x"34010004",
    14454 => x"4c250010", 14455 => x"34010001", 14456 => x"58610008",
    14457 => x"e0000002", 14458 => x"44850003", 14459 => x"58600004",
    14460 => x"e000000a", 14461 => x"28650004", 14462 => x"34010004",
    14463 => x"34a50001", 14464 => x"58650004", 14465 => x"4c250005",
    14466 => x"34010002", 14467 => x"58610008", 14468 => x"3441fe0c",
    14469 => x"5861000c", 14470 => x"78030001", 14471 => x"38638bdc",
    14472 => x"28650008", 14473 => x"44a00004", 14474 => x"34010001",
    14475 => x"5ca1001c", 14476 => x"e000000f", 14477 => x"44850005",
    14478 => x"28610004", 14479 => x"34210001", 14480 => x"58610004",
    14481 => x"e0000002", 14482 => x"58600004", 14483 => x"78030001",
    14484 => x"38638bdc", 14485 => x"28640004", 14486 => x"34010004",
    14487 => x"4c240010", 14488 => x"34010001", 14489 => x"58610008",
    14490 => x"e0000002", 14491 => x"44800003", 14492 => x"58600004",
    14493 => x"e000000a", 14494 => x"28640004", 14495 => x"34010004",
    14496 => x"34840001", 14497 => x"58640004", 14498 => x"4c240005",
    14499 => x"34010002", 14500 => x"58610008", 14501 => x"3441fe0c",
    14502 => x"5861000c", 14503 => x"3401251b", 14504 => x"4c220030",
    14505 => x"78020001", 14506 => x"38428bcc", 14507 => x"28440008",
    14508 => x"34010002", 14509 => x"3402ffff", 14510 => x"5c810031",
    14511 => x"78030001", 14512 => x"38638bdc", 14513 => x"28610008",
    14514 => x"5c24002d", 14515 => x"2862000c", 14516 => x"34011f3f",
    14517 => x"e0000002", 14518 => x"3442e0c0", 14519 => x"4841ffff",
    14520 => x"78030001", 14521 => x"38638bdc", 14522 => x"5862000c",
    14523 => x"78030001", 14524 => x"38638bcc", 14525 => x"2863000c",
    14526 => x"34011f3f", 14527 => x"e0000002", 14528 => x"3463e0c0",
    14529 => x"4861ffff", 14530 => x"78040001", 14531 => x"38848bcc",
    14532 => x"5883000c", 14533 => x"4c620003", 14534 => x"3444f060",
    14535 => x"e0000004", 14536 => x"34040000", 14537 => x"4c430002",
    14538 => x"34440fa0", 14539 => x"b4831800", 14540 => x"0062001f",
    14541 => x"b4431800", 14542 => x"14620001", 14543 => x"4c400003",
    14544 => x"34421f40", 14545 => x"e0000004", 14546 => x"34011f3f",
    14547 => x"4c220002", 14548 => x"3442e0c0", 14549 => x"59820000",
    14550 => x"34020001", 14551 => x"e0000008", 14552 => x"78010001",
    14553 => x"34420064", 14554 => x"38218bc8", 14555 => x"58220000",
    14556 => x"34010000", 14557 => x"f8000e94", 14558 => x"34020000",
    14559 => x"b8400800", 14560 => x"2b9d0004", 14561 => x"2b8b000c",
    14562 => x"2b8c0008", 14563 => x"379c000c", 14564 => x"c3a00000",
    14565 => x"379cfff8", 14566 => x"5b8b0008", 14567 => x"5b9d0004",
    14568 => x"78020001", 14569 => x"b8205800", 14570 => x"b8400800",
    14571 => x"382154b4", 14572 => x"fbfff893", 14573 => x"e0000003",
    14574 => x"34010064", 14575 => x"fbfffe55", 14576 => x"34010000",
    14577 => x"fbfff9e1", 14578 => x"4420fffc", 14579 => x"34010003",
    14580 => x"34020000", 14581 => x"34030001", 14582 => x"f8000da0",
    14583 => x"78020001", 14584 => x"b8400800", 14585 => x"382154cc",
    14586 => x"fbfff885", 14587 => x"e0000003", 14588 => x"34010064",
    14589 => x"fbfffe47", 14590 => x"34010000", 14591 => x"f8000e61",
    14592 => x"4420fffc", 14593 => x"78020001", 14594 => x"b8400800",
    14595 => x"38214adc", 14596 => x"fbfff87b", 14597 => x"78020001",
    14598 => x"b8400800", 14599 => x"382154dc", 14600 => x"fbfff877",
    14601 => x"fbffff34", 14602 => x"b9600800", 14603 => x"fbffff4a",
    14604 => x"4420fffe", 14605 => x"2b9d0004", 14606 => x"2b8b0008",
    14607 => x"379c0008", 14608 => x"c3a00000", 14609 => x"379cfff0",
    14610 => x"5b8b000c", 14611 => x"5b8c0008", 14612 => x"5b9d0004",
    14613 => x"b8405800", 14614 => x"34020003", 14615 => x"5c220020",
    14616 => x"fbffff25", 14617 => x"b9600800", 14618 => x"fbffff3b",
    14619 => x"4420fffe", 14620 => x"4c200002", 14621 => x"e000001a",
    14622 => x"37810010", 14623 => x"34020000", 14624 => x"f800036d",
    14625 => x"b8206000", 14626 => x"48010007", 14627 => x"29620000",
    14628 => x"2b810010", 14629 => x"3443ff38", 14630 => x"54610003",
    14631 => x"344200c8", 14632 => x"50410012", 14633 => x"34020001",
    14634 => x"b9600800", 14635 => x"f8000362", 14636 => x"78030001",
    14637 => x"b8206000", 14638 => x"29620000", 14639 => x"38635504",
    14640 => x"4c200003", 14641 => x"78030001", 14642 => x"386354fc",
    14643 => x"78010001", 14644 => x"3821550c", 14645 => x"fbfff84a",
    14646 => x"e0000004", 14647 => x"b9600800", 14648 => x"fbfffeee",
    14649 => x"b8206000", 14650 => x"29610000", 14651 => x"fbffef83",
    14652 => x"b9800800", 14653 => x"2b9d0004", 14654 => x"2b8b000c",
    14655 => x"2b8c0008", 14656 => x"379c0010", 14657 => x"c3a00000",
    14658 => x"379cfffc", 14659 => x"5b9d0004", 14660 => x"34010800",
    14661 => x"34020001", 14662 => x"fbfffaf2", 14663 => x"34010400",
    14664 => x"34020000", 14665 => x"fbfffaef", 14666 => x"34011000",
    14667 => x"34020000", 14668 => x"fbfffaec", 14669 => x"2b9d0004",
    14670 => x"379c0004", 14671 => x"c3a00000", 14672 => x"40230000",
    14673 => x"78020001", 14674 => x"40240001", 14675 => x"38428f98",
    14676 => x"28420000", 14677 => x"3c630008", 14678 => x"b8831800",
    14679 => x"58430010", 14680 => x"40240002", 14681 => x"40230003",
    14682 => x"3c840018", 14683 => x"3c630010", 14684 => x"b8832000",
    14685 => x"40230005", 14686 => x"b8832000", 14687 => x"40230004",
    14688 => x"3c630008", 14689 => x"b8830800", 14690 => x"58410014",
    14691 => x"c3a00000", 14692 => x"40230000", 14693 => x"40240003",
    14694 => x"78020001", 14695 => x"3c630018", 14696 => x"38428f98",
    14697 => x"b8831800", 14698 => x"40240001", 14699 => x"40210002",
    14700 => x"28420000", 14701 => x"3c840010", 14702 => x"3c210008",
    14703 => x"b8641800", 14704 => x"b8611800", 14705 => x"3401ff00",
    14706 => x"58430018", 14707 => x"a0611800", 14708 => x"34630001",
    14709 => x"58410020", 14710 => x"3801ea60", 14711 => x"5843001c",
    14712 => x"58410024", 14713 => x"78030001", 14714 => x"34210001",
    14715 => x"386357b0", 14716 => x"58410028", 14717 => x"34210001",
    14718 => x"5841002c", 14719 => x"28610000", 14720 => x"78030001",
    14721 => x"386357b4", 14722 => x"58410030", 14723 => x"38018cae",
    14724 => x"58410034", 14725 => x"28610000", 14726 => x"58410038",
    14727 => x"34011f40", 14728 => x"5841003c", 14729 => x"c3a00000",
    14730 => x"379cfff4", 14731 => x"5b8b000c", 14732 => x"5b8c0008",
    14733 => x"5b9d0004", 14734 => x"780b0001", 14735 => x"780c0001",
    14736 => x"396b7108", 14737 => x"398c7114", 14738 => x"e0000005",
    14739 => x"29620000", 14740 => x"b9600800", 14741 => x"356b000c",
    14742 => x"d8400000", 14743 => x"558bfffc", 14744 => x"2b9d0004",
    14745 => x"2b8b000c", 14746 => x"2b8c0008", 14747 => x"379c000c",
    14748 => x"c3a00000", 14749 => x"379cfff0", 14750 => x"5b8b0010",
    14751 => x"5b8c000c", 14752 => x"5b8d0008", 14753 => x"5b9d0004",
    14754 => x"780b0001", 14755 => x"780d0001", 14756 => x"340c0000",
    14757 => x"396b7108", 14758 => x"39ad7114", 14759 => x"e0000006",
    14760 => x"29620000", 14761 => x"b9600800", 14762 => x"356b000c",
    14763 => x"d8400000", 14764 => x"b5816000", 14765 => x"55abfffb",
    14766 => x"69810000", 14767 => x"2b9d0004", 14768 => x"2b8b0010",
    14769 => x"2b8c000c", 14770 => x"2b8d0008", 14771 => x"379c0010",
    14772 => x"c3a00000", 14773 => x"379cffec", 14774 => x"5b8b0014",
    14775 => x"5b8c0010", 14776 => x"5b8d000c", 14777 => x"5b8e0008",
    14778 => x"5b9d0004", 14779 => x"780b0001", 14780 => x"780d0001",
    14781 => x"b8207000", 14782 => x"396b7108", 14783 => x"39ad7114",
    14784 => x"e000000c", 14785 => x"296c0008", 14786 => x"e0000007",
    14787 => x"b9c01000", 14788 => x"f800124e", 14789 => x"5c200003",
    14790 => x"29810004", 14791 => x"e0000007", 14792 => x"358c0008",
    14793 => x"29810000", 14794 => x"5c20fff9", 14795 => x"356b000c",
    14796 => x"55abfff5", 14797 => x"78018000", 14798 => x"2b9d0004",
    14799 => x"2b8b0014", 14800 => x"2b8c0010", 14801 => x"2b8d000c",
    14802 => x"2b8e0008", 14803 => x"379c0014", 14804 => x"c3a00000",
    14805 => x"b8201800", 14806 => x"5c200008", 14807 => x"78010001",
    14808 => x"78020001", 14809 => x"38217108", 14810 => x"38427114",
    14811 => x"44220003", 14812 => x"28210008", 14813 => x"c3a00000",
    14814 => x"28620008", 14815 => x"34610008", 14816 => x"5c400016",
    14817 => x"78020001", 14818 => x"78040001", 14819 => x"38427108",
    14820 => x"38847114", 14821 => x"e000000f", 14822 => x"28410008",
    14823 => x"e000000a", 14824 => x"5c230008", 14825 => x"78030001",
    14826 => x"3442000c", 14827 => x"38637114", 14828 => x"34010000",
    14829 => x"50430009", 14830 => x"28410008", 14831 => x"c3a00000",
    14832 => x"34210008", 14833 => x"28250000", 14834 => x"5ca0fff6",
    14835 => x"3442000c", 14836 => x"5482fff2", 14837 => x"34010000",
    14838 => x"c3a00000", 14839 => x"379cffc8", 14840 => x"5b8b0038",
    14841 => x"5b8c0034", 14842 => x"5b8d0030", 14843 => x"5b8e002c",
    14844 => x"5b8f0028", 14845 => x"5b900024", 14846 => x"5b910020",
    14847 => x"5b92001c", 14848 => x"5b930018", 14849 => x"5b940014",
    14850 => x"5b950010", 14851 => x"5b96000c", 14852 => x"5b970008",
    14853 => x"5b9d0004", 14854 => x"b8207000", 14855 => x"34010000",
    14856 => x"b840b800", 14857 => x"78140001", 14858 => x"fbffffcb",
    14859 => x"78130001", 14860 => x"78120001", 14861 => x"78110001",
    14862 => x"78100001", 14863 => x"780f0001", 14864 => x"b8206800",
    14865 => x"34150000", 14866 => x"340b0000", 14867 => x"3a945740",
    14868 => x"3a734c00", 14869 => x"3a525538", 14870 => x"78168000",
    14871 => x"3a315314", 14872 => x"3a104458", 14873 => x"39ef530c",
    14874 => x"e0000028", 14875 => x"3562000f", 14876 => x"b5cb0800",
    14877 => x"4ae20006", 14878 => x"78020001", 14879 => x"38425530",
    14880 => x"fbfff751", 14881 => x"b5615800", 14882 => x"e0000021",
    14883 => x"29ac0004", 14884 => x"ba801800", 14885 => x"46a00002",
    14886 => x"ba601800", 14887 => x"29a40000", 14888 => x"ba401000",
    14889 => x"fbfff748", 14890 => x"b42b5800", 14891 => x"5d960005",
    14892 => x"b5cb0800", 14893 => x"b9e01000", 14894 => x"fbfff743",
    14895 => x"e000000e", 14896 => x"4d800006", 14897 => x"b5cb0800",
    14898 => x"ba001000", 14899 => x"fbfff73e", 14900 => x"c80c6000",
    14901 => x"b5615800", 14902 => x"2184ffff", 14903 => x"08842710",
    14904 => x"15830010", 14905 => x"b5cb0800", 14906 => x"00840010",
    14907 => x"ba201000", 14908 => x"fbfff735", 14909 => x"b42b5800",
    14910 => x"b9a00800", 14911 => x"fbffff96", 14912 => x"b8206800",
    14913 => x"36b50001", 14914 => x"5da0ffd9", 14915 => x"b9600800",
    14916 => x"2b9d0004", 14917 => x"2b8b0038", 14918 => x"2b8c0034",
    14919 => x"2b8d0030", 14920 => x"2b8e002c", 14921 => x"2b8f0028",
    14922 => x"2b900024", 14923 => x"2b910020", 14924 => x"2b92001c",
    14925 => x"2b930018", 14926 => x"2b940014", 14927 => x"2b950010",
    14928 => x"2b96000c", 14929 => x"2b970008", 14930 => x"379c0038",
    14931 => x"c3a00000", 14932 => x"379cffa8", 14933 => x"5b8b0008",
    14934 => x"5b9d0004", 14935 => x"378b000c", 14936 => x"b9600800",
    14937 => x"34020050", 14938 => x"fbffff9d", 14939 => x"78010001",
    14940 => x"b9601000", 14941 => x"3821461c", 14942 => x"fbfff721",
    14943 => x"34010000", 14944 => x"2b9d0004", 14945 => x"2b8b0008",
    14946 => x"379c0058", 14947 => x"c3a00000", 14948 => x"78010001",
    14949 => x"38218c38", 14950 => x"28210000", 14951 => x"28220008",
    14952 => x"2821000c", 14953 => x"202100ff", 14954 => x"c3a00000",
    14955 => x"78010001", 14956 => x"78030001", 14957 => x"386357b8",
    14958 => x"38218c38", 14959 => x"28210000", 14960 => x"28620000",
    14961 => x"78040001", 14962 => x"388457bc", 14963 => x"58220000",
    14964 => x"58200014", 14965 => x"28830000", 14966 => x"58200018",
    14967 => x"58200010", 14968 => x"58230000", 14969 => x"58220000",
    14970 => x"5820001c", 14971 => x"c3a00000", 14972 => x"78040001",
    14973 => x"34050002", 14974 => x"38848c38", 14975 => x"5c25000e",
    14976 => x"28810000", 14977 => x"1444001f", 14978 => x"20840007",
    14979 => x"b4831800", 14980 => x"f4832000", 14981 => x"00630003",
    14982 => x"b4821000", 14983 => x"3c42001d", 14984 => x"58200014",
    14985 => x"58200018", 14986 => x"b8431800", 14987 => x"58230010",
    14988 => x"e0000006", 14989 => x"28810000", 14990 => x"204200ff",
    14991 => x"58230014", 14992 => x"58220018", 14993 => x"58200010",
    14994 => x"78010001", 14995 => x"38218c38", 14996 => x"28210000",
    14997 => x"28220000", 14998 => x"38420004", 14999 => x"58220000",
    15000 => x"34010000", 15001 => x"c3a00000", 15002 => x"78050001",
    15003 => x"38a58c38", 15004 => x"28a50000", 15005 => x"202100ff",
    15006 => x"00630003", 15007 => x"58a20014", 15008 => x"58a10018",
    15009 => x"58a30010", 15010 => x"34010003", 15011 => x"5c810007",
    15012 => x"28a20000", 15013 => x"3401fff3", 15014 => x"a0410800",
    15015 => x"38210008", 15016 => x"58a10000", 15017 => x"c3a00000",
    15018 => x"34010001", 15019 => x"5c810007", 15020 => x"28a2001c",
    15021 => x"3401ffe7", 15022 => x"a0410800", 15023 => x"38210008",
    15024 => x"58a1001c", 15025 => x"c3a00000", 15026 => x"34010002",
    15027 => x"5c810006", 15028 => x"28a2001c", 15029 => x"3401ffe7",
    15030 => x"a0410800", 15031 => x"38210010", 15032 => x"58a1001c",
    15033 => x"c3a00000", 15034 => x"379cffe0", 15035 => x"5b8b0020",
    15036 => x"5b8c001c", 15037 => x"5b8d0018", 15038 => x"5b8e0014",
    15039 => x"5b8f0010", 15040 => x"5b90000c", 15041 => x"5b910008",
    15042 => x"5b9d0004", 15043 => x"b8206000", 15044 => x"78010001",
    15045 => x"382157a4", 15046 => x"282f0000", 15047 => x"780b0001",
    15048 => x"b8406800", 15049 => x"396b8c38", 15050 => x"fbffff9a",
    15051 => x"b8208800", 15052 => x"29610000", 15053 => x"b8408000",
    15054 => x"282e0004", 15055 => x"a1cf7000", 15056 => x"fbffff94",
    15057 => x"5c31fff9", 15058 => x"5c50fff8", 15059 => x"45800003",
    15060 => x"59810000", 15061 => x"59820004", 15062 => x"45a00003",
    15063 => x"3dc10003", 15064 => x"59a10000", 15065 => x"2b9d0004",
    15066 => x"2b8b0020", 15067 => x"2b8c001c", 15068 => x"2b8d0018",
    15069 => x"2b8e0014", 15070 => x"2b8f0010", 15071 => x"2b90000c",
    15072 => x"2b910008", 15073 => x"379c0020", 15074 => x"c3a00000",
    15075 => x"78010001", 15076 => x"38218c38", 15077 => x"28210000",
    15078 => x"28210000", 15079 => x"20210004", 15080 => x"64210000",
    15081 => x"c3a00000", 15082 => x"78020001", 15083 => x"38428c38",
    15084 => x"28420000", 15085 => x"2843001c", 15086 => x"44200003",
    15087 => x"38630006", 15088 => x"e0000003", 15089 => x"3401fff9",
    15090 => x"a0611800", 15091 => x"5843001c", 15092 => x"34010000",
    15093 => x"c3a00000", 15094 => x"379cffe0", 15095 => x"5b8b001c",
    15096 => x"5b8c0018", 15097 => x"5b8d0014", 15098 => x"5b8e0010",
    15099 => x"5b8f000c", 15100 => x"5b900008", 15101 => x"5b9d0004",
    15102 => x"b8205800", 15103 => x"78010001", 15104 => x"38218bec",
    15105 => x"b8406000", 15106 => x"40220000", 15107 => x"b8607000",
    15108 => x"b8807800", 15109 => x"b8a06800", 15110 => x"3401ffff",
    15111 => x"4440002b", 15112 => x"3d8c0001", 15113 => x"b9600800",
    15114 => x"fbfff93c", 15115 => x"218200fe", 15116 => x"b9600800",
    15117 => x"fbfff981", 15118 => x"01c20008", 15119 => x"b9600800",
    15120 => x"204200ff", 15121 => x"fbfff97d", 15122 => x"21c200ff",
    15123 => x"b9600800", 15124 => x"fbfff97a", 15125 => x"b9600800",
    15126 => x"fbfff944", 15127 => x"39820001", 15128 => x"b9600800",
    15129 => x"204200ff", 15130 => x"fbfff974", 15131 => x"340c0000",
    15132 => x"35aeffff", 15133 => x"37900023", 15134 => x"e0000009",
    15135 => x"b9600800", 15136 => x"ba001000", 15137 => x"34030000",
    15138 => x"fbfff9a9", 15139 => x"43820023", 15140 => x"b5ec0800",
    15141 => x"358c0001", 15142 => x"30220000", 15143 => x"55ccfff8",
    15144 => x"b9600800", 15145 => x"ba001000", 15146 => x"34030001",
    15147 => x"fbfff9a0", 15148 => x"43810023", 15149 => x"b5ee7000",
    15150 => x"31c10000", 15151 => x"b9600800", 15152 => x"fbfff946",
    15153 => x"b9a00800", 15154 => x"2b9d0004", 15155 => x"2b8b001c",
    15156 => x"2b8c0018", 15157 => x"2b8d0014", 15158 => x"2b8e0010",
    15159 => x"2b8f000c", 15160 => x"2b900008", 15161 => x"379c0020",
    15162 => x"c3a00000", 15163 => x"379cffe0", 15164 => x"5b8b0020",
    15165 => x"5b8c001c", 15166 => x"5b8d0018", 15167 => x"5b8e0014",
    15168 => x"5b8f0010", 15169 => x"5b90000c", 15170 => x"5b910008",
    15171 => x"5b9d0004", 15172 => x"b8205800", 15173 => x"78010001",
    15174 => x"38218bec", 15175 => x"b8606800", 15176 => x"40230000",
    15177 => x"3c4f0001", 15178 => x"b8808000", 15179 => x"b8a07000",
    15180 => x"3401ffff", 15181 => x"21ef00ff", 15182 => x"340c0000",
    15183 => x"5c60001f", 15184 => x"e0000020", 15185 => x"b9600800",
    15186 => x"fbfff8f4", 15187 => x"b9e01000", 15188 => x"b9600800",
    15189 => x"fbfff939", 15190 => x"01a20008", 15191 => x"b9600800",
    15192 => x"204200ff", 15193 => x"fbfff935", 15194 => x"21a200ff",
    15195 => x"b9600800", 15196 => x"fbfff932", 15197 => x"b60c1000",
    15198 => x"40420000", 15199 => x"b9600800", 15200 => x"35ad0001",
    15201 => x"fbfff92d", 15202 => x"b9600800", 15203 => x"fbfff913",
    15204 => x"b9600800", 15205 => x"fbfff8e1", 15206 => x"b9600800",
    15207 => x"b9e01000", 15208 => x"fbfff926", 15209 => x"b8208800",
    15210 => x"b9600800", 15211 => x"fbfff90b", 15212 => x"5e20fff8",
    15213 => x"358c0001", 15214 => x"55ccffe3", 15215 => x"b9c00800",
    15216 => x"2b9d0004", 15217 => x"2b8b0020", 15218 => x"2b8c001c",
    15219 => x"2b8d0018", 15220 => x"2b8e0014", 15221 => x"2b8f0010",
    15222 => x"2b90000c", 15223 => x"2b910008", 15224 => x"379c0020",
    15225 => x"c3a00000", 15226 => x"379cffec", 15227 => x"5b8b0014",
    15228 => x"5b8c0010", 15229 => x"5b8d000c", 15230 => x"5b8e0008",
    15231 => x"5b9d0004", 15232 => x"780d0001", 15233 => x"780c0001",
    15234 => x"39ad8bf0", 15235 => x"398c8bf4", 15236 => x"780b0001",
    15237 => x"59a10000", 15238 => x"59820000", 15239 => x"34030001",
    15240 => x"396b8bec", 15241 => x"202100ff", 15242 => x"204200ff",
    15243 => x"31630000", 15244 => x"fbfff99d", 15245 => x"b8207000",
    15246 => x"5c200006", 15247 => x"41a10003", 15248 => x"41820003",
    15249 => x"fbfff998", 15250 => x"5c2e0002", 15251 => x"31600000",
    15252 => x"2b9d0004", 15253 => x"2b8b0014", 15254 => x"2b8c0010",
    15255 => x"2b8d000c", 15256 => x"2b8e0008", 15257 => x"379c0014",
    15258 => x"c3a00000", 15259 => x"379cfff8", 15260 => x"5b8b0008",
    15261 => x"5b9d0004", 15262 => x"78010001", 15263 => x"78020001",
    15264 => x"38218bf0", 15265 => x"38428bf4", 15266 => x"40420003",
    15267 => x"780b0001", 15268 => x"40210003", 15269 => x"396b6eb0",
    15270 => x"34031004", 15271 => x"b9602000", 15272 => x"34050001",
    15273 => x"31600000", 15274 => x"fbffff91", 15275 => x"34030001",
    15276 => x"3402ffff", 15277 => x"5c230002", 15278 => x"41620000",
    15279 => x"b8400800", 15280 => x"2b9d0004", 15281 => x"2b8b0008",
    15282 => x"379c0008", 15283 => x"c3a00000", 15284 => x"379cffc4",
    15285 => x"5b8b001c", 15286 => x"5b8c0018", 15287 => x"5b8d0014",
    15288 => x"5b8e0010", 15289 => x"5b8f000c", 15290 => x"5b900008",
    15291 => x"5b9d0004", 15292 => x"b8205800", 15293 => x"206d00ff",
    15294 => x"34010002", 15295 => x"204c00ff", 15296 => x"3405fffc",
    15297 => x"55a10087", 15298 => x"78040001", 15299 => x"38846eb0",
    15300 => x"40820000", 15301 => x"340100ff", 15302 => x"5c41000d",
    15303 => x"78010001", 15304 => x"78020001", 15305 => x"38218bf0",
    15306 => x"38428bf4", 15307 => x"40420003", 15308 => x"40210003",
    15309 => x"34050001", 15310 => x"34031004", 15311 => x"fbffff27",
    15312 => x"34020001", 15313 => x"3405ffff", 15314 => x"5c220076",
    15315 => x"78010001", 15316 => x"38216eb0", 15317 => x"40230000",
    15318 => x"340200ff", 15319 => x"5c620002", 15320 => x"30200000",
    15321 => x"5d800021", 15322 => x"78010001", 15323 => x"38216eb0",
    15324 => x"40210000", 15325 => x"34050000", 15326 => x"442c006a",
    15327 => x"78010001", 15328 => x"78020001", 15329 => x"38218bf0",
    15330 => x"38428bf4", 15331 => x"09a3001d", 15332 => x"40420003",
    15333 => x"40210003", 15334 => x"3405001d", 15335 => x"34631005",
    15336 => x"b9602000", 15337 => x"fbffff0d", 15338 => x"3402001d",
    15339 => x"b9606000", 15340 => x"3405ffff", 15341 => x"5c22005b",
    15342 => x"3562001c", 15343 => x"34010000", 15344 => x"e0000005",
    15345 => x"41830000", 15346 => x"358c0001", 15347 => x"b4230800",
    15348 => x"202100ff", 15349 => x"5d82fffc", 15350 => x"4162001c",
    15351 => x"3405fffd", 15352 => x"5c410050", 15353 => x"e000004a",
    15354 => x"34010001", 15355 => x"5d810048", 15356 => x"780f0001",
    15357 => x"780e0001", 15358 => x"780d0001", 15359 => x"340c0000",
    15360 => x"39ef6eb0", 15361 => x"39ce8bf0", 15362 => x"39ad8bf4",
    15363 => x"37900020", 15364 => x"e0000015", 15365 => x"0983001d",
    15366 => x"41a20003", 15367 => x"41c10003", 15368 => x"34631005",
    15369 => x"ba002000", 15370 => x"3405001d", 15371 => x"fbfffeeb",
    15372 => x"3402001d", 15373 => x"5c22003a", 15374 => x"ba000800",
    15375 => x"b9601000", 15376 => x"34030010", 15377 => x"f8001084",
    15378 => x"5c200005", 15379 => x"78010001", 15380 => x"38215554",
    15381 => x"fbfff56a", 15382 => x"e0000005", 15383 => x"358c0001",
    15384 => x"218c00ff", 15385 => x"41e10000", 15386 => x"542cffeb",
    15387 => x"34010002", 15388 => x"3405fffe", 15389 => x"5581002b",
    15390 => x"3563001c", 15391 => x"b9600800", 15392 => x"34020000",
    15393 => x"e0000005", 15394 => x"40240000", 15395 => x"34210001",
    15396 => x"b4441000", 15397 => x"204200ff", 15398 => x"5c23fffc",
    15399 => x"780e0001", 15400 => x"780d0001", 15401 => x"3162001c",
    15402 => x"39ce8bf0", 15403 => x"39ad8bf4", 15404 => x"0983001d",
    15405 => x"41c10003", 15406 => x"41a20003", 15407 => x"b9602000",
    15408 => x"34631005", 15409 => x"3405001d", 15410 => x"780b0001",
    15411 => x"fbffff08", 15412 => x"396b6eb0", 15413 => x"41610000",
    15414 => x"542c000d", 15415 => x"78010001", 15416 => x"38215570",
    15417 => x"fbfff546", 15418 => x"41610000", 15419 => x"41a20003",
    15420 => x"34031004", 15421 => x"34210001", 15422 => x"31610000",
    15423 => x"41c10003", 15424 => x"b9602000", 15425 => x"34050001",
    15426 => x"fbfffef9", 15427 => x"78010001", 15428 => x"38216eb0",
    15429 => x"40250000", 15430 => x"e0000002", 15431 => x"3405ffff",
    15432 => x"b8a00800", 15433 => x"2b9d0004", 15434 => x"2b8b001c",
    15435 => x"2b8c0018", 15436 => x"2b8d0014", 15437 => x"2b8e0010",
    15438 => x"2b8f000c", 15439 => x"2b900008", 15440 => x"379c003c",
    15441 => x"c3a00000", 15442 => x"379cffcc", 15443 => x"5b8b0014",
    15444 => x"5b8c0010", 15445 => x"5b8d000c", 15446 => x"5b8e0008",
    15447 => x"5b9d0004", 15448 => x"340d0000", 15449 => x"b8205800",
    15450 => x"340c0001", 15451 => x"378e0018", 15452 => x"e0000027",
    15453 => x"b9c00800", 15454 => x"34020000", 15455 => x"b9a01800",
    15456 => x"fbffff54", 15457 => x"b8206000", 15458 => x"4c010023",
    15459 => x"b9c00800", 15460 => x"b9601000", 15461 => x"34030010",
    15462 => x"f800102f", 15463 => x"35ad0001", 15464 => x"5c20001b",
    15465 => x"2b81002c", 15466 => x"340c0001", 15467 => x"00220018",
    15468 => x"31610017", 15469 => x"31620014", 15470 => x"00220010",
    15471 => x"31620015", 15472 => x"00220008", 15473 => x"2b810030",
    15474 => x"31620016", 15475 => x"00220018", 15476 => x"3161001b",
    15477 => x"31620018", 15478 => x"00220010", 15479 => x"31620019",
    15480 => x"00220008", 15481 => x"2b810028", 15482 => x"3162001a",
    15483 => x"00220018", 15484 => x"31610013", 15485 => x"31620010",
    15486 => x"00220010", 15487 => x"31620011", 15488 => x"00220008",
    15489 => x"31620012", 15490 => x"e0000003", 15491 => x"498dffda",
    15492 => x"340c0000", 15493 => x"b9800800", 15494 => x"2b9d0004",
    15495 => x"2b8b0014", 15496 => x"2b8c0010", 15497 => x"2b8d000c",
    15498 => x"2b8e0008", 15499 => x"379c0034", 15500 => x"c3a00000",
    15501 => x"379cfff8", 15502 => x"5b8b0008", 15503 => x"5b9d0004",
    15504 => x"78030001", 15505 => x"b8205800", 15506 => x"204200ff",
    15507 => x"78010001", 15508 => x"38218bf0", 15509 => x"38638bf4",
    15510 => x"44400015", 15511 => x"29640000", 15512 => x"78028000",
    15513 => x"34050004", 15514 => x"b8821000", 15515 => x"59620000",
    15516 => x"40620003", 15517 => x"40210003", 15518 => x"34031000",
    15519 => x"b9602000", 15520 => x"fbfffe9b", 15521 => x"7c210004",
    15522 => x"78040001", 15523 => x"38845784", 15524 => x"c8011000",
    15525 => x"29630000", 15526 => x"28810000", 15527 => x"38420001",
    15528 => x"a0610800", 15529 => x"59610000", 15530 => x"e0000013",
    15531 => x"40620003", 15532 => x"40210003", 15533 => x"34031000",
    15534 => x"b9602000", 15535 => x"34050004", 15536 => x"fbfffe46",
    15537 => x"34030004", 15538 => x"3402ffff", 15539 => x"5c23000a",
    15540 => x"29610000", 15541 => x"34020000", 15542 => x"4c200007",
    15543 => x"78030001", 15544 => x"38635784", 15545 => x"28620000",
    15546 => x"a0220800", 15547 => x"59610000", 15548 => x"34020001",
    15549 => x"b8400800", 15550 => x"2b9d0004", 15551 => x"2b8b0008",
    15552 => x"379c0008", 15553 => x"c3a00000", 15554 => x"379cfff8",
    15555 => x"5b9d0004", 15556 => x"78010001", 15557 => x"78020001",
    15558 => x"38218bf0", 15559 => x"38428bf4", 15560 => x"40420003",
    15561 => x"40210003", 15562 => x"34031074", 15563 => x"3784000a",
    15564 => x"34050002", 15565 => x"0f80000a", 15566 => x"fbfffe6d",
    15567 => x"34030002", 15568 => x"3402ffff", 15569 => x"5c230002",
    15570 => x"2f82000a", 15571 => x"b8400800", 15572 => x"2b9d0004",
    15573 => x"379c0008", 15574 => x"c3a00000", 15575 => x"379cffcc",
    15576 => x"5b8b002c", 15577 => x"5b8c0028", 15578 => x"5b8d0024",
    15579 => x"5b8e0020", 15580 => x"5b8f001c", 15581 => x"5b900018",
    15582 => x"5b910014", 15583 => x"5b920010", 15584 => x"5b93000c",
    15585 => x"5b940008", 15586 => x"5b9d0004", 15587 => x"78030001",
    15588 => x"78020001", 15589 => x"38638bf0", 15590 => x"b8208800",
    15591 => x"38428bf4", 15592 => x"34010020", 15593 => x"33810037",
    15594 => x"40420003", 15595 => x"40610003", 15596 => x"37840034",
    15597 => x"34031074", 15598 => x"34050002", 15599 => x"fbfffe07",
    15600 => x"34020002", 15601 => x"340bffff", 15602 => x"5c220051",
    15603 => x"2f820034", 15604 => x"3801ffff", 15605 => x"5c410002",
    15606 => x"0f800034", 15607 => x"780d0001", 15608 => x"780c0001",
    15609 => x"340b0001", 15610 => x"39ad8bf0", 15611 => x"398c8bf4",
    15612 => x"37900037", 15613 => x"e0000023", 15614 => x"41b40003",
    15615 => x"41930003", 15616 => x"b9c00800", 15617 => x"34721076",
    15618 => x"f8000f64", 15619 => x"b8202800", 15620 => x"b9c02000",
    15621 => x"ba800800", 15622 => x"ba601000", 15623 => x"ba401800",
    15624 => x"fbfffe33", 15625 => x"b8207000", 15626 => x"29e10000",
    15627 => x"f8000f5b", 15628 => x"5dc10036", 15629 => x"29e10000",
    15630 => x"2f8e0034", 15631 => x"f8000f57", 15632 => x"b5c11800",
    15633 => x"41820003", 15634 => x"41a10003", 15635 => x"2063ffff",
    15636 => x"0f830034", 15637 => x"ba002000", 15638 => x"34631076",
    15639 => x"34050001", 15640 => x"fbfffe23", 15641 => x"34020001",
    15642 => x"5c220028", 15643 => x"2f810034", 15644 => x"356b0001",
    15645 => x"216b00ff", 15646 => x"34210001", 15647 => x"0f810034",
    15648 => x"3d6f0002", 15649 => x"2f830034", 15650 => x"b62f7800",
    15651 => x"29ee0000", 15652 => x"5dc0ffda", 15653 => x"3401000a",
    15654 => x"33810037", 15655 => x"41820003", 15656 => x"41a10003",
    15657 => x"34631075", 15658 => x"37840037", 15659 => x"34050001",
    15660 => x"fbfffe0f", 15661 => x"34020001", 15662 => x"340bffff",
    15663 => x"5c220014", 15664 => x"41a10003", 15665 => x"41820003",
    15666 => x"34031074", 15667 => x"37840034", 15668 => x"34050002",
    15669 => x"fbfffe06", 15670 => x"b8207000", 15671 => x"34010002",
    15672 => x"5dc1000b", 15673 => x"41a10003", 15674 => x"41820003",
    15675 => x"34031074", 15676 => x"37840032", 15677 => x"34050002",
    15678 => x"fbfffdb8", 15679 => x"e42e5800", 15680 => x"356bffff",
    15681 => x"e0000002", 15682 => x"340bffff", 15683 => x"b9600800",
    15684 => x"2b9d0004", 15685 => x"2b8b002c", 15686 => x"2b8c0028",
    15687 => x"2b8d0024", 15688 => x"2b8e0020", 15689 => x"2b8f001c",
    15690 => x"2b900018", 15691 => x"2b910014", 15692 => x"2b920010",
    15693 => x"2b93000c", 15694 => x"2b940008", 15695 => x"379c0034",
    15696 => x"c3a00000", 15697 => x"379cffe4", 15698 => x"5b8b0018",
    15699 => x"5b8c0014", 15700 => x"5b8d0010", 15701 => x"5b8e000c",
    15702 => x"5b8f0008", 15703 => x"5b9d0004", 15704 => x"78010001",
    15705 => x"78020001", 15706 => x"38218bf0", 15707 => x"38428bf4",
    15708 => x"40420003", 15709 => x"40210003", 15710 => x"34031074",
    15711 => x"3784001c", 15712 => x"34050002", 15713 => x"fbfffd95",
    15714 => x"34030002", 15715 => x"3402ffff", 15716 => x"5c230025",
    15717 => x"2f81001c", 15718 => x"3802fffd", 15719 => x"3421ffff",
    15720 => x"2021ffff", 15721 => x"50410005", 15722 => x"78010001",
    15723 => x"38214c84", 15724 => x"0f80001c", 15725 => x"fbfff412",
    15726 => x"780e0001", 15727 => x"780d0001", 15728 => x"780c0001",
    15729 => x"340b0000", 15730 => x"39ce8bf0", 15731 => x"39ad8bf4",
    15732 => x"378f001f", 15733 => x"398c4c80", 15734 => x"e000000e",
    15735 => x"41a20003", 15736 => x"41c10003", 15737 => x"35631076",
    15738 => x"b9e02000", 15739 => x"34050001", 15740 => x"fbfffd7a",
    15741 => x"34020001", 15742 => x"5c22000a", 15743 => x"4382001f",
    15744 => x"b9800800", 15745 => x"356b0001", 15746 => x"fbfff3fd",
    15747 => x"216bffff", 15748 => x"2f81001c", 15749 => x"542bfff2",
    15750 => x"34020000", 15751 => x"e0000002", 15752 => x"3402ffff",
    15753 => x"b8400800", 15754 => x"2b9d0004", 15755 => x"2b8b0018",
    15756 => x"2b8c0014", 15757 => x"2b8d0010", 15758 => x"2b8e000c",
    15759 => x"2b8f0008", 15760 => x"379c001c", 15761 => x"c3a00000",
    15762 => x"379cffdc", 15763 => x"5b8b0024", 15764 => x"5b8c0020",
    15765 => x"5b8d001c", 15766 => x"5b8e0018", 15767 => x"5b8f0014",
    15768 => x"5b900010", 15769 => x"5b91000c", 15770 => x"5b920008",
    15771 => x"5b9d0004", 15772 => x"206300ff", 15773 => x"b8208800",
    15774 => x"205200ff", 15775 => x"5c600012", 15776 => x"78040001",
    15777 => x"78030001", 15778 => x"38848bf0", 15779 => x"38638bf4",
    15780 => x"40620003", 15781 => x"40810003", 15782 => x"78040001",
    15783 => x"34031074", 15784 => x"38848bf8", 15785 => x"34050002",
    15786 => x"fbfffd4c", 15787 => x"34020002", 15788 => x"3403ffff",
    15789 => x"5c22002b", 15790 => x"78030001", 15791 => x"38638bfa",
    15792 => x"0c610000", 15793 => x"78040001", 15794 => x"38848bfa",
    15795 => x"78030001", 15796 => x"38638bf8", 15797 => x"2c820000",
    15798 => x"2c610000", 15799 => x"34030000", 15800 => x"3442fffe",
    15801 => x"5041001f", 15802 => x"780d0001", 15803 => x"780c0001",
    15804 => x"340b0000", 15805 => x"b8807000", 15806 => x"39ad8bf0",
    15807 => x"398c8bf4", 15808 => x"3410000a", 15809 => x"2dc30000",
    15810 => x"3461fffe", 15811 => x"54320012", 15812 => x"41820003",
    15813 => x"41a10003", 15814 => x"34640001", 15815 => x"b62b7800",
    15816 => x"0dc40000", 15817 => x"34631074", 15818 => x"b9e02000",
    15819 => x"34050001", 15820 => x"fbfffd2a", 15821 => x"34020001",
    15822 => x"5c220009", 15823 => x"41e10000", 15824 => x"356b0001",
    15825 => x"216b00ff", 15826 => x"5c30ffef", 15827 => x"b9601800",
    15828 => x"e0000004", 15829 => x"3403fffd", 15830 => x"e0000002",
    15831 => x"3403ffff", 15832 => x"b8600800", 15833 => x"2b9d0004",
    15834 => x"2b8b0024", 15835 => x"2b8c0020", 15836 => x"2b8d001c",
    15837 => x"2b8e0018", 15838 => x"2b8f0014", 15839 => x"2b900010",
    15840 => x"2b91000c", 15841 => x"2b920008", 15842 => x"379c0024",
    15843 => x"c3a00000", 15844 => x"379cfffc", 15845 => x"5b9d0004",
    15846 => x"78010001", 15847 => x"38215588", 15848 => x"fbfff397",
    15849 => x"3401ffff", 15850 => x"2b9d0004", 15851 => x"379c0004",
    15852 => x"c3a00000", 15853 => x"379cfff8", 15854 => x"5b8b0008",
    15855 => x"5b9d0004", 15856 => x"78010001", 15857 => x"b8405800",
    15858 => x"78020001", 15859 => x"38425b64", 15860 => x"382155ac",
    15861 => x"fbfff38a", 15862 => x"78020001", 15863 => x"78010001",
    15864 => x"38428ec0", 15865 => x"38218ed0", 15866 => x"34460090",
    15867 => x"34050022", 15868 => x"34040033", 15869 => x"28220004",
    15870 => x"204300ff", 15871 => x"7c670042", 15872 => x"7c630028",
    15873 => x"a0e31800", 15874 => x"5c60000b", 15875 => x"28230000",
    15876 => x"31650000", 15877 => x"31640001", 15878 => x"31630002",
    15879 => x"00430018", 15880 => x"31630003", 15881 => x"00430010",
    15882 => x"00420008", 15883 => x"31630004", 15884 => x"31620005",
    15885 => x"34210010", 15886 => x"5c26ffef", 15887 => x"34010000",
    15888 => x"2b9d0004", 15889 => x"2b8b0008", 15890 => x"379c0008",
    15891 => x"c3a00000", 15892 => x"379cffe8", 15893 => x"5b8b0018",
    15894 => x"5b8c0014", 15895 => x"5b8d0010", 15896 => x"5b8e000c",
    15897 => x"5b8f0008", 15898 => x"5b9d0004", 15899 => x"780b0001",
    15900 => x"b8207800", 15901 => x"b8407000", 15902 => x"340d0008",
    15903 => x"340c0001", 15904 => x"396b6eb4", 15905 => x"a18e1800",
    15906 => x"29640008", 15907 => x"7c620000", 15908 => x"b9e00800",
    15909 => x"35adffff", 15910 => x"d8800000", 15911 => x"3d8c0001",
    15912 => x"5da0fff9", 15913 => x"2b9d0004", 15914 => x"2b8b0018",
    15915 => x"2b8c0014", 15916 => x"2b8d0010", 15917 => x"2b8e000c",
    15918 => x"2b8f0008", 15919 => x"379c0018", 15920 => x"c3a00000",
    15921 => x"379cffe8", 15922 => x"5b8b0018", 15923 => x"5b8c0014",
    15924 => x"5b8d0010", 15925 => x"5b8e000c", 15926 => x"5b8f0008",
    15927 => x"5b9d0004", 15928 => x"780b0001", 15929 => x"b8207800",
    15930 => x"340e0008", 15931 => x"340c0000", 15932 => x"340d0001",
    15933 => x"396b6eb4", 15934 => x"29620004", 15935 => x"b9e00800",
    15936 => x"35ceffff", 15937 => x"d8400000", 15938 => x"7c220000",
    15939 => x"c8021000", 15940 => x"a1a21000", 15941 => x"b9826000",
    15942 => x"3dad0001", 15943 => x"5dc0fff7", 15944 => x"34010064",
    15945 => x"fbffe9a1", 15946 => x"b9800800", 15947 => x"2b9d0004",
    15948 => x"2b8b0018", 15949 => x"2b8c0014", 15950 => x"2b8d0010",
    15951 => x"2b8e000c", 15952 => x"2b8f0008", 15953 => x"379c0018",
    15954 => x"c3a00000", 15955 => x"379cffc0", 15956 => x"5b8b0040",
    15957 => x"5b8c003c", 15958 => x"5b8d0038", 15959 => x"5b8e0034",
    15960 => x"5b8f0030", 15961 => x"5b90002c", 15962 => x"5b910028",
    15963 => x"5b920024", 15964 => x"5b930020", 15965 => x"5b94001c",
    15966 => x"5b950018", 15967 => x"5b960014", 15968 => x"5b970010",
    15969 => x"5b98000c", 15970 => x"5b990008", 15971 => x"5b9d0004",
    15972 => x"34020000", 15973 => x"b8206000", 15974 => x"34030080",
    15975 => x"34210008", 15976 => x"780d0001", 15977 => x"f8000d47",
    15978 => x"39ad6eb4", 15979 => x"29a10000", 15980 => x"340f0000",
    15981 => x"44200061", 15982 => x"b9805800", 15983 => x"34120000",
    15984 => x"34110000", 15985 => x"78194000", 15986 => x"34160001",
    15987 => x"34180008", 15988 => x"596c0008", 15989 => x"45e00022",
    15990 => x"29610000", 15991 => x"78028000", 15992 => x"34030000",
    15993 => x"59610010", 15994 => x"29610004", 15995 => x"59610014",
    15996 => x"a0590800", 15997 => x"44200003", 15998 => x"78024000",
    15999 => x"34030000", 16000 => x"a0710800", 16001 => x"a0522800",
    16002 => x"b8a12800", 16003 => x"29640010", 16004 => x"29610014",
    16005 => x"5ca0000e", 16006 => x"a4603000", 16007 => x"a0260800",
    16008 => x"59610014", 16009 => x"00630001", 16010 => x"3c41001f",
    16011 => x"a4403800", 16012 => x"00420001", 16013 => x"a0872000",
    16014 => x"b8231800", 16015 => x"59640010", 16016 => x"b8430800",
    16017 => x"5c25ffeb", 16018 => x"e000003c", 16019 => x"b8821000",
    16020 => x"b8231800", 16021 => x"59620010", 16022 => x"59630014",
    16023 => x"35ee0001", 16024 => x"29a20000", 16025 => x"3dce0004",
    16026 => x"b9800800", 16027 => x"b58e7000", 16028 => x"d8400000",
    16029 => x"5c360031", 16030 => x"b9800800", 16031 => x"340200f0",
    16032 => x"fbffff74", 16033 => x"34140040", 16034 => x"34130000",
    16035 => x"34100001", 16036 => x"34120000", 16037 => x"34110000",
    16038 => x"29a20004", 16039 => x"b9800800", 16040 => x"29d70004",
    16041 => x"d8400000", 16042 => x"29a20004", 16043 => x"b820a800",
    16044 => x"b9800800", 16045 => x"a2f0b800", 16046 => x"d8400000",
    16047 => x"46a10008", 16048 => x"29a30008", 16049 => x"baa01000",
    16050 => x"7eb50000", 16051 => x"b9800800", 16052 => x"d8600000",
    16053 => x"5eb60011", 16054 => x"e0000007", 16055 => x"29a30008",
    16056 => x"b9800800", 16057 => x"bae01000", 16058 => x"d8600000",
    16059 => x"46e00009", 16060 => x"e000000a", 16061 => x"29c10000",
    16062 => x"b8330800", 16063 => x"59c10000", 16064 => x"29c10004",
    16065 => x"b8300800", 16066 => x"59c10004", 16067 => x"e0000003",
    16068 => x"ba539000", 16069 => x"ba308800", 16070 => x"3e010001",
    16071 => x"3e730001", 16072 => x"f6018000", 16073 => x"3694ffff",
    16074 => x"b6139800", 16075 => x"b8208000", 16076 => x"5e80ffda",
    16077 => x"e0000014", 16078 => x"b9e00800", 16079 => x"2b9d0004",
    16080 => x"2b8b0040", 16081 => x"2b8c003c", 16082 => x"2b8d0038",
    16083 => x"2b8e0034", 16084 => x"2b8f0030", 16085 => x"2b90002c",
    16086 => x"2b910028", 16087 => x"2b920024", 16088 => x"2b930020",
    16089 => x"2b94001c", 16090 => x"2b950018", 16091 => x"2b960014",
    16092 => x"2b970010", 16093 => x"2b98000c", 16094 => x"2b990008",
    16095 => x"379c0040", 16096 => x"c3a00000", 16097 => x"35ef0001",
    16098 => x"356b0010", 16099 => x"5df8ff91", 16100 => x"e3ffffea",
    16101 => x"379cfff0", 16102 => x"5b8b0010", 16103 => x"5b8c000c",
    16104 => x"5b8d0008", 16105 => x"5b9d0004", 16106 => x"b8205800",
    16107 => x"78010001", 16108 => x"38216eb4", 16109 => x"28220000",
    16110 => x"29610000", 16111 => x"340c0000", 16112 => x"340d0040",
    16113 => x"d8400000", 16114 => x"29610000", 16115 => x"34020055",
    16116 => x"fbffff20", 16117 => x"29610008", 16118 => x"2962000c",
    16119 => x"b9801800", 16120 => x"358c0008", 16121 => x"f8000b7c",
    16122 => x"29610000", 16123 => x"fbffff19", 16124 => x"5d8dfff9",
    16125 => x"2b9d0004", 16126 => x"2b8b0010", 16127 => x"2b8c000c",
    16128 => x"2b8d0008", 16129 => x"379c0010", 16130 => x"c3a00000",
    16131 => x"28210000", 16132 => x"78020001", 16133 => x"38428f48",
    16134 => x"28420000", 16135 => x"3c210008", 16136 => x"3821000a",
    16137 => x"58410000", 16138 => x"28410000", 16139 => x"20230008",
    16140 => x"5c60fffe", 16141 => x"20210001", 16142 => x"18210001",
    16143 => x"c3a00000", 16144 => x"28210000", 16145 => x"78020001",
    16146 => x"38428f48", 16147 => x"28420000", 16148 => x"3c210008",
    16149 => x"38210009", 16150 => x"58410000", 16151 => x"28410000",
    16152 => x"20230008", 16153 => x"5c60fffe", 16154 => x"20210001",
    16155 => x"c3a00000", 16156 => x"28210000", 16157 => x"78030001",
    16158 => x"38638f48", 16159 => x"3c210008", 16160 => x"28630000",
    16161 => x"7c420000", 16162 => x"38210008", 16163 => x"b8221000",
    16164 => x"58620000", 16165 => x"28610000", 16166 => x"20210008",
    16167 => x"5c20fffe", 16168 => x"c3a00000", 16169 => x"78010001",
    16170 => x"78030001", 16171 => x"38218f48", 16172 => x"386357c0",
    16173 => x"28210000", 16174 => x"28620000", 16175 => x"58220004",
    16176 => x"c3a00000", 16177 => x"379cffc4", 16178 => x"5b8b001c",
    16179 => x"5b8c0018", 16180 => x"5b8d0014", 16181 => x"5b8e0010",
    16182 => x"5b8f000c", 16183 => x"5b900008", 16184 => x"5b9d0004",
    16185 => x"b8206000", 16186 => x"28210000", 16187 => x"340bffff",
    16188 => x"4420002a", 16189 => x"29820004", 16190 => x"44400028",
    16191 => x"fbffe85f", 16192 => x"780e0001", 16193 => x"b8206800",
    16194 => x"340b0000", 16195 => x"3410001f", 16196 => x"378f0020",
    16197 => x"39ce55c8", 16198 => x"e000000b", 16199 => x"fbffe857",
    16200 => x"202400ff", 16201 => x"b56d1000", 16202 => x"b5eb0800",
    16203 => x"30240000", 16204 => x"b8401800", 16205 => x"b9c00800",
    16206 => x"b8802800", 16207 => x"fbfff230", 16208 => x"356b0001",
    16209 => x"29810004", 16210 => x"ee0b1800", 16211 => x"358c0004",
    16212 => x"7c220000", 16213 => x"a0621000", 16214 => x"5c40fff1",
    16215 => x"78010001", 16216 => x"b9602000", 16217 => x"b9a01000",
    16218 => x"b9e01800", 16219 => x"38218ec0", 16220 => x"f80001cc",
    16221 => x"b8206000", 16222 => x"b9601800", 16223 => x"78010001",
    16224 => x"fd8b5800", 16225 => x"382155ec", 16226 => x"b9a01000",
    16227 => x"b9802000", 16228 => x"fbfff21b", 16229 => x"c80b5800",
    16230 => x"b9600800", 16231 => x"2b9d0004", 16232 => x"2b8b001c",
    16233 => x"2b8c0018", 16234 => x"2b8d0014", 16235 => x"2b8e0010",
    16236 => x"2b8f000c", 16237 => x"2b900008", 16238 => x"379c003c",
    16239 => x"c3a00000", 16240 => x"379cffc8", 16241 => x"5b8b0018",
    16242 => x"5b8c0014", 16243 => x"5b8d0010", 16244 => x"5b8e000c",
    16245 => x"5b8f0008", 16246 => x"5b9d0004", 16247 => x"b8205800",
    16248 => x"28210000", 16249 => x"3405ffff", 16250 => x"4420002c",
    16251 => x"29620004", 16252 => x"4440002a", 16253 => x"fbffe821",
    16254 => x"b8207000", 16255 => x"29610004", 16256 => x"fbffe81e",
    16257 => x"b8205800", 16258 => x"34010020", 16259 => x"4c2b0002",
    16260 => x"340b0020", 16261 => x"378d001c", 16262 => x"78010001",
    16263 => x"b9602000", 16264 => x"b9c01000", 16265 => x"b9a01800",
    16266 => x"38218ec0", 16267 => x"f8000189", 16268 => x"b8206000",
    16269 => x"78010001", 16270 => x"b9601800", 16271 => x"3821560c",
    16272 => x"b9c01000", 16273 => x"b9802000", 16274 => x"fbfff1ed",
    16275 => x"e98b5800", 16276 => x"ec0c0800", 16277 => x"3405ffff",
    16278 => x"b9615800", 16279 => x"5d60000f", 16280 => x"b9a07800",
    16281 => x"780d0001", 16282 => x"39ad55c8", 16283 => x"b5eb0800",
    16284 => x"40240000", 16285 => x"b56e1000", 16286 => x"b9a00800",
    16287 => x"b8401800", 16288 => x"b8802800", 16289 => x"356b0001",
    16290 => x"fbfff1dd", 16291 => x"498bfff8", 16292 => x"fd8b2800",
    16293 => x"c8052800", 16294 => x"b8a00800", 16295 => x"2b9d0004",
    16296 => x"2b8b0018", 16297 => x"2b8c0014", 16298 => x"2b8d0010",
    16299 => x"2b8e000c", 16300 => x"2b8f0008", 16301 => x"379c0038",
    16302 => x"c3a00000", 16303 => x"379cffe4", 16304 => x"5b8b001c",
    16305 => x"5b8c0018", 16306 => x"5b8d0014", 16307 => x"5b8e0010",
    16308 => x"5b8f000c", 16309 => x"5b900008", 16310 => x"5b9d0004",
    16311 => x"780d0001", 16312 => x"39ad8ec0", 16313 => x"b9a00800",
    16314 => x"780b0001", 16315 => x"780f0001", 16316 => x"780e0001",
    16317 => x"fbfffe96", 16318 => x"396b8ed0", 16319 => x"340c0000",
    16320 => x"39ef562c", 16321 => x"39ce5644", 16322 => x"34100008",
    16323 => x"29630000", 16324 => x"29640004", 16325 => x"b8640800",
    16326 => x"44200010", 16327 => x"b9801000", 16328 => x"b9e00800",
    16329 => x"fbfff1b6", 16330 => x"3d810004", 16331 => x"34020000",
    16332 => x"34210008", 16333 => x"b5a10800", 16334 => x"f8000015",
    16335 => x"2023ffff", 16336 => x"08632710", 16337 => x"b8201000",
    16338 => x"14420010", 16339 => x"14630010", 16340 => x"b9c00800",
    16341 => x"fbfff1aa", 16342 => x"358c0001", 16343 => x"356b0010",
    16344 => x"5d90ffeb", 16345 => x"34010000", 16346 => x"2b9d0004",
    16347 => x"2b8b001c", 16348 => x"2b8c0018", 16349 => x"2b8d0014",
    16350 => x"2b8e0010", 16351 => x"2b8f000c", 16352 => x"2b900008",
    16353 => x"379c001c", 16354 => x"c3a00000", 16355 => x"379cffec",
    16356 => x"5b8b0014", 16357 => x"5b8c0010", 16358 => x"5b8d000c",
    16359 => x"5b8e0008", 16360 => x"5b9d0004", 16361 => x"402d000f",
    16362 => x"b8206000", 16363 => x"34010028", 16364 => x"b8407000",
    16365 => x"45a10005", 16366 => x"34010042", 16367 => x"45a10003",
    16368 => x"34010010", 16369 => x"5da10034", 16370 => x"21cb0002",
    16371 => x"5d60000f", 16372 => x"b9800800", 16373 => x"fbfffef0",
    16374 => x"29810000", 16375 => x"34020044", 16376 => x"21ce0001",
    16377 => x"fbfffe1b", 16378 => x"34010000", 16379 => x"5dcb002d",
    16380 => x"780b0001", 16381 => x"396b6eb4", 16382 => x"29620004",
    16383 => x"29810000", 16384 => x"d8400000", 16385 => x"4420fffd",
    16386 => x"b9800800", 16387 => x"fbfffee2", 16388 => x"29810000",
    16389 => x"780b0001", 16390 => x"340200be", 16391 => x"396b8bfc",
    16392 => x"fbfffe0c", 16393 => x"356e0008", 16394 => x"e0000005",
    16395 => x"29810000", 16396 => x"fbfffe25", 16397 => x"31610000",
    16398 => x"356b0001", 16399 => x"5d6efffc", 16400 => x"78020001",
    16401 => x"38428bfc", 16402 => x"40410001", 16403 => x"40430000",
    16404 => x"3c210008", 16405 => x"b8230800", 16406 => x"34030028",
    16407 => x"dc200800", 16408 => x"45a3000b", 16409 => x"34030042",
    16410 => x"45a30009", 16411 => x"34030010", 16412 => x"5da3000b",
    16413 => x"40420006", 16414 => x"3c21000f", 16415 => x"3c42000c",
    16416 => x"3421c000", 16417 => x"b8220800", 16418 => x"e0000006",
    16419 => x"3c21000c", 16420 => x"e0000004", 16421 => x"78018000",
    16422 => x"e0000002", 16423 => x"34010000", 16424 => x"2b9d0004",
    16425 => x"2b8b0014", 16426 => x"2b8c0010", 16427 => x"2b8d000c",
    16428 => x"2b8e0008", 16429 => x"379c0014", 16430 => x"c3a00000",
    16431 => x"379cfffc", 16432 => x"5b9d0004", 16433 => x"34030000",
    16434 => x"b8202000", 16435 => x"34090028", 16436 => x"34080042",
    16437 => x"34070010", 16438 => x"34060008", 16439 => x"40850017",
    16440 => x"44a90003", 16441 => x"44a80002", 16442 => x"5ca70006",
    16443 => x"3c630004", 16444 => x"34630008", 16445 => x"b4230800",
    16446 => x"fbffffa5", 16447 => x"e0000005", 16448 => x"34630001",
    16449 => x"34840010", 16450 => x"5c66fff5", 16451 => x"78018000",
    16452 => x"2b9d0004", 16453 => x"379c0004", 16454 => x"c3a00000",
    16455 => x"379cffe0", 16456 => x"5b8b0020", 16457 => x"5b8c001c",
    16458 => x"5b8d0018", 16459 => x"5b8e0014", 16460 => x"5b8f0010",
    16461 => x"5b90000c", 16462 => x"5b910008", 16463 => x"5b9d0004",
    16464 => x"b8205800", 16465 => x"b8408800", 16466 => x"b8608000",
    16467 => x"b8806000", 16468 => x"fbfffe91", 16469 => x"29610000",
    16470 => x"3402000f", 16471 => x"222e00ff", 16472 => x"fbfffdbc",
    16473 => x"29610000", 16474 => x"b9c01000", 16475 => x"2231ff00",
    16476 => x"fbfffdb8", 16477 => x"16310008", 16478 => x"29610000",
    16479 => x"ba201000", 16480 => x"340d0000", 16481 => x"fbfffdb3",
    16482 => x"e0000006", 16483 => x"b60d1000", 16484 => x"29610000",
    16485 => x"40420000", 16486 => x"35ad0001", 16487 => x"fbfffdad",
    16488 => x"498dfffb", 16489 => x"b9600800", 16490 => x"fbfffe7b",
    16491 => x"29610000", 16492 => x"340200aa", 16493 => x"fbfffda7",
    16494 => x"29610000", 16495 => x"fbfffdc2", 16496 => x"b8207800",
    16497 => x"5c2e0022", 16498 => x"29610000", 16499 => x"fbfffdbe",
    16500 => x"b8207000", 16501 => x"5c310020", 16502 => x"29610000",
    16503 => x"340d0000", 16504 => x"fbfffdb9", 16505 => x"b8208800",
    16506 => x"e0000007", 16507 => x"29610000", 16508 => x"fbfffdb5",
    16509 => x"b60d1000", 16510 => x"40420000", 16511 => x"5c220018",
    16512 => x"35ad0001", 16513 => x"498dfffa", 16514 => x"b9600800",
    16515 => x"fbfffe62", 16516 => x"29610000", 16517 => x"34020055",
    16518 => x"fbfffd8e", 16519 => x"29610000", 16520 => x"b9e01000",
    16521 => x"fbfffd8b", 16522 => x"29610000", 16523 => x"b9c01000",
    16524 => x"fbfffd88", 16525 => x"29610000", 16526 => x"ba201000",
    16527 => x"fbfffd85", 16528 => x"34012710", 16529 => x"fbffe759",
    16530 => x"e0000006", 16531 => x"340cffff", 16532 => x"e0000004",
    16533 => x"340cfffe", 16534 => x"e0000002", 16535 => x"340cfffd",
    16536 => x"b9800800", 16537 => x"2b9d0004", 16538 => x"2b8b0020",
    16539 => x"2b8c001c", 16540 => x"2b8d0018", 16541 => x"2b8e0014",
    16542 => x"2b8f0010", 16543 => x"2b90000c", 16544 => x"2b910008",
    16545 => x"379c0020", 16546 => x"c3a00000", 16547 => x"379cffe4",
    16548 => x"5b8b001c", 16549 => x"5b8c0018", 16550 => x"5b8d0014",
    16551 => x"5b8e0010", 16552 => x"5b8f000c", 16553 => x"5b900008",
    16554 => x"5b9d0004", 16555 => x"b8208000", 16556 => x"2041001f",
    16557 => x"b8405800", 16558 => x"b8607000", 16559 => x"b8806000",
    16560 => x"340d0000", 16561 => x"44200030", 16562 => x"3441ffff",
    16563 => x"b4240800", 16564 => x"1422001f", 16565 => x"b8807800",
    16566 => x"0042001b", 16567 => x"b4410800", 16568 => x"1562001f",
    16569 => x"14210005", 16570 => x"0042001b", 16571 => x"b44b1000",
    16572 => x"14420005", 16573 => x"4422000c", 16574 => x"78010001",
    16575 => x"382157c4", 16576 => x"28220000", 16577 => x"a1621000",
    16578 => x"4c400005", 16579 => x"3442ffff", 16580 => x"3401ffe0",
    16581 => x"b8411000", 16582 => x"34420001", 16583 => x"340f0020",
    16584 => x"c9e27800", 16585 => x"ba000800", 16586 => x"b9601000",
    16587 => x"b9c01800", 16588 => x"b9e02000", 16589 => x"fbffff7a",
    16590 => x"b8206800", 16591 => x"48010016", 16592 => x"b5cf7000",
    16593 => x"b56f5800", 16594 => x"c98f6000", 16595 => x"e000000e",
    16596 => x"b9802000", 16597 => x"4dec0002", 16598 => x"34040020",
    16599 => x"ba000800", 16600 => x"b9601000", 16601 => x"b9c01800",
    16602 => x"fbffff6d", 16603 => x"48010009", 16604 => x"b5a16800",
    16605 => x"35ce0020", 16606 => x"356b0020", 16607 => x"358cffe0",
    16608 => x"e0000002", 16609 => x"340f0020", 16610 => x"4980fff2",
    16611 => x"e0000002", 16612 => x"b8206800", 16613 => x"b9a00800",
    16614 => x"2b9d0004", 16615 => x"2b8b001c", 16616 => x"2b8c0018",
    16617 => x"2b8d0014", 16618 => x"2b8e0010", 16619 => x"2b8f000c",
    16620 => x"2b900008", 16621 => x"379c001c", 16622 => x"c3a00000",
    16623 => x"379cffec", 16624 => x"5b8b0014", 16625 => x"5b8c0010",
    16626 => x"5b8d000c", 16627 => x"5b8e0008", 16628 => x"5b9d0004",
    16629 => x"b8405800", 16630 => x"b8206000", 16631 => x"b8607000",
    16632 => x"b8806800", 16633 => x"fbfffdec", 16634 => x"29810000",
    16635 => x"340200f0", 16636 => x"fbfffd18", 16637 => x"29810000",
    16638 => x"216200ff", 16639 => x"fbfffd15", 16640 => x"2162ff00",
    16641 => x"29810000", 16642 => x"00420008", 16643 => x"340b0000",
    16644 => x"fbfffd10", 16645 => x"e0000006", 16646 => x"29810000",
    16647 => x"fbfffd2a", 16648 => x"b5cb1000", 16649 => x"30410000",
    16650 => x"356b0001", 16651 => x"49abfffb", 16652 => x"b9a00800",
    16653 => x"2b9d0004", 16654 => x"2b8b0014", 16655 => x"2b8c0010",
    16656 => x"2b8d000c", 16657 => x"2b8e0008", 16658 => x"379c0014",
    16659 => x"c3a00000", 16660 => x"379cfffc", 16661 => x"5b9d0004",
    16662 => x"34050000", 16663 => x"b8203000", 16664 => x"34080043",
    16665 => x"34070008", 16666 => x"40c90017", 16667 => x"5d280006",
    16668 => x"3ca50004", 16669 => x"34a50008", 16670 => x"b4250800",
    16671 => x"fbffffd0", 16672 => x"e0000005", 16673 => x"34a50001",
    16674 => x"34c60010", 16675 => x"5ca7fff7", 16676 => x"3401ffff",
    16677 => x"2b9d0004", 16678 => x"379c0004", 16679 => x"c3a00000",
    16680 => x"379cfffc", 16681 => x"5b9d0004", 16682 => x"34050000",
    16683 => x"b8203000", 16684 => x"34080043", 16685 => x"34070008",
    16686 => x"40c90017", 16687 => x"5d280006", 16688 => x"3ca50004",
    16689 => x"34a50008", 16690 => x"b4250800", 16691 => x"fbffff70",
    16692 => x"e0000005", 16693 => x"34a50001", 16694 => x"34c60010",
    16695 => x"5ca7fff7", 16696 => x"3401ffff", 16697 => x"2b9d0004",
    16698 => x"379c0004", 16699 => x"c3a00000", 16700 => x"379cfff4",
    16701 => x"5b8b000c", 16702 => x"5b8c0008", 16703 => x"5b9d0004",
    16704 => x"780b0001", 16705 => x"396b8c0c", 16706 => x"29610000",
    16707 => x"5c200009", 16708 => x"fbfff5fb", 16709 => x"78020001",
    16710 => x"342103e8", 16711 => x"38428c04", 16712 => x"58410000",
    16713 => x"29610000", 16714 => x"34210001", 16715 => x"59610000",
    16716 => x"780b0001", 16717 => x"396b8c08", 16718 => x"296c0000",
    16719 => x"fbfff5f0", 16720 => x"78020001", 16721 => x"38428c04",
    16722 => x"28440000", 16723 => x"c8242800", 16724 => x"34010000",
    16725 => x"48050018", 16726 => x"21830001", 16727 => x"78010001",
    16728 => x"3c650002", 16729 => x"38215b78", 16730 => x"b4250800",
    16731 => x"28210000", 16732 => x"b4242000", 16733 => x"29610000",
    16734 => x"58440000", 16735 => x"34020001", 16736 => x"34210001",
    16737 => x"59610000", 16738 => x"78010001", 16739 => x"38218ec0",
    16740 => x"44620003", 16741 => x"fbfffeca", 16742 => x"e0000006",
    16743 => x"34020002", 16744 => x"fbfffec7", 16745 => x"78020001",
    16746 => x"38426ec0", 16747 => x"58410004", 16748 => x"34010001",
    16749 => x"2b9d0004", 16750 => x"2b8b000c", 16751 => x"2b8c0008",
    16752 => x"379c000c", 16753 => x"c3a00000", 16754 => x"78010001",
    16755 => x"38218f74", 16756 => x"28220000", 16757 => x"78010001",
    16758 => x"38218f9c", 16759 => x"58220000", 16760 => x"340103c6",
    16761 => x"58410004", 16762 => x"c3a00000", 16763 => x"c3a00000",
    16764 => x"379cfff8", 16765 => x"5b8b0008", 16766 => x"5b9d0004",
    16767 => x"b8205800", 16768 => x"3401000a", 16769 => x"5d610003",
    16770 => x"3401000d", 16771 => x"fbfffff9", 16772 => x"78020001",
    16773 => x"38428f9c", 16774 => x"28420000", 16775 => x"28410000",
    16776 => x"20210001", 16777 => x"5c20fffe", 16778 => x"584b0008",
    16779 => x"2b9d0004", 16780 => x"2b8b0008", 16781 => x"379c0008",
    16782 => x"c3a00000", 16783 => x"379cfff4", 16784 => x"5b8b000c",
    16785 => x"5b8c0008", 16786 => x"5b9d0004", 16787 => x"b8206000",
    16788 => x"b8205800", 16789 => x"e0000004", 16790 => x"b8400800",
    16791 => x"356b0001", 16792 => x"fbffffe4", 16793 => x"41620000",
    16794 => x"5c40fffc", 16795 => x"c96c0800", 16796 => x"2b9d0004",
    16797 => x"2b8b000c", 16798 => x"2b8c0008", 16799 => x"379c000c",
    16800 => x"c3a00000", 16801 => x"78010001", 16802 => x"38218f9c",
    16803 => x"28220000", 16804 => x"3401ffff", 16805 => x"28430000",
    16806 => x"20630002", 16807 => x"44600003", 16808 => x"2841000c",
    16809 => x"202100ff", 16810 => x"c3a00000", 16811 => x"28250008",
    16812 => x"28240000", 16813 => x"28260004", 16814 => x"b4451800",
    16815 => x"88642000", 16816 => x"5822001c", 16817 => x"88461000",
    16818 => x"b4821000", 16819 => x"2824000c", 16820 => x"1442000c",
    16821 => x"b4442000", 16822 => x"28220014", 16823 => x"4c820005",
    16824 => x"28240010", 16825 => x"44800008", 16826 => x"4ca3000b",
    16827 => x"e0000006", 16828 => x"28220018", 16829 => x"4c440006",
    16830 => x"28240010", 16831 => x"44800002", 16832 => x"4c650005",
    16833 => x"58230008", 16834 => x"e0000003", 16835 => x"58230008",
    16836 => x"b8801000", 16837 => x"58220020", 16838 => x"b8400800",
    16839 => x"c3a00000", 16840 => x"2822000c", 16841 => x"58200008",
    16842 => x"58220020", 16843 => x"c3a00000", 16844 => x"379cfff8",
    16845 => x"5b8b0008", 16846 => x"5b9d0004", 16847 => x"b8205800",
    16848 => x"58200014", 16849 => x"b8400800", 16850 => x"f800093b",
    16851 => x"2963000c", 16852 => x"29620000", 16853 => x"4823000b",
    16854 => x"29610004", 16855 => x"4c410003", 16856 => x"34420001",
    16857 => x"59620000", 16858 => x"29620000", 16859 => x"5c410011",
    16860 => x"34010001", 16861 => x"59610014", 16862 => x"59610010",
    16863 => x"e000000e", 16864 => x"29610008", 16865 => x"4c220003",
    16866 => x"3442ffff", 16867 => x"59620000", 16868 => x"29620000",
    16869 => x"5c410007", 16870 => x"34010001", 16871 => x"59610014",
    16872 => x"59600000", 16873 => x"59600010", 16874 => x"3401ffff",
    16875 => x"e0000002", 16876 => x"29610010", 16877 => x"2b9d0004",
    16878 => x"2b8b0008", 16879 => x"379c0008", 16880 => x"c3a00000",
    16881 => x"58200010", 16882 => x"58200000", 16883 => x"58200014",
    16884 => x"c3a00000", 16885 => x"78030001", 16886 => x"38638f80",
    16887 => x"28640000", 16888 => x"48810013", 16889 => x"78030001",
    16890 => x"38638c20", 16891 => x"c8240800", 16892 => x"44400007",
    16893 => x"28620000", 16894 => x"34040001", 16895 => x"bc810800",
    16896 => x"28430028", 16897 => x"b8230800", 16898 => x"e0000007",
    16899 => x"28620000", 16900 => x"34040001", 16901 => x"bc810800",
    16902 => x"28430028", 16903 => x"a4200800", 16904 => x"a0230800",
    16905 => x"58410028", 16906 => x"c3a00000", 16907 => x"78030001",
    16908 => x"38638c20", 16909 => x"44400007", 16910 => x"28620000",
    16911 => x"34040001", 16912 => x"bc810800", 16913 => x"28430024",
    16914 => x"b8230800", 16915 => x"e0000007", 16916 => x"28620000",
    16917 => x"34040001", 16918 => x"bc810800", 16919 => x"28430024",
    16920 => x"a4200800", 16921 => x"a0230800", 16922 => x"58410024",
    16923 => x"c3a00000", 16924 => x"379cfff0", 16925 => x"5b8b0010",
    16926 => x"5b8c000c", 16927 => x"5b8d0008", 16928 => x"5b9d0004",
    16929 => x"b8406800", 16930 => x"b8606000", 16931 => x"34020000",
    16932 => x"34030028", 16933 => x"b8205800", 16934 => x"f800098a",
    16935 => x"b9600800", 16936 => x"b9a01000", 16937 => x"34030014",
    16938 => x"f8000908", 16939 => x"596c0014", 16940 => x"2b9d0004",
    16941 => x"2b8b0010", 16942 => x"2b8c000c", 16943 => x"2b8d0008",
    16944 => x"379c0010", 16945 => x"c3a00000", 16946 => x"b8201800",
    16947 => x"e0000004", 16948 => x"28840000", 16949 => x"34630008",
    16950 => x"44820006", 16951 => x"28610004", 16952 => x"b8602000",
    16953 => x"5c20fffb", 16954 => x"78010001", 16955 => x"38215660",
    16956 => x"c3a00000", 16957 => x"78020001", 16958 => x"38428c20",
    16959 => x"28420000", 16960 => x"b8201800", 16961 => x"34010000",
    16962 => x"28440008", 16963 => x"20840002", 16964 => x"4480000c",
    16965 => x"34040002", 16966 => x"58440008", 16967 => x"78060001",
    16968 => x"28420010", 16969 => x"38c657c8", 16970 => x"28c40000",
    16971 => x"3445ff9b", 16972 => x"54a40004", 16973 => x"08420064",
    16974 => x"34010001", 16975 => x"58620000", 16976 => x"c3a00000",
    16977 => x"379cfff0", 16978 => x"5b8b0010", 16979 => x"5b8c000c",
    16980 => x"5b8d0008", 16981 => x"5b9d0004", 16982 => x"780b0001",
    16983 => x"b8206000", 16984 => x"78010001", 16985 => x"396b8f80",
    16986 => x"38218f78", 16987 => x"28210000", 16988 => x"296d0000",
    16989 => x"b42d6800", 16990 => x"29810000", 16991 => x"b9a01000",
    16992 => x"f8000114", 16993 => x"29810004", 16994 => x"29630000",
    16995 => x"b9a01000", 16996 => x"f8000199", 16997 => x"5980000c",
    16998 => x"59800008", 16999 => x"2b9d0004", 17000 => x"2b8b0010",
    17001 => x"2b8c000c", 17002 => x"2b8d0008", 17003 => x"379c0010",
    17004 => x"c3a00000", 17005 => x"379cfff8", 17006 => x"5b8b0008",
    17007 => x"5b9d0004", 17008 => x"b8205800", 17009 => x"28210000",
    17010 => x"f800016c", 17011 => x"78010001", 17012 => x"38218c20",
    17013 => x"28210000", 17014 => x"34020001", 17015 => x"34030009",
    17016 => x"58220004", 17017 => x"5963000c", 17018 => x"78030001",
    17019 => x"386357cc", 17020 => x"59620008", 17021 => x"28620000",
    17022 => x"5822004c", 17023 => x"2b9d0004", 17024 => x"2b8b0008",
    17025 => x"379c0008", 17026 => x"c3a00000", 17027 => x"b8201000",
    17028 => x"28210000", 17029 => x"2823004c", 17030 => x"34010000",
    17031 => x"44600016", 17032 => x"28430004", 17033 => x"28630038",
    17034 => x"44600013", 17035 => x"78030001", 17036 => x"38638c20",
    17037 => x"28630000", 17038 => x"28640004", 17039 => x"20840004",
    17040 => x"4480000d", 17041 => x"28630004", 17042 => x"20630008",
    17043 => x"5c60000a", 17044 => x"2842000c", 17045 => x"3403000a",
    17046 => x"34010001", 17047 => x"54430006", 17048 => x"78010001",
    17049 => x"3c420002", 17050 => x"38215ba8", 17051 => x"b4220800",
    17052 => x"28210000", 17053 => x"c3a00000", 17054 => x"379cfff0",
    17055 => x"5b8b000c", 17056 => x"5b8c0008", 17057 => x"5b9d0004",
    17058 => x"2822000c", 17059 => x"b8205800", 17060 => x"34010009",
    17061 => x"3442ffff", 17062 => x"340c0000", 17063 => x"544100a5",
    17064 => x"78010001", 17065 => x"3c420002", 17066 => x"38215b80",
    17067 => x"b4220800", 17068 => x"28210000", 17069 => x"c0200000",
    17070 => x"78010001", 17071 => x"38218c20", 17072 => x"28210000",
    17073 => x"340c0000", 17074 => x"28220004", 17075 => x"20420008",
    17076 => x"5c400098", 17077 => x"28230004", 17078 => x"78028000",
    17079 => x"b8621000", 17080 => x"58220004", 17081 => x"3401000a",
    17082 => x"e0000090", 17083 => x"78010001", 17084 => x"38218c20",
    17085 => x"28210000", 17086 => x"78040001", 17087 => x"38845784",
    17088 => x"28230004", 17089 => x"28820000", 17090 => x"a0621000",
    17091 => x"58220004", 17092 => x"28220004", 17093 => x"20420008",
    17094 => x"5c400083", 17095 => x"28210004", 17096 => x"340c0001",
    17097 => x"20210004", 17098 => x"44220082", 17099 => x"596c000c",
    17100 => x"e0000080", 17101 => x"29610000", 17102 => x"340c0000",
    17103 => x"2821004c", 17104 => x"4420007c", 17105 => x"fbffbda1",
    17106 => x"29610004", 17107 => x"f8000151", 17108 => x"fbffbda7",
    17109 => x"34010008", 17110 => x"e0000074", 17111 => x"78010001",
    17112 => x"38218c20", 17113 => x"28210000", 17114 => x"34020002",
    17115 => x"340c0000", 17116 => x"58220008", 17117 => x"29610000",
    17118 => x"2821004c", 17119 => x"4420006d", 17120 => x"29610004",
    17121 => x"28210038", 17122 => x"4420006a", 17123 => x"78010001",
    17124 => x"38218c34", 17125 => x"28210000", 17126 => x"340300a2",
    17127 => x"58230000", 17128 => x"34030003", 17129 => x"58230010",
    17130 => x"34030001", 17131 => x"5823001c", 17132 => x"5962000c",
    17133 => x"e000005e", 17134 => x"78010001", 17135 => x"38218c34",
    17136 => x"28210000", 17137 => x"340c0000", 17138 => x"2822001c",
    17139 => x"20420001", 17140 => x"44400058", 17141 => x"34020002",
    17142 => x"5822001c", 17143 => x"fbfff448", 17144 => x"342107d0",
    17145 => x"59610010", 17146 => x"34010003", 17147 => x"e000004f",
    17148 => x"fbfff443", 17149 => x"29620010", 17150 => x"340c0000",
    17151 => x"c8220800", 17152 => x"4801004c", 17153 => x"34010007",
    17154 => x"5961000c", 17155 => x"5960001c", 17156 => x"e0000047",
    17157 => x"37810010", 17158 => x"fbffff37", 17159 => x"340c0000",
    17160 => x"44200044", 17161 => x"78030001", 17162 => x"386357d0",
    17163 => x"28620000", 17164 => x"2b810010", 17165 => x"f80007a4",
    17166 => x"3802c34f", 17167 => x"e8221000", 17168 => x"64210000",
    17169 => x"b8410800", 17170 => x"44200005", 17171 => x"34010064",
    17172 => x"59610014", 17173 => x"3401ff9c", 17174 => x"e0000003",
    17175 => x"59600014", 17176 => x"34010064", 17177 => x"59610018",
    17178 => x"34010004", 17179 => x"e000002f", 17180 => x"29610004",
    17181 => x"340c0000", 17182 => x"f80001df", 17183 => x"5c20002d",
    17184 => x"37810010", 17185 => x"fbffff1c", 17186 => x"442c002a",
    17187 => x"78040001", 17188 => x"388457d0", 17189 => x"2b810010",
    17190 => x"28820000", 17191 => x"f800078a", 17192 => x"29620014",
    17193 => x"5b810010", 17194 => x"44220009", 17195 => x"2961001c",
    17196 => x"29620018", 17197 => x"b4410800", 17198 => x"5961001c",
    17199 => x"29610004", 17200 => x"2962001c", 17201 => x"f80001aa",
    17202 => x"e0000019", 17203 => x"29620014", 17204 => x"340c0001",
    17205 => x"5c220017", 17206 => x"2961001c", 17207 => x"34217530",
    17208 => x"5961001c", 17209 => x"29610004", 17210 => x"2962001c",
    17211 => x"f80001a0", 17212 => x"34010005", 17213 => x"5961000c",
    17214 => x"e000000e", 17215 => x"29610004", 17216 => x"340c0000",
    17217 => x"f80001bc", 17218 => x"5c20000a", 17219 => x"34010006",
    17220 => x"e0000006", 17221 => x"b9600800", 17222 => x"fbffff3d",
    17223 => x"340c0000", 17224 => x"5c200004", 17225 => x"34010009",
    17226 => x"5961000c", 17227 => x"340c0001", 17228 => x"b9800800",
    17229 => x"2b9d0004", 17230 => x"2b8b000c", 17231 => x"2b8c0008",
    17232 => x"379c0010", 17233 => x"c3a00000", 17234 => x"78040001",
    17235 => x"64630000", 17236 => x"38848c20", 17237 => x"28850000",
    17238 => x"c8031800", 17239 => x"78048000", 17240 => x"78060001",
    17241 => x"a0641800", 17242 => x"38c657d4", 17243 => x"b4641800",
    17244 => x"28c40000", 17245 => x"3c210018", 17246 => x"a0441000",
    17247 => x"b8410800", 17248 => x"b8231800", 17249 => x"58a3004c",
    17250 => x"c3a00000", 17251 => x"78040001", 17252 => x"64630000",
    17253 => x"38848c20", 17254 => x"28850000", 17255 => x"c8031800",
    17256 => x"78048000", 17257 => x"78060001", 17258 => x"a0641800",
    17259 => x"38c657d4", 17260 => x"b4641800", 17261 => x"28c40000",
    17262 => x"3c210018", 17263 => x"a0441000", 17264 => x"b8410800",
    17265 => x"b8231800", 17266 => x"58a3004c", 17267 => x"c3a00000",
    17268 => x"34030005", 17269 => x"5823002c", 17270 => x"3803fffb",
    17271 => x"58230030", 17272 => x"3403ff6a", 17273 => x"5823001c",
    17274 => x"3403fffe", 17275 => x"58230018", 17276 => x"34030001",
    17277 => x"58230028", 17278 => x"340300c8", 17279 => x"58230048",
    17280 => x"34032710", 17281 => x"58230040", 17282 => x"34030064",
    17283 => x"58230044", 17284 => x"5822000c", 17285 => x"58200014",
    17286 => x"c3a00000", 17287 => x"379cfff0", 17288 => x"5b8b0010",
    17289 => x"5b8c000c", 17290 => x"5b8d0008", 17291 => x"5b9d0004",
    17292 => x"b8205800", 17293 => x"2821000c", 17294 => x"b8406800",
    17295 => x"340c0000", 17296 => x"5c610047", 17297 => x"34010022",
    17298 => x"34030000", 17299 => x"fbffffbf", 17300 => x"29620004",
    17301 => x"34010025", 17302 => x"34030000", 17303 => x"fbffffbb",
    17304 => x"29610008", 17305 => x"4c200004", 17306 => x"596d0004",
    17307 => x"596d0008", 17308 => x"e000003b", 17309 => x"4da10005",
    17310 => x"29620000", 17311 => x"78010040", 17312 => x"b4410800",
    17313 => x"59610000", 17314 => x"29630000", 17315 => x"78050001",
    17316 => x"29620004", 17317 => x"38a557d8", 17318 => x"28a10000",
    17319 => x"b5a32000", 17320 => x"c8826000", 17321 => x"482c0006",
    17322 => x"78050001", 17323 => x"38a557dc", 17324 => x"28a10000",
    17325 => x"49810002", 17326 => x"e0000002", 17327 => x"b8206000",
    17328 => x"78050001", 17329 => x"38a557e0", 17330 => x"28a10000",
    17331 => x"4c240006", 17332 => x"4c220005", 17333 => x"c8611800",
    17334 => x"c8410800", 17335 => x"59630000", 17336 => x"59610004",
    17337 => x"29610004", 17338 => x"b9801000", 17339 => x"596d0008",
    17340 => x"34214000", 17341 => x"59610004", 17342 => x"35610018",
    17343 => x"fbfffdec", 17344 => x"78030001", 17345 => x"38638c20",
    17346 => x"29620010", 17347 => x"b8206800", 17348 => x"28610000",
    17349 => x"34030000", 17350 => x"582d0040", 17351 => x"34410001",
    17352 => x"59610010", 17353 => x"34010026", 17354 => x"fbffff88",
    17355 => x"34010020", 17356 => x"b9a01000", 17357 => x"34030000",
    17358 => x"fbffff84", 17359 => x"b9801000", 17360 => x"34010021",
    17361 => x"34030001", 17362 => x"fbffff80", 17363 => x"b9801000",
    17364 => x"3561003c", 17365 => x"fbfffdf7", 17366 => x"7c2c0000",
    17367 => x"b9800800", 17368 => x"2b9d0004", 17369 => x"2b8b0010",
    17370 => x"2b8c000c", 17371 => x"2b8d0008", 17372 => x"379c0010",
    17373 => x"c3a00000", 17374 => x"379cfff8", 17375 => x"5b8b0008",
    17376 => x"5b9d0004", 17377 => x"b8205800", 17378 => x"2821002c",
    17379 => x"59600004", 17380 => x"59600000", 17381 => x"59610024",
    17382 => x"3401ffff", 17383 => x"59610008", 17384 => x"59600010",
    17385 => x"35610018", 17386 => x"fbfffdde", 17387 => x"3561003c",
    17388 => x"fbfffe05", 17389 => x"78020001", 17390 => x"35610054",
    17391 => x"34030010", 17392 => x"38425bd4", 17393 => x"fbfffe2b",
    17394 => x"2961000c", 17395 => x"34020001", 17396 => x"fbfffe01",
    17397 => x"34010024", 17398 => x"34020001", 17399 => x"34030001",
    17400 => x"fbffff5a", 17401 => x"2b9d0004", 17402 => x"2b8b0008",
    17403 => x"379c0008", 17404 => x"c3a00000", 17405 => x"379cfff8",
    17406 => x"5b8b0008", 17407 => x"5b9d0004", 17408 => x"b8205800",
    17409 => x"34010005", 17410 => x"59610018", 17411 => x"3801fffa",
    17412 => x"5961001c", 17413 => x"34010001", 17414 => x"59610014",
    17415 => x"34017530", 17416 => x"59610010", 17417 => x"3401fbb4",
    17418 => x"59610008", 17419 => x"3401ffe2", 17420 => x"59610004",
    17421 => x"340104b0", 17422 => x"59610034", 17423 => x"340103e8",
    17424 => x"5961002c", 17425 => x"34010064", 17426 => x"59610030",
    17427 => x"78010001", 17428 => x"38218f80", 17429 => x"28210000",
    17430 => x"59630074", 17431 => x"59620070", 17432 => x"c8611800",
    17433 => x"59630080", 17434 => x"35610004", 17435 => x"5960007c",
    17436 => x"59600084", 17437 => x"fbfffdab", 17438 => x"35610028",
    17439 => x"fbfffdd2", 17440 => x"2b9d0004", 17441 => x"2b8b0008",
    17442 => x"379c0008", 17443 => x"c3a00000", 17444 => x"379cfff8",
    17445 => x"5b8b0008", 17446 => x"5b9d0004", 17447 => x"b8205800",
    17448 => x"58200044", 17449 => x"58200040", 17450 => x"3401ffff",
    17451 => x"59610048", 17452 => x"5961004c", 17453 => x"59610050",
    17454 => x"59610054", 17455 => x"34010001", 17456 => x"59610084",
    17457 => x"59600058", 17458 => x"35610004", 17459 => x"5960005c",
    17460 => x"59600060", 17461 => x"59600068", 17462 => x"5960006c",
    17463 => x"59600078", 17464 => x"fbfffd90", 17465 => x"35610028",
    17466 => x"fbfffdb7", 17467 => x"29610070", 17468 => x"34020001",
    17469 => x"fbfffdb8", 17470 => x"29610074", 17471 => x"34020001",
    17472 => x"fbfffdb5", 17473 => x"34010004", 17474 => x"34020001",
    17475 => x"34030001", 17476 => x"fbffff1f", 17477 => x"2b9d0004",
    17478 => x"2b8b0008", 17479 => x"379c0008", 17480 => x"c3a00000",
    17481 => x"379cfff8", 17482 => x"5b8b0008", 17483 => x"5b9d0004",
    17484 => x"b8205800", 17485 => x"28210074", 17486 => x"34020000",
    17487 => x"fbfffda6", 17488 => x"59600084", 17489 => x"2b9d0004",
    17490 => x"2b8b0008", 17491 => x"379c0008", 17492 => x"c3a00000",
    17493 => x"379cfff0", 17494 => x"5b8b0010", 17495 => x"5b8c000c",
    17496 => x"5b8d0008", 17497 => x"5b9d0004", 17498 => x"28240084",
    17499 => x"b8205800", 17500 => x"34010001", 17501 => x"44800078",
    17502 => x"29610070", 17503 => x"5c610002", 17504 => x"59620048",
    17505 => x"29610074", 17506 => x"5c610002", 17507 => x"5962004c",
    17508 => x"29610048", 17509 => x"48010009", 17510 => x"29620050",
    17511 => x"48020006", 17512 => x"4c220005", 17513 => x"29630040",
    17514 => x"78020040", 17515 => x"b4621000", 17516 => x"59620040",
    17517 => x"59610050", 17518 => x"2961004c", 17519 => x"48010009",
    17520 => x"29620054", 17521 => x"48020006", 17522 => x"4c220005",
    17523 => x"29630044", 17524 => x"78020040", 17525 => x"b4621000",
    17526 => x"59620044", 17527 => x"59610054", 17528 => x"29630048",
    17529 => x"34010000", 17530 => x"4803005b", 17531 => x"2962004c",
    17532 => x"48020059", 17533 => x"296c0040", 17534 => x"29610038",
    17535 => x"b46c1800", 17536 => x"296c0044", 17537 => x"c8621000",
    17538 => x"c84c6000", 17539 => x"44200006", 17540 => x"218c3fff",
    17541 => x"21812000", 17542 => x"44200003", 17543 => x"3401c000",
    17544 => x"b9816000", 17545 => x"b9801000", 17546 => x"35610004",
    17547 => x"fbfffd20", 17548 => x"29620080", 17549 => x"78030001",
    17550 => x"38638c20", 17551 => x"2042000f", 17552 => x"b8206800",
    17553 => x"3c420010", 17554 => x"28610000", 17555 => x"21a3ffff",
    17556 => x"b8621000", 17557 => x"58220044", 17558 => x"29630040",
    17559 => x"29620048", 17560 => x"34010005", 17561 => x"b4621000",
    17562 => x"34030000", 17563 => x"fbfffec8", 17564 => x"29630044",
    17565 => x"2962004c", 17566 => x"34010002", 17567 => x"b4621000",
    17568 => x"34030000", 17569 => x"fbfffec2", 17570 => x"34010001",
    17571 => x"b9801000", 17572 => x"34030000", 17573 => x"fbfffebe",
    17574 => x"29620078", 17575 => x"34030000", 17576 => x"34410001",
    17577 => x"59610078", 17578 => x"34010006", 17579 => x"fbfffeb8",
    17580 => x"34010000", 17581 => x"b9a01000", 17582 => x"34030001",
    17583 => x"fbfffeb4", 17584 => x"78020001", 17585 => x"3401ffff",
    17586 => x"384257e4", 17587 => x"5961004c", 17588 => x"59610048",
    17589 => x"29630040", 17590 => x"28410000", 17591 => x"4c23000a",
    17592 => x"29620044", 17593 => x"4c220008", 17594 => x"78040001",
    17595 => x"388457e8", 17596 => x"28810000", 17597 => x"b4611800",
    17598 => x"b4410800", 17599 => x"59630040", 17600 => x"59610044",
    17601 => x"29610038", 17602 => x"4420000f", 17603 => x"2961006c",
    17604 => x"29620068", 17605 => x"4c220006", 17606 => x"34210001",
    17607 => x"5961006c", 17608 => x"29610040", 17609 => x"3421ffff",
    17610 => x"e0000006", 17611 => x"4c410006", 17612 => x"3421ffff",
    17613 => x"5961006c", 17614 => x"29610040", 17615 => x"34210001",
    17616 => x"59610040", 17617 => x"35610028", 17618 => x"b9801000",
    17619 => x"fbfffcf9", 17620 => x"7c210000", 17621 => x"2b9d0004",
    17622 => x"2b8b0010", 17623 => x"2b8c000c", 17624 => x"2b8d0008",
    17625 => x"379c0010", 17626 => x"c3a00000", 17627 => x"379cfff0",
    17628 => x"5b8b0008", 17629 => x"5b9d0004", 17630 => x"b8205800",
    17631 => x"1443001f", 17632 => x"3781000c", 17633 => x"4802000b",
    17634 => x"00440012", 17635 => x"3c63000e", 17636 => x"3c42000e",
    17637 => x"b8641800", 17638 => x"5b820010", 17639 => x"34021f40",
    17640 => x"5b83000c", 17641 => x"fbffc191", 17642 => x"2b820010",
    17643 => x"e0000009", 17644 => x"0842c000", 17645 => x"5b820010",
    17646 => x"1442001f", 17647 => x"5b82000c", 17648 => x"34021f40",
    17649 => x"fbffc189", 17650 => x"2b820010", 17651 => x"c8021000",
    17652 => x"0041001f", 17653 => x"b4221000", 17654 => x"14420001",
    17655 => x"34010000", 17656 => x"59620068", 17657 => x"2b9d0004",
    17658 => x"2b8b0008", 17659 => x"379c0010", 17660 => x"c3a00000",
    17661 => x"28220068", 17662 => x"2821006c", 17663 => x"fc410800",
    17664 => x"c3a00000", 17665 => x"58220004", 17666 => x"5820001c",
    17667 => x"58230008", 17668 => x"5820000c", 17669 => x"58200010",
    17670 => x"58200000", 17671 => x"c3a00000", 17672 => x"379cfffc",
    17673 => x"5b9d0004", 17674 => x"34020001", 17675 => x"58220000",
    17676 => x"58200014", 17677 => x"5820001c", 17678 => x"5820000c",
    17679 => x"58200010", 17680 => x"28210004", 17681 => x"fbfffce4",
    17682 => x"78010001", 17683 => x"38218f80", 17684 => x"28210000",
    17685 => x"34020001", 17686 => x"fbfffcdf", 17687 => x"2b9d0004",
    17688 => x"379c0004", 17689 => x"c3a00000", 17690 => x"379cffb0",
    17691 => x"5b8b0010", 17692 => x"5b8c000c", 17693 => x"5b8d0008",
    17694 => x"5b9d0004", 17695 => x"b8205800", 17696 => x"b8406000",
    17697 => x"b8606800", 17698 => x"37810014", 17699 => x"34020000",
    17700 => x"34030040", 17701 => x"f800068b", 17702 => x"3401c000",
    17703 => x"78040001", 17704 => x"5b810020", 17705 => x"38848f80",
    17706 => x"34014000", 17707 => x"5b810044", 17708 => x"28810000",
    17709 => x"5da10005", 17710 => x"78030001", 17711 => x"38636fbc",
    17712 => x"586c0000", 17713 => x"e0000027", 17714 => x"3dad0005",
    17715 => x"b56d5800", 17716 => x"29610000", 17717 => x"44200023",
    17718 => x"78030001", 17719 => x"38636fbc", 17720 => x"28610000",
    17721 => x"29620010", 17722 => x"c9810800", 17723 => x"20213fff",
    17724 => x"1423000c", 17725 => x"5c400007", 17726 => x"3c630002",
    17727 => x"5961000c", 17728 => x"34010001", 17729 => x"59630014",
    17730 => x"59610010", 17731 => x"e0000015", 17732 => x"2964000c",
    17733 => x"34420001", 17734 => x"b4240800", 17735 => x"29640014",
    17736 => x"b4641800", 17737 => x"3c630002", 17738 => x"37840050",
    17739 => x"b4831800", 17740 => x"2863ffc4", 17741 => x"59620010",
    17742 => x"b4230800", 17743 => x"29630008", 17744 => x"5961000c",
    17745 => x"5c430007", 17746 => x"f8000532", 17747 => x"59610018",
    17748 => x"34010001", 17749 => x"5961001c", 17750 => x"5960000c",
    17751 => x"59600010", 17752 => x"34010000", 17753 => x"2b9d0004",
    17754 => x"2b8b0010", 17755 => x"2b8c000c", 17756 => x"2b8d0008",
    17757 => x"379c0050", 17758 => x"c3a00000", 17759 => x"78030001",
    17760 => x"38638c20", 17761 => x"5c40000a", 17762 => x"34040001",
    17763 => x"28620000", 17764 => x"bc810800", 17765 => x"202100ff",
    17766 => x"28430020", 17767 => x"3c210010", 17768 => x"a4200800",
    17769 => x"a0230800", 17770 => x"e0000008", 17771 => x"28620000",
    17772 => x"34040001", 17773 => x"bc810800", 17774 => x"28430020",
    17775 => x"202100ff", 17776 => x"3c210010", 17777 => x"b8230800",
    17778 => x"58410020", 17779 => x"c3a00000", 17780 => x"379cfff8",
    17781 => x"5b8b0008", 17782 => x"5b9d0004", 17783 => x"34020001",
    17784 => x"44220009", 17785 => x"34020002", 17786 => x"4422000c",
    17787 => x"5c200017", 17788 => x"78010001", 17789 => x"38218c20",
    17790 => x"282b0000", 17791 => x"356b0018", 17792 => x"e000000a",
    17793 => x"78010001", 17794 => x"38218c20", 17795 => x"282b0000",
    17796 => x"356b0014", 17797 => x"e0000005", 17798 => x"78010001",
    17799 => x"38218c20", 17800 => x"282b0000", 17801 => x"356b001c",
    17802 => x"340107d0", 17803 => x"fbfff1b9", 17804 => x"78030001",
    17805 => x"386357a4", 17806 => x"29620000", 17807 => x"28610000",
    17808 => x"a0410800", 17809 => x"e0000002", 17810 => x"34010000",
    17811 => x"2b9d0004", 17812 => x"2b8b0008", 17813 => x"379c0008",
    17814 => x"c3a00000", 17815 => x"379cfff8", 17816 => x"5b8b0008",
    17817 => x"5b9d0004", 17818 => x"b8201800", 17819 => x"78010001",
    17820 => x"b8405800", 17821 => x"38218cf4", 17822 => x"44600007",
    17823 => x"3461ffff", 17824 => x"08210090", 17825 => x"78030001",
    17826 => x"38638c3c", 17827 => x"34210148", 17828 => x"b4230800",
    17829 => x"b9601000", 17830 => x"fbffff35", 17831 => x"78010001",
    17832 => x"38218c3c", 17833 => x"582b0018", 17834 => x"2b9d0004",
    17835 => x"2b8b0008", 17836 => x"379c0008", 17837 => x"c3a00000",
    17838 => x"379cffec", 17839 => x"5b8b0014", 17840 => x"5b8c0010",
    17841 => x"5b8d000c", 17842 => x"5b8e0008", 17843 => x"5b9d0004",
    17844 => x"780c0001", 17845 => x"780d0001", 17846 => x"b8207000",
    17847 => x"340b0000", 17848 => x"398c8f80", 17849 => x"39ad8c10",
    17850 => x"e000000a", 17851 => x"29a10000", 17852 => x"942b0800",
    17853 => x"20210001", 17854 => x"44200005", 17855 => x"35620013",
    17856 => x"3c420005", 17857 => x"b5c20800", 17858 => x"fbffff46",
    17859 => x"356b0001", 17860 => x"29810000", 17861 => x"482bfff6",
    17862 => x"2b9d0004", 17863 => x"2b8b0014", 17864 => x"2b8c0010",
    17865 => x"2b8d000c", 17866 => x"2b8e0008", 17867 => x"379c0014",
    17868 => x"c3a00000", 17869 => x"379cffbc", 17870 => x"5b8b0044",
    17871 => x"5b8c0040", 17872 => x"5b8d003c", 17873 => x"5b8e0038",
    17874 => x"5b8f0034", 17875 => x"5b900030", 17876 => x"5b91002c",
    17877 => x"5b920028", 17878 => x"5b930024", 17879 => x"5b940020",
    17880 => x"5b95001c", 17881 => x"5b960018", 17882 => x"5b970014",
    17883 => x"5b980010", 17884 => x"5b99000c", 17885 => x"5b9b0008",
    17886 => x"5b9d0004", 17887 => x"781b0001", 17888 => x"780b0001",
    17889 => x"78190001", 17890 => x"780d0001", 17891 => x"78110001",
    17892 => x"78100001", 17893 => x"780c0001", 17894 => x"78170001",
    17895 => x"780f0001", 17896 => x"3b7b8c20", 17897 => x"396b8c3c",
    17898 => x"34140009", 17899 => x"3b395be8", 17900 => x"34180001",
    17901 => x"34130003", 17902 => x"39ad8cd4", 17903 => x"34120008",
    17904 => x"3a318cf4", 17905 => x"3a108c58", 17906 => x"398c8f80",
    17907 => x"3af78e9c", 17908 => x"39ef8f78", 17909 => x"e0000079",
    17910 => x"2875007c", 17911 => x"780100ff", 17912 => x"3821ffff",
    17913 => x"02ae0018", 17914 => x"a2a1a800", 17915 => x"29610004",
    17916 => x"21ce007f", 17917 => x"3421ffff", 17918 => x"54340050",
    17919 => x"3c210002", 17920 => x"b7210800", 17921 => x"28210000",
    17922 => x"c0200000", 17923 => x"2961004c", 17924 => x"58610040",
    17925 => x"296100d4", 17926 => x"296200d0", 17927 => x"b4410800",
    17928 => x"0022001f", 17929 => x"b4410800", 17930 => x"14210001",
    17931 => x"34020001", 17932 => x"58610044", 17933 => x"29810000",
    17934 => x"fbfffbe7", 17935 => x"fbfff130", 17936 => x"34210032",
    17937 => x"59610008", 17938 => x"3401000a", 17939 => x"e0000011",
    17940 => x"29760008", 17941 => x"fbfff12a", 17942 => x"cac10800",
    17943 => x"4c200037", 17944 => x"29610000", 17945 => x"5c380003",
    17946 => x"59780004", 17947 => x"e0000033", 17948 => x"59730004",
    17949 => x"e0000031", 17950 => x"29810000", 17951 => x"34020000",
    17952 => x"fbfffbd5", 17953 => x"b9a00800", 17954 => x"fbfffc4b",
    17955 => x"34010002", 17956 => x"59610004", 17957 => x"e0000029",
    17958 => x"b9a00800", 17959 => x"fbfffc5c", 17960 => x"e0000012",
    17961 => x"ba000800", 17962 => x"fbfffdb4", 17963 => x"34010004",
    17964 => x"e3fffff8", 17965 => x"29610068", 17966 => x"44200020",
    17967 => x"2961006c", 17968 => x"4420001e", 17969 => x"29610000",
    17970 => x"5c330009", 17971 => x"34010005", 17972 => x"e3fffff0",
    17973 => x"ba200800", 17974 => x"fbfffdee", 17975 => x"34010006",
    17976 => x"e3ffffec", 17977 => x"296100f0", 17978 => x"44200014",
    17979 => x"b9600800", 17980 => x"fbffff72", 17981 => x"59720004",
    17982 => x"e0000010", 17983 => x"29610000", 17984 => x"5c380004",
    17985 => x"b9a00800", 17986 => x"fbfffc41", 17987 => x"44200007",
    17988 => x"29610068", 17989 => x"44200005", 17990 => x"29610000",
    17991 => x"5c330007", 17992 => x"296100f0", 17993 => x"5c200005",
    17994 => x"29610010", 17995 => x"34210001", 17996 => x"59610010",
    17997 => x"59740004", 17998 => x"ba000800", 17999 => x"baa01000",
    18000 => x"b9c01800", 18001 => x"fbfffd36", 18002 => x"29610068",
    18003 => x"4420001b", 18004 => x"ba200800", 18005 => x"baa01000",
    18006 => x"b9c01800", 18007 => x"fbfffdfe", 18008 => x"29610004",
    18009 => x"5c320015", 18010 => x"29610000", 18011 => x"34160000",
    18012 => x"5c33000c", 18013 => x"e0000008", 18014 => x"0ac10090",
    18015 => x"baa01000", 18016 => x"b9c01800", 18017 => x"34210148",
    18018 => x"b5610800", 18019 => x"fbfffdf2", 18020 => x"36d60001",
    18021 => x"29e10000", 18022 => x"3421ffff", 18023 => x"4836fff7",
    18024 => x"29810000", 18025 => x"49c10005", 18026 => x"bae00800",
    18027 => x"baa01000", 18028 => x"b9c01800", 18029 => x"fbfffead",
    18030 => x"2b630000", 18031 => x"78020002", 18032 => x"28610080",
    18033 => x"a0220800", 18034 => x"4420ff84", 18035 => x"29610014",
    18036 => x"34210001", 18037 => x"59610014", 18038 => x"34010001",
    18039 => x"d0410000", 18040 => x"2b9d0004", 18041 => x"2b8b0044",
    18042 => x"2b8c0040", 18043 => x"2b8d003c", 18044 => x"2b8e0038",
    18045 => x"2b8f0034", 18046 => x"2b900030", 18047 => x"2b91002c",
    18048 => x"2b920028", 18049 => x"2b930024", 18050 => x"2b940020",
    18051 => x"2b95001c", 18052 => x"2b960018", 18053 => x"2b970014",
    18054 => x"2b980010", 18055 => x"2b99000c", 18056 => x"2b9b0008",
    18057 => x"379c0044", 18058 => x"c3a00000", 18059 => x"78010001",
    18060 => x"38218c38", 18061 => x"28220000", 18062 => x"78030001",
    18063 => x"78010001", 18064 => x"38218c34", 18065 => x"386357ec",
    18066 => x"58220000", 18067 => x"28610000", 18068 => x"58410000",
    18069 => x"c3a00000", 18070 => x"379cffd4", 18071 => x"5b8b0028",
    18072 => x"5b8c0024", 18073 => x"5b8d0020", 18074 => x"5b8e001c",
    18075 => x"5b8f0018", 18076 => x"5b900014", 18077 => x"5b910010",
    18078 => x"5b92000c", 18079 => x"5b930008", 18080 => x"5b9d0004",
    18081 => x"b8205800", 18082 => x"b8408000", 18083 => x"b8609000",
    18084 => x"fbffb9ce", 18085 => x"78010001", 18086 => x"38218fac",
    18087 => x"28240000", 18088 => x"78010001", 18089 => x"38218c20",
    18090 => x"58240000", 18091 => x"78010001", 18092 => x"28850000",
    18093 => x"38218c38", 18094 => x"28210000", 18095 => x"78020001",
    18096 => x"38428c34", 18097 => x"00a60010", 18098 => x"58410000",
    18099 => x"78020001", 18100 => x"38428f80", 18101 => x"20c6003f",
    18102 => x"00a50018", 18103 => x"58460000", 18104 => x"78020001",
    18105 => x"38428f78", 18106 => x"20a50007", 18107 => x"58450000",
    18108 => x"78050001", 18109 => x"38a58c3c", 18110 => x"58ab0000",
    18111 => x"58a00010", 18112 => x"58800040", 18113 => x"58800044",
    18114 => x"58800000", 18115 => x"58800028", 18116 => x"58800024",
    18117 => x"58800004", 18118 => x"78030001", 18119 => x"58800020",
    18120 => x"340203e8", 18121 => x"386357b8", 18122 => x"58820048",
    18123 => x"28620000", 18124 => x"5820001c", 18125 => x"58220000",
    18126 => x"34010004", 18127 => x"5d610004", 18128 => x"34010007",
    18129 => x"58a10004", 18130 => x"e0000006", 18131 => x"34010009",
    18132 => x"58a10004", 18133 => x"34010003", 18134 => x"5d610002",
    18135 => x"ba003000", 18136 => x"78010001", 18137 => x"b8c01000",
    18138 => x"38218c58", 18139 => x"780d0001", 18140 => x"fbfffc98",
    18141 => x"39ad8f80", 18142 => x"29a30000", 18143 => x"78010001",
    18144 => x"38218cf4", 18145 => x"ba001000", 18146 => x"780f0001",
    18147 => x"780e0001", 18148 => x"fbfffd19", 18149 => x"340c0000",
    18150 => x"39ef8f78", 18151 => x"39ce8c3c", 18152 => x"34130001",
    18153 => x"e000000c", 18154 => x"09910090", 18155 => x"29a40000",
    18156 => x"ba001000", 18157 => x"36210148", 18158 => x"34840001",
    18159 => x"b48c1800", 18160 => x"b5c10800", 18161 => x"b5d18800",
    18162 => x"fbfffd0b", 18163 => x"358c0001", 18164 => x"5a330140",
    18165 => x"29e10000", 18166 => x"3421ffff", 18167 => x"482cfff3",
    18168 => x"34010002", 18169 => x"5d610006", 18170 => x"78010001",
    18171 => x"38218c34", 18172 => x"28210000", 18173 => x"34020006",
    18174 => x"5822001c", 18175 => x"780e0001", 18176 => x"780d0001",
    18177 => x"340c0000", 18178 => x"39ce8f80", 18179 => x"39ad8c3c",
    18180 => x"e0000008", 18181 => x"35810013", 18182 => x"3c210005",
    18183 => x"b9801000", 18184 => x"b5a10800", 18185 => x"34030200",
    18186 => x"fbfffdf7", 18187 => x"358c0001", 18188 => x"29c20000",
    18189 => x"484cfff8", 18190 => x"34010001", 18191 => x"5d610017",
    18192 => x"78010001", 18193 => x"38218c20", 18194 => x"28210000",
    18195 => x"28210004", 18196 => x"20210002", 18197 => x"44200021",
    18198 => x"78010001", 18199 => x"78040001", 18200 => x"38218c3c",
    18201 => x"38848c58", 18202 => x"58240098", 18203 => x"78040001",
    18204 => x"38848cf4", 18205 => x"5824009c", 18206 => x"78010001",
    18207 => x"38218f78", 18208 => x"28240000", 18209 => x"78010001",
    18210 => x"38218cd4", 18211 => x"b4441000", 18212 => x"ba401800",
    18213 => x"fbfffb2c", 18214 => x"78010001", 18215 => x"38218c20",
    18216 => x"28210000", 18217 => x"78020002", 18218 => x"e0000003",
    18219 => x"2823007c", 18220 => x"5b83002c", 18221 => x"28230080",
    18222 => x"a0621800", 18223 => x"4460fffc", 18224 => x"34020001",
    18225 => x"58220064", 18226 => x"28220028", 18227 => x"38420001",
    18228 => x"58220028", 18229 => x"fbffb946", 18230 => x"2b9d0004",
    18231 => x"2b8b0028", 18232 => x"2b8c0024", 18233 => x"2b8d0020",
    18234 => x"2b8e001c", 18235 => x"2b8f0018", 18236 => x"2b900014",
    18237 => x"2b910010", 18238 => x"2b92000c", 18239 => x"2b930008",
    18240 => x"379c002c", 18241 => x"c3a00000", 18242 => x"379cfffc",
    18243 => x"5b9d0004", 18244 => x"78020001", 18245 => x"38428c3c",
    18246 => x"28430004", 18247 => x"64240000", 18248 => x"7c630008",
    18249 => x"b8831800", 18250 => x"5c600006", 18251 => x"3421ffff",
    18252 => x"08210090", 18253 => x"34210148", 18254 => x"b4410800",
    18255 => x"fbfffcd5", 18256 => x"2b9d0004", 18257 => x"379c0004",
    18258 => x"c3a00000", 18259 => x"379cfffc", 18260 => x"5b9d0004",
    18261 => x"44200008", 18262 => x"3421ffff", 18263 => x"08210090",
    18264 => x"78020001", 18265 => x"38428c3c", 18266 => x"34210148",
    18267 => x"b4220800", 18268 => x"fbfffced", 18269 => x"2b9d0004",
    18270 => x"379c0004", 18271 => x"c3a00000", 18272 => x"78020001",
    18273 => x"b8201800", 18274 => x"38428c3c", 18275 => x"5c200004",
    18276 => x"28410004", 18277 => x"64210008", 18278 => x"c3a00000",
    18279 => x"28450004", 18280 => x"34040008", 18281 => x"34010000",
    18282 => x"5ca40006", 18283 => x"3463ffff", 18284 => x"08630090",
    18285 => x"b4431000", 18286 => x"28410180", 18287 => x"7c210000",
    18288 => x"c3a00000", 18289 => x"379cffe8", 18290 => x"5b8b0018",
    18291 => x"5b8c0014", 18292 => x"5b8d0010", 18293 => x"5b8e000c",
    18294 => x"5b8f0008", 18295 => x"5b9d0004", 18296 => x"3403ffff",
    18297 => x"b8407800", 18298 => x"5c230016", 18299 => x"34010000",
    18300 => x"780c0001", 18301 => x"780d0001", 18302 => x"fbfffe19",
    18303 => x"340b0000", 18304 => x"398c8f78", 18305 => x"39ad8c3c",
    18306 => x"340e0004", 18307 => x"e0000009", 18308 => x"09610090",
    18309 => x"b5a10800", 18310 => x"28210140", 18311 => x"5c2e0004",
    18312 => x"35610001", 18313 => x"b9e01000", 18314 => x"fbfffe0d",
    18315 => x"356b0001", 18316 => x"29810000", 18317 => x"3421ffff",
    18318 => x"482bfff6", 18319 => x"e0000002", 18320 => x"fbfffe07",
    18321 => x"2b9d0004", 18322 => x"2b8b0018", 18323 => x"2b8c0014",
    18324 => x"2b8d0010", 18325 => x"2b8e000c", 18326 => x"2b8f0008",
    18327 => x"379c0018", 18328 => x"c3a00000", 18329 => x"379cfff0",
    18330 => x"5b8b0010", 18331 => x"5b8c000c", 18332 => x"5b8d0008",
    18333 => x"5b9d0004", 18334 => x"780b0001", 18335 => x"b8406800",
    18336 => x"b8606000", 18337 => x"396b8cf4", 18338 => x"44200007",
    18339 => x"342bffff", 18340 => x"096b0090", 18341 => x"78010001",
    18342 => x"38218c3c", 18343 => x"356b0148", 18344 => x"b5615800",
    18345 => x"45a0000b", 18346 => x"2962006c", 18347 => x"34041f40",
    18348 => x"34030000", 18349 => x"3c420001", 18350 => x"1441001f",
    18351 => x"f80002ae", 18352 => x"3c210012", 18353 => x"0044000e",
    18354 => x"b8242000", 18355 => x"59a40000", 18356 => x"4580000b",
    18357 => x"29620068", 18358 => x"34030000", 18359 => x"34041f40",
    18360 => x"3c420001", 18361 => x"1441001f", 18362 => x"f80002a3",
    18363 => x"3c210012", 18364 => x"0042000e", 18365 => x"b8221000",
    18366 => x"59820000", 18367 => x"2b9d0004", 18368 => x"2b8b0010",
    18369 => x"2b8c000c", 18370 => x"2b8d0008", 18371 => x"379c0010",
    18372 => x"c3a00000", 18373 => x"379cfff0", 18374 => x"5b8b0010",
    18375 => x"5b8c000c", 18376 => x"5b8d0008", 18377 => x"5b9d0004",
    18378 => x"b8205800", 18379 => x"b8406800", 18380 => x"78010001",
    18381 => x"3d620005", 18382 => x"38218c3c", 18383 => x"b4220800",
    18384 => x"28240278", 18385 => x"b8606000", 18386 => x"4c800003",
    18387 => x"34844000", 18388 => x"e0000004", 18389 => x"34013fff",
    18390 => x"4c240002", 18391 => x"3484c000", 18392 => x"3c840001",
    18393 => x"34010000", 18394 => x"20823ffe", 18395 => x"34030000",
    18396 => x"34041f40", 18397 => x"f8000280", 18398 => x"3c210012",
    18399 => x"0044000e", 18400 => x"b8242000", 18401 => x"59a40000",
    18402 => x"4580000d", 18403 => x"78010001", 18404 => x"38218c10",
    18405 => x"35630013", 18406 => x"28220000", 18407 => x"3c630005",
    18408 => x"78010001", 18409 => x"38218c3c", 18410 => x"b4230800",
    18411 => x"28210004", 18412 => x"94410800", 18413 => x"20210001",
    18414 => x"59810000", 18415 => x"3d6b0005", 18416 => x"78020001",
    18417 => x"38428c3c", 18418 => x"b44b1000", 18419 => x"2841027c",
    18420 => x"2b9d0004", 18421 => x"2b8b0010", 18422 => x"2b8c000c",
    18423 => x"2b8d0008", 18424 => x"379c0010", 18425 => x"c3a00000",
    18426 => x"379cffec", 18427 => x"5b8b0014", 18428 => x"5b8c0010",
    18429 => x"5b9d000c", 18430 => x"780b0001", 18431 => x"396b8c3c",
    18432 => x"29610000", 18433 => x"4c010014", 18434 => x"296c0014",
    18435 => x"29620004", 18436 => x"78010001", 18437 => x"38215c10",
    18438 => x"fbfffa2c", 18439 => x"29640000", 18440 => x"b8201800",
    18441 => x"296500a4", 18442 => x"29660068", 18443 => x"296700f0",
    18444 => x"29680054", 18445 => x"296200dc", 18446 => x"29610010",
    18447 => x"5b820004", 18448 => x"5b810008", 18449 => x"78010001",
    18450 => x"3821566c", 18451 => x"b9801000", 18452 => x"fbffe96b",
    18453 => x"2b9d000c", 18454 => x"2b8b0014", 18455 => x"2b8c0010",
    18456 => x"379c0014", 18457 => x"c3a00000", 18458 => x"379cfffc",
    18459 => x"5b9d0004", 18460 => x"5c200004", 18461 => x"78010001",
    18462 => x"38218cf4", 18463 => x"e0000007", 18464 => x"3421ffff",
    18465 => x"08210090", 18466 => x"78020001", 18467 => x"38428c3c",
    18468 => x"34210148", 18469 => x"b4220800", 18470 => x"fbfffcd7",
    18471 => x"2b9d0004", 18472 => x"379c0004", 18473 => x"c3a00000",
    18474 => x"379cfff0", 18475 => x"5b8b0010", 18476 => x"5b8c000c",
    18477 => x"5b8d0008", 18478 => x"5b9d0004", 18479 => x"780d0001",
    18480 => x"780b0001", 18481 => x"b8206000", 18482 => x"39ad8c3c",
    18483 => x"396b8c10", 18484 => x"4440000d", 18485 => x"34020001",
    18486 => x"fbfff9bf", 18487 => x"35810013", 18488 => x"3c210005",
    18489 => x"b5a10800", 18490 => x"fbfffcce", 18491 => x"29610000",
    18492 => x"34020001", 18493 => x"bc4c6000", 18494 => x"b9816000",
    18495 => x"596c0000", 18496 => x"e000000a", 18497 => x"34030001",
    18498 => x"29640000", 18499 => x"bc611800", 18500 => x"a4601800",
    18501 => x"a0641800", 18502 => x"59630000", 18503 => x"29a30128",
    18504 => x"44230002", 18505 => x"fbfff9ac", 18506 => x"2b9d0004",
    18507 => x"2b8b0010", 18508 => x"2b8c000c", 18509 => x"2b8d0008",
    18510 => x"379c0010", 18511 => x"c3a00000", 18512 => x"08210090",
    18513 => x"78020001", 18514 => x"38428c3c", 18515 => x"b4411000",
    18516 => x"28410140", 18517 => x"28430140", 18518 => x"34020004",
    18519 => x"7c210001", 18520 => x"5c620002", 18521 => x"38210002",
    18522 => x"c3a00000", 18523 => x"4c200005", 18524 => x"78010001",
    18525 => x"38218c3c", 18526 => x"28210054", 18527 => x"c3a00000",
    18528 => x"78020001", 18529 => x"38428c3c", 18530 => x"5c200003",
    18531 => x"284100dc", 18532 => x"c3a00000", 18533 => x"3421ffff",
    18534 => x"08210090", 18535 => x"b4411000", 18536 => x"2841016c",
    18537 => x"c3a00000", 18538 => x"78030001", 18539 => x"38638c20",
    18540 => x"4c200007", 18541 => x"78010001", 18542 => x"38218c3c",
    18543 => x"58220054", 18544 => x"28610000", 18545 => x"58220040",
    18546 => x"c3a00000", 18547 => x"2024000f", 18548 => x"28630000",
    18549 => x"3c840010", 18550 => x"2045ffff", 18551 => x"b8a42000",
    18552 => x"58640044", 18553 => x"78030001", 18554 => x"38638c3c",
    18555 => x"5c200003", 18556 => x"586200dc", 18557 => x"c3a00000",
    18558 => x"3421ffff", 18559 => x"08210090", 18560 => x"b4611800",
    18561 => x"5862016c", 18562 => x"c3a00000", 18563 => x"379cffcc",
    18564 => x"5b8b0034", 18565 => x"5b8c0030", 18566 => x"5b8d002c",
    18567 => x"5b8e0028", 18568 => x"5b8f0024", 18569 => x"5b900020",
    18570 => x"5b91001c", 18571 => x"5b920018", 18572 => x"5b930014",
    18573 => x"5b940010", 18574 => x"5b95000c", 18575 => x"5b960008",
    18576 => x"5b9d0004", 18577 => x"78010001", 18578 => x"38218c3c",
    18579 => x"28220000", 18580 => x"34010001", 18581 => x"34140000",
    18582 => x"5c410005", 18583 => x"78010001", 18584 => x"38218cd4",
    18585 => x"fbfffa05", 18586 => x"b820a000", 18587 => x"78110001",
    18588 => x"780b0001", 18589 => x"780e0001", 18590 => x"340d0000",
    18591 => x"340c0001", 18592 => x"3a318f78", 18593 => x"396b8c3c",
    18594 => x"340f0001", 18595 => x"39ce8c20", 18596 => x"34120002",
    18597 => x"34160003", 18598 => x"34150004", 18599 => x"e0000047",
    18600 => x"3593ffff", 18601 => x"0a700090", 18602 => x"b5708000",
    18603 => x"2a010140", 18604 => x"442f000f", 18605 => x"29c10000",
    18606 => x"bdec1000", 18607 => x"28210020", 18608 => x"00210008",
    18609 => x"202100ff", 18610 => x"a0220800", 18611 => x"5c200008",
    18612 => x"b9800800", 18613 => x"fbfffe9e", 18614 => x"b9800800",
    18615 => x"34020000", 18616 => x"fbfffca7", 18617 => x"35ad0001",
    18618 => x"5a0f0140", 18619 => x"0a610090", 18620 => x"b5618000",
    18621 => x"2a020140", 18622 => x"44520014", 18623 => x"48520003",
    18624 => x"5c4f002d", 18625 => x"e0000004", 18626 => x"44560017",
    18627 => x"5c55002a", 18628 => x"e000001e", 18629 => x"296100f0",
    18630 => x"44200027", 18631 => x"29c10000", 18632 => x"bdec1000",
    18633 => x"28210020", 18634 => x"00210008", 18635 => x"202100ff",
    18636 => x"a0220800", 18637 => x"44200020", 18638 => x"b9800800",
    18639 => x"fbfffe73", 18640 => x"5a120140", 18641 => x"e000001b",
    18642 => x"2a010180", 18643 => x"4420001a", 18644 => x"29620018",
    18645 => x"b9800800", 18646 => x"fbfffcc1", 18647 => x"5a160140",
    18648 => x"e0000014", 18649 => x"34210148", 18650 => x"b5610800",
    18651 => x"fbfffc22", 18652 => x"5c200011", 18653 => x"b9800800",
    18654 => x"34020001", 18655 => x"fbfffc80", 18656 => x"5a150140",
    18657 => x"e000000b", 18658 => x"296100f0", 18659 => x"44200003",
    18660 => x"2a010180", 18661 => x"5c200008", 18662 => x"0a730090",
    18663 => x"b9800800", 18664 => x"34020000", 18665 => x"b5739800",
    18666 => x"fbfffc75", 18667 => x"5a6f0140", 18668 => x"35ad0001",
    18669 => x"358c0001", 18670 => x"2a210000", 18671 => x"482cffb9",
    18672 => x"29630000", 18673 => x"78020001", 18674 => x"38426fc4",
    18675 => x"5843000c", 18676 => x"29630014", 18677 => x"28410008",
    18678 => x"7dad0000", 18679 => x"58430010", 18680 => x"29630004",
    18681 => x"34210002", 18682 => x"b5b4a000", 18683 => x"58430014",
    18684 => x"296300a4", 18685 => x"58410008", 18686 => x"7e810000",
    18687 => x"58430018", 18688 => x"29630068", 18689 => x"5843001c",
    18690 => x"296300f0", 18691 => x"58430020", 18692 => x"29630054",
    18693 => x"58430024", 18694 => x"296300dc", 18695 => x"58430028",
    18696 => x"29630010", 18697 => x"5843002c", 18698 => x"2b9d0004",
    18699 => x"2b8b0034", 18700 => x"2b8c0030", 18701 => x"2b8d002c",
    18702 => x"2b8e0028", 18703 => x"2b8f0024", 18704 => x"2b900020",
    18705 => x"2b91001c", 18706 => x"2b920018", 18707 => x"2b930014",
    18708 => x"2b940010", 18709 => x"2b95000c", 18710 => x"2b960008",
    18711 => x"379c0034", 18712 => x"c3a00000", 18713 => x"379cfff8",
    18714 => x"5b8b0008", 18715 => x"5b9d0004", 18716 => x"fbffb756",
    18717 => x"34020000", 18718 => x"3401ffff", 18719 => x"fbffff4b",
    18720 => x"34010001", 18721 => x"fbfffc53", 18722 => x"380bffff",
    18723 => x"b9601000", 18724 => x"3401ffff", 18725 => x"fbffff45",
    18726 => x"34010001", 18727 => x"fbfffc4d", 18728 => x"34020000",
    18729 => x"34010000", 18730 => x"fbffff40", 18731 => x"34010000",
    18732 => x"fbfffc48", 18733 => x"b9601000", 18734 => x"34010000",
    18735 => x"fbffff3b", 18736 => x"34010000", 18737 => x"fbfffc43",
    18738 => x"34010002", 18739 => x"fbfffc41", 18740 => x"2b9d0004",
    18741 => x"2b8b0008", 18742 => x"379c0008", 18743 => x"c3a00000",
    18744 => x"379cfff0", 18745 => x"5b8b0010", 18746 => x"5b8c000c",
    18747 => x"5b8d0008", 18748 => x"5b9d0004", 18749 => x"78010001",
    18750 => x"780b0001", 18751 => x"38215744", 18752 => x"780c0001",
    18753 => x"396bf800", 18754 => x"282d0000", 18755 => x"398c5730",
    18756 => x"e0000005", 18757 => x"b9800800", 18758 => x"fbffe839",
    18759 => x"340103e8", 18760 => x"fbffedfc", 18761 => x"29610000",
    18762 => x"5c2dfffb", 18763 => x"2b9d0004", 18764 => x"2b8b0010",
    18765 => x"2b8c000c", 18766 => x"2b8d0008", 18767 => x"379c0010",
    18768 => x"c3a00000", 18769 => x"c3a00000", 18770 => x"379cfff8",
    18771 => x"5b8b0008", 18772 => x"5b9d0004", 18773 => x"28240014",
    18774 => x"b8201800", 18775 => x"b8403000", 18776 => x"44800015",
    18777 => x"28250010", 18778 => x"20a50002", 18779 => x"5ca00007",
    18780 => x"b4862000", 18781 => x"b8800800", 18782 => x"2b9d0004",
    18783 => x"2b8b0008", 18784 => x"379c0008", 18785 => x"c3a00000",
    18786 => x"346b0030", 18787 => x"b4861000", 18788 => x"b9600800",
    18789 => x"34030040", 18790 => x"f80001cc", 18791 => x"b9602000",
    18792 => x"b8800800", 18793 => x"2b9d0004", 18794 => x"2b8b0008",
    18795 => x"379c0008", 18796 => x"c3a00000", 18797 => x"28250010",
    18798 => x"20a70004", 18799 => x"5ce4ffeb", 18800 => x"2825001c",
    18801 => x"34040000", 18802 => x"44a7ffeb", 18803 => x"342b0030",
    18804 => x"34040040", 18805 => x"b9601800", 18806 => x"d8a00000",
    18807 => x"b9602000", 18808 => x"e3fffff0", 18809 => x"379cfff4",
    18810 => x"5b8b0008", 18811 => x"5b9d0004", 18812 => x"28220014",
    18813 => x"b8205800", 18814 => x"44400013", 18815 => x"2961000c",
    18816 => x"b4411000", 18817 => x"28430000", 18818 => x"78040001",
    18819 => x"388457f0", 18820 => x"28820000", 18821 => x"3401ffec",
    18822 => x"5c620007", 18823 => x"78020001", 18824 => x"38428c14",
    18825 => x"28430000", 18826 => x"34010000", 18827 => x"584b0000",
    18828 => x"5963007c", 18829 => x"2b9d0004", 18830 => x"2b8b0008",
    18831 => x"379c000c", 18832 => x"c3a00000", 18833 => x"28230010",
    18834 => x"20630004", 18835 => x"5c62ffec", 18836 => x"2825001c",
    18837 => x"2822000c", 18838 => x"3783000c", 18839 => x"34040004",
    18840 => x"d8a00000", 18841 => x"2b83000c", 18842 => x"e3ffffe8",
    18843 => x"379cfff0", 18844 => x"5b8b0010", 18845 => x"5b8c000c",
    18846 => x"5b8d0008", 18847 => x"5b9d0004", 18848 => x"b8205800",
    18849 => x"44400047", 18850 => x"2822000c", 18851 => x"58200080",
    18852 => x"582000b0", 18853 => x"58220090", 18854 => x"340c0000",
    18855 => x"b9600800", 18856 => x"fbffffaa", 18857 => x"59610028",
    18858 => x"4022003f", 18859 => x"5c400006", 18860 => x"78040001",
    18861 => x"388457f0", 18862 => x"28230000", 18863 => x"28820000",
    18864 => x"4462005d", 18865 => x"34010000", 18866 => x"45800030",
    18867 => x"3583ffff", 18868 => x"346c0028", 18869 => x"b58c0800",
    18870 => x"b4210800", 18871 => x"b5610800", 18872 => x"28220000",
    18873 => x"5c40000f", 18874 => x"34010000", 18875 => x"44620027",
    18876 => x"34620027", 18877 => x"b4421000", 18878 => x"b4421000",
    18879 => x"b5621000", 18880 => x"e0000002", 18881 => x"44610044",
    18882 => x"28410000", 18883 => x"3463ffff", 18884 => x"3442fffc",
    18885 => x"4420fffc", 18886 => x"596300b0", 18887 => x"346c0028",
    18888 => x"346d0024", 18889 => x"b5ad6800", 18890 => x"b5ad6800",
    18891 => x"b56d6800", 18892 => x"29a20000", 18893 => x"b9600800",
    18894 => x"b58c6000", 18895 => x"fbffff83", 18896 => x"b58c6000",
    18897 => x"b56c1000", 18898 => x"29a40000", 18899 => x"28430000",
    18900 => x"296c00b0", 18901 => x"34840040", 18902 => x"3463ffff",
    18903 => x"59610028", 18904 => x"59a40000", 18905 => x"58430000",
    18906 => x"35830020", 18907 => x"b4631800", 18908 => x"b4631800",
    18909 => x"b5631800", 18910 => x"2824000c", 18911 => x"28620000",
    18912 => x"b4441000", 18913 => x"59620074", 18914 => x"2b9d0004",
    18915 => x"2b8b0010", 18916 => x"2b8c000c", 18917 => x"2b8d0008",
    18918 => x"379c0010", 18919 => x"c3a00000", 18920 => x"28210028",
    18921 => x"296300b0", 18922 => x"34050002", 18923 => x"4024003f",
    18924 => x"eca32800", 18925 => x"64840002", 18926 => x"a0852000",
    18927 => x"4482ffc5", 18928 => x"34620020", 18929 => x"b4421000",
    18930 => x"b4421000", 18931 => x"b5621000", 18932 => x"28450000",
    18933 => x"34640025", 18934 => x"28220004", 18935 => x"b4842000",
    18936 => x"b4842000", 18937 => x"b4a21000", 18938 => x"b5642000",
    18939 => x"58820000", 18940 => x"2824000c", 18941 => x"34610021",
    18942 => x"b4210800", 18943 => x"b4210800", 18944 => x"b5610800",
    18945 => x"b4852800", 18946 => x"346c0001", 18947 => x"58250000",
    18948 => x"e3ffffa3", 18949 => x"34010000", 18950 => x"596000b0",
    18951 => x"2b9d0004", 18952 => x"2b8b0010", 18953 => x"2b8c000c",
    18954 => x"2b8d0008", 18955 => x"379c0010", 18956 => x"c3a00000",
    18957 => x"35820024", 18958 => x"b4421000", 18959 => x"b4421000",
    18960 => x"b5621800", 18961 => x"2c250004", 18962 => x"28640000",
    18963 => x"35820028", 18964 => x"b4421000", 18965 => x"b4421000",
    18966 => x"b5621000", 18967 => x"34a5ffff", 18968 => x"34840040",
    18969 => x"58450000", 18970 => x"58640000", 18971 => x"596c00b0",
    18972 => x"e3ffffbe", 18973 => x"379cffec", 18974 => x"5b8b0014",
    18975 => x"5b8c0010", 18976 => x"5b8d000c", 18977 => x"5b8e0008",
    18978 => x"5b9d0004", 18979 => x"b8406000", 18980 => x"34020001",
    18981 => x"b8205800", 18982 => x"b8607000", 18983 => x"b8806800",
    18984 => x"fbffff73", 18985 => x"b9600800", 18986 => x"34020000",
    18987 => x"fbffff70", 18988 => x"b8202800", 18989 => x"4420001e",
    18990 => x"28a10018", 18991 => x"5c2cfffa", 18992 => x"28a1001c",
    18993 => x"5c2efff8", 18994 => x"28a10020", 18995 => x"5c2dfff6",
    18996 => x"296100b0", 18997 => x"59650028", 18998 => x"28a2000c",
    18999 => x"34210020", 19000 => x"b4210800", 19001 => x"b4210800",
    19002 => x"b5610800", 19003 => x"28230000", 19004 => x"34010000",
    19005 => x"b4431800", 19006 => x"59630074", 19007 => x"28a30014",
    19008 => x"59600078", 19009 => x"34630001", 19010 => x"c8621000",
    19011 => x"59620070", 19012 => x"2b9d0004", 19013 => x"2b8b0014",
    19014 => x"2b8c0010", 19015 => x"2b8d000c", 19016 => x"2b8e0008",
    19017 => x"379c0014", 19018 => x"c3a00000", 19019 => x"3401fffe",
    19020 => x"e3fffff8", 19021 => x"379cfff8", 19022 => x"5b8b0008",
    19023 => x"5b9d0004", 19024 => x"b8205800", 19025 => x"fbffffcc",
    19026 => x"4c200005", 19027 => x"2b9d0004", 19028 => x"2b8b0008",
    19029 => x"379c0008", 19030 => x"c3a00000", 19031 => x"29610074",
    19032 => x"59600028", 19033 => x"2b9d0004", 19034 => x"2b8b0008",
    19035 => x"379c0008", 19036 => x"c3a00000", 19037 => x"2045ffff",
    19038 => x"00460010", 19039 => x"2088ffff", 19040 => x"00890010",
    19041 => x"89053800", 19042 => x"89064000", 19043 => x"89252800",
    19044 => x"00ea0010", 19045 => x"89263000", 19046 => x"b5052800",
    19047 => x"b4aa2800", 19048 => x"50a80003", 19049 => x"78080001",
    19050 => x"b4c83000", 19051 => x"88431000", 19052 => x"88812000",
    19053 => x"00a10010", 19054 => x"3ca50010", 19055 => x"b4c13000",
    19056 => x"20e7ffff", 19057 => x"b4440800", 19058 => x"b4260800",
    19059 => x"b4a71000", 19060 => x"c3a00000", 19061 => x"44600008",
    19062 => x"34040020", 19063 => x"c8832000", 19064 => x"48800006",
    19065 => x"c8041000", 19066 => x"34030000", 19067 => x"80221000",
    19068 => x"b8600800", 19069 => x"c3a00000", 19070 => x"bc242000",
    19071 => x"80431000", 19072 => x"80231800", 19073 => x"b8821000",
    19074 => x"b8600800", 19075 => x"e3fffffa", 19076 => x"379cfff8",
    19077 => x"5b8b0008", 19078 => x"5b9d0004", 19079 => x"44400022",
    19080 => x"b8412000", 19081 => x"3403000f", 19082 => x"5483000b",
    19083 => x"78030001", 19084 => x"38635c68", 19085 => x"3c210004",
    19086 => x"b4621000", 19087 => x"b4410800", 19088 => x"40210000",
    19089 => x"2b9d0004", 19090 => x"2b8b0008", 19091 => x"379c0008",
    19092 => x"c3a00000", 19093 => x"340b0000", 19094 => x"4c200003",
    19095 => x"c8010800", 19096 => x"340b0001", 19097 => x"4c400003",
    19098 => x"c8021000", 19099 => x"196b0001", 19100 => x"90c01800",
    19101 => x"20630002", 19102 => x"44600008", 19103 => x"8c220800",
    19104 => x"45600002", 19105 => x"c8010800", 19106 => x"2b9d0004",
    19107 => x"2b8b0008", 19108 => x"379c0008", 19109 => x"c3a00000",
    19110 => x"34030000", 19111 => x"f800004a", 19112 => x"e3fffff8",
    19113 => x"90000800", 19114 => x"20210001", 19115 => x"3c210001",
    19116 => x"d0010000", 19117 => x"90e00800", 19118 => x"bba0f000",
    19119 => x"342100a0", 19120 => x"c0200000", 19121 => x"379cfff8",
    19122 => x"5b8b0008", 19123 => x"5b9d0004", 19124 => x"44400015",
    19125 => x"340b0000", 19126 => x"4c200003", 19127 => x"c8010800",
    19128 => x"340b0001", 19129 => x"1443001f", 19130 => x"90c02000",
    19131 => x"98621000", 19132 => x"20840002", 19133 => x"c8431000",
    19134 => x"44800008", 19135 => x"c4220800", 19136 => x"45600002",
    19137 => x"c8010800", 19138 => x"2b9d0004", 19139 => x"2b8b0008",
    19140 => x"379c0008", 19141 => x"c3a00000", 19142 => x"34030001",
    19143 => x"f800002a", 19144 => x"e3fffff8", 19145 => x"90000800",
    19146 => x"20210001", 19147 => x"3c210001", 19148 => x"d0010000",
    19149 => x"90e00800", 19150 => x"bba0f000", 19151 => x"342100a0",
    19152 => x"c0200000", 19153 => x"379cfffc", 19154 => x"5b9d0004",
    19155 => x"44400006", 19156 => x"34030000", 19157 => x"f800001c",
    19158 => x"2b9d0004", 19159 => x"379c0004", 19160 => x"c3a00000",
    19161 => x"90000800", 19162 => x"20210001", 19163 => x"3c210001",
    19164 => x"d0010000", 19165 => x"90e00800", 19166 => x"bba0f000",
    19167 => x"342100a0", 19168 => x"c0200000", 19169 => x"379cfffc",
    19170 => x"5b9d0004", 19171 => x"44400006", 19172 => x"34030001",
    19173 => x"f800000c", 19174 => x"2b9d0004", 19175 => x"379c0004",
    19176 => x"c3a00000", 19177 => x"90000800", 19178 => x"20210001",
    19179 => x"3c210001", 19180 => x"d0010000", 19181 => x"90e00800",
    19182 => x"bba0f000", 19183 => x"342100a0", 19184 => x"c0200000",
    19185 => x"f4222000", 19186 => x"44800018", 19187 => x"34040001",
    19188 => x"4c40000b", 19189 => x"34050000", 19190 => x"54410003",
    19191 => x"c8220800", 19192 => x"b8a42800", 19193 => x"00840001",
    19194 => x"00420001", 19195 => x"5c80fffb", 19196 => x"5c600002",
    19197 => x"b8a00800", 19198 => x"c3a00000", 19199 => x"3c420001",
    19200 => x"3c840001", 19201 => x"f4222800", 19202 => x"7c860000",
    19203 => x"a0c52800", 19204 => x"44a00002", 19205 => x"4c40fffa",
    19206 => x"34050000", 19207 => x"4480fff5", 19208 => x"34050000",
    19209 => x"e3ffffed", 19210 => x"34040001", 19211 => x"34050000",
    19212 => x"e3ffffea", 19213 => x"1422001f", 19214 => x"98410800",
    19215 => x"c8220800", 19216 => x"c3a00000", 19217 => x"34060003",
    19218 => x"b8202000", 19219 => x"b8402800", 19220 => x"50c3000c",
    19221 => x"b8413000", 19222 => x"20c60003", 19223 => x"5cc0000b",
    19224 => x"34010003", 19225 => x"28860000", 19226 => x"28a20000",
    19227 => x"5cc20005", 19228 => x"3463fffc", 19229 => x"34840004",
    19230 => x"34a50004", 19231 => x"5461fffa", 19232 => x"34010000",
    19233 => x"4460000e", 19234 => x"40860000", 19235 => x"40a10000",
    19236 => x"3462ffff", 19237 => x"44c10006", 19238 => x"e000000a",
    19239 => x"40860000", 19240 => x"40a10000", 19241 => x"3442ffff",
    19242 => x"5cc10006", 19243 => x"34840001", 19244 => x"34a50001",
    19245 => x"5c40fffa", 19246 => x"34010000", 19247 => x"c3a00000",
    19248 => x"c8c10800", 19249 => x"c3a00000", 19250 => x"3404000f",
    19251 => x"b8203800", 19252 => x"b8403000", 19253 => x"5083002d",
    19254 => x"b8412000", 19255 => x"20840003", 19256 => x"5c80002b",
    19257 => x"b8402000", 19258 => x"b8202800", 19259 => x"b8603000",
    19260 => x"3407000f", 19261 => x"28880000", 19262 => x"34c6fff0",
    19263 => x"58a80000", 19264 => x"28880004", 19265 => x"58a80004",
    19266 => x"28880008", 19267 => x"58a80008", 19268 => x"2888000c",
    19269 => x"34840010", 19270 => x"58a8000c", 19271 => x"34a50010",
    19272 => x"54c7fff5", 19273 => x"3463fff0", 19274 => x"00660004",
    19275 => x"2063000f", 19276 => x"34c60001", 19277 => x"3cc60004",
    19278 => x"b4263800", 19279 => x"b4463000", 19280 => x"34020003",
    19281 => x"50430011", 19282 => x"34020000", 19283 => x"34080003",
    19284 => x"b4c22000", 19285 => x"28850000", 19286 => x"b4e22000",
    19287 => x"34420004", 19288 => x"58850000", 19289 => x"c8622000",
    19290 => x"5488fffa", 19291 => x"3463fffc", 19292 => x"00620002",
    19293 => x"20630003", 19294 => x"34420001", 19295 => x"3c420002",
    19296 => x"b4e23800", 19297 => x"b4c23000", 19298 => x"44600008",
    19299 => x"34020000", 19300 => x"b4c22000", 19301 => x"40850000",
    19302 => x"b4e22000", 19303 => x"34420001", 19304 => x"30850000",
    19305 => x"5c43fffb", 19306 => x"c3a00000", 19307 => x"b8203800",
    19308 => x"b8403000", 19309 => x"5041000c", 19310 => x"b4432000",
    19311 => x"5024000a", 19312 => x"4460003f", 19313 => x"b4231000",
    19314 => x"3484ffff", 19315 => x"40850000", 19316 => x"3442ffff",
    19317 => x"3463ffff", 19318 => x"30450000", 19319 => x"5c60fffb",
    19320 => x"c3a00000", 19321 => x"3404000f", 19322 => x"5083002d",
    19323 => x"b8412000", 19324 => x"20840003", 19325 => x"5c80002b",
    19326 => x"b8402000", 19327 => x"b8202800", 19328 => x"b8603000",
    19329 => x"3407000f", 19330 => x"28880000", 19331 => x"34c6fff0",
    19332 => x"58a80000", 19333 => x"28880004", 19334 => x"58a80004",
    19335 => x"28880008", 19336 => x"58a80008", 19337 => x"2888000c",
    19338 => x"34840010", 19339 => x"58a8000c", 19340 => x"34a50010",
    19341 => x"54c7fff5", 19342 => x"3463fff0", 19343 => x"00660004",
    19344 => x"2063000f", 19345 => x"34c60001", 19346 => x"3cc60004",
    19347 => x"b4263800", 19348 => x"b4463000", 19349 => x"34020003",
    19350 => x"50430011", 19351 => x"34020000", 19352 => x"34080003",
    19353 => x"b4c22000", 19354 => x"28850000", 19355 => x"b4e22000",
    19356 => x"34420004", 19357 => x"58850000", 19358 => x"c8622000",
    19359 => x"5488fffa", 19360 => x"3463fffc", 19361 => x"00620002",
    19362 => x"20630003", 19363 => x"34420001", 19364 => x"3c420002",
    19365 => x"b4e23800", 19366 => x"b4c23000", 19367 => x"44600008",
    19368 => x"34020000", 19369 => x"b4c22000", 19370 => x"40850000",
    19371 => x"b4e22000", 19372 => x"34420001", 19373 => x"30850000",
    19374 => x"5c43fffb", 19375 => x"c3a00000", 19376 => x"20250003",
    19377 => x"b8202000", 19378 => x"44a0000b", 19379 => x"4460002c",
    19380 => x"3463ffff", 19381 => x"204600ff", 19382 => x"e0000003",
    19383 => x"44600028", 19384 => x"3463ffff", 19385 => x"30860000",
    19386 => x"34840001", 19387 => x"20850003", 19388 => x"5ca0fffb",
    19389 => x"34050003", 19390 => x"50a3001a", 19391 => x"204500ff",
    19392 => x"3ca60008", 19393 => x"340a000f", 19394 => x"b8c52800",
    19395 => x"3ca60010", 19396 => x"b8804000", 19397 => x"b8c53000",
    19398 => x"b8603800", 19399 => x"b8802800", 19400 => x"3409000f",
    19401 => x"546a0017", 19402 => x"34040000", 19403 => x"34070003",
    19404 => x"b5042800", 19405 => x"34840004", 19406 => x"58a60000",
    19407 => x"c8642800", 19408 => x"54a7fffc", 19409 => x"3463fffc",
    19410 => x"00640002", 19411 => x"20630003", 19412 => x"34840001",
    19413 => x"3c840002", 19414 => x"b5044000", 19415 => x"b9002000",
    19416 => x"44600007", 19417 => x"204200ff", 19418 => x"34050000",
    19419 => x"b4853000", 19420 => x"30c20000", 19421 => x"34a50001",
    19422 => x"5c65fffd", 19423 => x"c3a00000", 19424 => x"58a60000",
    19425 => x"58a60004", 19426 => x"58a60008", 19427 => x"58a6000c",
    19428 => x"34e7fff0", 19429 => x"34a50010", 19430 => x"54e9fffa",
    19431 => x"3463fff0", 19432 => x"00680004", 19433 => x"2063000f",
    19434 => x"35080001", 19435 => x"3d080004", 19436 => x"b4884000",
    19437 => x"34040003", 19438 => x"5464ffdc", 19439 => x"b9002000",
    19440 => x"e3ffffe8", 19441 => x"78030001", 19442 => x"38636fc0",
    19443 => x"28670000", 19444 => x"b8204800", 19445 => x"34030000",
    19446 => x"34060001", 19447 => x"e0000009", 19448 => x"40840000",
    19449 => x"b4e44000", 19450 => x"41080001", 19451 => x"21080003",
    19452 => x"45060012", 19453 => x"c8a40800", 19454 => x"5c200013",
    19455 => x"44810012", 19456 => x"b5232800", 19457 => x"40a50000",
    19458 => x"b4432000", 19459 => x"34630001", 19460 => x"b4e54000",
    19461 => x"41080001", 19462 => x"21080003", 19463 => x"5d06fff1",
    19464 => x"40840000", 19465 => x"34a50020", 19466 => x"b4e44000",
    19467 => x"41080001", 19468 => x"21080003", 19469 => x"5d06fff0",
    19470 => x"34840020", 19471 => x"c8a40800", 19472 => x"4420ffef",
    19473 => x"c3a00000", 19474 => x"b8411800", 19475 => x"20630003",
    19476 => x"5c60001d", 19477 => x"b8202000", 19478 => x"28430000",
    19479 => x"28210000", 19480 => x"5c230018", 19481 => x"78030001",
    19482 => x"38635d68", 19483 => x"28670000", 19484 => x"78030001",
    19485 => x"38635d6c", 19486 => x"28660000", 19487 => x"a4201800",
    19488 => x"b4270800", 19489 => x"a0231800", 19490 => x"a0661800",
    19491 => x"34010000", 19492 => x"44600003", 19493 => x"e000001c",
    19494 => x"5c600019", 19495 => x"34840004", 19496 => x"28810000",
    19497 => x"34420004", 19498 => x"28480000", 19499 => x"b4272800",
    19500 => x"a4201800", 19501 => x"a0a31800", 19502 => x"a0661800",
    19503 => x"4428fff7", 19504 => x"b8800800", 19505 => x"40230000",
    19506 => x"5c600006", 19507 => x"e0000009", 19508 => x"34210001",
    19509 => x"40230000", 19510 => x"34420001", 19511 => x"44600005",
    19512 => x"40440000", 19513 => x"4464fffb", 19514 => x"c8640800",
    19515 => x"c3a00000", 19516 => x"40440000", 19517 => x"c8640800",
    19518 => x"c3a00000", 19519 => x"34010000", 19520 => x"c3a00000",
    19521 => x"c3a00000", 19522 => x"b8412800", 19523 => x"20a50003",
    19524 => x"b8403800", 19525 => x"b8202000", 19526 => x"5ca00018",
    19527 => x"78040001", 19528 => x"38845d68", 19529 => x"28430000",
    19530 => x"28880000", 19531 => x"78040001", 19532 => x"38845d6c",
    19533 => x"28870000", 19534 => x"a4603000", 19535 => x"b4682000",
    19536 => x"a0c43000", 19537 => x"a0c73000", 19538 => x"b8202000",
    19539 => x"5cc5000a", 19540 => x"58830000", 19541 => x"34420004",
    19542 => x"28430000", 19543 => x"34840004", 19544 => x"a4603000",
    19545 => x"b4682800", 19546 => x"a0c52800", 19547 => x"a0a72800",
    19548 => x"44a0fff8", 19549 => x"b8403800", 19550 => x"34030000",
    19551 => x"b4e32800", 19552 => x"40a50000", 19553 => x"b4833000",
    19554 => x"34630001", 19555 => x"30c50000", 19556 => x"5ca0fffb",
    19557 => x"c3a00000", 19558 => x"20220003", 19559 => x"4440002c",
    19560 => x"40230000", 19561 => x"34020000", 19562 => x"44600027",
    19563 => x"b8201000", 19564 => x"e0000003", 19565 => x"40430000",
    19566 => x"44600022", 19567 => x"34420001", 19568 => x"20430003",
    19569 => x"5c60fffc", 19570 => x"78040001", 19571 => x"38845d68",
    19572 => x"28430000", 19573 => x"28860000", 19574 => x"78040001",
    19575 => x"38845d6c", 19576 => x"28850000", 19577 => x"a4602000",
    19578 => x"b4661800", 19579 => x"a0641800", 19580 => x"a0651800",
    19581 => x"5c600011", 19582 => x"34420004", 19583 => x"28430000",
    19584 => x"b4662000", 19585 => x"a4601800", 19586 => x"a0831800",
    19587 => x"a0651800", 19588 => x"5c60000a", 19589 => x"34420004",
    19590 => x"28430000", 19591 => x"b4662000", 19592 => x"a4601800",
    19593 => x"a0831800", 19594 => x"a0651800", 19595 => x"4460fff3",
    19596 => x"e0000002", 19597 => x"34420001", 19598 => x"40430000",
    19599 => x"5c60fffe", 19600 => x"c8411000", 19601 => x"b8400800",
    19602 => x"c3a00000", 19603 => x"b8201000", 19604 => x"e3ffffde",
    19605 => x"34060000", 19606 => x"44600017", 19607 => x"b8413800",
    19608 => x"20e70003", 19609 => x"3464ffff", 19610 => x"44e00015",
    19611 => x"40230000", 19612 => x"40450000", 19613 => x"5c65000f",
    19614 => x"34060000", 19615 => x"4480000e", 19616 => x"34210001",
    19617 => x"34420001", 19618 => x"5c600004", 19619 => x"e000000a",
    19620 => x"44800033", 19621 => x"44600032", 19622 => x"40230000",
    19623 => x"40450000", 19624 => x"3484ffff", 19625 => x"34210001",
    19626 => x"34420001", 19627 => x"4465fff9", 19628 => x"c8653000",
    19629 => x"b8c00800", 19630 => x"c3a00000", 19631 => x"b8202800",
    19632 => x"34010003", 19633 => x"b8402000", 19634 => x"50230028",
    19635 => x"28a10000", 19636 => x"28420000", 19637 => x"5c220025",
    19638 => x"3463fffc", 19639 => x"b8e03000", 19640 => x"4460fff5",
    19641 => x"78020001", 19642 => x"38425d68", 19643 => x"28490000",
    19644 => x"78020001", 19645 => x"38425d6c", 19646 => x"28480000",
    19647 => x"a4201000", 19648 => x"b4290800", 19649 => x"a0220800",
    19650 => x"a0280800", 19651 => x"34070003", 19652 => x"5c20ffe9",
    19653 => x"34a50004", 19654 => x"34840004", 19655 => x"54670006",
    19656 => x"b8a00800", 19657 => x"b8801000", 19658 => x"44600014",
    19659 => x"3464ffff", 19660 => x"e3ffffcf", 19661 => x"28a10000",
    19662 => x"288a0000", 19663 => x"b4293000", 19664 => x"a4201000",
    19665 => x"a0c21000", 19666 => x"a0481000", 19667 => x"5c2a0007",
    19668 => x"3463fffc", 19669 => x"44600002", 19670 => x"4440ffef",
    19671 => x"34060000", 19672 => x"b8c00800", 19673 => x"c3a00000",
    19674 => x"b8801000", 19675 => x"b8a00800", 19676 => x"3464ffff",
    19677 => x"e3ffffbe", 19678 => x"40a30000", 19679 => x"40850000",
    19680 => x"c8653000", 19681 => x"e3ffffcc", 19682 => x"b8412000",
    19683 => x"20840003", 19684 => x"74650003", 19685 => x"64840000",
    19686 => x"b8403000", 19687 => x"a0852000", 19688 => x"b8202800",
    19689 => x"44800015", 19690 => x"78040001", 19691 => x"38845d68",
    19692 => x"28890000", 19693 => x"78040001", 19694 => x"38845d6c",
    19695 => x"28880000", 19696 => x"340a0003", 19697 => x"e0000006",
    19698 => x"58a40000", 19699 => x"3463fffc", 19700 => x"34a50004",
    19701 => x"34420004", 19702 => x"51430007", 19703 => x"28440000",
    19704 => x"a4803800", 19705 => x"b4893000", 19706 => x"a0e63000",
    19707 => x"a0c83000", 19708 => x"44c0fff6", 19709 => x"b8403000",
    19710 => x"44600014", 19711 => x"40c20000", 19712 => x"3463ffff",
    19713 => x"34a40001", 19714 => x"30a20000", 19715 => x"44400009",
    19716 => x"34c20001", 19717 => x"4460000e", 19718 => x"40450000",
    19719 => x"3463ffff", 19720 => x"34420001", 19721 => x"30850000",
    19722 => x"34840001", 19723 => x"5ca0fffa", 19724 => x"34020000",
    19725 => x"44600007", 19726 => x"b4822800", 19727 => x"30a00000",
    19728 => x"34420001", 19729 => x"5c62fffd", 19730 => x"c3a00000",
    19731 => x"c3a00000", 19732 => x"c3a00000", 19733 => x"34030000",
    19734 => x"4440000c", 19735 => x"40240000", 19736 => x"4480000a",
    19737 => x"3442ffff", 19738 => x"b8201800", 19739 => x"e0000004",
    19740 => x"40640000", 19741 => x"3442ffff", 19742 => x"44800003",
    19743 => x"34630001", 19744 => x"5c40fffc", 19745 => x"c8611800",
    19746 => x"b8600800", 19747 => x"c3a00000", 19748 => x"57522043",
    19749 => x"6f72653a", 19750 => x"20737461", 19751 => x"7274696e",
    19752 => x"67207570", 19753 => x"2e2e2e0a", 19754 => x"00000000",
    19755 => x"556e6162", 19756 => x"6c652074", 19757 => x"6f206465",
    19758 => x"7465726d", 19759 => x"696e6520", 19760 => x"4d414320",
    19761 => x"61646472", 19762 => x"6573730a", 19763 => x"00000000",
    19764 => x"4c6f6361", 19765 => x"6c204d41", 19766 => x"43206164",
    19767 => x"64726573", 19768 => x"733a2025", 19769 => x"3032783a",
    19770 => x"25303278", 19771 => x"3a253032", 19772 => x"783a2530",
    19773 => x"32783a25", 19774 => x"3032783a", 19775 => x"25303278",
    19776 => x"0a000000", 19777 => x"73706c6c", 19778 => x"2d626800",
    19779 => x"7368656c", 19780 => x"6c2b6775", 19781 => x"69000000",
    19782 => x"70747000", 19783 => x"75707469", 19784 => x"6d650000",
    19785 => x"63686563", 19786 => x"6b2d6c69", 19787 => x"6e6b0000",
    19788 => x"69646c65", 19789 => x"00000000", 19790 => x"64696167",
    19791 => x"2d66736d", 19792 => x"2d312d25", 19793 => x"733a2025",
    19794 => x"3039642e", 19795 => x"25303364", 19796 => x"3a200000",
    19797 => x"454e5445", 19798 => x"52202573", 19799 => x"2c207061",
    19800 => x"636b6574", 19801 => x"206c656e", 19802 => x"2025690a",
    19803 => x"00000000", 19804 => x"25733a20", 19805 => x"7265656e",
    19806 => x"74657220", 19807 => x"696e2025", 19808 => x"69206d73",
    19809 => x"0a000000", 19810 => x"4c454156", 19811 => x"45202573",
    19812 => x"20286e65", 19813 => x"78743a20", 19814 => x"25336929",
    19815 => x"0a0a0000", 19816 => x"52454356", 19817 => x"20253032",
    19818 => x"64206279", 19819 => x"74657320", 19820 => x"61742025",
    19821 => x"642e2530", 19822 => x"39642028", 19823 => x"74797065",
    19824 => x"2025782c", 19825 => x"20257329", 19826 => x"0a000000",
    19827 => x"66736d20", 19828 => x"666f7220", 19829 => x"25733a20",
    19830 => x"4572726f", 19831 => x"72202569", 19832 => x"20696e20",
    19833 => x"25730a00", 19834 => x"66736d3a", 19835 => x"20556e6b",
    19836 => x"6e6f776e", 19837 => x"20737461", 19838 => x"74652066",
    19839 => x"6f722070", 19840 => x"6f727420", 19841 => x"25730a00",
    19842 => x"70707369", 19843 => x"00000000", 19844 => x"25732d25",
    19845 => x"692d2573", 19846 => x"3a200000", 19847 => x"25733a20",
    19848 => x"6572726f", 19849 => x"72207061", 19850 => x"7273696e",
    19851 => x"67202225", 19852 => x"73220a00", 19853 => x"64696167",
    19854 => x"2d636f6e", 19855 => x"66696700", 19856 => x"64696167",
    19857 => x"2d657874", 19858 => x"656e7369", 19859 => x"6f6e0000",
    19860 => x"64696167", 19861 => x"2d626d63", 19862 => x"00000000",
    19863 => x"64696167", 19864 => x"2d736572", 19865 => x"766f0000",
    19866 => x"64696167", 19867 => x"2d667261", 19868 => x"6d657300",
    19869 => x"64696167", 19870 => x"2d74696d", 19871 => x"65000000",
    19872 => x"64696167", 19873 => x"2d66736d", 19874 => x"00000000",
    19875 => x"50505369", 19876 => x"20666f72", 19877 => x"20575250",
    19878 => x"432e2043", 19879 => x"6f6d6d69", 19880 => x"74202573",
    19881 => x"2c206275", 19882 => x"696c7420", 19883 => x"6f6e204e",
    19884 => x"6f762033", 19885 => x"30203230", 19886 => x"31360a00",
    19887 => x"70707369", 19888 => x"2d763230", 19889 => x"31342e30",
    19890 => x"372d3139", 19891 => x"362d6763", 19892 => x"39336437",
    19893 => x"31300000", 19894 => x"50545020", 19895 => x"73746172",
    19896 => x"740a0000", 19897 => x"50545020", 19898 => x"73746f70",
    19899 => x"0a000000", 19900 => x"4c6f636b", 19901 => x"696e6720",
    19902 => x"504c4c00", 19903 => x"0a4c6f63", 19904 => x"6b207469",
    19905 => x"6d656f75", 19906 => x"742e0000", 19907 => x"2e000000",
    19908 => x"77723100", 19909 => x"25732573", 19910 => x"25303278",
    19911 => x"2d253032", 19912 => x"782d2530", 19913 => x"32782d25",
    19914 => x"3032782d", 19915 => x"25303278", 19916 => x"2d253032",
    19917 => x"782d2530", 19918 => x"32782d25", 19919 => x"3032782d",
    19920 => x"25303278", 19921 => x"2d253032", 19922 => x"780a0000",
    19923 => x"25732573", 19924 => x"25732028", 19925 => x"73697a65",
    19926 => x"20256929", 19927 => x"0a000000", 19928 => x"25732573",
    19929 => x"00000000", 19930 => x"25303278", 19931 => x"00000000",
    19932 => x"25735645", 19933 => x"5253494f", 19934 => x"4e3a2075",
    19935 => x"6e737570", 19936 => x"706f7274", 19937 => x"65642028",
    19938 => x"2569290a", 19939 => x"00000000", 19940 => x"25735645",
    19941 => x"5253494f", 19942 => x"4e3a2025", 19943 => x"69202874",
    19944 => x"79706520", 19945 => x"25692c20", 19946 => x"6c656e20",
    19947 => x"25692c20", 19948 => x"646f6d61", 19949 => x"696e2025",
    19950 => x"69290a00", 19951 => x"2573464c", 19952 => x"4147533a",
    19953 => x"20307825", 19954 => x"30347820", 19955 => x"28636f72",
    19956 => x"72656374", 19957 => x"696f6e20", 19958 => x"2530386c",
    19959 => x"75290a00", 19960 => x"504f5254", 19961 => x"3a200000",
    19962 => x"25735245", 19963 => x"53543a20", 19964 => x"73657120",
    19965 => x"25692c20", 19966 => x"6374726c", 19967 => x"2025692c",
    19968 => x"206c6f67", 19969 => x"2d696e74", 19970 => x"65727661",
    19971 => x"6c202569", 19972 => x"0a000000", 19973 => x"25734d45",
    19974 => x"53534147", 19975 => x"453a2028", 19976 => x"45292053",
    19977 => x"594e430a", 19978 => x"00000000", 19979 => x"25732573",
    19980 => x"256c752e", 19981 => x"25303969", 19982 => x"0a000000",
    19983 => x"4d53472d", 19984 => x"53594e43", 19985 => x"3a200000",
    19986 => x"25734d45", 19987 => x"53534147", 19988 => x"453a2028",
    19989 => x"45292044", 19990 => x"454c4159", 19991 => x"5f524551",
    19992 => x"0a000000", 19993 => x"4d53472d", 19994 => x"44454c41",
    19995 => x"595f5245", 19996 => x"513a2000", 19997 => x"25734d45",
    19998 => x"53534147", 19999 => x"453a2028", 20000 => x"47292046",
    20001 => x"4f4c4c4f", 20002 => x"575f5550", 20003 => x"0a000000",
    20004 => x"4d53472d", 20005 => x"464f4c4c", 20006 => x"4f575f55",
    20007 => x"503a2000", 20008 => x"25734d45", 20009 => x"53534147",
    20010 => x"453a2028", 20011 => x"47292044", 20012 => x"454c4159",
    20013 => x"5f524553", 20014 => x"500a0000", 20015 => x"4d53472d",
    20016 => x"44454c41", 20017 => x"595f5245", 20018 => x"53503a20",
    20019 => x"00000000", 20020 => x"25734d45", 20021 => x"53534147",
    20022 => x"453a2028", 20023 => x"47292041", 20024 => x"4e4e4f55",
    20025 => x"4e43450a", 20026 => x"00000000", 20027 => x"4d53472d",
    20028 => x"414e4e4f", 20029 => x"554e4345", 20030 => x"3a207374",
    20031 => x"616d7020", 20032 => x"00000000", 20033 => x"25732573",
    20034 => x"25303278", 20035 => x"2d253032", 20036 => x"782d2530",
    20037 => x"34780a00", 20038 => x"4d53472d", 20039 => x"414e4e4f",
    20040 => x"554e4345", 20041 => x"3a206772", 20042 => x"616e646d",
    20043 => x"61737465", 20044 => x"722d7175", 20045 => x"616c6974",
    20046 => x"79200000", 20047 => x"25734d53", 20048 => x"472d414e",
    20049 => x"4e4f554e", 20050 => x"43453a20", 20051 => x"6772616e",
    20052 => x"646d6173", 20053 => x"7465722d", 20054 => x"7072696f",
    20055 => x"20256920", 20056 => x"25690a00", 20057 => x"25732573",
    20058 => x"25303278", 20059 => x"2d253032", 20060 => x"782d2530",
    20061 => x"32782d25", 20062 => x"3032782d", 20063 => x"25303278",
    20064 => x"2d253032", 20065 => x"782d2530", 20066 => x"32782d25",
    20067 => x"3032780a", 20068 => x"00000000", 20069 => x"4d53472d",
    20070 => x"414e4e4f", 20071 => x"554e4345", 20072 => x"3a206772",
    20073 => x"616e646d", 20074 => x"61737465", 20075 => x"722d6964",
    20076 => x"20000000", 20077 => x"25734d45", 20078 => x"53534147",
    20079 => x"453a2028", 20080 => x"47292053", 20081 => x"49474e41",
    20082 => x"4c494e47", 20083 => x"0a000000", 20084 => x"4d53472d",
    20085 => x"5349474e", 20086 => x"414c494e", 20087 => x"473a2074",
    20088 => x"61726765", 20089 => x"742d706f", 20090 => x"72742000",
    20091 => x"2573544c", 20092 => x"563a2074", 20093 => x"6f6f2073",
    20094 => x"686f7274", 20095 => x"20282569", 20096 => x"202d2025",
    20097 => x"69203d20", 20098 => x"2569290a", 20099 => x"00000000",
    20100 => x"2573544c", 20101 => x"563a2074", 20102 => x"79706520",
    20103 => x"25303478", 20104 => x"206c656e", 20105 => x"20256920",
    20106 => x"6f756920", 20107 => x"25303278", 20108 => x"3a253032",
    20109 => x"783a2530", 20110 => x"32782073", 20111 => x"75622025",
    20112 => x"3032783a", 20113 => x"25303278", 20114 => x"3a253032",
    20115 => x"780a0000", 20116 => x"2573544c", 20117 => x"563a2074",
    20118 => x"6f6f2073", 20119 => x"686f7274", 20120 => x"20286578",
    20121 => x"70656374", 20122 => x"65642025", 20123 => x"692c2074",
    20124 => x"6f74616c", 20125 => x"20256929", 20126 => x"0a000000",
    20127 => x"544c563a", 20128 => x"20000000", 20129 => x"746c762d",
    20130 => x"636f6e74", 20131 => x"656e7400", 20132 => x"44554d50",
    20133 => x"3a200000", 20134 => x"7061796c", 20135 => x"6f616400",
    20136 => x"20696e76", 20137 => x"616c6964", 20138 => x"00000000",
    20139 => x"25735449", 20140 => x"4d453a20", 20141 => x"28256c69",
    20142 => x"202d2030", 20143 => x"78256c78", 20144 => x"2920256c",
    20145 => x"692e2530", 20146 => x"366c6925", 20147 => x"730a0000",
    20148 => x"2573564c", 20149 => x"414e2025", 20150 => x"690a0000",
    20151 => x"25734554", 20152 => x"483a2025", 20153 => x"30347820",
    20154 => x"28253032", 20155 => x"783a2530", 20156 => x"32783a25",
    20157 => x"3032783a", 20158 => x"25303278", 20159 => x"3a253032",
    20160 => x"783a2530", 20161 => x"3278202d", 20162 => x"3e202530",
    20163 => x"32783a25", 20164 => x"3032783a", 20165 => x"25303278",
    20166 => x"3a253032", 20167 => x"783a2530", 20168 => x"32783a25",
    20169 => x"30327829", 20170 => x"0a000000", 20171 => x"25734950",
    20172 => x"3a202569", 20173 => x"20282569", 20174 => x"2e25692e",
    20175 => x"25692e25", 20176 => x"69202d3e", 20177 => x"2025692e",
    20178 => x"25692e25", 20179 => x"692e2569", 20180 => x"29206c65",
    20181 => x"6e202569", 20182 => x"0a000000", 20183 => x"25735544",
    20184 => x"503a2028", 20185 => x"2569202d", 20186 => x"3e202569",
    20187 => x"29206c65", 20188 => x"6e202569", 20189 => x"0a000000",
    20190 => x"25733a20", 20191 => x"256c690a", 20192 => x"00000000",
    20193 => x"5761726e", 20194 => x"696e673a", 20195 => x"2025733a",
    20196 => x"2063616e", 20197 => x"206e6f74", 20198 => x"2061646a",
    20199 => x"75737420", 20200 => x"66726571", 20201 => x"5f707062",
    20202 => x"20256c69", 20203 => x"0a000000", 20204 => x"25733a20",
    20205 => x"25396c75", 20206 => x"2e253039", 20207 => x"6c690a00",
    20208 => x"25733a20", 20209 => x"736e743d", 20210 => x"25642c20",
    20211 => x"7365633d", 20212 => x"25642c20", 20213 => x"6e736563",
    20214 => x"3d25640a", 20215 => x"00000000", 20216 => x"73656e64",
    20217 => x"3a200000", 20218 => x"72656376", 20219 => x"3a200000",
    20220 => x"696e6974", 20221 => x"69616c69", 20222 => x"7a696e67",
    20223 => x"00000000", 20224 => x"6661756c", 20225 => x"74790000",
    20226 => x"64697361", 20227 => x"626c6564", 20228 => x"00000000",
    20229 => x"6c697374", 20230 => x"656e696e", 20231 => x"67000000",
    20232 => x"756e6361", 20233 => x"6c696272", 20234 => x"61746564",
    20235 => x"00000000", 20236 => x"736c6176", 20237 => x"65000000",
    20238 => x"756e6361", 20239 => x"6c696272", 20240 => x"61746564",
    20241 => x"2f77722d", 20242 => x"70726573", 20243 => x"656e7400",
    20244 => x"6d617374", 20245 => x"65722f77", 20246 => x"722d6d2d",
    20247 => x"6c6f636b", 20248 => x"00000000", 20249 => x"756e6361",
    20250 => x"6c696272", 20251 => x"61746564", 20252 => x"2f77722d",
    20253 => x"732d6c6f", 20254 => x"636b0000", 20255 => x"756e6361",
    20256 => x"6c696272", 20257 => x"61746564", 20258 => x"2f77722d",
    20259 => x"6c6f636b", 20260 => x"65640000", 20261 => x"77722d63",
    20262 => x"616c6962", 20263 => x"72617469", 20264 => x"6f6e0000",
    20265 => x"77722d63", 20266 => x"616c6962", 20267 => x"72617465",
    20268 => x"64000000", 20269 => x"77722d72", 20270 => x"6573702d",
    20271 => x"63616c69", 20272 => x"622d7265", 20273 => x"71000000",
    20274 => x"77722d6c", 20275 => x"696e6b2d", 20276 => x"6f6e0000",
    20277 => x"686f6f6b", 20278 => x"3a202573", 20279 => x"0a000000",
    20280 => x"5432206f", 20281 => x"72205433", 20282 => x"20696e63",
    20283 => x"6f727265", 20284 => x"63742c20", 20285 => x"64697363",
    20286 => x"61726469", 20287 => x"6e672074", 20288 => x"75706c65",
    20289 => x"0a000000", 20290 => x"48616e64", 20291 => x"7368616b",
    20292 => x"65206661", 20293 => x"696c7572", 20294 => x"653a206e",
    20295 => x"6f77206e", 20296 => x"6f6e2d77", 20297 => x"72202573",
    20298 => x"0a000000", 20299 => x"52657472", 20300 => x"79206f6e",
    20301 => x"2074696d", 20302 => x"656f7574", 20303 => x"0a000000",
    20304 => x"25733a20", 20305 => x"73756273", 20306 => x"74617465",
    20307 => x"2025690a", 20308 => x"00000000", 20309 => x"54783d3e",
    20310 => x"3e736361", 20311 => x"6c656450", 20312 => x"69636f73",
    20313 => x"65636f6e", 20314 => x"64732e6d", 20315 => x"7362203d",
    20316 => x"20307825", 20317 => x"780a0000", 20318 => x"54783d3e",
    20319 => x"3e736361", 20320 => x"6c656450", 20321 => x"69636f73",
    20322 => x"65636f6e", 20323 => x"64732e6c", 20324 => x"7362203d",
    20325 => x"20307825", 20326 => x"780a0000", 20327 => x"52782066",
    20328 => x"69786564", 20329 => x"2064656c", 20330 => x"6179203d",
    20331 => x"2025640a", 20332 => x"00000000", 20333 => x"52783d3e",
    20334 => x"3e736361", 20335 => x"6c656450", 20336 => x"69636f73",
    20337 => x"65636f6e", 20338 => x"64732e6d", 20339 => x"7362203d",
    20340 => x"20307825", 20341 => x"780a0000", 20342 => x"52783d3e",
    20343 => x"3e736361", 20344 => x"6c656450", 20345 => x"69636f73",
    20346 => x"65636f6e", 20347 => x"64732e6c", 20348 => x"7362203d",
    20349 => x"20307825", 20350 => x"780a0000", 20351 => x"4552524f",
    20352 => x"523a204e", 20353 => x"65772063", 20354 => x"6c617373",
    20355 => x"2025690a", 20356 => x"00000000", 20357 => x"4255473a",
    20358 => x"20547279", 20359 => x"696e6720", 20360 => x"746f2073",
    20361 => x"656e6420", 20362 => x"696e7661", 20363 => x"6c696420",
    20364 => x"77725f6d", 20365 => x"7367206d", 20366 => x"6f64653d",
    20367 => x"25782069", 20368 => x"643d2578", 20369 => x"00000000",
    20370 => x"68616e64", 20371 => x"6c652053", 20372 => x"69676e61",
    20373 => x"6c696e67", 20374 => x"206d7367", 20375 => x"2c206661",
    20376 => x"696c6564", 20377 => x"2c205468", 20378 => x"69732069",
    20379 => x"73206e6f", 20380 => x"74206f72", 20381 => x"67616e69",
    20382 => x"7a617469", 20383 => x"6f6e2065", 20384 => x"7874656e",
    20385 => x"73696f6e", 20386 => x"20544c56", 20387 => x"203d2030",
    20388 => x"7825780a", 20389 => x"00000000", 20390 => x"68616e64",
    20391 => x"6c652053", 20392 => x"69676e61", 20393 => x"6c696e67",
    20394 => x"206d7367", 20395 => x"2c206661", 20396 => x"696c6564",
    20397 => x"2c206e6f", 20398 => x"74204345", 20399 => x"524e2773",
    20400 => x"204f5549", 20401 => x"203d2030", 20402 => x"7825780a",
    20403 => x"00000000", 20404 => x"68616e64", 20405 => x"6c652053",
    20406 => x"69676e61", 20407 => x"6c696e67", 20408 => x"206d7367",
    20409 => x"2c206661", 20410 => x"696c6564", 20411 => x"2c206e6f",
    20412 => x"74205768", 20413 => x"69746520", 20414 => x"52616262",
    20415 => x"6974206d", 20416 => x"61676963", 20417 => x"206e756d",
    20418 => x"62657220", 20419 => x"3d203078", 20420 => x"25780a00",
    20421 => x"68616e64", 20422 => x"6c652053", 20423 => x"69676e61",
    20424 => x"6c696e67", 20425 => x"206d7367", 20426 => x"2c206661",
    20427 => x"696c6564", 20428 => x"2c206e6f", 20429 => x"74207375",
    20430 => x"70706f72", 20431 => x"74656420", 20432 => x"76657273",
    20433 => x"696f6e20", 20434 => x"6e756d62", 20435 => x"6572203d",
    20436 => x"20307825", 20437 => x"780a0000", 20438 => x"25732825",
    20439 => x"6429204d", 20440 => x"65737361", 20441 => x"67652063",
    20442 => x"616e2774", 20443 => x"20626520", 20444 => x"73656e74",
    20445 => x"0a000000", 20446 => x"53454e54", 20447 => x"20253032",
    20448 => x"64206279", 20449 => x"74657320", 20450 => x"61742025",
    20451 => x"642e2530", 20452 => x"39642028", 20453 => x"2573290a",
    20454 => x"00000000", 20455 => x"556e696e", 20456 => x"69746961",
    20457 => x"6c697a65", 20458 => x"64000000", 20459 => x"20287761",
    20460 => x"69742066", 20461 => x"6f722068", 20462 => x"77290000",
    20463 => x"4552524f", 20464 => x"523a2025", 20465 => x"733a2054",
    20466 => x"696d6573", 20467 => x"74616d70", 20468 => x"73496e63",
    20469 => x"6f727265", 20470 => x"63743a20", 20471 => x"25642025",
    20472 => x"64202564", 20473 => x"2025640a", 20474 => x"00000000",
    20475 => x"2573203d", 20476 => x"2025643a", 20477 => x"25643a25",
    20478 => x"640a0000", 20479 => x"73657276", 20480 => x"6f3a7431",
    20481 => x"00000000", 20482 => x"73657276", 20483 => x"6f3a7432",
    20484 => x"00000000", 20485 => x"73657276", 20486 => x"6f3a7433",
    20487 => x"00000000", 20488 => x"73657276", 20489 => x"6f3a7434",
    20490 => x"00000000", 20491 => x"2d3e6d64", 20492 => x"656c6179",
    20493 => x"00000000", 20494 => x"504c4c20", 20495 => x"4f75744f",
    20496 => x"664c6f63", 20497 => x"6b2c2073", 20498 => x"686f756c",
    20499 => x"64207265", 20500 => x"73746172", 20501 => x"74207379",
    20502 => x"6e630a00", 20503 => x"73657276", 20504 => x"6f3a6275",
    20505 => x"73790a00", 20506 => x"6f666673", 20507 => x"65745f68",
    20508 => x"773a2025", 20509 => x"6c692e25", 20510 => x"30396c69",
    20511 => x"20282b25", 20512 => x"6c69290a", 20513 => x"00000000",
    20514 => x"77725f73", 20515 => x"6572766f", 20516 => x"20737461",
    20517 => x"74653a20", 20518 => x"25732573", 20519 => x"0a000000",
    20520 => x"6f6c6473", 20521 => x"65747020", 20522 => x"25692c20",
    20523 => x"6f666673", 20524 => x"65742025", 20525 => x"693a2530",
    20526 => x"34690a00", 20527 => x"61646a75", 20528 => x"73742070",
    20529 => x"68617365", 20530 => x"2025690a", 20531 => x"00000000",
    20532 => x"53594e43", 20533 => x"5f4e5345", 20534 => x"43000000",
    20535 => x"53594e43", 20536 => x"5f534543", 20537 => x"00000000",
    20538 => x"53594e43", 20539 => x"5f504841", 20540 => x"53450000",
    20541 => x"54524143", 20542 => x"4b5f5048", 20543 => x"41534500",
    20544 => x"57414954", 20545 => x"5f4f4646", 20546 => x"5345545f",
    20547 => x"53544142", 20548 => x"4c450000", 20549 => x"7072652d",
    20550 => x"6d617374", 20551 => x"65720000", 20552 => x"70617373",
    20553 => x"69766500", 20554 => x"25733a20", 20555 => x"63616e27",
    20556 => x"7420696e", 20557 => x"69742065", 20558 => x"7874656e",
    20559 => x"73696f6e", 20560 => x"0a000000", 20561 => x"636c6f63",
    20562 => x"6b20636c", 20563 => x"61737320", 20564 => x"3d202564",
    20565 => x"0a000000", 20566 => x"636c6f63", 20567 => x"6b206163",
    20568 => x"63757261", 20569 => x"6379203d", 20570 => x"2025640a",
    20571 => x"00000000", 20572 => x"70705f73", 20573 => x"6c617665",
    20574 => x"203a2044", 20575 => x"656c6179", 20576 => x"20526573",
    20577 => x"7020646f", 20578 => x"65736e27", 20579 => x"74206d61",
    20580 => x"74636820", 20581 => x"44656c61", 20582 => x"79205265",
    20583 => x"710a0000", 20584 => x"4e657720", 20585 => x"666f7265",
    20586 => x"69676e20", 20587 => x"4d617374", 20588 => x"65722025",
    20589 => x"69206164", 20590 => x"6465640a", 20591 => x"00000000",
    20592 => x"4552524f", 20593 => x"523a2025", 20594 => x"733a2046",
    20595 => x"6f6c6c6f", 20596 => x"77207570", 20597 => x"206d6573",
    20598 => x"73616765", 20599 => x"20697320", 20600 => x"6e6f7420",
    20601 => x"66726f6d", 20602 => x"20637572", 20603 => x"72656e74",
    20604 => x"20706172", 20605 => x"656e740a", 20606 => x"00000000",
    20607 => x"4552524f", 20608 => x"523a2025", 20609 => x"733a2053",
    20610 => x"6c617665", 20611 => x"20776173", 20612 => x"206e6f74",
    20613 => x"20776169", 20614 => x"74696e67", 20615 => x"20612066",
    20616 => x"6f6c6c6f", 20617 => x"77207570", 20618 => x"206d6573",
    20619 => x"73616765", 20620 => x"0a000000", 20621 => x"4552524f",
    20622 => x"523a2025", 20623 => x"733a2053", 20624 => x"65717565",
    20625 => x"6e636549", 20626 => x"44202564", 20627 => x"20646f65",
    20628 => x"736e2774", 20629 => x"206d6174", 20630 => x"6368206c",
    20631 => x"61737420", 20632 => x"53796e63", 20633 => x"206d6573",
    20634 => x"73616765", 20635 => x"2025640a", 20636 => x"00000000",
    20637 => x"416e6e6f", 20638 => x"756e6365", 20639 => x"206d6573",
    20640 => x"73616765", 20641 => x"2066726f", 20642 => x"6d20616e",
    20643 => x"6f746865", 20644 => x"7220666f", 20645 => x"72656967",
    20646 => x"6e206d61", 20647 => x"73746572", 20648 => x"0a000000",
    20649 => x"25733a25", 20650 => x"693a2045", 20651 => x"72726f72",
    20652 => x"20310a00", 20653 => x"25733a25", 20654 => x"693a2045",
    20655 => x"72726f72", 20656 => x"20320a00", 20657 => x"42657374",
    20658 => x"20666f72", 20659 => x"6569676e", 20660 => x"206d6173",
    20661 => x"74657220", 20662 => x"69732025", 20663 => x"692f2569",
    20664 => x"0a000000", 20665 => x"25733a20", 20666 => x"6572726f",
    20667 => x"720a0000", 20668 => x"25733a20", 20669 => x"70617373",
    20670 => x"6976650a", 20671 => x"00000000", 20672 => x"25733a20",
    20673 => x"6d617374", 20674 => x"65720a00", 20675 => x"4e657720",
    20676 => x"55544320", 20677 => x"6f666673", 20678 => x"65743a20",
    20679 => x"25690a00", 20680 => x"25733a20", 20681 => x"736c6176",
    20682 => x"650a0000", 20683 => x"73796e63", 20684 => x"00000000",
    20685 => x"64656c61", 20686 => x"795f7265", 20687 => x"71000000",
    20688 => x"7064656c", 20689 => x"61795f72", 20690 => x"65710000",
    20691 => x"7064656c", 20692 => x"61795f72", 20693 => x"65737000",
    20694 => x"64656c61", 20695 => x"795f7265", 20696 => x"73700000",
    20697 => x"7064656c", 20698 => x"61795f72", 20699 => x"6573705f",
    20700 => x"666f6c6c", 20701 => x"6f775f75", 20702 => x"70000000",
    20703 => x"616e6e6f", 20704 => x"756e6365", 20705 => x"00000000",
    20706 => x"7369676e", 20707 => x"616c696e", 20708 => x"67000000",
    20709 => x"6d616e61", 20710 => x"67656d65", 20711 => x"6e740000",
    20712 => x"4552524f", 20713 => x"523a2042", 20714 => x"55473a20",
    20715 => x"25732064", 20716 => x"6f65736e", 20717 => x"27742073",
    20718 => x"7570706f", 20719 => x"7274206e", 20720 => x"65676174",
    20721 => x"69766573", 20722 => x"0a000000", 20723 => x"4552524f",
    20724 => x"523a204e", 20725 => x"65676174", 20726 => x"69766520",
    20727 => x"76616c75", 20728 => x"65206361", 20729 => x"6e6e6f74",
    20730 => x"20626520", 20731 => x"636f6e76", 20732 => x"65727465",
    20733 => x"6420696e", 20734 => x"746f2074", 20735 => x"696d6573",
    20736 => x"74616d70", 20737 => x"0a000000", 20738 => x"4552524f",
    20739 => x"523a2074", 20740 => x"6f5f5469", 20741 => x"6d65496e",
    20742 => x"7465726e", 20743 => x"616c3a20", 20744 => x"7365636f",
    20745 => x"6e647320", 20746 => x"6669656c", 20747 => x"64206973",
    20748 => x"20686967", 20749 => x"68657220", 20750 => x"7468616e",
    20751 => x"20736967", 20752 => x"6e656420", 20753 => x"696e7465",
    20754 => x"67657220", 20755 => x"28333262", 20756 => x"69747329",
    20757 => x"0a000000", 20758 => x"2d000000", 20759 => x"25732564",
    20760 => x"2e253039", 20761 => x"64000000", 20762 => x"6572726f",
    20763 => x"7220696e", 20764 => x"20745f6f", 20765 => x"70732d3e",
    20766 => x"73657276", 20767 => x"6f5f696e", 20768 => x"69740000",
    20769 => x"496e6974", 20770 => x"69616c69", 20771 => x"7a65643a",
    20772 => x"206f6273", 20773 => x"5f647269", 20774 => x"66742025",
    20775 => x"6c6c690a", 20776 => x"00000000", 20777 => x"636f7272",
    20778 => x"65637469", 20779 => x"6f6e2066", 20780 => x"69656c64",
    20781 => x"20313a20", 20782 => x"25730a00", 20783 => x"64697363",
    20784 => x"61726420", 20785 => x"54332f54", 20786 => x"343a2077",
    20787 => x"65206d69", 20788 => x"73732054", 20789 => x"312f5432",
    20790 => x"0a000000", 20791 => x"636f7272", 20792 => x"65637469",
    20793 => x"6f6e2066", 20794 => x"69656c64", 20795 => x"20323a20",
    20796 => x"25730a00", 20797 => x"54313a20", 20798 => x"25730a00",
    20799 => x"54323a20", 20800 => x"25730a00", 20801 => x"54333a20",
    20802 => x"25730a00", 20803 => x"54343a20", 20804 => x"25730a00",
    20805 => x"4d617374", 20806 => x"65722074", 20807 => x"6f20736c",
    20808 => x"6176653a", 20809 => x"2025730a", 20810 => x"00000000",
    20811 => x"536c6176", 20812 => x"6520746f", 20813 => x"206d6173",
    20814 => x"7465723a", 20815 => x"2025730a", 20816 => x"00000000",
    20817 => x"6d65616e", 20818 => x"50617468", 20819 => x"44656c61",
    20820 => x"793a2025", 20821 => x"730a0000", 20822 => x"73657276",
    20823 => x"6f206162", 20824 => x"6f727465", 20825 => x"642c2064",
    20826 => x"656c6179", 20827 => x"20677265", 20828 => x"61746572",
    20829 => x"20746861", 20830 => x"6e203120", 20831 => x"7365636f",
    20832 => x"6e640a00", 20833 => x"73657276", 20834 => x"6f206162",
    20835 => x"6f727465", 20836 => x"642c2064", 20837 => x"656c6179",
    20838 => x"20256420", 20839 => x"6f722025", 20840 => x"64206772",
    20841 => x"65617465", 20842 => x"72207468", 20843 => x"616e2063",
    20844 => x"6f6e6669", 20845 => x"67757265", 20846 => x"64206d61",
    20847 => x"78696d75", 20848 => x"6d202564", 20849 => x"0a000000",
    20850 => x"5472696d", 20851 => x"20746f6f", 20852 => x"2d6c6f6e",
    20853 => x"67206d70", 20854 => x"643a2025", 20855 => x"690a0000",
    20856 => x"41667465", 20857 => x"72206176", 20858 => x"67282569",
    20859 => x"292c206d", 20860 => x"65616e50", 20861 => x"61746844",
    20862 => x"656c6179", 20863 => x"3a202569", 20864 => x"0a000000",
    20865 => x"4f666673", 20866 => x"65742066", 20867 => x"726f6d20",
    20868 => x"6d617374", 20869 => x"65723a20", 20870 => x"20202020",
    20871 => x"25730a00", 20872 => x"73657276", 20873 => x"6f206162",
    20874 => x"6f727465", 20875 => x"642c206f", 20876 => x"66667365",
    20877 => x"74206772", 20878 => x"65617465", 20879 => x"72207468",
    20880 => x"616e2031", 20881 => x"20736563", 20882 => x"6f6e640a",
    20883 => x"00000000", 20884 => x"73657276", 20885 => x"6f206162",
    20886 => x"6f727465", 20887 => x"642c206f", 20888 => x"66667365",
    20889 => x"74206772", 20890 => x"65617465", 20891 => x"72207468",
    20892 => x"616e2063", 20893 => x"6f6e6669", 20894 => x"67757265",
    20895 => x"64206d61", 20896 => x"78696d75", 20897 => x"6d202564",
    20898 => x"0a000000", 20899 => x"4f627365", 20900 => x"72766564",
    20901 => x"20647269", 20902 => x"66743a20", 20903 => x"2539690a",
    20904 => x"00000000", 20905 => x"74696d65", 20906 => x"6f757420",
    20907 => x"65787069", 20908 => x"7265643a", 20909 => x"2025730a",
    20910 => x"00000000", 20911 => x"50505f54", 20912 => x"4f5f4445",
    20913 => x"4c415952", 20914 => x"45510000", 20915 => x"50505f54",
    20916 => x"4f5f5359", 20917 => x"4e430000", 20918 => x"50505f54",
    20919 => x"4f5f414e", 20920 => x"4e5f5245", 20921 => x"43454950",
    20922 => x"54000000", 20923 => x"50505f54", 20924 => x"4f5f414e",
    20925 => x"4e5f494e", 20926 => x"54455256", 20927 => x"414c0000",
    20928 => x"50505f54", 20929 => x"4f5f4641", 20930 => x"554c5459",
    20931 => x"00000000", 20932 => x"50505f54", 20933 => x"4f5f4558",
    20934 => x"545f3000", 20935 => x"50505f54", 20936 => x"4f5f4558",
    20937 => x"545f3100", 20938 => x"50505f54", 20939 => x"4f5f4558",
    20940 => x"545f3200", 20941 => x"536c6176", 20942 => x"65204f6e",
    20943 => x"6c792c20", 20944 => x"636c6f63", 20945 => x"6b20636c",
    20946 => x"61737320", 20947 => x"73657420", 20948 => x"746f2032",
    20949 => x"35350a00", 20950 => x"25750000", 20951 => x"25752575",
    20952 => x"00000000", 20953 => x"6c6e6b3a", 20954 => x"25642072",
    20955 => x"783a2564", 20956 => x"2074783a", 20957 => x"25642000",
    20958 => x"6c6f636b", 20959 => x"3a256420", 20960 => x"00000000",
    20961 => x"7074703a", 20962 => x"25732000", 20963 => x"73763a25",
    20964 => x"64200000", 20965 => x"73733a27", 20966 => x"25732720",
    20967 => x"00000000", 20968 => x"6175783a", 20969 => x"25782000",
    20970 => x"7365633a", 20971 => x"2564206e", 20972 => x"7365633a",
    20973 => x"25642000", 20974 => x"6d753a25", 20975 => x"73200000",
    20976 => x"646d733a", 20977 => x"25732000", 20978 => x"6474786d",
    20979 => x"3a256420", 20980 => x"6472786d", 20981 => x"3a256420",
    20982 => x"00000000", 20983 => x"64747873", 20984 => x"3a256420",
    20985 => x"64727873", 20986 => x"3a256420", 20987 => x"00000000",
    20988 => x"6173796d", 20989 => x"3a256420", 20990 => x"00000000",
    20991 => x"63727474", 20992 => x"3a257320", 20993 => x"00000000",
    20994 => x"636b6f3a", 20995 => x"25642000", 20996 => x"73657470",
    20997 => x"3a256420", 20998 => x"00000000", 20999 => x"75636e74",
    21000 => x"3a256420", 21001 => x"00000000", 21002 => x"68643a25",
    21003 => x"64206d64", 21004 => x"3a256420", 21005 => x"61643a25",
    21006 => x"64200000", 21007 => x"70636200", 21008 => x"74656d70",
    21009 => x"3a202564", 21010 => x"2e253034", 21011 => x"64204300",
    21012 => x"0a0a5054", 21013 => x"50207374", 21014 => x"61747573",
    21015 => x"3a200000", 21016 => x"25730000", 21017 => x"0a0a5379",
    21018 => x"6e632069", 21019 => x"6e666f20", 21020 => x"6e6f7420",
    21021 => x"76616c69", 21022 => x"640a0a00", 21023 => x"0a0a5379",
    21024 => x"6e636872", 21025 => x"6f6e697a", 21026 => x"6174696f",
    21027 => x"6e207374", 21028 => x"61747573", 21029 => x"3a0a0a00",
    21030 => x"57522050", 21031 => x"54502043", 21032 => x"6f726520",
    21033 => x"53796e63", 21034 => x"204d6f6e", 21035 => x"69746f72",
    21036 => x"20762031", 21037 => x"2e300000", 21038 => x"45736320",
    21039 => x"3d206578", 21040 => x"69740000", 21041 => x"0a0a5441",
    21042 => x"49205469", 21043 => x"6d653a20", 21044 => x"20202020",
    21045 => x"20202020", 21046 => x"20202020", 21047 => x"20202020",
    21048 => x"20000000", 21049 => x"0a0a4c69", 21050 => x"6e6b2073",
    21051 => x"74617475", 21052 => x"733a0000", 21053 => x"25733a20",
    21054 => x"00000000", 21055 => x"77727531", 21056 => x"00000000",
    21057 => x"4c696e6b", 21058 => x"20757020", 21059 => x"20200000",
    21060 => x"4c696e6b", 21061 => x"20646f77", 21062 => x"6e200000",
    21063 => x"2852583a", 21064 => x"2025642c", 21065 => x"2054583a",
    21066 => x"20256429", 21067 => x"2c206d6f", 21068 => x"64653a20",
    21069 => x"00000000", 21070 => x"5752204f", 21071 => x"66660000",
    21072 => x"436c6f63", 21073 => x"6b206f66", 21074 => x"66736574",
    21075 => x"3a202020", 21076 => x"20202020", 21077 => x"20202020",
    21078 => x"20202020", 21079 => x"20200000", 21080 => x"2532692e",
    21081 => x"25303969", 21082 => x"20730000", 21083 => x"25396920",
    21084 => x"6e730000", 21085 => x"0a4f6e65", 21086 => x"2d776179",
    21087 => x"2064656c", 21088 => x"61792061", 21089 => x"76657261",
    21090 => x"6765643a", 21091 => x"20202020", 21092 => x"20202000",
    21093 => x"0a4f6273", 21094 => x"65727665", 21095 => x"64206472",
    21096 => x"6966743a", 21097 => x"20202020", 21098 => x"20202020",
    21099 => x"20202020", 21100 => x"20202000", 21101 => x"5752204d",
    21102 => x"61737465", 21103 => x"72202000", 21104 => x"57522053",
    21105 => x"6c617665", 21106 => x"20202000", 21107 => x"57522055",
    21108 => x"6e6b6e6f", 21109 => x"776e2020", 21110 => x"20000000",
    21111 => x"4c6f636b", 21112 => x"65642020", 21113 => x"00000000",
    21114 => x"4e6f4c6f", 21115 => x"636b2020", 21116 => x"00000000",
    21117 => x"43616c69", 21118 => x"62726174", 21119 => x"65642020",
    21120 => x"00000000", 21121 => x"556e6361", 21122 => x"6c696272",
    21123 => x"61746564", 21124 => x"20200000", 21125 => x"0a495076",
    21126 => x"343a2000", 21127 => x"424f4f54", 21128 => x"50207275",
    21129 => x"6e6e696e", 21130 => x"67000000", 21131 => x"25732028",
    21132 => x"66726f6d", 21133 => x"20626f6f", 21134 => x"74702900",
    21135 => x"25732028", 21136 => x"73746174", 21137 => x"69632061",
    21138 => x"73736967", 21139 => x"6e6d656e", 21140 => x"74290000",
    21141 => x"53657276", 21142 => x"6f207374", 21143 => x"6174653a",
    21144 => x"20202020", 21145 => x"20202020", 21146 => x"20202020",
    21147 => x"20202000", 21148 => x"50686173", 21149 => x"65207472",
    21150 => x"61636b69", 21151 => x"6e673a20", 21152 => x"20202020",
    21153 => x"20202020", 21154 => x"20202000", 21155 => x"4f4e0a00",
    21156 => x"4f46460a", 21157 => x"00000000", 21158 => x"41757820",
    21159 => x"636c6f63", 21160 => x"6b207374", 21161 => x"61747573",
    21162 => x"3a202020", 21163 => x"20202020", 21164 => x"20202000",
    21165 => x"656e6162", 21166 => x"6c656400", 21167 => x"2c206c6f",
    21168 => x"636b6564", 21169 => x"00000000", 21170 => x"0a54696d",
    21171 => x"696e6720", 21172 => x"70617261", 21173 => x"6d657465",
    21174 => x"72733a0a", 21175 => x"0a000000", 21176 => x"526f756e",
    21177 => x"642d7472", 21178 => x"69702074", 21179 => x"696d6520",
    21180 => x"286d7529", 21181 => x"3a202020", 21182 => x"20000000",
    21183 => x"25732070", 21184 => x"730a0000", 21185 => x"4d617374",
    21186 => x"65722d73", 21187 => x"6c617665", 21188 => x"2064656c",
    21189 => x"61793a20", 21190 => x"20202020", 21191 => x"20000000",
    21192 => x"4d617374", 21193 => x"65722050", 21194 => x"48592064",
    21195 => x"656c6179", 21196 => x"733a2020", 21197 => x"20202020",
    21198 => x"20000000", 21199 => x"54583a20", 21200 => x"25642070",
    21201 => x"732c2052", 21202 => x"583a2025", 21203 => x"64207073",
    21204 => x"0a000000", 21205 => x"536c6176", 21206 => x"65205048",
    21207 => x"59206465", 21208 => x"6c617973", 21209 => x"3a202020",
    21210 => x"20202020", 21211 => x"20000000", 21212 => x"546f7461",
    21213 => x"6c206c69", 21214 => x"6e6b2061", 21215 => x"73796d6d",
    21216 => x"65747279", 21217 => x"3a202020", 21218 => x"20000000",
    21219 => x"25396420", 21220 => x"70730a00", 21221 => x"4361626c",
    21222 => x"65207274", 21223 => x"74206465", 21224 => x"6c61793a",
    21225 => x"20202020", 21226 => x"20202020", 21227 => x"20000000",
    21228 => x"436c6f63", 21229 => x"6b206f66", 21230 => x"66736574",
    21231 => x"3a202020", 21232 => x"20202020", 21233 => x"20202020",
    21234 => x"20000000", 21235 => x"50686173", 21236 => x"65207365",
    21237 => x"74706f69", 21238 => x"6e743a20", 21239 => x"20202020",
    21240 => x"20202020", 21241 => x"20000000", 21242 => x"536b6577",
    21243 => x"3a202020", 21244 => x"20202020", 21245 => x"20202020",
    21246 => x"20202020", 21247 => x"20202020", 21248 => x"20000000",
    21249 => x"55706461", 21250 => x"74652063", 21251 => x"6f756e74",
    21252 => x"65723a20", 21253 => x"20202020", 21254 => x"20202020",
    21255 => x"20000000", 21256 => x"2539640a", 21257 => x"00000000",
    21258 => x"2d2d0000", 21259 => x"756e6b6e", 21260 => x"6f776e00",
    21261 => x"73746174", 21262 => x"73000000", 21263 => x"1b5b3125",
    21264 => x"63000000", 21265 => x"436f6d6d", 21266 => x"616e6420",
    21267 => x"22257322", 21268 => x"3a206572", 21269 => x"726f7220",
    21270 => x"25640a00", 21271 => x"556e7265", 21272 => x"636f676e",
    21273 => x"697a6564", 21274 => x"20636f6d", 21275 => x"6d616e64",
    21276 => x"20222573", 21277 => x"222e0a00", 21278 => x"77726323",
    21279 => x"20000000", 21280 => x"25630000", 21281 => x"456d7074",
    21282 => x"7920696e", 21283 => x"69742073", 21284 => x"63726970",
    21285 => x"742e2e2e", 21286 => x"0a000000", 21287 => x"65786563",
    21288 => x"7574696e", 21289 => x"673a2025", 21290 => x"730a0000",
    21291 => x"57522043", 21292 => x"6f726520", 21293 => x"6275696c",
    21294 => x"643a2025", 21295 => x"7325730a", 21296 => x"00000000",
    21297 => x"2028756e", 21298 => x"73757070", 21299 => x"6f727465",
    21300 => x"64206465", 21301 => x"76656c6f", 21302 => x"70657220",
    21303 => x"6275696c", 21304 => x"64290000", 21305 => x"4275696c",
    21306 => x"743a2025", 21307 => x"73202573", 21308 => x"20627920",
    21309 => x"25730a00", 21310 => x"4275696c", 21311 => x"7420666f",
    21312 => x"72202564", 21313 => x"206b4220", 21314 => x"52414d2c",
    21315 => x"20737461", 21316 => x"636b2069", 21317 => x"73202564",
    21318 => x"20627974", 21319 => x"65730a00", 21320 => x"5741524e",
    21321 => x"494e473a", 21322 => x"20686172", 21323 => x"64776172",
    21324 => x"65207361", 21325 => x"79732025", 21326 => x"696b4220",
    21327 => x"3c3d2052", 21328 => x"414d203c", 21329 => x"2025696b",
    21330 => x"420a0000", 21331 => x"76657200", 21332 => x"73746172",
    21333 => x"74000000", 21334 => x"73746f70", 21335 => x"00000000",
    21336 => x"676d0000", 21337 => x"6d6f6465", 21338 => x"00000000",
    21339 => x"6772616e", 21340 => x"646d6173", 21341 => x"74657200",
    21342 => x"41766169", 21343 => x"6c61626c", 21344 => x"6520636f",
    21345 => x"6d6d616e", 21346 => x"64733a0a", 21347 => x"00000000",
    21348 => x"20202573", 21349 => x"0a000000", 21350 => x"68656c70",
    21351 => x"00000000", 21352 => x"25303278", 21353 => x"3a253032",
    21354 => x"783a2530", 21355 => x"32783a25", 21356 => x"3032783a",
    21357 => x"25303278", 21358 => x"3a253032", 21359 => x"78000000",
    21360 => x"67657400", 21361 => x"67657470", 21362 => x"00000000",
    21363 => x"73657400", 21364 => x"73657470", 21365 => x"00000000",
    21366 => x"4d41432d", 21367 => x"61646472", 21368 => x"6573733a",
    21369 => x"2025730a", 21370 => x"00000000", 21371 => x"6d616300",
    21372 => x"72657365", 21373 => x"74000000", 21374 => x"20697465",
    21375 => x"72617469", 21376 => x"6f6e7320", 21377 => x"20202020",
    21378 => x"7365636f", 21379 => x"6e64732e", 21380 => x"6d696372",
    21381 => x"6f732020", 21382 => x"20206e61", 21383 => x"6d650a00",
    21384 => x"20202539", 21385 => x"6c692020", 21386 => x"2025396c",
    21387 => x"692e2530", 21388 => x"366c6920", 21389 => x"2025730a",
    21390 => x"00000000", 21391 => x"70730000", 21392 => x"55736167",
    21393 => x"653a2072", 21394 => x"65667265", 21395 => x"7368203c",
    21396 => x"7365636f", 21397 => x"6e64733e", 21398 => x"0a000000",
    21399 => x"72656672", 21400 => x"65736800", 21401 => x"73746174",
    21402 => x"69737469", 21403 => x"6373206e", 21404 => x"6f77206f",
    21405 => x"66660a00", 21406 => x"62747300", 21407 => x"6f666600",
    21408 => x"73746174", 21409 => x"00000000", 21410 => x"57726f6e",
    21411 => x"67207061", 21412 => x"72616d65", 21413 => x"7465720a",
    21414 => x"00000000", 21415 => x"65726173", 21416 => x"65000000",
    21417 => x"436f756c", 21418 => x"64206e6f", 21419 => x"74206572",
    21420 => x"61736520", 21421 => x"44420a00", 21422 => x"61646400",
    21423 => x"53465020", 21424 => x"44422069", 21425 => x"73206675",
    21426 => x"6c6c0a00", 21427 => x"49324320", 21428 => x"6572726f",
    21429 => x"720a0000", 21430 => x"53465020", 21431 => x"64617461",
    21432 => x"62617365", 21433 => x"20657272", 21434 => x"6f722028",
    21435 => x"2564290a", 21436 => x"00000000", 21437 => x"25642053",
    21438 => x"46507320", 21439 => x"696e2044", 21440 => x"420a0000",
    21441 => x"73686f77", 21442 => x"00000000", 21443 => x"53465020",
    21444 => x"64617461", 21445 => x"62617365", 21446 => x"20656d70",
    21447 => x"74790a00", 21448 => x"25643a20", 21449 => x"504e3a00",
    21450 => x"20645478", 21451 => x"3a202538", 21452 => x"64206452",
    21453 => x"783a2025", 21454 => x"38642061", 21455 => x"6c706861",
    21456 => x"3a202538", 21457 => x"640a0000", 21458 => x"6d617463",
    21459 => x"68000000", 21460 => x"4e6f2053", 21461 => x"46502e0a",
    21462 => x"00000000", 21463 => x"53465020", 21464 => x"72656164",
    21465 => x"20657272", 21466 => x"6f720a00", 21467 => x"436f756c",
    21468 => x"64206e6f", 21469 => x"74206d61", 21470 => x"74636820",
    21471 => x"746f2044", 21472 => x"420a0000", 21473 => x"53465020",
    21474 => x"6d617463", 21475 => x"6865642c", 21476 => x"20645478",
    21477 => x"3d256420", 21478 => x"6452783d", 21479 => x"25642061",
    21480 => x"6c706861", 21481 => x"3d25640a", 21482 => x"00000000",
    21483 => x"656e6100", 21484 => x"73667000", 21485 => x"696e6974",
    21486 => x"00000000", 21487 => x"636c0000", 21488 => x"73707300",
    21489 => x"67707300", 21490 => x"25642025", 21491 => x"640a0000",
    21492 => x"73646163", 21493 => x"00000000", 21494 => x"67646163",
    21495 => x"00000000", 21496 => x"63686563", 21497 => x"6b76636f",
    21498 => x"00000000", 21499 => x"706c6c00", 21500 => x"666f7263",
    21501 => x"65000000", 21502 => x"466f756e", 21503 => x"64207068",
    21504 => x"61736520", 21505 => x"7472616e", 21506 => x"73697469",
    21507 => x"6f6e2069", 21508 => x"6e204545", 21509 => x"50524f4d",
    21510 => x"3a202564", 21511 => x"70730a00", 21512 => x"4d656173",
    21513 => x"7572696e", 21514 => x"67207432", 21515 => x"2f743420",
    21516 => x"70686173", 21517 => x"65207472", 21518 => x"616e7369",
    21519 => x"74696f6e", 21520 => x"2e2e2e0a", 21521 => x"00000000",
    21522 => x"63616c69", 21523 => x"62726174", 21524 => x"696f6e00",
    21525 => x"73657473", 21526 => x"65630000", 21527 => x"7365746e",
    21528 => x"73656300", 21529 => x"72617700", 21530 => x"2573202b",
    21531 => x"2564206e", 21532 => x"616e6f73", 21533 => x"65636f6e",
    21534 => x"64732e0a", 21535 => x"00000000", 21536 => x"74696d65",
    21537 => x"00000000", 21538 => x"67756900", 21539 => x"73646200",
    21540 => x"4f4e0000", 21541 => x"4f464600", 21542 => x"656e6162",
    21543 => x"6c650000", 21544 => x"64697361", 21545 => x"626c6500",
    21546 => x"70686173", 21547 => x"65207472", 21548 => x"61636b69",
    21549 => x"6e672025", 21550 => x"730a0000", 21551 => x"70747261",
    21552 => x"636b0000", 21553 => x"25642e25", 21554 => x"642e2564",
    21555 => x"2e256400", 21556 => x"49502d61", 21557 => x"64647265",
    21558 => x"73733a20", 21559 => x"696e2074", 21560 => x"7261696e",
    21561 => x"696e670a", 21562 => x"00000000", 21563 => x"49502d61",
    21564 => x"64647265", 21565 => x"73733a20", 21566 => x"25732028",
    21567 => x"66726f6d", 21568 => x"20626f6f", 21569 => x"7470290a",
    21570 => x"00000000", 21571 => x"49502d61", 21572 => x"64647265",
    21573 => x"73733a20", 21574 => x"25732028", 21575 => x"73746174",
    21576 => x"69632061", 21577 => x"73736967", 21578 => x"6e6d656e",
    21579 => x"74290a00", 21580 => x"69700000", 21581 => x"50505349",
    21582 => x"20766572", 21583 => x"626f7369", 21584 => x"74793a20",
    21585 => x"2530386c", 21586 => x"780a0000", 21587 => x"76657262",
    21588 => x"6f736500", 21589 => x"436f756c", 21590 => x"64206e6f",
    21591 => x"74206572", 21592 => x"61736520", 21593 => x"696e6974",
    21594 => x"20736372", 21595 => x"6970740a", 21596 => x"00000000",
    21597 => x"436f756c", 21598 => x"64206e6f", 21599 => x"74206164",
    21600 => x"64207468", 21601 => x"6520636f", 21602 => x"6d6d616e",
    21603 => x"640a0000", 21604 => x"4f4b2e0a", 21605 => x"00000000",
    21606 => x"626f6f74", 21607 => x"00000000", 21608 => x"25732c20",
    21609 => x"25732025", 21610 => x"642c2025", 21611 => x"642c2025",
    21612 => x"3032643a", 21613 => x"25303264", 21614 => x"3a253032",
    21615 => x"64000000", 21616 => x"25732025", 21617 => x"32642025",
    21618 => x"3032643a", 21619 => x"25303264", 21620 => x"3a253032",
    21621 => x"64000000", 21622 => x"2534642d", 21623 => x"25303264",
    21624 => x"2d253032", 21625 => x"642d2530", 21626 => x"32643a25",
    21627 => x"3032643a", 21628 => x"25303264", 21629 => x"00000000",
    21630 => x"1b5b3025", 21631 => x"643b3325", 21632 => x"646d0000",
    21633 => x"1b5b6d00", 21634 => x"1b5b2564", 21635 => x"3b256466",
    21636 => x"00000000", 21637 => x"1b5b324a", 21638 => x"1b5b313b",
    21639 => x"31480000", 21640 => x"53756e00", 21641 => x"4d6f6e00",
    21642 => x"54756500", 21643 => x"57656400", 21644 => x"54687500",
    21645 => x"46726900", 21646 => x"53617400", 21647 => x"4a616e00",
    21648 => x"46656200", 21649 => x"4d617200", 21650 => x"41707200",
    21651 => x"4d617900", 21652 => x"4a756e00", 21653 => x"4a756c00",
    21654 => x"41756700", 21655 => x"53657000", 21656 => x"4f637400",
    21657 => x"4e6f7600", 21658 => x"44656300", 21659 => x"4c6f6f70",
    21660 => x"73207065", 21661 => x"72206a69", 21662 => x"6666793a",
    21663 => x"2025690a", 21664 => x"00000000", 21665 => x"25733a20",
    21666 => x"6e6f2073", 21667 => x"6f636b65", 21668 => x"7420736c",
    21669 => x"6f747320", 21670 => x"6c656674", 21671 => x"0a000000",
    21672 => x"77723000", 21673 => x"6e65742d", 21674 => x"62680000",
    21675 => x"69707634", 21676 => x"00000000", 21677 => x"61727000",
    21678 => x"44697363", 21679 => x"6f766572", 21680 => x"65642049",
    21681 => x"50206164", 21682 => x"64726573", 21683 => x"73202825",
    21684 => x"642e2564", 21685 => x"2e25642e", 21686 => x"25642921",
    21687 => x"0a000000", 21688 => x"534e4d50", 21689 => x"3a205346",
    21690 => x"50207570", 21691 => x"64617465", 21692 => x"6420696e",
    21693 => x"206d656d", 21694 => x"6f72792c", 21695 => x"20726573",
    21696 => x"74617274", 21697 => x"20505450", 21698 => x"0a000000",
    21699 => x"494e5641", 21700 => x"4c494400", 21701 => x"25642e25",
    21702 => x"30346400", 21703 => x"736e6d70", 21704 => x"00000000",
    21705 => x"4e6f7620", 21706 => x"33302032", 21707 => x"30313620",
    21708 => x"32303a35", 21709 => x"393a3538", 21710 => x"00000000",
    21711 => x"30313233", 21712 => x"34353637", 21713 => x"38396162",
    21714 => x"63646566", 21715 => x"00000000", 21716 => x"49443a20",
    21717 => x"25780a00", 21718 => x"6e6f2070", 21719 => x"66696c74",
    21720 => x"65722072", 21721 => x"756c652d", 21722 => x"73657421",
    21723 => x"0a000000", 21724 => x"7066696c", 21725 => x"7465723a",
    21726 => x"2077726f", 21727 => x"6e67206d", 21728 => x"61676963",
    21729 => x"206e756d", 21730 => x"62657220", 21731 => x"28676f74",
    21732 => x"20307825", 21733 => x"78290a00", 21734 => x"7066696c",
    21735 => x"7465723a", 21736 => x"2077726f", 21737 => x"6e672072",
    21738 => x"756c652d", 21739 => x"7365742c", 21740 => x"2063616e",
    21741 => x"27742061", 21742 => x"70706c79", 21743 => x"0a000000",
    21744 => x"696e7661", 21745 => x"6c696420", 21746 => x"64657363",
    21747 => x"72697074", 21748 => x"6f722040", 21749 => x"2578203d",
    21750 => x"2025780a", 21751 => x"00000000", 21752 => x"5761726e",
    21753 => x"696e673a", 21754 => x"20747820", 21755 => x"6e6f7420",
    21756 => x"7465726d", 21757 => x"696e6174", 21758 => x"65642069",
    21759 => x"6e66696e", 21760 => x"69746520", 21761 => x"6d63723d",
    21762 => x"30782578", 21763 => x"0a000000", 21764 => x"5761726e",
    21765 => x"696e673a", 21766 => x"20747820", 21767 => x"74696d65",
    21768 => x"7374616d", 21769 => x"70206e65", 21770 => x"76657220",
    21771 => x"62656361", 21772 => x"6d652061", 21773 => x"7661696c",
    21774 => x"61626c65", 21775 => x"0a000000", 21776 => x"64657620",
    21777 => x"20307825", 21778 => x"30386c78", 21779 => x"20402025",
    21780 => x"30366c78", 21781 => x"2c202573", 21782 => x"0a000000",
    21783 => x"66706761", 21784 => x"2d617265", 21785 => x"61000000",
    21786 => x"4572726f", 21787 => x"72202564", 21788 => x"20776869",
    21789 => x"6c652072", 21790 => x"65616469", 21791 => x"6e672074",
    21792 => x"32347020", 21793 => x"66726f6d", 21794 => x"2073746f",
    21795 => x"72616765", 21796 => x"0a000000", 21797 => x"74323470",
    21798 => x"20726561", 21799 => x"64206672", 21800 => x"6f6d2073",
    21801 => x"746f7261", 21802 => x"67653a20", 21803 => x"25642070",
    21804 => x"730a0000", 21805 => x"57616974", 21806 => x"696e6720",
    21807 => x"666f7220", 21808 => x"6c696e6b", 21809 => x"2e2e2e0a",
    21810 => x"00000000", 21811 => x"4c6f636b", 21812 => x"696e6720",
    21813 => x"504c4c2e", 21814 => x"2e2e0a00", 21815 => x"43616c69",
    21816 => x"62726174", 21817 => x"696e6720", 21818 => x"52582074",
    21819 => x"696d6573", 21820 => x"74616d70", 21821 => x"65722e2e",
    21822 => x"2e0a0000", 21823 => x"4661696c", 21824 => x"65640000",
    21825 => x"53756363", 21826 => x"65737300", 21827 => x"57726f74",
    21828 => x"65206e65", 21829 => x"77207432", 21830 => x"34702076",
    21831 => x"616c7565", 21832 => x"3a202564", 21833 => x"20707320",
    21834 => x"28257329", 21835 => x"0a000000", 21836 => x"20454e4f",
    21837 => x"53504300", 21838 => x"25732573", 21839 => x"3a000000",
    21840 => x"74656d70", 21841 => x"00000000", 21842 => x"74656d70",
    21843 => x"65726174", 21844 => x"75726500", 21845 => x"55706461",
    21846 => x"74652065", 21847 => x"78697374", 21848 => x"696e6720",
    21849 => x"53465020", 21850 => x"656e7472", 21851 => x"790a0000",
    21852 => x"41646469", 21853 => x"6e67206e", 21854 => x"65772053",
    21855 => x"46502065", 21856 => x"6e747279", 21857 => x"0a000000",
    21858 => x"43616e27", 21859 => x"74207361", 21860 => x"76652070",
    21861 => x"65727369", 21862 => x"7374656e", 21863 => x"74204d41",
    21864 => x"43206164", 21865 => x"64726573", 21866 => x"730a0000",
    21867 => x"25733a20", 21868 => x"5573696e", 21869 => x"67205731",
    21870 => x"20736572", 21871 => x"69616c20", 21872 => x"6e756d62",
    21873 => x"65720a00", 21874 => x"6f666673", 21875 => x"65742025",
    21876 => x"34692028", 21877 => x"30782530", 21878 => x"3378293a",
    21879 => x"20253369", 21880 => x"20283078", 21881 => x"25303278",
    21882 => x"290a0000", 21883 => x"77726974", 21884 => x"65283078",
    21885 => x"25782c20", 21886 => x"2569293a", 21887 => x"20726573",
    21888 => x"756c7420", 21889 => x"3d202569", 21890 => x"0a000000",
    21891 => x"72656164", 21892 => x"28307825", 21893 => x"782c2025",
    21894 => x"69293a20", 21895 => x"72657375", 21896 => x"6c74203d",
    21897 => x"2025690a", 21898 => x"00000000", 21899 => x"64657669",
    21900 => x"63652025", 21901 => x"693a2025", 21902 => x"30387825",
    21903 => x"3038780a", 21904 => x"00000000", 21905 => x"74656d70",
    21906 => x"3a202564", 21907 => x"2e253034", 21908 => x"640a0000",
    21909 => x"77310000", 21910 => x"77317200", 21911 => x"77317700",
    21912 => x"3c756e6b", 21913 => x"6e6f776e", 21914 => x"3e000000",
    21915 => x"736f6674", 21916 => x"706c6c3a", 21917 => x"20697271",
    21918 => x"73202564", 21919 => x"20736571", 21920 => x"20257320",
    21921 => x"6d6f6465", 21922 => x"20256420", 21923 => x"616c6967",
    21924 => x"6e6d656e", 21925 => x"745f7374", 21926 => x"61746520",
    21927 => x"25642048", 21928 => x"4c256420", 21929 => x"4d4c2564",
    21930 => x"2048593d", 21931 => x"2564204d", 21932 => x"593d2564",
    21933 => x"2044656c", 21934 => x"436e743d", 21935 => x"25640a00",
    21936 => x"73746172", 21937 => x"742d6578", 21938 => x"74000000",
    21939 => x"77616974", 21940 => x"2d657874", 21941 => x"00000000",
    21942 => x"73746172", 21943 => x"742d6865", 21944 => x"6c706572",
    21945 => x"00000000", 21946 => x"77616974", 21947 => x"2d68656c",
    21948 => x"70657200", 21949 => x"73746172", 21950 => x"742d6d61",
    21951 => x"696e0000", 21952 => x"77616974", 21953 => x"2d6d6169",
    21954 => x"6e000000", 21955 => x"72656164", 21956 => x"79000000",
    21957 => x"636c6561", 21958 => x"722d6461", 21959 => x"63730000",
    21960 => x"77616974", 21961 => x"2d636c65", 21962 => x"61722d64",
    21963 => x"61637300", 21964 => x"53746163", 21965 => x"6b206f76",
    21966 => x"6572666c", 21967 => x"6f77210a", 21968 => x"00000000",
    21969 => x"badc0ffe", 21970 => x"3b9aca00", 21971 => x"000f4240",
    21972 => x"00080030", 21973 => x"d4a51000", 21974 => x"3b9ac9ff",
    21975 => x"c4653600", 21976 => x"7ffffffe", 21977 => x"80000001",
    21978 => x"fff06000", 21979 => x"0007d000", 21980 => x"41c64e6d",
    21981 => x"00010043", 21982 => x"00010044", 21983 => x"00015180",
    21984 => x"83aa7e80", 21985 => x"7fffffff", 21986 => x"00062000",
    21987 => x"005ee000", 21988 => x"01000001", 21989 => x"11223344",
    21990 => x"e0001fff", 21991 => x"111ee000", 21992 => x"01554000",
    21993 => x"0fffffff", 21994 => x"059682f0", 21995 => x"0ee6b27f",
    21996 => x"c0a80001", 21997 => x"4b002f40", 21998 => x"01312d02",
    21999 => x"01312d0a", 22000 => x"003d0137", 22001 => x"8000001f",
    22002 => x"009895b6", 22003 => x"c4000001", 22004 => x"000186a0",
    22005 => x"00ffffff", 22006 => x"fffdb610", 22007 => x"000249f0",
    22008 => x"05f5e100", 22009 => x"0bebc200", 22010 => x"fa0a1f00",
    22011 => x"01312d03", 22012 => x"5344422d", 22013 => x"011b1900",
    22014 => x"00000000", 22015 => x"70705f64", 22016 => x"6961675f",
    22017 => x"70617273", 22018 => x"65000000", 22019 => x"00000000",
    22020 => x"00013634", 22021 => x"00013640", 22022 => x"00013650",
    22023 => x"0001365c", 22024 => x"00013668", 22025 => x"00013674",
    22026 => x"00013680", 22027 => x"000014dc", 22028 => x"0000154c",
    22029 => x"00001804", 22030 => x"00001804", 22031 => x"00001804",
    22032 => x"00001804", 22033 => x"00001804", 22034 => x"00001804",
    22035 => x"000015c8", 22036 => x"00001638", 22037 => x"00001804",
    22038 => x"000016cc", 22039 => x"000017d8", 22040 => x"77727063",
    22041 => x"5f74696d", 22042 => x"655f6164", 22043 => x"6a757374",
    22044 => x"5f6f6666", 22045 => x"73657400", 22046 => x"77727063",
    22047 => x"5f74696d", 22048 => x"655f6164", 22049 => x"6a757374",
    22050 => x"00000000", 22051 => x"77727063", 22052 => x"5f74696d",
    22053 => x"655f7365", 22054 => x"74000000", 22055 => x"77727063",
    22056 => x"5f74696d", 22057 => x"655f6765", 22058 => x"74000000",
    22059 => x"77727063", 22060 => x"5f6e6574", 22061 => x"5f73656e",
    22062 => x"64000000", 22063 => x"77725f75", 22064 => x"6e706163",
    22065 => x"6b5f616e", 22066 => x"6e6f756e", 22067 => x"63650000",
    22068 => x"77725f70", 22069 => x"61636b5f", 22070 => x"616e6e6f",
    22071 => x"756e6365", 22072 => x"00000000", 22073 => x"77725f68",
    22074 => x"616e646c", 22075 => x"655f666f", 22076 => x"6c6c6f77",
    22077 => x"75700000", 22078 => x"77725f68", 22079 => x"616e646c",
    22080 => x"655f616e", 22081 => x"6e6f756e", 22082 => x"63650000",
    22083 => x"77725f65", 22084 => x"78656375", 22085 => x"74655f73",
    22086 => x"6c617665", 22087 => x"00000000", 22088 => x"77725f73",
    22089 => x"31000000", 22090 => x"77725f68", 22091 => x"616e646c",
    22092 => x"655f7265", 22093 => x"73700000", 22094 => x"77725f6e",
    22095 => x"65775f73", 22096 => x"6c617665", 22097 => x"00000000",
    22098 => x"77725f6d", 22099 => x"61737465", 22100 => x"725f6d73",
    22101 => x"67000000", 22102 => x"77725f6c", 22103 => x"69737465",
    22104 => x"6e696e67", 22105 => x"00000000", 22106 => x"77725f6f",
    22107 => x"70656e00", 22108 => x"77725f69", 22109 => x"6e697400",
    22110 => x"00002ddc", 22111 => x"00002e04", 22112 => x"00002e24",
    22113 => x"00002e94", 22114 => x"00002eb4", 22115 => x"00002ed0",
    22116 => x"00002ef0", 22117 => x"00002f7c", 22118 => x"00002f9c",
    22119 => x"77725f63", 22120 => x"616c6962", 22121 => x"72617469",
    22122 => x"6f6e0000", 22123 => x"00004420", 22124 => x"00004408",
    22125 => x"00004448", 22126 => x"00004554", 22127 => x"0000449c",
    22128 => x"00013f9c", 22129 => x"000140d0", 22130 => x"000140dc",
    22131 => x"000140e8", 22132 => x"000140f4", 22133 => x"00014100",
    22134 => x"77725f73", 22135 => x"6572766f", 22136 => x"5f757064",
    22137 => x"61746500", 22138 => x"70705f69", 22139 => x"6e697469",
    22140 => x"616c697a", 22141 => x"696e6700", 22142 => x"73745f63",
    22143 => x"6f6d5f73", 22144 => x"6c617665", 22145 => x"5f68616e",
    22146 => x"646c655f", 22147 => x"666f6c6c", 22148 => x"6f777570",
    22149 => x"00000000", 22150 => x"626d635f", 22151 => x"64617461",
    22152 => x"7365745f", 22153 => x"636d7000", 22154 => x"626d635f",
    22155 => x"73746174", 22156 => x"655f6465", 22157 => x"63697369",
    22158 => x"6f6e0000", 22159 => x"63466965", 22160 => x"6c645f74",
    22161 => x"6f5f5469", 22162 => x"6d65496e", 22163 => x"7465726e",
    22164 => x"616c0000", 22165 => x"00014c2c", 22166 => x"00014d6c",
    22167 => x"00014118", 22168 => x"00013c30", 22169 => x"0000001f",
    22170 => x"0000001c", 22171 => x"0000001f", 22172 => x"0000001e",
    22173 => x"0000001f", 22174 => x"0000001e", 22175 => x"0000001f",
    22176 => x"0000001f", 22177 => x"0000001e", 22178 => x"0000001f",
    22179 => x"0000001e", 22180 => x"0000001f", 22181 => x"0000001f",
    22182 => x"0000001d", 22183 => x"0000001f", 22184 => x"0000001e",
    22185 => x"0000001f", 22186 => x"0000001e", 22187 => x"0000001f",
    22188 => x"0000001f", 22189 => x"0000001e", 22190 => x"0000001f",
    22191 => x"0000001e", 22192 => x"0000001f", 22193 => x"00015220",
    22194 => x"00015224", 22195 => x"00015228", 22196 => x"0001522c",
    22197 => x"00015230", 22198 => x"00015234", 22199 => x"00015238",
    22200 => x"0001523c", 22201 => x"00015240", 22202 => x"00015244",
    22203 => x"00015248", 22204 => x"0001524c", 22205 => x"00015250",
    22206 => x"00015254", 22207 => x"00015258", 22208 => x"0001525c",
    22209 => x"00015260", 22210 => x"00015264", 22211 => x"00015268",
    22212 => x"70747064", 22213 => x"5f6e6574", 22214 => x"69665f63",
    22215 => x"72656174", 22216 => x"655f736f", 22217 => x"636b6574",
    22218 => x"00000000", 22219 => x"0000b614", 22220 => x"0000b624",
    22221 => x"0000b688", 22222 => x"0000b688", 22223 => x"0000b634",
    22224 => x"0000b688", 22225 => x"0000b688", 22226 => x"30ff0201",
    22227 => x"fa040670", 22228 => x"75626c69", 22229 => x"63fdff02",
    22230 => x"f90201fc", 22231 => x"0201fb30", 22232 => x"ff30ff06",
    22233 => x"6765745f", 22234 => x"70657273", 22235 => x"69737465",
    22236 => x"6e745f6d", 22237 => x"61630000", 22238 => x"000000c8",
    22239 => x"000039d0", 22240 => x"00010b34", 22241 => x"00010bb8",
    22242 => x"00010bf0", 22243 => x"00010c70", 22244 => x"00010cfc",
    22245 => x"00010d14", 22246 => x"00010c14", 22247 => x"00010b5c",
    22248 => x"00010ab8", 22249 => x"00010aec", 22250 => x"00000000",
    22251 => x"00000000", 22252 => x"00000000", 22253 => x"00000000",
    22254 => x"00000001", 22255 => x"00000001", 22256 => x"00000001",
    22257 => x"00000001", 22258 => x"00000000", 22259 => x"00000000",
    22260 => x"00000000", 22261 => x"0000ece8", 22262 => x"0000ece8",
    22263 => x"00000000", 22264 => x"0000d9d0", 22265 => x"00000000",
    22266 => x"00011878", 22267 => x"00011898", 22268 => x"000118a4",
    22269 => x"000118b4", 22270 => x"000118d4", 22271 => x"000118e4",
    22272 => x"00011938", 22273 => x"000118fc", 22274 => x"0001180c",
    22275 => x"00011850", 22276 => x"00000001", 22277 => x"000156c0",
    22278 => x"00000002", 22279 => x"000156cc", 22280 => x"00000003",
    22281 => x"000156d8", 22282 => x"00000004", 22283 => x"000156e8",
    22284 => x"00000005", 22285 => x"000156f4", 22286 => x"00000006",
    22287 => x"00015700", 22288 => x"00000007", 22289 => x"00013c08",
    22290 => x"00000008", 22291 => x"0001570c", 22292 => x"00000009",
    22293 => x"00015714", 22294 => x"0000000a", 22295 => x"00015720",
    22296 => x"00000000", 22297 => x"00000000", 22298 => x"00000000",
    22299 => x"00000000", 22300 => x"00000000", 22301 => x"00000000",
    22302 => x"00010000", 22303 => x"00000000", 22304 => x"00000000",
    22305 => x"00000000", 22306 => x"00020100", 22307 => x"00000000",
    22308 => x"00000000", 22309 => x"00000000", 22310 => x"00030101",
    22311 => x"00000000", 22312 => x"00000000", 22313 => x"00000000",
    22314 => x"00040201", 22315 => x"01000000", 22316 => x"00000000",
    22317 => x"00000000", 22318 => x"00050201", 22319 => x"01010000",
    22320 => x"00000000", 22321 => x"00000000", 22322 => x"00060302",
    22323 => x"01010100", 22324 => x"00000000", 22325 => x"00000000",
    22326 => x"00070302", 22327 => x"01010101", 22328 => x"00000000",
    22329 => x"00000000", 22330 => x"00080402", 22331 => x"02010101",
    22332 => x"01000000", 22333 => x"00000000", 22334 => x"00090403",
    22335 => x"02010101", 22336 => x"01010000", 22337 => x"00000000",
    22338 => x"000a0503", 22339 => x"02020101", 22340 => x"01010100",
    22341 => x"00000000", 22342 => x"000b0503", 22343 => x"02020101",
    22344 => x"01010101", 22345 => x"00000000", 22346 => x"000c0604",
    22347 => x"03020201", 22348 => x"01010101", 22349 => x"01000000",
    22350 => x"000d0604", 22351 => x"03020201", 22352 => x"01010101",
    22353 => x"01010000", 22354 => x"000e0704", 22355 => x"03020202",
    22356 => x"01010101", 22357 => x"01010100", 22358 => x"000f0705",
    22359 => x"03030202", 22360 => x"01010101", 22361 => x"01010101",
    22362 => x"fefefeff", 22363 => x"80808080", 22364 => x"00202020",
    22365 => x"20202020", 22366 => x"20202828", 22367 => x"28282820",
    22368 => x"20202020", 22369 => x"20202020", 22370 => x"20202020",
    22371 => x"20202020", 22372 => x"20881010", 22373 => x"10101010",
    22374 => x"10101010", 22375 => x"10101010", 22376 => x"10040404",
    22377 => x"04040404", 22378 => x"04040410", 22379 => x"10101010",
    22380 => x"10104141", 22381 => x"41414141", 22382 => x"01010101",
    22383 => x"01010101", 22384 => x"01010101", 22385 => x"01010101",
    22386 => x"01010101", 22387 => x"10101010", 22388 => x"10104242",
    22389 => x"42424242", 22390 => x"02020202", 22391 => x"02020202",
    22392 => x"02020202", 22393 => x"02020202", 22394 => x"02020202",
    22395 => x"10101010", 22396 => x"20000000", 22397 => x"00000000",
    22398 => x"00000000", 22399 => x"00000000", 22400 => x"00000000",
    22401 => x"00000000", 22402 => x"00000000", 22403 => x"00000000",
    22404 => x"00000000", 22405 => x"00000000", 22406 => x"00000000",
    22407 => x"00000000", 22408 => x"00000000", 22409 => x"00000000",
    22410 => x"00000000", 22411 => x"00000000", 22412 => x"00000000",
    22413 => x"00000000", 22414 => x"00000000", 22415 => x"00000000",
    22416 => x"00000000", 22417 => x"00000000", 22418 => x"00000000",
    22419 => x"00000000", 22420 => x"00000000", 22421 => x"00000000",
    22422 => x"00000000", 22423 => x"00000000", 22424 => x"00000000",
    22425 => x"00000000", 22426 => x"00000000", 22427 => x"00000000",
    22428 => x"00000000", 22429 => x"00000000", 22430 => x"00016ff8",
    22431 => x"00017018", 22432 => x"00017028", 22433 => x"00017038",
    22434 => x"000003e8", 22435 => x"00000001", 22436 => x"00000955",
    22437 => x"ffffffff", 22438 => x"00000000", 22439 => x"00000000",
    22440 => x"00000000", 22441 => x"00000000", 22442 => x"00000000",
    22443 => x"00000000", 22444 => x"00000000", 22445 => x"00000000",
    22446 => x"0001620c", 22447 => x"0001632c", 22448 => x"00016310",
    22449 => x"00017290", 22450 => x"00017310", 22451 => x"00000000",
    22452 => x"00000000", 22453 => x"00000000", 22454 => x"00000000",
    22455 => x"00000000", 22456 => x"00000000", 22457 => x"00000000",
    22458 => x"00000000", 22459 => x"00000000", 22460 => x"00000000",
    22461 => x"00000000", 22462 => x"00000000", 22463 => x"00000000",
    22464 => x"00000000", 22465 => x"00000000", 22466 => x"00000000",
    22467 => x"00000000", 22468 => x"00000000", 22469 => x"00000000",
    22470 => x"00000000", 22471 => x"00000000", 22472 => x"00000000",
    22473 => x"00000000", 22474 => x"00000000", 22475 => x"00000000",
    22476 => x"00000000", 22477 => x"00000000", 22478 => x"00000000",
    22479 => x"00000000", 22480 => x"00000000", 22481 => x"00000000",
    22482 => x"00000000", 22483 => x"00000000", 22484 => x"00000000",
    22485 => x"00000000", 22486 => x"00000000", 22487 => x"00000000",
    22488 => x"00000000", 22489 => x"00000000", 22490 => x"00000000",
    22491 => x"00000000", 22492 => x"00000000", 22493 => x"00000000",
    22494 => x"00000000", 22495 => x"00000000", 22496 => x"00000000",
    22497 => x"00000000", 22498 => x"00000000", 22499 => x"00000000",
    22500 => x"00000000", 22501 => x"00000000", 22502 => x"00000000",
    22503 => x"00000000", 22504 => x"00000000", 22505 => x"00000000",
    22506 => x"00000000", 22507 => x"00000000", 22508 => x"00000000",
    22509 => x"00000000", 22510 => x"00000000", 22511 => x"00000000",
    22512 => x"00000000", 22513 => x"00000000", 22514 => x"00000000",
    22515 => x"00000000", 22516 => x"00000000", 22517 => x"00000000",
    22518 => x"00000000", 22519 => x"00000000", 22520 => x"00000000",
    22521 => x"00000000", 22522 => x"00000000", 22523 => x"00000000",
    22524 => x"00000000", 22525 => x"00000000", 22526 => x"00000000",
    22527 => x"00000000", 22528 => x"00000000", 22529 => x"00000000",
    22530 => x"00000000", 22531 => x"00000000", 22532 => x"00000000",
    22533 => x"00000000", 22534 => x"00000000", 22535 => x"00000000",
    22536 => x"00000000", 22537 => x"00000000", 22538 => x"00000000",
    22539 => x"00000000", 22540 => x"00000000", 22541 => x"00000000",
    22542 => x"00000000", 22543 => x"00000000", 22544 => x"00000000",
    22545 => x"00000000", 22546 => x"00000000", 22547 => x"00000000",
    22548 => x"00000000", 22549 => x"00000000", 22550 => x"00000000",
    22551 => x"00000000", 22552 => x"00000000", 22553 => x"00000000",
    22554 => x"00000000", 22555 => x"00000000", 22556 => x"00000000",
    22557 => x"00000000", 22558 => x"00000000", 22559 => x"00000000",
    22560 => x"00000000", 22561 => x"00000000", 22562 => x"00000000",
    22563 => x"00000000", 22564 => x"00000000", 22565 => x"00000000",
    22566 => x"00000000", 22567 => x"00000000", 22568 => x"00000000",
    22569 => x"00000000", 22570 => x"00000000", 22571 => x"00000000",
    22572 => x"00000000", 22573 => x"00000000", 22574 => x"00000000",
    22575 => x"00000000", 22576 => x"00000000", 22577 => x"00000000",
    22578 => x"00000000", 22579 => x"00000000", 22580 => x"00000000",
    22581 => x"00000000", 22582 => x"00000000", 22583 => x"00000000",
    22584 => x"00000000", 22585 => x"00000000", 22586 => x"00000000",
    22587 => x"00000000", 22588 => x"00000000", 22589 => x"00000000",
    22590 => x"00000000", 22591 => x"00000000", 22592 => x"00000000",
    22593 => x"00000000", 22594 => x"00000000", 22595 => x"00000000",
    22596 => x"00000000", 22597 => x"00000000", 22598 => x"00000000",
    22599 => x"00000000", 22600 => x"00000000", 22601 => x"00000000",
    22602 => x"00000000", 22603 => x"00000000", 22604 => x"00000000",
    22605 => x"00000000", 22606 => x"00000000", 22607 => x"00000000",
    22608 => x"00000000", 22609 => x"00000000", 22610 => x"00000000",
    22611 => x"00000000", 22612 => x"00000000", 22613 => x"00000000",
    22614 => x"00000000", 22615 => x"00000000", 22616 => x"00016254",
    22617 => x"00000000", 22618 => x"00000000", 22619 => x"00000000",
    22620 => x"00000000", 22621 => x"00000000", 22622 => x"00000000",
    22623 => x"00000000", 22624 => x"00000000", 22625 => x"00000000",
    22626 => x"00000000", 22627 => x"00000000", 22628 => x"00000000",
    22629 => x"00000000", 22630 => x"00000000", 22631 => x"00000000",
    22632 => x"00000000", 22633 => x"00000000", 22634 => x"00000000",
    22635 => x"00000000", 22636 => x"00000000", 22637 => x"00000000",
    22638 => x"00000000", 22639 => x"00000000", 22640 => x"00000000",
    22641 => x"00000000", 22642 => x"00013710", 22643 => x"00013710",
    22644 => x"00000000", 22645 => x"00000001", 22646 => x"00000000",
    22647 => x"00000000", 22648 => x"00000000", 22649 => x"00000000",
    22650 => x"00000000", 22651 => x"00000000", 22652 => x"00000000",
    22653 => x"00000000", 22654 => x"00000000", 22655 => x"00000000",
    22656 => x"00000000", 22657 => x"00000000", 22658 => x"00000000",
    22659 => x"00015e98", 22660 => x"00017390", 22661 => x"00000000",
    22662 => x"000173d0", 22663 => x"000173ec", 22664 => x"0001741c",
    22665 => x"0001743c", 22666 => x"00000000", 22667 => x"00000000",
    22668 => x"00000000", 22669 => x"00000000", 22670 => x"00000000",
    22671 => x"00000000", 22672 => x"00000000", 22673 => x"00000000",
    22674 => x"00000000", 22675 => x"00017460", 22676 => x"000003e8",
    22677 => x"00000000", 22678 => x"00000000", 22679 => x"00000000",
    22680 => x"00000000", 22681 => x"00016268", 22682 => x"000162d4",
    22683 => x"00000000", 22684 => x"00000000", 22685 => x"00000000",
    22686 => x"00000000", 22687 => x"00000000", 22688 => x"00000000",
    22689 => x"00000000", 22690 => x"00000000", 22691 => x"00000000",
    22692 => x"00000000", 22693 => x"00000000", 22694 => x"00000000",
    22695 => x"00000000", 22696 => x"00000000", 22697 => x"00000000",
    22698 => x"00000000", 22699 => x"00000000", 22700 => x"00000000",
    22701 => x"00000000", 22702 => x"00000000", 22703 => x"00000000",
    22704 => x"00000000", 22705 => x"00000000", 22706 => x"00000000",
    22707 => x"00000000", 22708 => x"00000000", 22709 => x"00000a58",
    22710 => x"00000a8c", 22711 => x"00000b0c", 22712 => x"00000b14",
    22713 => x"00000b6c", 22714 => x"00000b98", 22715 => x"00000bf0",
    22716 => x"00000c14", 22717 => x"00000cd8", 22718 => x"00000ce0",
    22719 => x"00000ce8", 22720 => x"00000d4c", 22721 => x"00000d68",
    22722 => x"00000b38", 22723 => x"00000000", 22724 => x"00001c8c",
    22725 => x"00001c10", 22726 => x"00001bb4", 22727 => x"00001b5c",
    22728 => x"00000000", 22729 => x"00000000", 22730 => x"00001b2c",
    22731 => x"00001f18", 22732 => x"00001ef8", 22733 => x"00001e28",
    22734 => x"00001d0c", 22735 => x"00000000", 22736 => x"00000000",
    22737 => x"00000000", 22738 => x"00000000", 22739 => x"00000000",
    22740 => x"00000000", 22741 => x"00000000", 22742 => x"00000000",
    22743 => x"00000000", 22744 => x"00000000", 22745 => x"00000000",
    22746 => x"00000200", 22747 => x"00000000", 22748 => x"00017570",
    22749 => x"00000001", 22750 => x"00013bf0", 22751 => x"00004748",
    22752 => x"00000002", 22753 => x"00013c00", 22754 => x"00004914",
    22755 => x"00000003", 22756 => x"00013c08", 22757 => x"000049d0",
    22758 => x"00000004", 22759 => x"00013c14", 22760 => x"000049e0",
    22761 => x"00000006", 22762 => x"00014118", 22763 => x"00004b8c",
    22764 => x"00000008", 22765 => x"00013c20", 22766 => x"00004ecc",
    22767 => x"00000009", 22768 => x"00013c30", 22769 => x"00004f40",
    22770 => x"00000064", 22771 => x"00013c38", 22772 => x"00002814",
    22773 => x"00000066", 22774 => x"00013c50", 22775 => x"0000298c",
    22776 => x"00000065", 22777 => x"00013c64", 22778 => x"00002ab8",
    22779 => x"00000067", 22780 => x"00013c7c", 22781 => x"00002bbc",
    22782 => x"00000068", 22783 => x"00013c94", 22784 => x"00002ce8",
    22785 => x"00000069", 22786 => x"00013ca4", 22787 => x"00003004",
    22788 => x"0000006a", 22789 => x"00013cb4", 22790 => x"00003118",
    22791 => x"0000006b", 22792 => x"00013cc8", 22793 => x"0000329c",
    22794 => x"00000000", 22795 => x"00000000", 22796 => x"00000000",
    22797 => x"00000001", 22798 => x"00013bf0", 22799 => x"00004748",
    22800 => x"00000002", 22801 => x"00013c00", 22802 => x"00004914",
    22803 => x"00000003", 22804 => x"00013c08", 22805 => x"000049d0",
    22806 => x"00000004", 22807 => x"00013c14", 22808 => x"000049e0",
    22809 => x"00000005", 22810 => x"00014114", 22811 => x"00004af8",
    22812 => x"00000006", 22813 => x"00014118", 22814 => x"00004b8c",
    22815 => x"00000007", 22816 => x"00014120", 22817 => x"00004e08",
    22818 => x"00000008", 22819 => x"00013c20", 22820 => x"00004ecc",
    22821 => x"00000009", 22822 => x"00013c30", 22823 => x"00004f40",
    22824 => x"00000000", 22825 => x"00000000", 22826 => x"00000000",
    22827 => x"00002218", 22828 => x"00002138", 22829 => x"00000000",
    22830 => x"000020f0", 22831 => x"000025b0", 22832 => x"00002568",
    22833 => x"0000247c", 22834 => x"00002060", 22835 => x"00001fd4",
    22836 => x"00002404", 22837 => x"0000238c", 22838 => x"00002324",
    22839 => x"000022b8", 22840 => x"00000001", 22841 => x"0001432c",
    22842 => x"00014334", 22843 => x"00014340", 22844 => x"0001434c",
    22845 => x"00000000", 22846 => x"00000000", 22847 => x"00000000",
    22848 => x"00000000", 22849 => x"00014370", 22850 => x"00014358",
    22851 => x"00014364", 22852 => x"0001437c", 22853 => x"00014388",
    22854 => x"00014394", 22855 => x"00000000", 22856 => x"00000000",
    22857 => x"000146bc", 22858 => x"000146cc", 22859 => x"000146d8",
    22860 => x"000146ec", 22861 => x"00014700", 22862 => x"00014710",
    22863 => x"0001471c", 22864 => x"00014728", 22865 => x"bbfef060",
    22866 => x"00000000", 22867 => x"00000000", 22868 => x"00000000",
    22869 => x"00000000", 22870 => x"00000000", 22871 => x"00000000",
    22872 => x"00000000", 22873 => x"00000000", 22874 => x"00000000",
    22875 => x"00000000", 22876 => x"00000000", 22877 => x"00000000",
    22878 => x"00000001", 22879 => x"00000000", 22880 => x"000a03e8",
    22881 => x"00060100", 22882 => x"80800000", 22883 => x"00000000",
    22884 => x"00015e98", 22885 => x"00000000", 22886 => x"00000000",
    22887 => x"00000000", 22888 => x"00000000", 22889 => x"00000000",
    22890 => x"00000000", 22891 => x"00000000", 22892 => x"00000000",
    22893 => x"00000000", 22894 => x"00000000", 22895 => x"00000200",
    22896 => x"00000000", 22897 => x"00017a9c", 22898 => x"00000000",
    22899 => x"00000000", 22900 => x"00000000", 22901 => x"00000000",
    22902 => x"00000000", 22903 => x"00000000", 22904 => x"00000000",
    22905 => x"00000000", 22906 => x"00000000", 22907 => x"00000000",
    22908 => x"00000060", 22909 => x"00000000", 22910 => x"00017c9c",
    22911 => x"00000000", 22912 => x"00000000", 22913 => x"00000000",
    22914 => x"00000000", 22915 => x"00000000", 22916 => x"00000000",
    22917 => x"00000000", 22918 => x"00000000", 22919 => x"00000000",
    22920 => x"00000000", 22921 => x"00000080", 22922 => x"00000000",
    22923 => x"00017cfc", 22924 => x"00000000", 22925 => x"00000000",
    22926 => x"00000000", 22927 => x"00000000", 22928 => x"00000000",
    22929 => x"00000000", 22930 => x"00000000", 22931 => x"00000000",
    22932 => x"00000000", 22933 => x"00000000", 22934 => x"00000080",
    22935 => x"00000000", 22936 => x"00017d80", 22937 => x"63757465",
    22938 => x"00000000", 22939 => x"00000000", 22940 => x"00000000",
    22941 => x"00000000", 22942 => x"00000000", 22943 => x"00000000",
    22944 => x"00000000", 22945 => x"00016748", 22946 => x"0000bb64",
    22947 => x"00016754", 22948 => x"09000000", 22949 => x"000167b8",
    22950 => x"0000bb64", 22951 => x"000167c4", 22952 => x"09000000",
    22953 => x"00016814", 22954 => x"0000b954", 22955 => x"00016820",
    22956 => x"0a000000", 22957 => x"0001685c", 22958 => x"0000bb64",
    22959 => x"00016868", 22960 => x"09000000", 22961 => x"00016930",
    22962 => x"0000bb64", 22963 => x"0001693c", 22964 => x"09000000",
    22965 => x"00016aa4", 22966 => x"0000bb64", 22967 => x"00016ab0",
    22968 => x"09000000", 22969 => x"00016b3c", 22970 => x"0000bb64",
    22971 => x"00016b48", 22972 => x"09000000", 22973 => x"00016bc0",
    22974 => x"0000b954", 22975 => x"00016bcc", 22976 => x"0a000000",
    22977 => x"00000000", 22978 => x"00000000", 22979 => x"00000000",
    22980 => x"00000000", 22981 => x"00000000", 22982 => x"00000000",
    22983 => x"00000000", 22984 => x"00000000", 22985 => x"00000000",
    22986 => x"00000000", 22987 => x"00000000", 22988 => x"00000000",
    22989 => x"00000000", 22990 => x"00000000", 22991 => x"00000100",
    22992 => x"00000000", 22993 => x"00017e28", 22994 => x"2b060104",
    22995 => x"01606501", 22996 => x"01000000", 22997 => x"00016c30",
    22998 => x"0000c0e0", 22999 => x"00000000", 23000 => x"00016664",
    23001 => x"02040020", 23002 => x"00016c34", 23003 => x"0000c0b4",
    23004 => x"00000000", 23005 => x"00015e78", 23006 => x"02040004",
    23007 => x"00016c38", 23008 => x"0000c0b4", 23009 => x"00000000",
    23010 => x"00015e84", 23011 => x"02040004", 23012 => x"00016c3c",
    23013 => x"0000c0b4", 23014 => x"00000000", 23015 => x"00016c40",
    23016 => x"02040004", 23017 => x"00000000", 23018 => x"00000000",
    23019 => x"00000000", 23020 => x"00000000", 23021 => x"00000000",
    23022 => x"2b060104", 23023 => x"01606501", 23024 => x"02000000",
    23025 => x"00016c44", 23026 => x"0000c478", 23027 => x"00000000",
    23028 => x"00000004", 23029 => x"02460001", 23030 => x"00016c48",
    23031 => x"0000c478", 23032 => x"00000000", 23033 => x"00000005",
    23034 => x"02040001", 23035 => x"00016c4c", 23036 => x"0000c478",
    23037 => x"00000000", 23038 => x"00000002", 23039 => x"02430001",
    23040 => x"00000000", 23041 => x"00000000", 23042 => x"00000000",
    23043 => x"00000000", 23044 => x"00000000", 23045 => x"2b060104",
    23046 => x"01606501", 23047 => x"03010000", 23048 => x"00016c50",
    23049 => x"0000c348", 23050 => x"00000000", 23051 => x"00000000",
    23052 => x"01040001", 23053 => x"00016c54", 23054 => x"0000c348",
    23055 => x"00000000", 23056 => x"00000000", 23057 => x"01040001",
    23058 => x"00000000", 23059 => x"00000000", 23060 => x"00000000",
    23061 => x"00000000", 23062 => x"00000000", 23063 => x"2b060104",
    23064 => x"01606501", 23065 => x"04000000", 23066 => x"00016c58",
    23067 => x"0000c0e0", 23068 => x"00000000", 23069 => x"00016fd0",
    23070 => x"02020004", 23071 => x"00016c5c", 23072 => x"0000c0e0",
    23073 => x"00000000", 23074 => x"00016fd4", 23075 => x"02410004",
    23076 => x"00016c60", 23077 => x"0000c0e0", 23078 => x"00000000",
    23079 => x"00016fd8", 23080 => x"02020004", 23081 => x"00016c64",
    23082 => x"0000c0e0", 23083 => x"00000000", 23084 => x"00016fdc",
    23085 => x"02020004", 23086 => x"00016c68", 23087 => x"0000c0e0",
    23088 => x"00000000", 23089 => x"00016fe0", 23090 => x"02410004",
    23091 => x"00016c6c", 23092 => x"0000c0e0", 23093 => x"00000000",
    23094 => x"00016fe4", 23095 => x"02410004", 23096 => x"00016c70",
    23097 => x"0000c0e0", 23098 => x"00000000", 23099 => x"00016fe8",
    23100 => x"02020004", 23101 => x"00016c74", 23102 => x"0000c0e0",
    23103 => x"00000000", 23104 => x"00016fec", 23105 => x"02020004",
    23106 => x"00016c78", 23107 => x"0000c0e0", 23108 => x"00000000",
    23109 => x"00016ff0", 23110 => x"02410004", 23111 => x"00000000",
    23112 => x"00000000", 23113 => x"00000000", 23114 => x"00000000",
    23115 => x"00000000", 23116 => x"2b060104", 23117 => x"01606501",
    23118 => x"05000000", 23119 => x"00016c7c", 23120 => x"0000c0b4",
    23121 => x"00000000", 23122 => x"00017e04", 23123 => x"02021404",
    23124 => x"00016c80", 23125 => x"0000c028", 23126 => x"00000000",
    23127 => x"00017e04", 23128 => x"0202e808", 23129 => x"00016c84",
    23130 => x"0000c028", 23131 => x"00000000", 23132 => x"00017e04",
    23133 => x"0202e008", 23134 => x"00016c88", 23135 => x"0000c0b4",
    23136 => x"00000000", 23137 => x"00017e04", 23138 => x"0246a008",
    23139 => x"00016c8c", 23140 => x"0000c0b4", 23141 => x"00000000",
    23142 => x"00017e04", 23143 => x"0241b804", 23144 => x"00016c90",
    23145 => x"0000bf28", 23146 => x"00000000", 23147 => x"00000001",
    23148 => x"02460001", 23149 => x"00016c94", 23150 => x"0000c0b4",
    23151 => x"00000000", 23152 => x"00017e04", 23153 => x"02021804",
    23154 => x"00016c98", 23155 => x"0000c0b4", 23156 => x"00000000",
    23157 => x"00017e04", 23158 => x"02021c04", 23159 => x"00016c9c",
    23160 => x"0000c0b4", 23161 => x"00000000", 23162 => x"00017e04",
    23163 => x"02022004", 23164 => x"00016ca0", 23165 => x"0000c0b4",
    23166 => x"00000000", 23167 => x"00017e04", 23168 => x"02022404",
    23169 => x"00016ca4", 23170 => x"0000c0b4", 23171 => x"00000000",
    23172 => x"00017e04", 23173 => x"0241f004", 23174 => x"00016ca8",
    23175 => x"0000c0b4", 23176 => x"00000000", 23177 => x"00017e04",
    23178 => x"0241f404", 23179 => x"00016cac", 23180 => x"0000c0b4",
    23181 => x"00000000", 23182 => x"00017e04", 23183 => x"0241f804",
    23184 => x"00016cb0", 23185 => x"0000bf28", 23186 => x"00000000",
    23187 => x"00000002", 23188 => x"02460001", 23189 => x"00016cb4",
    23190 => x"0000c0e0", 23191 => x"00000000", 23192 => x"00016204",
    23193 => x"02410004", 23194 => x"00016cb8", 23195 => x"0000c0e0",
    23196 => x"00000000", 23197 => x"00016208", 23198 => x"02410004",
    23199 => x"00016cbc", 23200 => x"0000c0b4", 23201 => x"00000000",
    23202 => x"00017e04", 23203 => x"02022804", 23204 => x"00000000",
    23205 => x"00000000", 23206 => x"00000000", 23207 => x"00000000",
    23208 => x"00000000", 23209 => x"2b060104", 23210 => x"01606501",
    23211 => x"06000000", 23212 => x"00016cc0", 23213 => x"0000c0e0",
    23214 => x"0000c168", 23215 => x"00017f28", 23216 => x"02020004",
    23217 => x"00016cc4", 23218 => x"0000c0e0", 23219 => x"0000c1c8",
    23220 => x"00017f2c", 23221 => x"02020004", 23222 => x"00016cc8",
    23223 => x"0000c0e0", 23224 => x"0000b930", 23225 => x"00017e08",
    23226 => x"02040010", 23227 => x"00016ccc", 23228 => x"0000c0e0",
    23229 => x"0000b930", 23230 => x"00017e1c", 23231 => x"02020004",
    23232 => x"00016cd0", 23233 => x"0000c0e0", 23234 => x"0000b930",
    23235 => x"00017e20", 23236 => x"02020004", 23237 => x"00016cd4",
    23238 => x"0000c0e0", 23239 => x"0000b930", 23240 => x"00017e18",
    23241 => x"02020004", 23242 => x"00000000", 23243 => x"00000000",
    23244 => x"00000000", 23245 => x"00000000", 23246 => x"00000000",
    23247 => x"2b060104", 23248 => x"01606501", 23249 => x"07000000",
    23250 => x"00016cd8", 23251 => x"0000c108", 23252 => x"00000000",
    23253 => x"00000001", 23254 => x"02020001", 23255 => x"00016cdc",
    23256 => x"0000c0e0", 23257 => x"00000000", 23258 => x"00018c24",
    23259 => x"02040010", 23260 => x"00016ce0", 23261 => x"0000c0e0",
    23262 => x"00000000", 23263 => x"00018bc0", 23264 => x"02020004",
    23265 => x"00016ce4", 23266 => x"0000c0e0", 23267 => x"00000000",
    23268 => x"00018f6c", 23269 => x"02410004", 23270 => x"00016ce8",
    23271 => x"0000c0e0", 23272 => x"00000000", 23273 => x"00018f70",
    23274 => x"02410004", 23275 => x"00000000", 23276 => x"00000000",
    23277 => x"00000000", 23278 => x"00000000", 23279 => x"00000000",
    23280 => x"2b060104", 23281 => x"01606501", 23282 => x"08010000",
    23283 => x"00016cec", 23284 => x"0000bdf8", 23285 => x"00000000",
    23286 => x"00000000", 23287 => x"01040001", 23288 => x"00016cf0",
    23289 => x"0000bdf8", 23290 => x"00000000", 23291 => x"00000000",
    23292 => x"01020001", 23293 => x"00016cf4", 23294 => x"0000bdf8",
    23295 => x"00000000", 23296 => x"00000000", 23297 => x"01020001",
    23298 => x"00016cf8", 23299 => x"0000bdf8", 23300 => x"00000000",
    23301 => x"00000000", 23302 => x"01020001", 23303 => x"00000000",
    23304 => x"00000000", 23305 => x"00000000", 23306 => x"00000000",
    23307 => x"00000000", 23308 => x"01000000", 23309 => x"02000000",
    23310 => x"03000000", 23311 => x"04000000", 23312 => x"00015324",
    23313 => x"01000000", 23314 => x"02000000", 23315 => x"03000000",
    23316 => x"02000000", 23317 => x"03000000", 23318 => x"01000000",
    23319 => x"02000000", 23320 => x"03000000", 23321 => x"04000000",
    23322 => x"05000000", 23323 => x"06000000", 23324 => x"07000000",
    23325 => x"08000000", 23326 => x"09000000", 23327 => x"05000000",
    23328 => x"08000000", 23329 => x"09000000", 23330 => x"0a000000",
    23331 => x"0c000000", 23332 => x"0d000000", 23333 => x"0e000000",
    23334 => x"0f000000", 23335 => x"10000000", 23336 => x"11000000",
    23337 => x"12000000", 23338 => x"13000000", 23339 => x"14000000",
    23340 => x"16000000", 23341 => x"17000000", 23342 => x"18000000",
    23343 => x"1a000000", 23344 => x"01000000", 23345 => x"02000000",
    23346 => x"03000000", 23347 => x"04000000", 23348 => x"05000000",
    23349 => x"06000000", 23350 => x"01000000", 23351 => x"02000000",
    23352 => x"03000000", 23353 => x"04000000", 23354 => x"05000000",
    23355 => x"02000000", 23356 => x"03000000", 23357 => x"04000000",
    23358 => x"05000000", 23359 => x"00016ed0", 23360 => x"00016fbc",
    23361 => x"00000000", 23362 => x"00000000", 23363 => x"00000004",
    23364 => x"00000008", 23365 => x"00000100", 23366 => x"00000200",
    23367 => x"046362a0", 23368 => x"00018fa4", 23369 => x"00000000",
    23370 => x"00000000", 23371 => x"0000ce42", 23372 => x"ab28633a",
    23373 => x"00000000", 23374 => x"00018c18", 23375 => x"00000000",
    23376 => x"00000000", 23377 => x"0000ce42", 23378 => x"650c2d4f",
    23379 => x"00000000", 23380 => x"00018fac", 23381 => x"00000000",
    23382 => x"00000000", 23383 => x"0000ce42", 23384 => x"65158dc0",
    23385 => x"00000000", 23386 => x"00018c38", 23387 => x"00000000",
    23388 => x"00000000", 23389 => x"0000ce42", 23390 => x"de0d8ced",
    23391 => x"00000000", 23392 => x"00018fa8", 23393 => x"00000000",
    23394 => x"00000000", 23395 => x"0000ce42", 23396 => x"ff07fc47",
    23397 => x"00000000", 23398 => x"00018f74", 23399 => x"00000000",
    23400 => x"00000000", 23401 => x"0000ce42", 23402 => x"e2d13d04",
    23403 => x"00000000", 23404 => x"00018f48", 23405 => x"00000000",
    23406 => x"00000000", 23407 => x"0000ce42", 23408 => x"779c5443",
    23409 => x"00000000", 23410 => x"00018fa0", 23411 => x"00000000",
    23412 => x"00000000", 23413 => x"00000651", 23414 => x"68202b22",
    23415 => x"00000000", 23416 => x"00018f98", 23417 => x"00000000",
    23418 => x"00000000", 23419 => x"00001103", 23420 => x"c0413599",
    23421 => x"00000000", 23422 => x"0001545c", 23423 => x"00000000",
    23424 => x"00000001", 23425 => x"00030000", 23426 => x"00000004",
    23427 => x"00000000", 23428 => x"00000000", 23429 => x"00000000",
    23430 => x"00000000", 23431 => x"00000000", 23432 => x"00000000",
    23433 => x"00000000", 23434 => x"00000000", 23435 => x"00000000",
    23436 => x"00000000", 23437 => x"00000000", 23438 => x"00000000",
    23439 => x"00000000", 23440 => x"00000000", 23441 => x"00000000",
    23442 => x"00000000", 23443 => x"00000000", 23444 => x"00000000",
    23445 => x"00000000", 23446 => x"00000000", 23447 => x"00000000",
    23448 => x"00000000", 23449 => x"00000000", 23450 => x"00000000",
    23451 => x"00000000", 23452 => x"00000000", 23453 => x"00000000",
    23454 => x"00000000", 23455 => x"00000000", 23456 => x"00000000",
    23457 => x"00000000", 23458 => x"00000000", 23459 => x"00000000",
    23460 => x"00000000", 23461 => x"00000000", 23462 => x"00000000",
    23463 => x"00000000", 23464 => x"00000000", 23465 => x"00000000",
    23466 => x"00000000", 23467 => x"00000000", 23468 => x"ff000000",
    23469 => x"0000fc0c", 23470 => x"0000fc40", 23471 => x"0000fc70",
    23472 => x"0001483c", 23473 => x"80000000", 23474 => x"00000000",
    23475 => x"00000000", 23476 => x"44332211", 23477 => x"00000000",
    23478 => x"04000000", 23479 => x"138046e2", 23480 => x"01000000",
    23481 => x"9000cfea", 23482 => x"01000000", 23483 => x"108157f3",
    23484 => x"01000000", 23485 => x"0be0ffff", 23486 => x"01000000",
    23487 => x"88e0ffff", 23488 => x"01000000", 23489 => x"08e1ffff",
    23490 => x"01000000", 23491 => x"1b0020e0", 23492 => x"01000000",
    23493 => x"9800c0eb", 23494 => x"01000000", 23495 => x"6b2130e0",
    23496 => x"01000000", 23497 => x"69610de0", 23498 => x"01000000",
    23499 => x"10a38900", 23500 => x"04000000", 23501 => x"33e31ef1",
    23502 => x"01000000", 23503 => x"31c35ff9", 23504 => x"01000000",
    23505 => x"2b0300e1", 23506 => x"01000000", 23507 => x"43c300e1",
    23508 => x"01000000", 23509 => x"79411400", 23510 => x"04000000",
    23511 => x"cb250060", 23512 => x"00000000", 23513 => x"d3250260",
    23514 => x"00000000", 23515 => x"81c88001", 23516 => x"04000000",
    23517 => x"c02fc100", 23518 => x"04000000", 23519 => x"50ea8101",
    23520 => x"04000000", 23521 => x"5b090080", 23522 => x"01000000",
    23523 => x"59092080", 23524 => x"01000000", 23525 => x"c86a8101",
    23526 => x"04000000", 23527 => x"63097afd", 23528 => x"01000000",
    23529 => x"e88a8101", 23530 => x"04000000", 23531 => x"fc8a8101",
    23532 => x"04000000", 23533 => x"00000000", 23534 => x"08000000",
    23535 => x"ffffffff", 23536 => x"00015d70", 23537 => x"5b1157a7",
    23538 => x"00000003", 23539 => x"00000000", 23540 => x"00000000",
    23541 => x"00000000", 23542 => x"00000000", 23543 => x"00000000",
    23544 => x"00000000", 23545 => x"00000000", 23546 => x"00000000",
    23547 => x"00000000", 23548 => x"00000000", 23549 => x"00000000",
    23550 => x"77727063", 23551 => x"2d76332e", 23552 => x"302d3238",
    23553 => x"342d6764", 23554 => x"31613339", 23555 => x"61302d64",
    23556 => x"69727479", 23557 => x"00000000", 23558 => x"4e6f7620",
    23559 => x"33302032", 23560 => x"30313600", 23561 => x"00000000",
    23562 => x"32313a31", 23563 => x"323a3137", 23564 => x"00000000",
    23565 => x"00000000", 23566 => x"686f6e67", 23567 => x"6d696e67",
    23568 => x"00000000", 23569 => x"00000000", 23570 => x"00000000",
    23571 => x"00000000", 23572 => x"00000000", 23573 => x"00000000",
    23574 => x"00014d4c", 23575 => x"00008880", 23576 => x"00013518",
    23577 => x"00008940", 23578 => x"00014d64", 23579 => x"000089a0",
    23580 => x"00014d98", 23581 => x"00008a3c", 23582 => x"00014dec",
    23583 => x"00008b54", 23584 => x"00014e3c", 23585 => x"00008c64",
    23586 => x"00014e5c", 23587 => x"00008d44", 23588 => x"00014e80",
    23589 => x"00008da4", 23590 => x"00014fb0", 23591 => x"00008ea8",
    23592 => x"00014fec", 23593 => x"00009240", 23594 => x"00015048",
    23595 => x"000094a8", 23596 => x"00015080", 23597 => x"00009580",
    23598 => x"00015088", 23599 => x"000096e0", 23600 => x"0001508c",
    23601 => x"000096f8", 23602 => x"000150bc", 23603 => x"00009714",
    23604 => x"00015130", 23605 => x"00009864", 23606 => x"0001514c",
    23607 => x"00009954", 23608 => x"00014fb4", 23609 => x"0000999c",
    23610 => x"00015540", 23611 => x"0000e950", 23612 => x"00015654",
    23613 => x"0000febc", 23614 => x"00015658", 23615 => x"0000fdc0",
    23616 => x"0001565c", 23617 => x"0000fcc4", 23618 => x"000104f0",
    23619 => x"00000000", 23620 => x"00016ec0", 23621 => x"00013530",
    23622 => x"00000000", 23623 => x"00000214", 23624 => x"00000000",
    23625 => x"00000000", 23626 => x"00000000", 23627 => x"00000000",
    23628 => x"00013504", 23629 => x"00000000", 23630 => x"00000000",
    23631 => x"0001220c", 23632 => x"00000000", 23633 => x"00000000",
    23634 => x"00000000", 23635 => x"0001350c", 23636 => x"00000000",
    23637 => x"000087d4", 23638 => x"000004f8", 23639 => x"00000000",
    23640 => x"00000000", 23641 => x"00000000", 23642 => x"00013518",
    23643 => x"00000000", 23644 => x"00000000", 23645 => x"000010e8",
    23646 => x"00000000", 23647 => x"00000000", 23648 => x"00000000",
    23649 => x"0001351c", 23650 => x"00000000", 23651 => x"000004d4",
    23652 => x"00000468", 23653 => x"00000000", 23654 => x"00000000",
    23655 => x"00000000", 23656 => x"00013524", 23657 => x"00000000",
    23658 => x"00000000", 23659 => x"00000378", 23660 => x"00000000",
    23661 => x"00000000", 23662 => x"00000000", 23663 => x"00014c34",
    23664 => x"00000000", 23665 => x"00000000", 23666 => x"00007678",
    23667 => x"00000000", 23668 => x"00000000", 23669 => x"00000000",
    23670 => x"000152a4", 23671 => x"00018f88", 23672 => x"00000000",
    23673 => x"0000a0d8", 23674 => x"00000000", 23675 => x"00000000",
    23676 => x"00000000", 23677 => x"000152ac", 23678 => x"00018f88",
    23679 => x"0000a848", 23680 => x"0000a8f8", 23681 => x"00000000",
    23682 => x"00000000", 23683 => x"00000000", 23684 => x"000152b4",
    23685 => x"00018f88", 23686 => x"0000ae04", 23687 => x"0000ac78",
    23688 => x"00000000", 23689 => x"00000000", 23690 => x"00000000",
    23691 => x"0001531c", 23692 => x"00018f88", 23693 => x"0000c524",
    23694 => x"0000b54c", 23695 => x"00000000", 23696 => x"00000000",
    23697 => x"00000000", 23698 => x"00015548", 23699 => x"00000000",
    23700 => x"0000e628", 23701 => x"0000e674", 23702 => x"00000000",
    23703 => x"00000000", 23704 => x"00000000", 23705 => x"00000000",
    23706 => x"00000000", 23707 => x"00000000", 23708 => x"00000000",
    23709 => x"00000000", 23710 => x"00000000", 23711 => x"00000000",
    23712 => x"00000000", 23713 => x"00000000", 23714 => x"00000000",
    23715 => x"00000000", 23716 => x"00000000", 23717 => x"00000000",
    23718 => x"00000000", 23719 => x"00000000", 23720 => x"00000000",
    23721 => x"00000000", 23722 => x"00000000", 23723 => x"00000000",
    23724 => x"00000000", 23725 => x"00000000", 23726 => x"00000000",
    23727 => x"00000000", 23728 => x"00000000", 23729 => x"00000000",
    23730 => x"00000000", 23731 => x"00000000", 23732 => x"00000000",
    23733 => x"00000000", 23734 => x"00000000", 23735 => x"00000000",
    23736 => x"00000000", 23737 => x"00000000", 23738 => x"00000000",
    23739 => x"00000000", 23740 => x"00000000", 23741 => x"00000000",
    23742 => x"00000000", 23743 => x"00000000", 23744 => x"00000000",
    23745 => x"00000000", 23746 => x"00000000", 23747 => x"00000000",
    23748 => x"00000000", 23749 => x"00000000", 23750 => x"00000000",
    23751 => x"00000000", 23752 => x"00000000", 23753 => x"00000000",
    23754 => x"00000000", 23755 => x"00000000", 23756 => x"00000000",
    23757 => x"00000000", 23758 => x"00000000", 23759 => x"00000000",
    23760 => x"00000000", 23761 => x"00000000", 23762 => x"00000000",
    23763 => x"00000000", 23764 => x"00000000", 23765 => x"00000000",
    23766 => x"00000000", 23767 => x"00000000", 23768 => x"00000000",
    23769 => x"00000000", 23770 => x"00000000", 23771 => x"00000000",
    23772 => x"00000000", 23773 => x"00000000", 23774 => x"00000000",
    23775 => x"00000000", 23776 => x"00000000", 23777 => x"00000000",
    23778 => x"00000000", 23779 => x"00000000", 23780 => x"00000000",
    23781 => x"00000000", 23782 => x"00000000", 23783 => x"00000000",
    23784 => x"00000000", 23785 => x"00000000", 23786 => x"00000000",
    23787 => x"00000000", 23788 => x"00000000", 23789 => x"00000000",
    23790 => x"00000000", 23791 => x"00000000", 23792 => x"00000000",
    23793 => x"00000000", 23794 => x"00000000", 23795 => x"00000000",
    23796 => x"00000000", 23797 => x"00000000", 23798 => x"00000000",
    23799 => x"00000000", 23800 => x"00000000", 23801 => x"00000000",
    23802 => x"00000000", 23803 => x"00000000", 23804 => x"00000000",
    23805 => x"00000000", 23806 => x"00000000", 23807 => x"00000000",
    23808 => x"00000000", 23809 => x"00000000", 23810 => x"00000000",
    23811 => x"00000000", 23812 => x"00000000", 23813 => x"00000000",
    23814 => x"00000000", 23815 => x"00000000", 23816 => x"00000000",
    23817 => x"00000000", 23818 => x"00000000", 23819 => x"00000000",
    23820 => x"00000000", 23821 => x"00000000", 23822 => x"00000000",
    23823 => x"00000000", 23824 => x"00000000", 23825 => x"00000000",
    23826 => x"00000000", 23827 => x"00000000", 23828 => x"00000000",
    23829 => x"00000000", 23830 => x"00000000", 23831 => x"00000000",
    23832 => x"00000000", 23833 => x"00000000", 23834 => x"00000000",
    23835 => x"00000000", 23836 => x"00000000", 23837 => x"00000000",
    23838 => x"00000000", 23839 => x"00000000", 23840 => x"00000000",
    23841 => x"00000000", 23842 => x"00000000", 23843 => x"00000000",
    23844 => x"00000000", 23845 => x"00000000", 23846 => x"00000000",
    23847 => x"00000000", 23848 => x"00000000", 23849 => x"00000000",
    23850 => x"00000000", 23851 => x"00000000", 23852 => x"00000000",
    23853 => x"00000000", 23854 => x"00000000", 23855 => x"00000000",
    23856 => x"00000000", 23857 => x"00000000", 23858 => x"00000000",
    23859 => x"00000000", 23860 => x"00000000", 23861 => x"00000000",
    23862 => x"00000000", 23863 => x"00000000", 23864 => x"00000000",
    23865 => x"00000000", 23866 => x"00000000", 23867 => x"00000000",
    23868 => x"00000000", 23869 => x"00000000", 23870 => x"00000000",
    23871 => x"00000000", 23872 => x"00000000", 23873 => x"00000000",
    23874 => x"00000000", 23875 => x"00000000", 23876 => x"00000000",
    23877 => x"00000000", 23878 => x"00000000", 23879 => x"00000000",
    23880 => x"00000000", 23881 => x"00000000", 23882 => x"00000000",
    23883 => x"00000000", 23884 => x"00000000", 23885 => x"00000000",
    23886 => x"00000000", 23887 => x"00000000", 23888 => x"00000000",
    23889 => x"00000000", 23890 => x"00000000", 23891 => x"00000000",
    23892 => x"00000000", 23893 => x"00000000", 23894 => x"00000000",
    23895 => x"00000000", 23896 => x"00000000", 23897 => x"00000000",
    23898 => x"00000000", 23899 => x"00000000", 23900 => x"00000000",
    23901 => x"00000000", 23902 => x"00000000", 23903 => x"00000000",
    23904 => x"00000000", 23905 => x"00000000", 23906 => x"00000000",
    23907 => x"00000000", 23908 => x"00000000", 23909 => x"00000000",
    23910 => x"00000000", 23911 => x"00000000", 23912 => x"00000000",
    23913 => x"00000000", 23914 => x"00000000", 23915 => x"00000000",
    23916 => x"00000000", 23917 => x"00000000", 23918 => x"00000000",
    23919 => x"00000000", 23920 => x"00000000", 23921 => x"00000000",
    23922 => x"00000000", 23923 => x"00000000", 23924 => x"00000000",
    23925 => x"00000000", 23926 => x"00000000", 23927 => x"00000000",
    23928 => x"00000000", 23929 => x"00000000", 23930 => x"00000000",
    23931 => x"00000000", 23932 => x"00000000", 23933 => x"00000000",
    23934 => x"00000000", 23935 => x"00000000", 23936 => x"00000000",
    23937 => x"00000000", 23938 => x"00000000", 23939 => x"00000000",
    23940 => x"00000000", 23941 => x"00000000", 23942 => x"00000000",
    23943 => x"00000000", 23944 => x"00000000", 23945 => x"00000000",
    23946 => x"00000000", 23947 => x"00000000", 23948 => x"00000000",
    23949 => x"00000000", 23950 => x"00000000", 23951 => x"00000000",
    23952 => x"00000000", 23953 => x"00000000", 23954 => x"00000000",
    23955 => x"00000000", 23956 => x"00000000", 23957 => x"00000000",
    23958 => x"00000000", 23959 => x"00000000", 23960 => x"00000000",
    23961 => x"00000000", 23962 => x"00000000", 23963 => x"00000000",
    23964 => x"00000000", 23965 => x"00000000", 23966 => x"00000000",
    23967 => x"00000000", 23968 => x"00000000", 23969 => x"00000000",
    23970 => x"00000000", 23971 => x"00000000", 23972 => x"00000000",
    23973 => x"00000000", 23974 => x"00000000", 23975 => x"00000000",
    23976 => x"00000000", 23977 => x"00000000", 23978 => x"00000000",
    23979 => x"00000000", 23980 => x"00000000", 23981 => x"00000000",
    23982 => x"00000000", 23983 => x"00000000", 23984 => x"00000000",
    23985 => x"00000000", 23986 => x"00000000", 23987 => x"00000000",
    23988 => x"00000000", 23989 => x"00000000", 23990 => x"00000000",
    23991 => x"00000000", 23992 => x"00000000", 23993 => x"00000000",
    23994 => x"00000000", 23995 => x"00000000", 23996 => x"00000000",
    23997 => x"00000000", 23998 => x"00000000", 23999 => x"00000000",
    24000 => x"00000000", 24001 => x"00000000", 24002 => x"00000000",
    24003 => x"00000000", 24004 => x"00000000", 24005 => x"00000000",
    24006 => x"00000000", 24007 => x"00000000", 24008 => x"00000000",
    24009 => x"00000000", 24010 => x"00000000", 24011 => x"00000000",
    24012 => x"00000000", 24013 => x"00000000", 24014 => x"00000000",
    24015 => x"00000000", 24016 => x"00000000", 24017 => x"00000000",
    24018 => x"00000000", 24019 => x"00000000", 24020 => x"00000000",
    24021 => x"00000000", 24022 => x"00000000", 24023 => x"00000000",
    24024 => x"00000000", 24025 => x"00000000", 24026 => x"00000000",
    24027 => x"00000000", 24028 => x"00000000", 24029 => x"00000000",
    24030 => x"00000000", 24031 => x"00000000", 24032 => x"00000000",
    24033 => x"00000000", 24034 => x"00000000", 24035 => x"00000000",
    24036 => x"00000000", 24037 => x"00000000", 24038 => x"00000000",
    24039 => x"00000000", 24040 => x"00000000", 24041 => x"00000000",
    24042 => x"00000000", 24043 => x"00000000", 24044 => x"00000000",
    24045 => x"00000000", 24046 => x"00000000", 24047 => x"00000000",
    24048 => x"00000000", 24049 => x"00000000", 24050 => x"00000000",
    24051 => x"00000000", 24052 => x"00000000", 24053 => x"00000000",
    24054 => x"00000000", 24055 => x"00000000", 24056 => x"00000000",
    24057 => x"00000000", 24058 => x"00000000", 24059 => x"00000000",
    24060 => x"00000000", 24061 => x"00000000", 24062 => x"00000000",
    24063 => x"00000000", 24064 => x"00000000", 24065 => x"00000000",
    24066 => x"00000000", 24067 => x"00000000", 24068 => x"00000000",
    24069 => x"00000000", 24070 => x"00000000", 24071 => x"00000000",
    24072 => x"00000000", 24073 => x"00000000", 24074 => x"00000000",
    24075 => x"00000000", 24076 => x"00000000", 24077 => x"00000000",
    24078 => x"00000000", 24079 => x"00000000", 24080 => x"00000000",
    24081 => x"00000000", 24082 => x"00000000", 24083 => x"00000000",
    24084 => x"00000000", 24085 => x"00000000", 24086 => x"00000000",
    24087 => x"00000000", 24088 => x"00000000", 24089 => x"00000000",
    24090 => x"00000000", 24091 => x"00000000", 24092 => x"00000000",
    24093 => x"00000000", 24094 => x"00000000", 24095 => x"00000000",
    24096 => x"00000000", 24097 => x"00000000", 24098 => x"00000000",
    24099 => x"00000000", 24100 => x"00000000", 24101 => x"00000000",
    24102 => x"00000000", 24103 => x"00000000", 24104 => x"00000000",
    24105 => x"00000000", 24106 => x"00000000", 24107 => x"00000000",
    24108 => x"00000000", 24109 => x"00000000", 24110 => x"00000000",
    24111 => x"00000000", 24112 => x"00000000", 24113 => x"00000000",
    24114 => x"00000000", 24115 => x"00000000", 24116 => x"00000000",
    24117 => x"00000000", 24118 => x"00000000", 24119 => x"00000000",
    24120 => x"00000000", 24121 => x"00000000", 24122 => x"00000000",
    24123 => x"00000000", 24124 => x"00000000", 24125 => x"00000000",
    24126 => x"00000000", 24127 => x"00000000", 24128 => x"00000000",
    24129 => x"00000000", 24130 => x"00000000", 24131 => x"00000000",
    24132 => x"00000000", 24133 => x"00000000", 24134 => x"00000000",
    24135 => x"00000000", 24136 => x"00000000", 24137 => x"00000000",
    24138 => x"00000000", 24139 => x"00000000", 24140 => x"00000000",
    24141 => x"00000000", 24142 => x"00000000", 24143 => x"00000000",
    24144 => x"00000000", 24145 => x"00000000", 24146 => x"00000000",
    24147 => x"00000000", 24148 => x"00000000", 24149 => x"00000000",
    24150 => x"00000000", 24151 => x"00000000", 24152 => x"00000000",
    24153 => x"00000000", 24154 => x"00000000", 24155 => x"00000000",
    24156 => x"00000000", 24157 => x"00000000", 24158 => x"00000000",
    24159 => x"00000000", 24160 => x"00000000", 24161 => x"00000000",
    24162 => x"00000000", 24163 => x"00000000", 24164 => x"00000000",
    24165 => x"00000000", 24166 => x"00000000", 24167 => x"00000000",
    24168 => x"00000000", 24169 => x"00000000", 24170 => x"00000000",
    24171 => x"00000000", 24172 => x"00000000", 24173 => x"00000000",
    24174 => x"00000000", 24175 => x"00000000", 24176 => x"00000000",
    24177 => x"00000000", 24178 => x"00000000", 24179 => x"00000000",
    24180 => x"00000000", 24181 => x"00000000", 24182 => x"00000000",
    24183 => x"00000000", 24184 => x"00000000", 24185 => x"00000000",
    24186 => x"00000000", 24187 => x"00000000", 24188 => x"00000000",
    24189 => x"00000000", 24190 => x"00000000", 24191 => x"00000000",
    24192 => x"00000000", 24193 => x"00000000", 24194 => x"00000000",
    24195 => x"00000000", 24196 => x"00000000", 24197 => x"00000000",
    24198 => x"00000000", 24199 => x"00000000", 24200 => x"00000000",
    24201 => x"00000000", 24202 => x"00000000", 24203 => x"00000000",
    24204 => x"00000000", 24205 => x"00000000", 24206 => x"00000000",
    24207 => x"00000000", 24208 => x"00000000", 24209 => x"00000000",
    24210 => x"00000000", 24211 => x"00000000", 24212 => x"00000000",
    24213 => x"00000000", 24214 => x"00000000", 24215 => x"00000000",
    24216 => x"00000000", 24217 => x"00000000", 24218 => x"00000000",
    24219 => x"00000000", 24220 => x"00000000", 24221 => x"00000000",
    24222 => x"00000000", 24223 => x"00000000", 24224 => x"00000000",
    24225 => x"00000000", 24226 => x"00000000", 24227 => x"00000000",
    24228 => x"00000000", 24229 => x"00000000", 24230 => x"00000000",
    24231 => x"00000000", 24232 => x"00000000", 24233 => x"00000000",
    24234 => x"00000000", 24235 => x"00000000", 24236 => x"00000000",
    24237 => x"00000000", 24238 => x"00000000", 24239 => x"00000000",
    24240 => x"00000000", 24241 => x"00000000", 24242 => x"00000000",
    24243 => x"00000000", 24244 => x"00000000", 24245 => x"00000000",
    24246 => x"00000000", 24247 => x"00000000", 24248 => x"00000000",
    24249 => x"00000000", 24250 => x"00000000", 24251 => x"00000000",
    24252 => x"00000000", 24253 => x"00000000", 24254 => x"00000000",
    24255 => x"00000000", 24256 => x"00000000", 24257 => x"00000000",
    24258 => x"00000000", 24259 => x"00000000", 24260 => x"00000000",
    24261 => x"00000000", 24262 => x"00000000", 24263 => x"00000000",
    24264 => x"00000000", 24265 => x"00000000", 24266 => x"00000000",
    24267 => x"00000000", 24268 => x"00000000", 24269 => x"00000000",
    24270 => x"00000000", 24271 => x"00000000", 24272 => x"00000000",
    24273 => x"00000000", 24274 => x"00000000", 24275 => x"00000000",
    24276 => x"00000000", 24277 => x"00000000", 24278 => x"00000000",
    24279 => x"00000000", 24280 => x"00000000", 24281 => x"00000000",
    24282 => x"00000000", 24283 => x"00000000", 24284 => x"00000000",
    24285 => x"00000000", 24286 => x"00000000", 24287 => x"00000000",
    24288 => x"00000000", 24289 => x"00000000", 24290 => x"00000000",
    24291 => x"00000000", 24292 => x"00000000", 24293 => x"00000000",
    24294 => x"00000000", 24295 => x"00000000", 24296 => x"00000000",
    24297 => x"00000000", 24298 => x"00000000", 24299 => x"00000000",
    24300 => x"00000000", 24301 => x"00000000", 24302 => x"00000000",
    24303 => x"00000000", 24304 => x"00000000", 24305 => x"00000000",
    24306 => x"00000000", 24307 => x"00000000", 24308 => x"00000000",
    24309 => x"00000000", 24310 => x"00000000", 24311 => x"00000000",
    24312 => x"00000000", 24313 => x"00000000", 24314 => x"00000000",
    24315 => x"00000000", 24316 => x"00000000", 24317 => x"00000000",
    24318 => x"00000000", 24319 => x"00000000", 24320 => x"00000000",
    24321 => x"00000000", 24322 => x"00000000", 24323 => x"00000000",
    24324 => x"00000000", 24325 => x"00000000", 24326 => x"00000000",
    24327 => x"00000000", 24328 => x"00000000", 24329 => x"00000000",
    24330 => x"00000000", 24331 => x"00000000", 24332 => x"00000000",
    24333 => x"00000000", 24334 => x"00000000", 24335 => x"00000000",
    24336 => x"00000000", 24337 => x"00000000", 24338 => x"00000000",
    24339 => x"00000000", 24340 => x"00000000", 24341 => x"00000000",
    24342 => x"00000000", 24343 => x"00000000", 24344 => x"00000000",
    24345 => x"00000000", 24346 => x"00000000", 24347 => x"00000000",
    24348 => x"00000000", 24349 => x"00000000", 24350 => x"00000000",
    24351 => x"00000000", 24352 => x"00000000", 24353 => x"00000000",
    24354 => x"00000000", 24355 => x"00000000", 24356 => x"00000000",
    24357 => x"00000000", 24358 => x"00000000", 24359 => x"00000000",
    24360 => x"00000000", 24361 => x"00000000", 24362 => x"00000000",
    24363 => x"00000000", 24364 => x"00000000", 24365 => x"00000000",
    24366 => x"00000000", 24367 => x"00000000", 24368 => x"00000000",
    24369 => x"00000000", 24370 => x"00000000", 24371 => x"00000000",
    24372 => x"00000000", 24373 => x"00000000", 24374 => x"00000000",
    24375 => x"00000000", 24376 => x"00000000", 24377 => x"00000000",
    24378 => x"00000000", 24379 => x"00000000", 24380 => x"00000000",
    24381 => x"00000000", 24382 => x"00000000", 24383 => x"00000000",
    24384 => x"00000000", 24385 => x"00000000", 24386 => x"00000000",
    24387 => x"00000000", 24388 => x"00000000", 24389 => x"00000000",
    24390 => x"00000000", 24391 => x"00000000", 24392 => x"00000000",
    24393 => x"00000000", 24394 => x"00000000", 24395 => x"00000000",
    24396 => x"00000000", 24397 => x"00000000", 24398 => x"00000000",
    24399 => x"00000000", 24400 => x"00000000", 24401 => x"00000000",
    24402 => x"00000000", 24403 => x"00000000", 24404 => x"00000000",
    24405 => x"00000000", 24406 => x"00000000", 24407 => x"00000000",
    24408 => x"00000000", 24409 => x"00000000", 24410 => x"00000000",
    24411 => x"00000000", 24412 => x"00000000", 24413 => x"00000000",
    24414 => x"00000000", 24415 => x"00000000", 24416 => x"00000000",
    24417 => x"00000000", 24418 => x"00000000", 24419 => x"00000000",
    24420 => x"00000000", 24421 => x"00000000", 24422 => x"00000000",
    24423 => x"00000000", 24424 => x"00000000", 24425 => x"00000000",
    24426 => x"00000000", 24427 => x"00000000", 24428 => x"00000000",
    24429 => x"00000000", 24430 => x"00000000", 24431 => x"00000000",
    24432 => x"00000000", 24433 => x"00000000", 24434 => x"00000000",
    24435 => x"00000000", 24436 => x"00000000", 24437 => x"00000000",
    24438 => x"00000000", 24439 => x"00000000", 24440 => x"00000000",
    24441 => x"00000000", 24442 => x"00000000", 24443 => x"00000000",
    24444 => x"00000000", 24445 => x"00000000", 24446 => x"00000000",
    24447 => x"00000000", 24448 => x"00000000", 24449 => x"00000000",
    24450 => x"00000000", 24451 => x"00000000", 24452 => x"00000000",
    24453 => x"00000000", 24454 => x"00000000", 24455 => x"00000000",
    24456 => x"00000000", 24457 => x"00000000", 24458 => x"00000000",
    24459 => x"00000000", 24460 => x"00000000", 24461 => x"00000000",
    24462 => x"00000000", 24463 => x"00000000", 24464 => x"00000000",
    24465 => x"00000000", 24466 => x"00000000", 24467 => x"00000000",
    24468 => x"00000000", 24469 => x"00000000", 24470 => x"00000000",
    24471 => x"00000000", 24472 => x"00000000", 24473 => x"00000000",
    24474 => x"00000000", 24475 => x"00000000", 24476 => x"00000000",
    24477 => x"00000000", 24478 => x"00000000", 24479 => x"00000000",
    24480 => x"00000000", 24481 => x"00000000", 24482 => x"00000000",
    24483 => x"00000000", 24484 => x"00000000", 24485 => x"00000000",
    24486 => x"00000000", 24487 => x"00000000", 24488 => x"00000000",
    24489 => x"00000000", 24490 => x"00000000", 24491 => x"00000000",
    24492 => x"00000000", 24493 => x"00000000", 24494 => x"00000000",
    24495 => x"00000000", 24496 => x"00000000", 24497 => x"00000000",
    24498 => x"00000000", 24499 => x"00000000", 24500 => x"00000000",
    24501 => x"00000000", 24502 => x"00000000", 24503 => x"00000000",
    24504 => x"00000000", 24505 => x"00000000", 24506 => x"00000000",
    24507 => x"00000000", 24508 => x"00000000", 24509 => x"00000000",
    24510 => x"00000000", 24511 => x"00000000", 24512 => x"00000000",
    24513 => x"00000000", 24514 => x"00000000", 24515 => x"00000000",
    24516 => x"00000000", 24517 => x"00000000", 24518 => x"00000000",
    24519 => x"00000000", 24520 => x"00000000", 24521 => x"00000000",
    24522 => x"00000000", 24523 => x"00000000", 24524 => x"00000000",
    24525 => x"00000000", 24526 => x"00000000", 24527 => x"00000000",
    24528 => x"00000000", 24529 => x"00000000", 24530 => x"00000000",
    24531 => x"00000000", 24532 => x"00000000", 24533 => x"00000000",
    24534 => x"00000000", 24535 => x"00000000", 24536 => x"00000000",
    24537 => x"00000000", 24538 => x"00000000", 24539 => x"00000000",
    24540 => x"00000000", 24541 => x"00000000", 24542 => x"00000000",
    24543 => x"00000000", 24544 => x"00000000", 24545 => x"00000000",
    24546 => x"00000000", 24547 => x"00000000", 24548 => x"00000000",
    24549 => x"00000000", 24550 => x"00000000", 24551 => x"00000000",
    24552 => x"00000000", 24553 => x"00000000", 24554 => x"00000000",
    24555 => x"00000000", 24556 => x"00000000", 24557 => x"00000000",
    24558 => x"00000000", 24559 => x"00000000", 24560 => x"00000000",
    24561 => x"00000000", 24562 => x"00000000", 24563 => x"00000000",
    24564 => x"00000000", 24565 => x"00000000", 24566 => x"00000000",
    24567 => x"00000000", 24568 => x"00000000", 24569 => x"00000000",
    24570 => x"00000000", 24571 => x"00000000", 24572 => x"00000000",
    24573 => x"00000000", 24574 => x"00000000", 24575 => x"00000000",
    24576 => x"00000000", 24577 => x"00000000", 24578 => x"00000000",
    24579 => x"00000000", 24580 => x"00000000", 24581 => x"00000000",
    24582 => x"00000000", 24583 => x"00000000", 24584 => x"00000000",
    24585 => x"00000000", 24586 => x"00000000", 24587 => x"00000000",
    24588 => x"00000000", 24589 => x"00000000", 24590 => x"00000000",
    24591 => x"00000000", 24592 => x"00000000", 24593 => x"00000000",
    24594 => x"00000000", 24595 => x"00000000", 24596 => x"00000000",
    24597 => x"00000000", 24598 => x"00000000", 24599 => x"00000000",
    24600 => x"00000000", 24601 => x"00000000", 24602 => x"00000000",
    24603 => x"00000000", 24604 => x"00000000", 24605 => x"00000000",
    24606 => x"00000000", 24607 => x"00000000", 24608 => x"00000000",
    24609 => x"00000000", 24610 => x"00000000", 24611 => x"00000000",
    24612 => x"00000000", 24613 => x"00000000", 24614 => x"00000000",
    24615 => x"00000000", 24616 => x"00000000", 24617 => x"00000000",
    24618 => x"00000000", 24619 => x"00000000", 24620 => x"00000000",
    24621 => x"00000000", 24622 => x"00000000", 24623 => x"00000000",
    24624 => x"00000000", 24625 => x"00000000", 24626 => x"00000000",
    24627 => x"00000000", 24628 => x"00000000", 24629 => x"00000000",
    24630 => x"00000000", 24631 => x"00000000", 24632 => x"00000000",
    24633 => x"00000000", 24634 => x"00000000", 24635 => x"00000000",
    24636 => x"00000000", 24637 => x"00000000", 24638 => x"00000000",
    24639 => x"00000000", 24640 => x"00000000", 24641 => x"00000000",
    24642 => x"00000000", 24643 => x"00000000", 24644 => x"00000000",
    24645 => x"00000000", 24646 => x"00000000", 24647 => x"00000000",
    24648 => x"00000000", 24649 => x"00000000", 24650 => x"00000000",
    24651 => x"00000000", 24652 => x"00000000", 24653 => x"00000000",
    24654 => x"00000000", 24655 => x"00000000", 24656 => x"00000000",
    24657 => x"00000000", 24658 => x"00000000", 24659 => x"00000000",
    24660 => x"00000000", 24661 => x"00000000", 24662 => x"00000000",
    24663 => x"00000000", 24664 => x"00000000", 24665 => x"00000000",
    24666 => x"00000000", 24667 => x"00000000", 24668 => x"00000000",
    24669 => x"00000000", 24670 => x"00000000", 24671 => x"00000000",
    24672 => x"00000000", 24673 => x"00000000", 24674 => x"00000000",
    24675 => x"00000000", 24676 => x"00000000", 24677 => x"00000000",
    24678 => x"00000000", 24679 => x"00000000", 24680 => x"00000000",
    24681 => x"00000000", 24682 => x"00000000", 24683 => x"00000000",
    24684 => x"00000000", 24685 => x"00000000", 24686 => x"00000000",
    24687 => x"00000000", 24688 => x"00000000", 24689 => x"00000000",
    24690 => x"00000000", 24691 => x"00000000", 24692 => x"00000000",
    24693 => x"00000000", 24694 => x"00000000", 24695 => x"00000000",
    24696 => x"00000000", 24697 => x"00000000", 24698 => x"00000000",
    24699 => x"00000000", 24700 => x"00000000", 24701 => x"00000000",
    24702 => x"00000000", 24703 => x"00000000", 24704 => x"00000000",
    24705 => x"00000000", 24706 => x"00000000", 24707 => x"00000000",
    24708 => x"00000000", 24709 => x"00000000", 24710 => x"00000000",
    24711 => x"00000000", 24712 => x"00000000", 24713 => x"00000000",
    24714 => x"00000000", 24715 => x"00000000", 24716 => x"00000000",
    24717 => x"00000000", 24718 => x"00000000", 24719 => x"00000000",
    24720 => x"00000000", 24721 => x"00000000", 24722 => x"00000000",
    24723 => x"00000000", 24724 => x"00000000", 24725 => x"00000000",
    24726 => x"00000000", 24727 => x"00000000", 24728 => x"00000000",
    24729 => x"00000000", 24730 => x"00000000", 24731 => x"00000000",
    24732 => x"00000000", 24733 => x"00000000", 24734 => x"00000000",
    24735 => x"00000000", 24736 => x"00000000", 24737 => x"00000000",
    24738 => x"00000000", 24739 => x"00000000", 24740 => x"00000000",
    24741 => x"00000000", 24742 => x"00000000", 24743 => x"00000000",
    24744 => x"00000000", 24745 => x"00000000", 24746 => x"00000000",
    24747 => x"00000000", 24748 => x"00000000", 24749 => x"00000000",
    24750 => x"00000000", 24751 => x"00000000", 24752 => x"00000000",
    24753 => x"00000000", 24754 => x"00000000", 24755 => x"00000000",
    24756 => x"00000000", 24757 => x"00000000", 24758 => x"00000000",
    24759 => x"00000000", 24760 => x"00000000", 24761 => x"00000000",
    24762 => x"00000000", 24763 => x"00000000", 24764 => x"00000000",
    24765 => x"00000000", 24766 => x"00000000", 24767 => x"00000000",
    24768 => x"00000000", 24769 => x"00000000", 24770 => x"00000000",
    24771 => x"00000000", 24772 => x"00000000", 24773 => x"00000000",
    24774 => x"00000000", 24775 => x"00000000", 24776 => x"00000000",
    24777 => x"00000000", 24778 => x"00000000", 24779 => x"00000000",
    24780 => x"00000000", 24781 => x"00000000", 24782 => x"00000000",
    24783 => x"00000000", 24784 => x"00000000", 24785 => x"00000000",
    24786 => x"00000000", 24787 => x"00000000", 24788 => x"00000000",
    24789 => x"00000000", 24790 => x"00000000", 24791 => x"00000000",
    24792 => x"00000000", 24793 => x"00000000", 24794 => x"00000000",
    24795 => x"00000000", 24796 => x"00000000", 24797 => x"00000000",
    24798 => x"00000000", 24799 => x"00000000", 24800 => x"00000000",
    24801 => x"00000000", 24802 => x"00000000", 24803 => x"00000000",
    24804 => x"00000000", 24805 => x"00000000", 24806 => x"00000000",
    24807 => x"00000000", 24808 => x"00000000", 24809 => x"00000000",
    24810 => x"00000000", 24811 => x"00000000", 24812 => x"00000000",
    24813 => x"00000000", 24814 => x"00000000", 24815 => x"00000000",
    24816 => x"00000000", 24817 => x"00000000", 24818 => x"00000000",
    24819 => x"00000000", 24820 => x"00000000", 24821 => x"00000000",
    24822 => x"00000000", 24823 => x"00000000", 24824 => x"00000000",
    24825 => x"00000000", 24826 => x"00000000", 24827 => x"00000000",
    24828 => x"00000000", 24829 => x"00000000", 24830 => x"00000000",
    24831 => x"00000000", 24832 => x"00000000", 24833 => x"00000000",
    24834 => x"00000000", 24835 => x"00000000", 24836 => x"00000000",
    24837 => x"00000000", 24838 => x"00000000", 24839 => x"00000000",
    24840 => x"00000000", 24841 => x"00000000", 24842 => x"00000000",
    24843 => x"00000000", 24844 => x"00000000", 24845 => x"00000000",
    24846 => x"00000000", 24847 => x"00000000", 24848 => x"00000000",
    24849 => x"00000000", 24850 => x"00000000", 24851 => x"00000000",
    24852 => x"00000000", 24853 => x"00000000", 24854 => x"00000000",
    24855 => x"00000000", 24856 => x"00000000", 24857 => x"00000000",
    24858 => x"00000000", 24859 => x"00000000", 24860 => x"00000000",
    24861 => x"00000000", 24862 => x"00000000", 24863 => x"00000000",
    24864 => x"00000000", 24865 => x"00000000", 24866 => x"00000000",
    24867 => x"00000000", 24868 => x"00000000", 24869 => x"00000000",
    24870 => x"00000000", 24871 => x"00000000", 24872 => x"00000000",
    24873 => x"00000000", 24874 => x"00000000", 24875 => x"00000000",
    24876 => x"00000000", 24877 => x"00000000", 24878 => x"00000000",
    24879 => x"00000000", 24880 => x"00000000", 24881 => x"00000000",
    24882 => x"00000000", 24883 => x"00000000", 24884 => x"00000000",
    24885 => x"00000000", 24886 => x"00000000", 24887 => x"00000000",
    24888 => x"00000000", 24889 => x"00000000", 24890 => x"00000000",
    24891 => x"00000000", 24892 => x"00000000", 24893 => x"00000000",
    24894 => x"00000000", 24895 => x"00000000", 24896 => x"00000000",
    24897 => x"00000000", 24898 => x"00000000", 24899 => x"00000000",
    24900 => x"00000000", 24901 => x"00000000", 24902 => x"00000000",
    24903 => x"00000000", 24904 => x"00000000", 24905 => x"00000000",
    24906 => x"00000000", 24907 => x"00000000", 24908 => x"00000000",
    24909 => x"00000000", 24910 => x"00000000", 24911 => x"00000000",
    24912 => x"00000000", 24913 => x"00000000", 24914 => x"00000000",
    24915 => x"00000000", 24916 => x"00000000", 24917 => x"00000000",
    24918 => x"00000000", 24919 => x"00000000", 24920 => x"00000000",
    24921 => x"00000000", 24922 => x"00000000", 24923 => x"00000000",
    24924 => x"00000000", 24925 => x"00000000", 24926 => x"00000000",
    24927 => x"00000000", 24928 => x"00000000", 24929 => x"00000000",
    24930 => x"00000000", 24931 => x"00000000", 24932 => x"00000000",
    24933 => x"00000000", 24934 => x"00000000", 24935 => x"00000000",
    24936 => x"00000000", 24937 => x"00000000", 24938 => x"00000000",
    24939 => x"00000000", 24940 => x"00000000", 24941 => x"00000000",
    24942 => x"00000000", 24943 => x"00000000", 24944 => x"00000000",
    24945 => x"00000000", 24946 => x"00000000", 24947 => x"00000000",
    24948 => x"00000000", 24949 => x"00000000", 24950 => x"00000000",
    24951 => x"00000000", 24952 => x"00000000", 24953 => x"00000000",
    24954 => x"00000000", 24955 => x"00000000", 24956 => x"00000000",
    24957 => x"00000000", 24958 => x"00000000", 24959 => x"00000000",
    24960 => x"00000000", 24961 => x"00000000", 24962 => x"00000000",
    24963 => x"00000000", 24964 => x"00000000", 24965 => x"00000000",
    24966 => x"00000000", 24967 => x"00000000", 24968 => x"00000000",
    24969 => x"00000000", 24970 => x"00000000", 24971 => x"00000000",
    24972 => x"00000000", 24973 => x"00000000", 24974 => x"00000000",
    24975 => x"00000000", 24976 => x"00000000", 24977 => x"00000000",
    24978 => x"00000000", 24979 => x"00000000", 24980 => x"00000000",
    24981 => x"00000000", 24982 => x"00000000", 24983 => x"00000000",
    24984 => x"00000000", 24985 => x"00000000", 24986 => x"00000000",
    24987 => x"00000000", 24988 => x"00000000", 24989 => x"00000000",
    24990 => x"00000000", 24991 => x"00000000", 24992 => x"00000000",
    24993 => x"00000000", 24994 => x"00000000", 24995 => x"00000000",
    24996 => x"00000000", 24997 => x"00000000", 24998 => x"00000000",
    24999 => x"00000000", 25000 => x"00000000", 25001 => x"00000000",
    25002 => x"00000000", 25003 => x"00000000", 25004 => x"00000000",
    25005 => x"00000000", 25006 => x"00000000", 25007 => x"00000000",
    25008 => x"00000000", 25009 => x"00000000", 25010 => x"00000000",
    25011 => x"00000000", 25012 => x"00000000", 25013 => x"00000000",
    25014 => x"00000000", 25015 => x"00000000", 25016 => x"00000000",
    25017 => x"00000000", 25018 => x"00000000", 25019 => x"00000000",
    25020 => x"00000000", 25021 => x"00000000", 25022 => x"00000000",
    25023 => x"00000000", 25024 => x"00000000", 25025 => x"00000000",
    25026 => x"00000000", 25027 => x"00000000", 25028 => x"00000000",
    25029 => x"00000000", 25030 => x"00000000", 25031 => x"00000000",
    25032 => x"00000000", 25033 => x"00000000", 25034 => x"00000000",
    25035 => x"00000000", 25036 => x"00000000", 25037 => x"00000000",
    25038 => x"00000000", 25039 => x"00000000", 25040 => x"00000000",
    25041 => x"00000000", 25042 => x"00000000", 25043 => x"00000000",
    25044 => x"00000000", 25045 => x"00000000", 25046 => x"00000000",
    25047 => x"00000000", 25048 => x"00000000", 25049 => x"00000000",
    25050 => x"00000000", 25051 => x"00000000", 25052 => x"00000000",
    25053 => x"00000000", 25054 => x"00000000", 25055 => x"00000000",
    25056 => x"00000000", 25057 => x"00000000", 25058 => x"00000000",
    25059 => x"00000000", 25060 => x"00000000", 25061 => x"00000000",
    25062 => x"00000000", 25063 => x"00000000", 25064 => x"00000000",
    25065 => x"00000000", 25066 => x"00000000", 25067 => x"00000000",
    25068 => x"00000000", 25069 => x"00000000", 25070 => x"00000000",
    25071 => x"00000000", 25072 => x"00000000", 25073 => x"00000000",
    25074 => x"00000000", 25075 => x"00000000", 25076 => x"00000000",
    25077 => x"00000000", 25078 => x"00000000", 25079 => x"00000000",
    25080 => x"00000000", 25081 => x"00000000", 25082 => x"00000000",
    25083 => x"00000000", 25084 => x"00000000", 25085 => x"00000000",
    25086 => x"00000000", 25087 => x"00000000", 25088 => x"00000000",
    25089 => x"00000000", 25090 => x"00000000", 25091 => x"00000000",
    25092 => x"00000000", 25093 => x"00000000", 25094 => x"00000000",
    25095 => x"00000000", 25096 => x"00000000", 25097 => x"00000000",
    25098 => x"00000000", 25099 => x"00000000", 25100 => x"00000000",
    25101 => x"00000000", 25102 => x"00000000", 25103 => x"00000000",
    25104 => x"00000000", 25105 => x"00000000", 25106 => x"00000000",
    25107 => x"00000000", 25108 => x"00000000", 25109 => x"00000000",
    25110 => x"00000000", 25111 => x"00000000", 25112 => x"00000000",
    25113 => x"00000000", 25114 => x"00000000", 25115 => x"00000000",
    25116 => x"00000000", 25117 => x"00000000", 25118 => x"00000000",
    25119 => x"00000000", 25120 => x"00000000", 25121 => x"00000000",
    25122 => x"00000000", 25123 => x"00000000", 25124 => x"00000000",
    25125 => x"00000000", 25126 => x"00000000", 25127 => x"00000000",
    25128 => x"00000000", 25129 => x"00000000", 25130 => x"00000000",
    25131 => x"00000000", 25132 => x"00000000", 25133 => x"00000000",
    25134 => x"00000000", 25135 => x"00000000", 25136 => x"00000000",
    25137 => x"00000000", 25138 => x"00000000", 25139 => x"00000000",
    25140 => x"00000000", 25141 => x"00000000", 25142 => x"00000000",
    25143 => x"00000000", 25144 => x"00000000", 25145 => x"00000000",
    25146 => x"00000000", 25147 => x"00000000", 25148 => x"00000000",
    25149 => x"00000000", 25150 => x"00000000", 25151 => x"00000000",
    25152 => x"00000000", 25153 => x"00000000", 25154 => x"00000000",
    25155 => x"00000000", 25156 => x"00000000", 25157 => x"00000000",
    25158 => x"00000000", 25159 => x"00000000", 25160 => x"00000000",
    25161 => x"00000000", 25162 => x"00000000", 25163 => x"00000000",
    25164 => x"00000000", 25165 => x"00000000", 25166 => x"00000000",
    25167 => x"00000000", 25168 => x"00000000", 25169 => x"00000000",
    25170 => x"00000000", 25171 => x"00000000", 25172 => x"00000000",
    25173 => x"00000000", 25174 => x"00000000", 25175 => x"00000000",
    25176 => x"00000000", 25177 => x"00000000", 25178 => x"00000000",
    25179 => x"00000000", 25180 => x"00000000", 25181 => x"00000000",
    25182 => x"00000000", 25183 => x"00000000", 25184 => x"00000000",
    25185 => x"00000000", 25186 => x"00000000", 25187 => x"00000000",
    25188 => x"00000000", 25189 => x"00000000", 25190 => x"00000000",
    25191 => x"00000000", 25192 => x"00000000", 25193 => x"00000000",
    25194 => x"00000000", 25195 => x"00000000", 25196 => x"00000000",
    25197 => x"00000000", 25198 => x"00000000", 25199 => x"00000000",
    25200 => x"00000000", 25201 => x"00000000", 25202 => x"00000000",
    25203 => x"00000000", 25204 => x"00000000", 25205 => x"00000000",
    25206 => x"00000000", 25207 => x"00000000", 25208 => x"00000000",
    25209 => x"00000000", 25210 => x"00000000", 25211 => x"00000000",
    25212 => x"00000000", 25213 => x"00000000", 25214 => x"00000000",
    25215 => x"00000000", 25216 => x"00000000", 25217 => x"00000000",
    25218 => x"00000000", 25219 => x"00000000", 25220 => x"00000000",
    25221 => x"00000000", 25222 => x"00000000", 25223 => x"00000000",
    25224 => x"00000000", 25225 => x"00000000", 25226 => x"00000000",
    25227 => x"00000000", 25228 => x"00000000", 25229 => x"00000000",
    25230 => x"00000000", 25231 => x"00000000", 25232 => x"00000000",
    25233 => x"00000000", 25234 => x"00000000", 25235 => x"00000000",
    25236 => x"00000000", 25237 => x"00000000", 25238 => x"00000000",
    25239 => x"00000000", 25240 => x"00000000", 25241 => x"00000000",
    25242 => x"00000000", 25243 => x"00000000", 25244 => x"00000000",
    25245 => x"00000000", 25246 => x"00000000", 25247 => x"00000000",
    25248 => x"00000000", 25249 => x"00000000", 25250 => x"00000000",
    25251 => x"00000000", 25252 => x"00000000", 25253 => x"00000000",
    25254 => x"00000000", 25255 => x"00000000", 25256 => x"00000000",
    25257 => x"00000000", 25258 => x"00000000", 25259 => x"00000000",
    25260 => x"00000000", 25261 => x"00000000", 25262 => x"00000000",
    25263 => x"00000000", 25264 => x"00000000", 25265 => x"00000000",
    25266 => x"00000000", 25267 => x"00000000", 25268 => x"00000000",
    25269 => x"00000000", 25270 => x"00000000", 25271 => x"00000000",
    25272 => x"00000000", 25273 => x"00000000", 25274 => x"00000000",
    25275 => x"00000000", 25276 => x"00000000", 25277 => x"00000000",
    25278 => x"00000000", 25279 => x"00000000", 25280 => x"00000000",
    25281 => x"00000000", 25282 => x"00000000", 25283 => x"00000000",
    25284 => x"00000000", 25285 => x"00000000", 25286 => x"00000000",
    25287 => x"00000000", 25288 => x"00000000", 25289 => x"00000000",
    25290 => x"00000000", 25291 => x"00000000", 25292 => x"00000000",
    25293 => x"00000000", 25294 => x"00000000", 25295 => x"00000000",
    25296 => x"00000000", 25297 => x"00000000", 25298 => x"00000000",
    25299 => x"00000000", 25300 => x"00000000", 25301 => x"00000000",
    25302 => x"00000000", 25303 => x"00000000", 25304 => x"00000000",
    25305 => x"00000000", 25306 => x"00000000", 25307 => x"00000000",
    25308 => x"00000000", 25309 => x"00000000", 25310 => x"00000000",
    25311 => x"00000000", 25312 => x"00000000", 25313 => x"00000000",
    25314 => x"00000000", 25315 => x"00000000", 25316 => x"00000000",
    25317 => x"00000000", 25318 => x"00000000", 25319 => x"00000000",
    25320 => x"00000000", 25321 => x"00000000", 25322 => x"00000000",
    25323 => x"00000000", 25324 => x"00000000", 25325 => x"00000000",
    25326 => x"00000000", 25327 => x"00000000", 25328 => x"00000000",
    25329 => x"00000000", 25330 => x"00000000", 25331 => x"00000000",
    25332 => x"00000000", 25333 => x"00000000", 25334 => x"00000000",
    25335 => x"00000000", 25336 => x"00000000", 25337 => x"00000000",
    25338 => x"00000000", 25339 => x"00000000", 25340 => x"00000000",
    25341 => x"00000000", 25342 => x"00000000", 25343 => x"00000000",
    25344 => x"00000000", 25345 => x"00000000", 25346 => x"00000000",
    25347 => x"00000000", 25348 => x"00000000", 25349 => x"00000000",
    25350 => x"00000000", 25351 => x"00000000", 25352 => x"00000000",
    25353 => x"00000000", 25354 => x"00000000", 25355 => x"00000000",
    25356 => x"00000000", 25357 => x"00000000", 25358 => x"00000000",
    25359 => x"00000000", 25360 => x"00000000", 25361 => x"00000000",
    25362 => x"00000000", 25363 => x"00000000", 25364 => x"00000000",
    25365 => x"00000000", 25366 => x"00000000", 25367 => x"00000000",
    25368 => x"00000000", 25369 => x"00000000", 25370 => x"00000000",
    25371 => x"00000000", 25372 => x"00000000", 25373 => x"00000000",
    25374 => x"00000000", 25375 => x"00000000", 25376 => x"00000000",
    25377 => x"00000000", 25378 => x"00000000", 25379 => x"00000000",
    25380 => x"00000000", 25381 => x"00000000", 25382 => x"00000000",
    25383 => x"00000000", 25384 => x"00000000", 25385 => x"00000000",
    25386 => x"00000000", 25387 => x"00000000", 25388 => x"00000000",
    25389 => x"00000000", 25390 => x"00000000", 25391 => x"00000000",
    25392 => x"00000000", 25393 => x"00000000", 25394 => x"00000000",
    25395 => x"00000000", 25396 => x"00000000", 25397 => x"00000000",
    25398 => x"00000000", 25399 => x"00000000", 25400 => x"00000000",
    25401 => x"00000000", 25402 => x"00000000", 25403 => x"00000000",
    25404 => x"00000000", 25405 => x"00000000", 25406 => x"00000000",
    25407 => x"00000000", 25408 => x"00000000", 25409 => x"00000000",
    25410 => x"00000000", 25411 => x"00000000", 25412 => x"00000000",
    25413 => x"00000000", 25414 => x"00000000", 25415 => x"00000000",
    25416 => x"00000000", 25417 => x"00000000", 25418 => x"00000000",
    25419 => x"00000000", 25420 => x"00000000", 25421 => x"00000000",
    25422 => x"00000000", 25423 => x"00000000", 25424 => x"00000000",
    25425 => x"00000000", 25426 => x"00000000", 25427 => x"00000000",
    25428 => x"00000000", 25429 => x"00000000", 25430 => x"00000000",
    25431 => x"00000000", 25432 => x"00000000", 25433 => x"00000000",
    25434 => x"00000000", 25435 => x"00000000", 25436 => x"00000000",
    25437 => x"00000000", 25438 => x"00000000", 25439 => x"00000000",
    25440 => x"00000000", 25441 => x"00000000", 25442 => x"00000000",
    25443 => x"00000000", 25444 => x"00000000", 25445 => x"00000000",
    25446 => x"00000000", 25447 => x"00000000", 25448 => x"00000000",
    25449 => x"00000000", 25450 => x"00000000", 25451 => x"00000000",
    25452 => x"00000000", 25453 => x"00000000", 25454 => x"00000000",
    25455 => x"00000000", 25456 => x"00000000", 25457 => x"00000000",
    25458 => x"00000000", 25459 => x"00000000", 25460 => x"00000000",
    25461 => x"00000000", 25462 => x"00000000", 25463 => x"00000000",
    25464 => x"00000000", 25465 => x"00000000", 25466 => x"00000000",
    25467 => x"00000000", 25468 => x"00000000", 25469 => x"00000000",
    25470 => x"00000000", 25471 => x"00000000", 25472 => x"00000000",
    25473 => x"00000000", 25474 => x"00000000", 25475 => x"00000000",
    25476 => x"00000000", 25477 => x"00000000", 25478 => x"00000000",
    25479 => x"00000000", 25480 => x"00000000", 25481 => x"00000000",
    25482 => x"00000000", 25483 => x"00000000", 25484 => x"00000000",
    25485 => x"00000000", 25486 => x"00000000", 25487 => x"00000000",
    25488 => x"00000000", 25489 => x"00000000", 25490 => x"00000000",
    25491 => x"00000000", 25492 => x"00000000", 25493 => x"00000000",
    25494 => x"00000000", 25495 => x"00000000", 25496 => x"00000000",
    25497 => x"00000000", 25498 => x"00000000", 25499 => x"00000000",
    25500 => x"00000000", 25501 => x"00000000", 25502 => x"00000000",
    25503 => x"00000000", 25504 => x"00000000", 25505 => x"00000000",
    25506 => x"00000000", 25507 => x"00000000", 25508 => x"00000000",
    25509 => x"00000000", 25510 => x"00000000", 25511 => x"00000000",
    25512 => x"00000000", 25513 => x"00000000", 25514 => x"00000000",
    25515 => x"00000000", 25516 => x"00000000", 25517 => x"00000000",
    25518 => x"00000000", 25519 => x"00000000", 25520 => x"00000000",
    25521 => x"00000000", 25522 => x"00000000", 25523 => x"00000000",
    25524 => x"00000000", 25525 => x"00000000", 25526 => x"00000000",
    25527 => x"00000000", 25528 => x"00000000", 25529 => x"00000000",
    25530 => x"00000000", 25531 => x"00000000", 25532 => x"00000000",
    25533 => x"00000000", 25534 => x"00000000", 25535 => x"00000000",
    25536 => x"00000000", 25537 => x"00000000", 25538 => x"00000000",
    25539 => x"00000000", 25540 => x"00000000", 25541 => x"00000000",
    25542 => x"00000000", 25543 => x"00000000", 25544 => x"00000000",
    25545 => x"00000000", 25546 => x"00000000", 25547 => x"00000000",
    25548 => x"00000000", 25549 => x"00000000", 25550 => x"00000000",
    25551 => x"00000000", 25552 => x"00000000", 25553 => x"00000000",
    25554 => x"00000000", 25555 => x"00000000", 25556 => x"00000000",
    25557 => x"00000000", 25558 => x"00000000", 25559 => x"00000000",
    25560 => x"00000000", 25561 => x"00000000", 25562 => x"00000000",
    25563 => x"00000000", 25564 => x"00000000", 25565 => x"00000000",
    25566 => x"00000000", 25567 => x"00000000", 25568 => x"00000000",
    25569 => x"00000000", 25570 => x"00000000", 25571 => x"00000000",
    25572 => x"00000000", 25573 => x"00000000", 25574 => x"00000000",
    25575 => x"00000000", 25576 => x"00000000", 25577 => x"00000000",
    25578 => x"00000000", 25579 => x"00000000", 25580 => x"00000000",
    25581 => x"00000000", 25582 => x"00000000", 25583 => x"00000000",
    25584 => x"00000000", 25585 => x"00000000", 25586 => x"00000000",
    25587 => x"00000000", 25588 => x"00000000", 25589 => x"00000000",
    25590 => x"00000000", 25591 => x"00000000", 25592 => x"00000000",
    25593 => x"00000000", 25594 => x"00000000", 25595 => x"00000000",
    25596 => x"00000000", 25597 => x"00000000", 25598 => x"00000000",
    25599 => x"00000000", 25600 => x"00000000", 25601 => x"00000000",
    25602 => x"00000000", 25603 => x"00000000", 25604 => x"00000000",
    25605 => x"00000000", 25606 => x"00000000", 25607 => x"00000000",
    25608 => x"00000000", 25609 => x"00000000", 25610 => x"00000000",
    25611 => x"00000000", 25612 => x"00000000", 25613 => x"00000000",
    25614 => x"00000000", 25615 => x"00000000", 25616 => x"00000000",
    25617 => x"00000000", 25618 => x"00000000", 25619 => x"00000000",
    25620 => x"00000000", 25621 => x"00000000", 25622 => x"00000000",
    25623 => x"00000000", 25624 => x"00000000", 25625 => x"00000000",
    25626 => x"00000000", 25627 => x"00000000", 25628 => x"00000000",
    25629 => x"00000000", 25630 => x"00000000", 25631 => x"00000000",
    25632 => x"00000000", 25633 => x"00000000", 25634 => x"00000000",
    25635 => x"00000000", 25636 => x"00000000", 25637 => x"00000000",
    25638 => x"00000000", 25639 => x"00000000", 25640 => x"00000000",
    25641 => x"00000000", 25642 => x"00000000", 25643 => x"00000000",
    25644 => x"00000000", 25645 => x"00000000", 25646 => x"00000000",
    25647 => x"00000000", 25648 => x"00000000", 25649 => x"00000000",
    25650 => x"00000000", 25651 => x"00000000", 25652 => x"00000000",
    25653 => x"00000000", 25654 => x"00000000", 25655 => x"00000000",
    25656 => x"00000000", 25657 => x"00000000", 25658 => x"00000000",
    25659 => x"00000000", 25660 => x"00000000", 25661 => x"00000000",
    25662 => x"00000000", 25663 => x"00000000", 25664 => x"00000000",
    25665 => x"00000000", 25666 => x"00000000", 25667 => x"00000000",
    25668 => x"00000000", 25669 => x"00000000", 25670 => x"00000000",
    25671 => x"00000000", 25672 => x"00000000", 25673 => x"00000000",
    25674 => x"00000000", 25675 => x"00000000", 25676 => x"00000000",
    25677 => x"00000000", 25678 => x"00000000", 25679 => x"00000000",
    25680 => x"00000000", 25681 => x"00000000", 25682 => x"00000000",
    25683 => x"00000000", 25684 => x"00000000", 25685 => x"00000000",
    25686 => x"00000000", 25687 => x"00000000", 25688 => x"00000000",
    25689 => x"00000000", 25690 => x"00000000", 25691 => x"00000000",
    25692 => x"00000000", 25693 => x"00000000", 25694 => x"00000000",
    25695 => x"00000000", 25696 => x"00000000", 25697 => x"00000000",
    25698 => x"00000000", 25699 => x"00000000", 25700 => x"00000000",
    25701 => x"00000000", 25702 => x"00000000", 25703 => x"00000000",
    25704 => x"00000000", 25705 => x"00000000", 25706 => x"00000000",
    25707 => x"00000000", 25708 => x"00000000", 25709 => x"00000000",
    25710 => x"00000000", 25711 => x"00000000", 25712 => x"00000000",
    25713 => x"00000000", 25714 => x"00000000", 25715 => x"00000000",
    25716 => x"00000000", 25717 => x"00000000", 25718 => x"00000000",
    25719 => x"00000000", 25720 => x"00000000", 25721 => x"00000000",
    25722 => x"00000000", 25723 => x"00000000", 25724 => x"00000000",
    25725 => x"00000000", 25726 => x"00000000", 25727 => x"00000000",
    25728 => x"00000000", 25729 => x"00000000", 25730 => x"00000000",
    25731 => x"00000000", 25732 => x"00000000", 25733 => x"00000000",
    25734 => x"00000000", 25735 => x"00000000", 25736 => x"00000000",
    25737 => x"00000000", 25738 => x"00000000", 25739 => x"00000000",
    25740 => x"00000000", 25741 => x"00000000", 25742 => x"00000000",
    25743 => x"00000000", 25744 => x"00000000", 25745 => x"00000000",
    25746 => x"00000000", 25747 => x"00000000", 25748 => x"00000000",
    25749 => x"00000000", 25750 => x"00000000", 25751 => x"00000000",
    25752 => x"00000000", 25753 => x"00000000", 25754 => x"00000000",
    25755 => x"00000000", 25756 => x"00000000", 25757 => x"00000000",
    25758 => x"00000000", 25759 => x"00000000", 25760 => x"00000000",
    25761 => x"00000000", 25762 => x"00000000", 25763 => x"00000000",
    25764 => x"00000000", 25765 => x"00000000", 25766 => x"00000000",
    25767 => x"00000000", 25768 => x"00000000", 25769 => x"00000000",
    25770 => x"00000000", 25771 => x"00000000", 25772 => x"00000000",
    25773 => x"00000000", 25774 => x"00000000", 25775 => x"00000000",
    25776 => x"00000000", 25777 => x"00000000", 25778 => x"00000000",
    25779 => x"00000000", 25780 => x"00000000", 25781 => x"00000000",
    25782 => x"00000000", 25783 => x"00000000", 25784 => x"00000000",
    25785 => x"00000000", 25786 => x"00000000", 25787 => x"00000000",
    25788 => x"00000000", 25789 => x"00000000", 25790 => x"00000000",
    25791 => x"00000000", 25792 => x"00000000", 25793 => x"00000000",
    25794 => x"00000000", 25795 => x"00000000", 25796 => x"00000000",
    25797 => x"00000000", 25798 => x"00000000", 25799 => x"00000000",
    25800 => x"00000000", 25801 => x"00000000", 25802 => x"00000000",
    25803 => x"00000000", 25804 => x"00000000", 25805 => x"00000000",
    25806 => x"00000000", 25807 => x"00000000", 25808 => x"00000000",
    25809 => x"00000000", 25810 => x"00000000", 25811 => x"00000000",
    25812 => x"00000000", 25813 => x"00000000", 25814 => x"00000000",
    25815 => x"00000000", 25816 => x"00000000", 25817 => x"00000000",
    25818 => x"00000000", 25819 => x"00000000", 25820 => x"00000000",
    25821 => x"00000000", 25822 => x"00000000", 25823 => x"00000000",
    25824 => x"00000000", 25825 => x"00000000", 25826 => x"00000000",
    25827 => x"00000000", 25828 => x"00000000", 25829 => x"00000000",
    25830 => x"00000000", 25831 => x"00000000", 25832 => x"00000000",
    25833 => x"00000000", 25834 => x"00000000", 25835 => x"00000000",
    25836 => x"00000000", 25837 => x"00000000", 25838 => x"00000000",
    25839 => x"00000000", 25840 => x"00000000", 25841 => x"00000000",
    25842 => x"00000000", 25843 => x"00000000", 25844 => x"00000000",
    25845 => x"00000000", 25846 => x"00000000", 25847 => x"00000000",
    25848 => x"00000000", 25849 => x"00000000", 25850 => x"00000000",
    25851 => x"00000000", 25852 => x"00000000", 25853 => x"00000000",
    25854 => x"00000000", 25855 => x"00000000", 25856 => x"00000000",
    25857 => x"00000000", 25858 => x"00000000", 25859 => x"00000000",
    25860 => x"00000000", 25861 => x"00000000", 25862 => x"00000000",
    25863 => x"00000000", 25864 => x"00000000", 25865 => x"00000000",
    25866 => x"00000000", 25867 => x"00000000", 25868 => x"00000000",
    25869 => x"00000000", 25870 => x"00000000", 25871 => x"00000000",
    25872 => x"00000000", 25873 => x"00000000", 25874 => x"00000000",
    25875 => x"00000000", 25876 => x"00000000", 25877 => x"00000000",
    25878 => x"00000000", 25879 => x"00000000", 25880 => x"00000000",
    25881 => x"00000000", 25882 => x"00000000", 25883 => x"00000000",
    25884 => x"00000000", 25885 => x"00000000", 25886 => x"00000000",
    25887 => x"00000000", 25888 => x"00000000", 25889 => x"00000000",
    25890 => x"00000000", 25891 => x"00000000", 25892 => x"00000000",
    25893 => x"00000000", 25894 => x"00000000", 25895 => x"00000000",
    25896 => x"00000000", 25897 => x"00000000", 25898 => x"00000000",
    25899 => x"00000000", 25900 => x"00000000", 25901 => x"00000000",
    25902 => x"00000000", 25903 => x"00000000", 25904 => x"00000000",
    25905 => x"00000000", 25906 => x"00000000", 25907 => x"00000000",
    25908 => x"00000000", 25909 => x"00000000", 25910 => x"00000000",
    25911 => x"00000000", 25912 => x"00000000", 25913 => x"00000000",
    25914 => x"00000000", 25915 => x"00000000", 25916 => x"00000000",
    25917 => x"00000000", 25918 => x"00000000", 25919 => x"00000000",
    25920 => x"00000000", 25921 => x"00000000", 25922 => x"00000000",
    25923 => x"00000000", 25924 => x"00000000", 25925 => x"00000000",
    25926 => x"00000000", 25927 => x"00000000", 25928 => x"00000000",
    25929 => x"00000000", 25930 => x"00000000", 25931 => x"00000000",
    25932 => x"00000000", 25933 => x"00000000", 25934 => x"00000000",
    25935 => x"00000000", 25936 => x"00000000", 25937 => x"00000000",
    25938 => x"00000000", 25939 => x"00000000", 25940 => x"00000000",
    25941 => x"00000000", 25942 => x"00000000", 25943 => x"00000000",
    25944 => x"00000000", 25945 => x"00000000", 25946 => x"00000000",
    25947 => x"00000000", 25948 => x"00000000", 25949 => x"00000000",
    25950 => x"00000000", 25951 => x"00000000", 25952 => x"00000000",
    25953 => x"00000000", 25954 => x"00000000", 25955 => x"00000000",
    25956 => x"00000000", 25957 => x"00000000", 25958 => x"00000000",
    25959 => x"00000000", 25960 => x"00000000", 25961 => x"00000000",
    25962 => x"00000000", 25963 => x"00000000", 25964 => x"00000000",
    25965 => x"00000000", 25966 => x"00000000", 25967 => x"00000000",
    25968 => x"00000000", 25969 => x"00000000", 25970 => x"00000000",
    25971 => x"00000000", 25972 => x"00000000", 25973 => x"00000000",
    25974 => x"00000000", 25975 => x"00000000", 25976 => x"00000000",
    25977 => x"00000000", 25978 => x"00000000", 25979 => x"00000000",
    25980 => x"00000000", 25981 => x"00000000", 25982 => x"00000000",
    25983 => x"00000000", 25984 => x"00000000", 25985 => x"00000000",
    25986 => x"00000000", 25987 => x"00000000", 25988 => x"00000000",
    25989 => x"00000000", 25990 => x"00000000", 25991 => x"00000000",
    25992 => x"00000000", 25993 => x"00000000", 25994 => x"00000000",
    25995 => x"00000000", 25996 => x"00000000", 25997 => x"00000000",
    25998 => x"00000000", 25999 => x"00000000", 26000 => x"00000000",
    26001 => x"00000000", 26002 => x"00000000", 26003 => x"00000000",
    26004 => x"00000000", 26005 => x"00000000", 26006 => x"00000000",
    26007 => x"00000000", 26008 => x"00000000", 26009 => x"00000000",
    26010 => x"00000000", 26011 => x"00000000", 26012 => x"00000000",
    26013 => x"00000000", 26014 => x"00000000", 26015 => x"00000000",
    26016 => x"00000000", 26017 => x"00000000", 26018 => x"00000000",
    26019 => x"00000000", 26020 => x"00000000", 26021 => x"00000000",
    26022 => x"00000000", 26023 => x"00000000", 26024 => x"00000000",
    26025 => x"00000000", 26026 => x"00000000", 26027 => x"00000000",
    26028 => x"00000000", 26029 => x"00000000", 26030 => x"00000000",
    26031 => x"00000000", 26032 => x"00000000", 26033 => x"00000000",
    26034 => x"00000000", 26035 => x"00000000", 26036 => x"00000000",
    26037 => x"00000000", 26038 => x"00000000", 26039 => x"00000000",
    26040 => x"00000000", 26041 => x"00000000", 26042 => x"00000000",
    26043 => x"00000000", 26044 => x"00000000", 26045 => x"00000000",
    26046 => x"00000000", 26047 => x"00000000", 26048 => x"00000000",
    26049 => x"00000000", 26050 => x"00000000", 26051 => x"00000000",
    26052 => x"00000000", 26053 => x"00000000", 26054 => x"00000000",
    26055 => x"00000000", 26056 => x"00000000", 26057 => x"00000000",
    26058 => x"00000000", 26059 => x"00000000", 26060 => x"00000000",
    26061 => x"00000000", 26062 => x"00000000", 26063 => x"00000000",
    26064 => x"00000000", 26065 => x"00000000", 26066 => x"00000000",
    26067 => x"00000000", 26068 => x"00000000", 26069 => x"00000000",
    26070 => x"00000000", 26071 => x"00000000", 26072 => x"00000000",
    26073 => x"00000000", 26074 => x"00000000", 26075 => x"00000000",
    26076 => x"00000000", 26077 => x"00000000", 26078 => x"00000000",
    26079 => x"00000000", 26080 => x"00000000", 26081 => x"00000000",
    26082 => x"00000000", 26083 => x"00000000", 26084 => x"00000000",
    26085 => x"00000000", 26086 => x"00000000", 26087 => x"00000000",
    26088 => x"00000000", 26089 => x"00000000", 26090 => x"00000000",
    26091 => x"00000000", 26092 => x"00000000", 26093 => x"00000000",
    26094 => x"00000000", 26095 => x"00000000", 26096 => x"00000000",
    26097 => x"00000000", 26098 => x"00000000", 26099 => x"00000000",
    26100 => x"00000000", 26101 => x"00000000", 26102 => x"00000000",
    26103 => x"00000000", 26104 => x"00000000", 26105 => x"00000000",
    26106 => x"00000000", 26107 => x"00000000", 26108 => x"00000000",
    26109 => x"00000000", 26110 => x"00000000", 26111 => x"00000000",
    26112 => x"00000000", 26113 => x"00000000", 26114 => x"00000000",
    26115 => x"00000000", 26116 => x"00000000", 26117 => x"00000000",
    26118 => x"00000000", 26119 => x"00000000", 26120 => x"00000000",
    26121 => x"00000000", 26122 => x"00000000", 26123 => x"00000000",
    26124 => x"00000000", 26125 => x"00000000", 26126 => x"00000000",
    26127 => x"00000000", 26128 => x"00000000", 26129 => x"00000000",
    26130 => x"00000000", 26131 => x"00000000", 26132 => x"00000000",
    26133 => x"00000000", 26134 => x"00000000", 26135 => x"00000000",
    26136 => x"00000000", 26137 => x"00000000", 26138 => x"00000000",
    26139 => x"00000000", 26140 => x"00000000", 26141 => x"00000000",
    26142 => x"00000000", 26143 => x"00000000", 26144 => x"00000000",
    26145 => x"00000000", 26146 => x"00000000", 26147 => x"00000000",
    26148 => x"00000000", 26149 => x"00000000", 26150 => x"00000000",
    26151 => x"00000000", 26152 => x"00000000", 26153 => x"00000000",
    26154 => x"00000000", 26155 => x"00000000", 26156 => x"00000000",
    26157 => x"00000000", 26158 => x"00000000", 26159 => x"00000000",
    26160 => x"00000000", 26161 => x"00000000", 26162 => x"00000000",
    26163 => x"00000000", 26164 => x"00000000", 26165 => x"00000000",
    26166 => x"00000000", 26167 => x"00000000", 26168 => x"00000000",
    26169 => x"00000000", 26170 => x"00000000", 26171 => x"00000000",
    26172 => x"00000000", 26173 => x"00000000", 26174 => x"00000000",
    26175 => x"00000000", 26176 => x"00000000", 26177 => x"00000000",
    26178 => x"00000000", 26179 => x"00000000", 26180 => x"00000000",
    26181 => x"00000000", 26182 => x"00000000", 26183 => x"00000000",
    26184 => x"00000000", 26185 => x"00000000", 26186 => x"00000000",
    26187 => x"00000000", 26188 => x"00000000", 26189 => x"00000000",
    26190 => x"00000000", 26191 => x"00000000", 26192 => x"00000000",
    26193 => x"00000000", 26194 => x"00000000", 26195 => x"00000000",
    26196 => x"00000000", 26197 => x"00000000", 26198 => x"00000000",
    26199 => x"00000000", 26200 => x"00000000", 26201 => x"00000000",
    26202 => x"00000000", 26203 => x"00000000", 26204 => x"00000000",
    26205 => x"00000000", 26206 => x"00000000", 26207 => x"00000000",
    26208 => x"00000000", 26209 => x"00000000", 26210 => x"00000000",
    26211 => x"00000000", 26212 => x"00000000", 26213 => x"00000000",
    26214 => x"00000000", 26215 => x"00000000", 26216 => x"00000000",
    26217 => x"00000000", 26218 => x"00000000", 26219 => x"00000000",
    26220 => x"00000000", 26221 => x"00000000", 26222 => x"00000000",
    26223 => x"00000000", 26224 => x"00000000", 26225 => x"00000000",
    26226 => x"00000000", 26227 => x"00000000", 26228 => x"00000000",
    26229 => x"00000000", 26230 => x"00000000", 26231 => x"00000000",
    26232 => x"00000000", 26233 => x"00000000", 26234 => x"00000000",
    26235 => x"00000000", 26236 => x"00000000", 26237 => x"00000000",
    26238 => x"00000000", 26239 => x"00000000", 26240 => x"00000000",
    26241 => x"00000000", 26242 => x"00000000", 26243 => x"00000000",
    26244 => x"00000000", 26245 => x"00000000", 26246 => x"00000000",
    26247 => x"00000000", 26248 => x"00000000", 26249 => x"00000000",
    26250 => x"00000000", 26251 => x"00000000", 26252 => x"00000000",
    26253 => x"00000000", 26254 => x"00000000", 26255 => x"00000000",
    26256 => x"00000000", 26257 => x"00000000", 26258 => x"00000000",
    26259 => x"00000000", 26260 => x"00000000", 26261 => x"00000000",
    26262 => x"00000000", 26263 => x"00000000", 26264 => x"00000000",
    26265 => x"00000000", 26266 => x"00000000", 26267 => x"00000000",
    26268 => x"00000000", 26269 => x"00000000", 26270 => x"00000000",
    26271 => x"00000000", 26272 => x"00000000", 26273 => x"00000000",
    26274 => x"00000000", 26275 => x"00000000", 26276 => x"00000000",
    26277 => x"00000000", 26278 => x"00000000", 26279 => x"00000000",
    26280 => x"00000000", 26281 => x"00000000", 26282 => x"00000000",
    26283 => x"00000000", 26284 => x"00000000", 26285 => x"00000000",
    26286 => x"00000000", 26287 => x"00000000", 26288 => x"00000000",
    26289 => x"00000000", 26290 => x"00000000", 26291 => x"00000000",
    26292 => x"00000000", 26293 => x"00000000", 26294 => x"00000000",
    26295 => x"00000000", 26296 => x"00000000", 26297 => x"00000000",
    26298 => x"00000000", 26299 => x"00000000", 26300 => x"00000000",
    26301 => x"00000000", 26302 => x"00000000", 26303 => x"00000000",
    26304 => x"00000000", 26305 => x"00000000", 26306 => x"00000000",
    26307 => x"00000000", 26308 => x"00000000", 26309 => x"00000000",
    26310 => x"00000000", 26311 => x"00000000", 26312 => x"00000000",
    26313 => x"00000000", 26314 => x"00000000", 26315 => x"00000000",
    26316 => x"00000000", 26317 => x"00000000", 26318 => x"00000000",
    26319 => x"00000000", 26320 => x"00000000", 26321 => x"00000000",
    26322 => x"00000000", 26323 => x"00000000", 26324 => x"00000000",
    26325 => x"00000000", 26326 => x"00000000", 26327 => x"00000000",
    26328 => x"00000000", 26329 => x"00000000", 26330 => x"00000000",
    26331 => x"00000000", 26332 => x"00000000", 26333 => x"00000000",
    26334 => x"00000000", 26335 => x"00000000", 26336 => x"00000000",
    26337 => x"00000000", 26338 => x"00000000", 26339 => x"00000000",
    26340 => x"00000000", 26341 => x"00000000", 26342 => x"00000000",
    26343 => x"00000000", 26344 => x"00000000", 26345 => x"00000000",
    26346 => x"00000000", 26347 => x"00000000", 26348 => x"00000000",
    26349 => x"00000000", 26350 => x"00000000", 26351 => x"00000000",
    26352 => x"00000000", 26353 => x"00000000", 26354 => x"00000000",
    26355 => x"00000000", 26356 => x"00000000", 26357 => x"00000000",
    26358 => x"00000000", 26359 => x"00000000", 26360 => x"00000000",
    26361 => x"00000000", 26362 => x"00000000", 26363 => x"00000000",
    26364 => x"00000000", 26365 => x"00000000", 26366 => x"00000000",
    26367 => x"00000000", 26368 => x"00000000", 26369 => x"00000000",
    26370 => x"00000000", 26371 => x"00000000", 26372 => x"00000000",
    26373 => x"00000000", 26374 => x"00000000", 26375 => x"00000000",
    26376 => x"00000000", 26377 => x"00000000", 26378 => x"00000000",
    26379 => x"00000000", 26380 => x"00000000", 26381 => x"00000000",
    26382 => x"00000000", 26383 => x"00000000", 26384 => x"00000000",
    26385 => x"00000000", 26386 => x"00000000", 26387 => x"00000000",
    26388 => x"00000000", 26389 => x"00000000", 26390 => x"00000000",
    26391 => x"00000000", 26392 => x"00000000", 26393 => x"00000000",
    26394 => x"00000000", 26395 => x"00000000", 26396 => x"00000000",
    26397 => x"00000000", 26398 => x"00000000", 26399 => x"00000000",
    26400 => x"00000000", 26401 => x"00000000", 26402 => x"00000000",
    26403 => x"00000000", 26404 => x"00000000", 26405 => x"00000000",
    26406 => x"00000000", 26407 => x"00000000", 26408 => x"00000000",
    26409 => x"00000000", 26410 => x"00000000", 26411 => x"00000000",
    26412 => x"00000000", 26413 => x"00000000", 26414 => x"00000000",
    26415 => x"00000000", 26416 => x"00000000", 26417 => x"00000000",
    26418 => x"00000000", 26419 => x"00000000", 26420 => x"00000000",
    26421 => x"00000000", 26422 => x"00000000", 26423 => x"00000000",
    26424 => x"00000000", 26425 => x"00000000", 26426 => x"00000000",
    26427 => x"00000000", 26428 => x"00000000", 26429 => x"00000000",
    26430 => x"00000000", 26431 => x"00000000", 26432 => x"00000000",
    26433 => x"00000000", 26434 => x"00000000", 26435 => x"00000000",
    26436 => x"00000000", 26437 => x"00000000", 26438 => x"00000000",
    26439 => x"00000000", 26440 => x"00000000", 26441 => x"00000000",
    26442 => x"00000000", 26443 => x"00000000", 26444 => x"00000000",
    26445 => x"00000000", 26446 => x"00000000", 26447 => x"00000000",
    26448 => x"00000000", 26449 => x"00000000", 26450 => x"00000000",
    26451 => x"00000000", 26452 => x"00000000", 26453 => x"00000000",
    26454 => x"00000000", 26455 => x"00000000", 26456 => x"00000000",
    26457 => x"00000000", 26458 => x"00000000", 26459 => x"00000000",
    26460 => x"00000000", 26461 => x"00000000", 26462 => x"00000000",
    26463 => x"00000000", 26464 => x"00000000", 26465 => x"00000000",
    26466 => x"00000000", 26467 => x"00000000", 26468 => x"00000000",
    26469 => x"00000000", 26470 => x"00000000", 26471 => x"00000000",
    26472 => x"00000000", 26473 => x"00000000", 26474 => x"00000000",
    26475 => x"00000000", 26476 => x"00000000", 26477 => x"00000000",
    26478 => x"00000000", 26479 => x"00000000", 26480 => x"00000000",
    26481 => x"00000000", 26482 => x"00000000", 26483 => x"00000000",
    26484 => x"00000000", 26485 => x"00000000", 26486 => x"00000000",
    26487 => x"00000000", 26488 => x"00000000", 26489 => x"00000000",
    26490 => x"00000000", 26491 => x"00000000", 26492 => x"00000000",
    26493 => x"00000000", 26494 => x"00000000", 26495 => x"00000000",
    26496 => x"00000000", 26497 => x"00000000", 26498 => x"00000000",
    26499 => x"00000000", 26500 => x"00000000", 26501 => x"00000000",
    26502 => x"00000000", 26503 => x"00000000", 26504 => x"00000000",
    26505 => x"00000000", 26506 => x"00000000", 26507 => x"00000000",
    26508 => x"00000000", 26509 => x"00000000", 26510 => x"00000000",
    26511 => x"00000000", 26512 => x"00000000", 26513 => x"00000000",
    26514 => x"00000000", 26515 => x"00000000", 26516 => x"00000000",
    26517 => x"00000000", 26518 => x"00000000", 26519 => x"00000000",
    26520 => x"00000000", 26521 => x"00000000", 26522 => x"00000000",
    26523 => x"00000000", 26524 => x"00000000", 26525 => x"00000000",
    26526 => x"00000000", 26527 => x"00000000", 26528 => x"00000000",
    26529 => x"00000000", 26530 => x"00000000", 26531 => x"00000000",
    26532 => x"00000000", 26533 => x"00000000", 26534 => x"00000000",
    26535 => x"00000000", 26536 => x"00000000", 26537 => x"00000000",
    26538 => x"00000000", 26539 => x"00000000", 26540 => x"00000000",
    26541 => x"00000000", 26542 => x"00000000", 26543 => x"00000000",
    26544 => x"00000000", 26545 => x"00000000", 26546 => x"00000000",
    26547 => x"00000000", 26548 => x"00000000", 26549 => x"00000000",
    26550 => x"00000000", 26551 => x"00000000", 26552 => x"00000000",
    26553 => x"00000000", 26554 => x"00000000", 26555 => x"00000000",
    26556 => x"00000000", 26557 => x"00000000", 26558 => x"00000000",
    26559 => x"00000000", 26560 => x"00000000", 26561 => x"00000000",
    26562 => x"00000000", 26563 => x"00000000", 26564 => x"00000000",
    26565 => x"00000000", 26566 => x"00000000", 26567 => x"00000000",
    26568 => x"00000000", 26569 => x"00000000", 26570 => x"00000000",
    26571 => x"00000000", 26572 => x"00000000", 26573 => x"00000000",
    26574 => x"00000000", 26575 => x"00000000", 26576 => x"00000000",
    26577 => x"00000000", 26578 => x"00000000", 26579 => x"00000000",
    26580 => x"00000000", 26581 => x"00000000", 26582 => x"00000000",
    26583 => x"00000000", 26584 => x"00000000", 26585 => x"00000000",
    26586 => x"00000000", 26587 => x"00000000", 26588 => x"00000000",
    26589 => x"00000000", 26590 => x"00000000", 26591 => x"00000000",
    26592 => x"00000000", 26593 => x"00000000", 26594 => x"00000000",
    26595 => x"00000000", 26596 => x"00000000", 26597 => x"00000000",
    26598 => x"00000000", 26599 => x"00000000", 26600 => x"00000000",
    26601 => x"00000000", 26602 => x"00000000", 26603 => x"00000000",
    26604 => x"00000000", 26605 => x"00000000", 26606 => x"00000000",
    26607 => x"00000000", 26608 => x"00000000", 26609 => x"00000000",
    26610 => x"00000000", 26611 => x"00000000", 26612 => x"00000000",
    26613 => x"00000000", 26614 => x"00000000", 26615 => x"00000000",
    26616 => x"00000000", 26617 => x"00000000", 26618 => x"00000000",
    26619 => x"00000000", 26620 => x"00000000", 26621 => x"00000000",
    26622 => x"00000000", 26623 => x"00000000", 26624 => x"00000000",
    26625 => x"00000000", 26626 => x"00000000", 26627 => x"00000000",
    26628 => x"00000000", 26629 => x"00000000", 26630 => x"00000000",
    26631 => x"00000000", 26632 => x"00000000", 26633 => x"00000000",
    26634 => x"00000000", 26635 => x"00000000", 26636 => x"00000000",
    26637 => x"00000000", 26638 => x"00000000", 26639 => x"00000000",
    26640 => x"00000000", 26641 => x"00000000", 26642 => x"00000000",
    26643 => x"00000000", 26644 => x"00000000", 26645 => x"00000000",
    26646 => x"00000000", 26647 => x"00000000", 26648 => x"00000000",
    26649 => x"00000000", 26650 => x"00000000", 26651 => x"00000000",
    26652 => x"00000000", 26653 => x"00000000", 26654 => x"00000000",
    26655 => x"00000000", 26656 => x"00000000", 26657 => x"00000000",
    26658 => x"00000000", 26659 => x"00000000", 26660 => x"00000000",
    26661 => x"00000000", 26662 => x"00000000", 26663 => x"00000000",
    26664 => x"00000000", 26665 => x"00000000", 26666 => x"00000000",
    26667 => x"00000000", 26668 => x"00000000", 26669 => x"00000000",
    26670 => x"00000000", 26671 => x"00000000", 26672 => x"00000000",
    26673 => x"00000000", 26674 => x"00000000", 26675 => x"00000000",
    26676 => x"00000000", 26677 => x"00000000", 26678 => x"00000000",
    26679 => x"00000000", 26680 => x"00000000", 26681 => x"00000000",
    26682 => x"00000000", 26683 => x"00000000", 26684 => x"00000000",
    26685 => x"00000000", 26686 => x"00000000", 26687 => x"00000000",
    26688 => x"00000000", 26689 => x"00000000", 26690 => x"00000000",
    26691 => x"00000000", 26692 => x"00000000", 26693 => x"00000000",
    26694 => x"00000000", 26695 => x"00000000", 26696 => x"00000000",
    26697 => x"00000000", 26698 => x"00000000", 26699 => x"00000000",
    26700 => x"00000000", 26701 => x"00000000", 26702 => x"00000000",
    26703 => x"00000000", 26704 => x"00000000", 26705 => x"00000000",
    26706 => x"00000000", 26707 => x"00000000", 26708 => x"00000000",
    26709 => x"00000000", 26710 => x"00000000", 26711 => x"00000000",
    26712 => x"00000000", 26713 => x"00000000", 26714 => x"00000000",
    26715 => x"00000000", 26716 => x"00000000", 26717 => x"00000000",
    26718 => x"00000000", 26719 => x"00000000", 26720 => x"00000000",
    26721 => x"00000000", 26722 => x"00000000", 26723 => x"00000000",
    26724 => x"00000000", 26725 => x"00000000", 26726 => x"00000000",
    26727 => x"00000000", 26728 => x"00000000", 26729 => x"00000000",
    26730 => x"00000000", 26731 => x"00000000", 26732 => x"00000000",
    26733 => x"00000000", 26734 => x"00000000", 26735 => x"00000000",
    26736 => x"00000000", 26737 => x"00000000", 26738 => x"00000000",
    26739 => x"00000000", 26740 => x"00000000", 26741 => x"00000000",
    26742 => x"00000000", 26743 => x"00000000", 26744 => x"00000000",
    26745 => x"00000000", 26746 => x"00000000", 26747 => x"00000000",
    26748 => x"00000000", 26749 => x"00000000", 26750 => x"00000000",
    26751 => x"00000000", 26752 => x"00000000", 26753 => x"00000000",
    26754 => x"00000000", 26755 => x"00000000", 26756 => x"00000000",
    26757 => x"00000000", 26758 => x"00000000", 26759 => x"00000000",
    26760 => x"00000000", 26761 => x"00000000", 26762 => x"00000000",
    26763 => x"00000000", 26764 => x"00000000", 26765 => x"00000000",
    26766 => x"00000000", 26767 => x"00000000", 26768 => x"00000000",
    26769 => x"00000000", 26770 => x"00000000", 26771 => x"00000000",
    26772 => x"00000000", 26773 => x"00000000", 26774 => x"00000000",
    26775 => x"00000000", 26776 => x"00000000", 26777 => x"00000000",
    26778 => x"00000000", 26779 => x"00000000", 26780 => x"00000000",
    26781 => x"00000000", 26782 => x"00000000", 26783 => x"00000000",
    26784 => x"00000000", 26785 => x"00000000", 26786 => x"00000000",
    26787 => x"00000000", 26788 => x"00000000", 26789 => x"00000000",
    26790 => x"00000000", 26791 => x"00000000", 26792 => x"00000000",
    26793 => x"00000000", 26794 => x"00000000", 26795 => x"00000000",
    26796 => x"00000000", 26797 => x"00000000", 26798 => x"00000000",
    26799 => x"00000000", 26800 => x"00000000", 26801 => x"00000000",
    26802 => x"00000000", 26803 => x"00000000", 26804 => x"00000000",
    26805 => x"00000000", 26806 => x"00000000", 26807 => x"00000000",
    26808 => x"00000000", 26809 => x"00000000", 26810 => x"00000000",
    26811 => x"00000000", 26812 => x"00000000", 26813 => x"00000000",
    26814 => x"00000000", 26815 => x"00000000", 26816 => x"00000000",
    26817 => x"00000000", 26818 => x"00000000", 26819 => x"00000000",
    26820 => x"00000000", 26821 => x"00000000", 26822 => x"00000000",
    26823 => x"00000000", 26824 => x"00000000", 26825 => x"00000000",
    26826 => x"00000000", 26827 => x"00000000", 26828 => x"00000000",
    26829 => x"00000000", 26830 => x"00000000", 26831 => x"00000000",
    26832 => x"00000000", 26833 => x"00000000", 26834 => x"00000000",
    26835 => x"00000000", 26836 => x"00000000", 26837 => x"00000000",
    26838 => x"00000000", 26839 => x"00000000", 26840 => x"00000000",
    26841 => x"00000000", 26842 => x"00000000", 26843 => x"00000000",
    26844 => x"00000000", 26845 => x"00000000", 26846 => x"00000000",
    26847 => x"00000000", 26848 => x"00000000", 26849 => x"00000000",
    26850 => x"00000000", 26851 => x"00000000", 26852 => x"00000000",
    26853 => x"00000000", 26854 => x"00000000", 26855 => x"00000000",
    26856 => x"00000000", 26857 => x"00000000", 26858 => x"00000000",
    26859 => x"00000000", 26860 => x"00000000", 26861 => x"00000000",
    26862 => x"00000000", 26863 => x"00000000", 26864 => x"00000000",
    26865 => x"00000000", 26866 => x"00000000", 26867 => x"00000000",
    26868 => x"00000000", 26869 => x"00000000", 26870 => x"00000000",
    26871 => x"00000000", 26872 => x"00000000", 26873 => x"00000000",
    26874 => x"00000000", 26875 => x"00000000", 26876 => x"00000000",
    26877 => x"00000000", 26878 => x"00000000", 26879 => x"00000000",
    26880 => x"00000000", 26881 => x"00000000", 26882 => x"00000000",
    26883 => x"00000000", 26884 => x"00000000", 26885 => x"00000000",
    26886 => x"00000000", 26887 => x"00000000", 26888 => x"00000000",
    26889 => x"00000000", 26890 => x"00000000", 26891 => x"00000000",
    26892 => x"00000000", 26893 => x"00000000", 26894 => x"00000000",
    26895 => x"00000000", 26896 => x"00000000", 26897 => x"00000000",
    26898 => x"00000000", 26899 => x"00000000", 26900 => x"00000000",
    26901 => x"00000000", 26902 => x"00000000", 26903 => x"00000000",
    26904 => x"00000000", 26905 => x"00000000", 26906 => x"00000000",
    26907 => x"00000000", 26908 => x"00000000", 26909 => x"00000000",
    26910 => x"00000000", 26911 => x"00000000", 26912 => x"00000000",
    26913 => x"00000000", 26914 => x"00000000", 26915 => x"00000000",
    26916 => x"00000000", 26917 => x"00000000", 26918 => x"00000000",
    26919 => x"00000000", 26920 => x"00000000", 26921 => x"00000000",
    26922 => x"00000000", 26923 => x"00000000", 26924 => x"00000000",
    26925 => x"00000000", 26926 => x"00000000", 26927 => x"00000000",
    26928 => x"00000000", 26929 => x"00000000", 26930 => x"00000000",
    26931 => x"00000000", 26932 => x"00000000", 26933 => x"00000000",
    26934 => x"00000000", 26935 => x"00000000", 26936 => x"00000000",
    26937 => x"00000000", 26938 => x"00000000", 26939 => x"00000000",
    26940 => x"00000000", 26941 => x"00000000", 26942 => x"00000000",
    26943 => x"00000000", 26944 => x"00000000", 26945 => x"00000000",
    26946 => x"00000000", 26947 => x"00000000", 26948 => x"00000000",
    26949 => x"00000000", 26950 => x"00000000", 26951 => x"00000000",
    26952 => x"00000000", 26953 => x"00000000", 26954 => x"00000000",
    26955 => x"00000000", 26956 => x"00000000", 26957 => x"00000000",
    26958 => x"00000000", 26959 => x"00000000", 26960 => x"00000000",
    26961 => x"00000000", 26962 => x"00000000", 26963 => x"00000000",
    26964 => x"00000000", 26965 => x"00000000", 26966 => x"00000000",
    26967 => x"00000000", 26968 => x"00000000", 26969 => x"00000000",
    26970 => x"00000000", 26971 => x"00000000", 26972 => x"00000000",
    26973 => x"00000000", 26974 => x"00000000", 26975 => x"00000000",
    26976 => x"00000000", 26977 => x"00000000", 26978 => x"00000000",
    26979 => x"00000000", 26980 => x"00000000", 26981 => x"00000000",
    26982 => x"00000000", 26983 => x"00000000", 26984 => x"00000000",
    26985 => x"00000000", 26986 => x"00000000", 26987 => x"00000000",
    26988 => x"00000000", 26989 => x"00000000", 26990 => x"00000000",
    26991 => x"00000000", 26992 => x"00000000", 26993 => x"00000000",
    26994 => x"00000000", 26995 => x"00000000", 26996 => x"00000000",
    26997 => x"00000000", 26998 => x"00000000", 26999 => x"00000000",
    27000 => x"00000000", 27001 => x"00000000", 27002 => x"00000000",
    27003 => x"00000000", 27004 => x"00000000", 27005 => x"00000000",
    27006 => x"00000000", 27007 => x"00000000", 27008 => x"00000000",
    27009 => x"00000000", 27010 => x"00000000", 27011 => x"00000000",
    27012 => x"00000000", 27013 => x"00000000", 27014 => x"00000000",
    27015 => x"00000000", 27016 => x"00000000", 27017 => x"00000000",
    27018 => x"00000000", 27019 => x"00000000", 27020 => x"00000000",
    27021 => x"00000000", 27022 => x"00000000", 27023 => x"00000000",
    27024 => x"00000000", 27025 => x"00000000", 27026 => x"00000000",
    27027 => x"00000000", 27028 => x"00000000", 27029 => x"00000000",
    27030 => x"00000000", 27031 => x"00000000", 27032 => x"00000000",
    27033 => x"00000000", 27034 => x"00000000", 27035 => x"00000000",
    27036 => x"00000000", 27037 => x"00000000", 27038 => x"00000000",
    27039 => x"00000000", 27040 => x"00000000", 27041 => x"00000000",
    27042 => x"00000000", 27043 => x"00000000", 27044 => x"00000000",
    27045 => x"00000000", 27046 => x"00000000", 27047 => x"00000000",
    27048 => x"00000000", 27049 => x"00000000", 27050 => x"00000000",
    27051 => x"00000000", 27052 => x"00000000", 27053 => x"00000000",
    27054 => x"00000000", 27055 => x"00000000", 27056 => x"00000000",
    27057 => x"00000000", 27058 => x"00000000", 27059 => x"00000000",
    27060 => x"00000000", 27061 => x"00000000", 27062 => x"00000000",
    27063 => x"00000000", 27064 => x"00000000", 27065 => x"00000000",
    27066 => x"00000000", 27067 => x"00000000", 27068 => x"00000000",
    27069 => x"00000000", 27070 => x"00000000", 27071 => x"00000000",
    27072 => x"00000000", 27073 => x"00000000", 27074 => x"00000000",
    27075 => x"00000000", 27076 => x"00000000", 27077 => x"00000000",
    27078 => x"00000000", 27079 => x"00000000", 27080 => x"00000000",
    27081 => x"00000000", 27082 => x"00000000", 27083 => x"00000000",
    27084 => x"00000000", 27085 => x"00000000", 27086 => x"00000000",
    27087 => x"00000000", 27088 => x"00000000", 27089 => x"00000000",
    27090 => x"00000000", 27091 => x"00000000", 27092 => x"00000000",
    27093 => x"00000000", 27094 => x"00000000", 27095 => x"00000000",
    27096 => x"00000000", 27097 => x"00000000", 27098 => x"00000000",
    27099 => x"00000000", 27100 => x"00000000", 27101 => x"00000000",
    27102 => x"00000000", 27103 => x"00000000", 27104 => x"00000000",
    27105 => x"00000000", 27106 => x"00000000", 27107 => x"00000000",
    27108 => x"00000000", 27109 => x"00000000", 27110 => x"00000000",
    27111 => x"00000000", 27112 => x"00000000", 27113 => x"00000000",
    27114 => x"00000000", 27115 => x"00000000", 27116 => x"00000000",
    27117 => x"00000000", 27118 => x"00000000", 27119 => x"00000000",
    27120 => x"00000000", 27121 => x"00000000", 27122 => x"00000000",
    27123 => x"00000000", 27124 => x"00000000", 27125 => x"00000000",
    27126 => x"00000000", 27127 => x"00000000", 27128 => x"00000000",
    27129 => x"00000000", 27130 => x"00000000", 27131 => x"00000000",
    27132 => x"00000000", 27133 => x"00000000", 27134 => x"00000000",
    27135 => x"00000000", 27136 => x"00000000", 27137 => x"00000000",
    27138 => x"00000000", 27139 => x"00000000", 27140 => x"00000000",
    27141 => x"00000000", 27142 => x"00000000", 27143 => x"00000000",
    27144 => x"00000000", 27145 => x"00000000", 27146 => x"00000000",
    27147 => x"00000000", 27148 => x"00000000", 27149 => x"00000000",
    27150 => x"00000000", 27151 => x"00000000", 27152 => x"00000000",
    27153 => x"00000000", 27154 => x"00000000", 27155 => x"00000000",
    27156 => x"00000000", 27157 => x"00000000", 27158 => x"00000000",
    27159 => x"00000000", 27160 => x"00000000", 27161 => x"00000000",
    27162 => x"00000000", 27163 => x"00000000", 27164 => x"00000000",
    27165 => x"00000000", 27166 => x"00000000", 27167 => x"00000000",
    27168 => x"00000000", 27169 => x"00000000", 27170 => x"00000000",
    27171 => x"00000000", 27172 => x"00000000", 27173 => x"00000000",
    27174 => x"00000000", 27175 => x"00000000", 27176 => x"00000000",
    27177 => x"00000000", 27178 => x"00000000", 27179 => x"00000000",
    27180 => x"00000000", 27181 => x"00000000", 27182 => x"00000000",
    27183 => x"00000000", 27184 => x"00000000", 27185 => x"00000000",
    27186 => x"00000000", 27187 => x"00000000", 27188 => x"00000000",
    27189 => x"00000000", 27190 => x"00000000", 27191 => x"00000000",
    27192 => x"00000000", 27193 => x"00000000", 27194 => x"00000000",
    27195 => x"00000000", 27196 => x"00000000", 27197 => x"00000000",
    27198 => x"00000000", 27199 => x"00000000", 27200 => x"00000000",
    27201 => x"00000000", 27202 => x"00000000", 27203 => x"00000000",
    27204 => x"00000000", 27205 => x"00000000", 27206 => x"00000000",
    27207 => x"00000000", 27208 => x"00000000", 27209 => x"00000000",
    27210 => x"00000000", 27211 => x"00000000", 27212 => x"00000000",
    27213 => x"00000000", 27214 => x"00000000", 27215 => x"00000000",
    27216 => x"00000000", 27217 => x"00000000", 27218 => x"00000000",
    27219 => x"00000000", 27220 => x"00000000", 27221 => x"00000000",
    27222 => x"00000000", 27223 => x"00000000", 27224 => x"00000000",
    27225 => x"00000000", 27226 => x"00000000", 27227 => x"00000000",
    27228 => x"00000000", 27229 => x"00000000", 27230 => x"00000000",
    27231 => x"00000000", 27232 => x"00000000", 27233 => x"00000000",
    27234 => x"00000000", 27235 => x"00000000", 27236 => x"00000000",
    27237 => x"00000000", 27238 => x"00000000", 27239 => x"00000000",
    27240 => x"00000000", 27241 => x"00000000", 27242 => x"00000000",
    27243 => x"00000000", 27244 => x"00000000", 27245 => x"00000000",
    27246 => x"00000000", 27247 => x"00000000", 27248 => x"00000000",
    27249 => x"00000000", 27250 => x"00000000", 27251 => x"00000000",
    27252 => x"00000000", 27253 => x"00000000", 27254 => x"00000000",
    27255 => x"00000000", 27256 => x"00000000", 27257 => x"00000000",
    27258 => x"00000000", 27259 => x"00000000", 27260 => x"00000000",
    27261 => x"00000000", 27262 => x"00000000", 27263 => x"00000000",
    27264 => x"00000000", 27265 => x"00000000", 27266 => x"00000000",
    27267 => x"00000000", 27268 => x"00000000", 27269 => x"00000000",
    27270 => x"00000000", 27271 => x"00000000", 27272 => x"00000000",
    27273 => x"00000000", 27274 => x"00000000", 27275 => x"00000000",
    27276 => x"00000000", 27277 => x"00000000", 27278 => x"00000000",
    27279 => x"00000000", 27280 => x"00000000", 27281 => x"00000000",
    27282 => x"00000000", 27283 => x"00000000", 27284 => x"00000000",
    27285 => x"00000000", 27286 => x"00000000", 27287 => x"00000000",
    27288 => x"00000000", 27289 => x"00000000", 27290 => x"00000000",
    27291 => x"00000000", 27292 => x"00000000", 27293 => x"00000000",
    27294 => x"00000000", 27295 => x"00000000", 27296 => x"00000000",
    27297 => x"00000000", 27298 => x"00000000", 27299 => x"00000000",
    27300 => x"00000000", 27301 => x"00000000", 27302 => x"00000000",
    27303 => x"00000000", 27304 => x"00000000", 27305 => x"00000000",
    27306 => x"00000000", 27307 => x"00000000", 27308 => x"00000000",
    27309 => x"00000000", 27310 => x"00000000", 27311 => x"00000000",
    27312 => x"00000000", 27313 => x"00000000", 27314 => x"00000000",
    27315 => x"00000000", 27316 => x"00000000", 27317 => x"00000000",
    27318 => x"00000000", 27319 => x"00000000", 27320 => x"00000000",
    27321 => x"00000000", 27322 => x"00000000", 27323 => x"00000000",
    27324 => x"00000000", 27325 => x"00000000", 27326 => x"00000000",
    27327 => x"00000000", 27328 => x"00000000", 27329 => x"00000000",
    27330 => x"00000000", 27331 => x"00000000", 27332 => x"00000000",
    27333 => x"00000000", 27334 => x"00000000", 27335 => x"00000000",
    27336 => x"00000000", 27337 => x"00000000", 27338 => x"00000000",
    27339 => x"00000000", 27340 => x"00000000", 27341 => x"00000000",
    27342 => x"00000000", 27343 => x"00000000", 27344 => x"00000000",
    27345 => x"00000000", 27346 => x"00000000", 27347 => x"00000000",
    27348 => x"00000000", 27349 => x"00000000", 27350 => x"00000000",
    27351 => x"00000000", 27352 => x"00000000", 27353 => x"00000000",
    27354 => x"00000000", 27355 => x"00000000", 27356 => x"00000000",
    27357 => x"00000000", 27358 => x"00000000", 27359 => x"00000000",
    27360 => x"00000000", 27361 => x"00000000", 27362 => x"00000000",
    27363 => x"00000000", 27364 => x"00000000", 27365 => x"00000000",
    27366 => x"00000000", 27367 => x"00000000", 27368 => x"00000000",
    27369 => x"00000000", 27370 => x"00000000", 27371 => x"00000000",
    27372 => x"00000000", 27373 => x"00000000", 27374 => x"00000000",
    27375 => x"00000000", 27376 => x"00000000", 27377 => x"00000000",
    27378 => x"00000000", 27379 => x"00000000", 27380 => x"00000000",
    27381 => x"00000000", 27382 => x"00000000", 27383 => x"00000000",
    27384 => x"00000000", 27385 => x"00000000", 27386 => x"00000000",
    27387 => x"00000000", 27388 => x"00000000", 27389 => x"00000000",
    27390 => x"00000000", 27391 => x"00000000", 27392 => x"00000000",
    27393 => x"00000000", 27394 => x"00000000", 27395 => x"00000000",
    27396 => x"00000000", 27397 => x"00000000", 27398 => x"00000000",
    27399 => x"00000000", 27400 => x"00000000", 27401 => x"00000000",
    27402 => x"00000000", 27403 => x"00000000", 27404 => x"00000000",
    27405 => x"00000000", 27406 => x"00000000", 27407 => x"00000000",
    27408 => x"00000000", 27409 => x"00000000", 27410 => x"00000000",
    27411 => x"00000000", 27412 => x"00000000", 27413 => x"00000000",
    27414 => x"00000000", 27415 => x"00000000", 27416 => x"00000000",
    27417 => x"00000000", 27418 => x"00000000", 27419 => x"00000000",
    27420 => x"00000000", 27421 => x"00000000", 27422 => x"00000000",
    27423 => x"00000000", 27424 => x"00000000", 27425 => x"00000000",
    27426 => x"00000000", 27427 => x"00000000", 27428 => x"00000000",
    27429 => x"00000000", 27430 => x"00000000", 27431 => x"00000000",
    27432 => x"00000000", 27433 => x"00000000", 27434 => x"00000000",
    27435 => x"00000000", 27436 => x"00000000", 27437 => x"00000000",
    27438 => x"00000000", 27439 => x"00000000", 27440 => x"00000000",
    27441 => x"00000000", 27442 => x"00000000", 27443 => x"00000000",
    27444 => x"00000000", 27445 => x"00000000", 27446 => x"00000000",
    27447 => x"00000000", 27448 => x"00000000", 27449 => x"00000000",
    27450 => x"00000000", 27451 => x"00000000", 27452 => x"00000000",
    27453 => x"00000000", 27454 => x"00000000", 27455 => x"00000000",
    27456 => x"00000000", 27457 => x"00000000", 27458 => x"00000000",
    27459 => x"00000000", 27460 => x"00000000", 27461 => x"00000000",
    27462 => x"00000000", 27463 => x"00000000", 27464 => x"00000000",
    27465 => x"00000000", 27466 => x"00000000", 27467 => x"00000000",
    27468 => x"00000000", 27469 => x"00000000", 27470 => x"00000000",
    27471 => x"00000000", 27472 => x"00000000", 27473 => x"00000000",
    27474 => x"00000000", 27475 => x"00000000", 27476 => x"00000000",
    27477 => x"00000000", 27478 => x"00000000", 27479 => x"00000000",
    27480 => x"00000000", 27481 => x"00000000", 27482 => x"00000000",
    27483 => x"00000000", 27484 => x"00000000", 27485 => x"00000000",
    27486 => x"00000000", 27487 => x"00000000", 27488 => x"00000000",
    27489 => x"00000000", 27490 => x"00000000", 27491 => x"00000000",
    27492 => x"00000000", 27493 => x"00000000", 27494 => x"00000000",
    27495 => x"00000000", 27496 => x"00000000", 27497 => x"00000000",
    27498 => x"00000000", 27499 => x"00000000", 27500 => x"00000000",
    27501 => x"00000000", 27502 => x"00000000", 27503 => x"00000000",
    27504 => x"00000000", 27505 => x"00000000", 27506 => x"00000000",
    27507 => x"00000000", 27508 => x"00000000", 27509 => x"00000000",
    27510 => x"00000000", 27511 => x"00000000", 27512 => x"00000000",
    27513 => x"00000000", 27514 => x"00000000", 27515 => x"00000000",
    27516 => x"00000000", 27517 => x"00000000", 27518 => x"00000000",
    27519 => x"00000000", 27520 => x"00000000", 27521 => x"00000000",
    27522 => x"00000000", 27523 => x"00000000", 27524 => x"00000000",
    27525 => x"00000000", 27526 => x"00000000", 27527 => x"00000000",
    27528 => x"00000000", 27529 => x"00000000", 27530 => x"00000000",
    27531 => x"00000000", 27532 => x"00000000", 27533 => x"00000000",
    27534 => x"00000000", 27535 => x"00000000", 27536 => x"00000000",
    27537 => x"00000000", 27538 => x"00000000", 27539 => x"00000000",
    27540 => x"00000000", 27541 => x"00000000", 27542 => x"00000000",
    27543 => x"00000000", 27544 => x"00000000", 27545 => x"00000000",
    27546 => x"00000000", 27547 => x"00000000", 27548 => x"00000000",
    27549 => x"00000000", 27550 => x"00000000", 27551 => x"00000000",
    27552 => x"00000000", 27553 => x"00000000", 27554 => x"00000000",
    27555 => x"00000000", 27556 => x"00000000", 27557 => x"00000000",
    27558 => x"00000000", 27559 => x"00000000", 27560 => x"00000000",
    27561 => x"00000000", 27562 => x"00000000", 27563 => x"00000000",
    27564 => x"00000000", 27565 => x"00000000", 27566 => x"00000000",
    27567 => x"00000000", 27568 => x"00000000", 27569 => x"00000000",
    27570 => x"00000000", 27571 => x"00000000", 27572 => x"00000000",
    27573 => x"00000000", 27574 => x"00000000", 27575 => x"00000000",
    27576 => x"00000000", 27577 => x"00000000", 27578 => x"00000000",
    27579 => x"00000000", 27580 => x"00000000", 27581 => x"00000000",
    27582 => x"00000000", 27583 => x"00000000", 27584 => x"00000000",
    27585 => x"00000000", 27586 => x"00000000", 27587 => x"00000000",
    27588 => x"00000000", 27589 => x"00000000", 27590 => x"00000000",
    27591 => x"00000000", 27592 => x"00000000", 27593 => x"00000000",
    27594 => x"00000000", 27595 => x"00000000", 27596 => x"00000000",
    27597 => x"00000000", 27598 => x"00000000", 27599 => x"00000000",
    27600 => x"00000000", 27601 => x"00000000", 27602 => x"00000000",
    27603 => x"00000000", 27604 => x"00000000", 27605 => x"00000000",
    27606 => x"00000000", 27607 => x"00000000", 27608 => x"00000000",
    27609 => x"00000000", 27610 => x"00000000", 27611 => x"00000000",
    27612 => x"00000000", 27613 => x"00000000", 27614 => x"00000000",
    27615 => x"00000000", 27616 => x"00000000", 27617 => x"00000000",
    27618 => x"00000000", 27619 => x"00000000", 27620 => x"00000000",
    27621 => x"00000000", 27622 => x"00000000", 27623 => x"00000000",
    27624 => x"00000000", 27625 => x"00000000", 27626 => x"00000000",
    27627 => x"00000000", 27628 => x"00000000", 27629 => x"00000000",
    27630 => x"00000000", 27631 => x"00000000", 27632 => x"00000000",
    27633 => x"00000000", 27634 => x"00000000", 27635 => x"00000000",
    27636 => x"00000000", 27637 => x"00000000", 27638 => x"00000000",
    27639 => x"00000000", 27640 => x"00000000", 27641 => x"00000000",
    27642 => x"00000000", 27643 => x"00000000", 27644 => x"00000000",
    27645 => x"00000000", 27646 => x"00000000", 27647 => x"00000000",
    27648 => x"00000000", 27649 => x"00000000", 27650 => x"00000000",
    27651 => x"00000000", 27652 => x"00000000", 27653 => x"00000000",
    27654 => x"00000000", 27655 => x"00000000", 27656 => x"00000000",
    27657 => x"00000000", 27658 => x"00000000", 27659 => x"00000000",
    27660 => x"00000000", 27661 => x"00000000", 27662 => x"00000000",
    27663 => x"00000000", 27664 => x"00000000", 27665 => x"00000000",
    27666 => x"00000000", 27667 => x"00000000", 27668 => x"00000000",
    27669 => x"00000000", 27670 => x"00000000", 27671 => x"00000000",
    27672 => x"00000000", 27673 => x"00000000", 27674 => x"00000000",
    27675 => x"00000000", 27676 => x"00000000", 27677 => x"00000000",
    27678 => x"00000000", 27679 => x"00000000", 27680 => x"00000000",
    27681 => x"00000000", 27682 => x"00000000", 27683 => x"00000000",
    27684 => x"00000000", 27685 => x"00000000", 27686 => x"00000000",
    27687 => x"00000000", 27688 => x"00000000", 27689 => x"00000000",
    27690 => x"00000000", 27691 => x"00000000", 27692 => x"00000000",
    27693 => x"00000000", 27694 => x"00000000", 27695 => x"00000000",
    27696 => x"00000000", 27697 => x"00000000", 27698 => x"00000000",
    27699 => x"00000000", 27700 => x"00000000", 27701 => x"00000000",
    27702 => x"00000000", 27703 => x"00000000", 27704 => x"00000000",
    27705 => x"00000000", 27706 => x"00000000", 27707 => x"00000000",
    27708 => x"00000000", 27709 => x"00000000", 27710 => x"00000000",
    27711 => x"00000000", 27712 => x"00000000", 27713 => x"00000000",
    27714 => x"00000000", 27715 => x"00000000", 27716 => x"00000000",
    27717 => x"00000000", 27718 => x"00000000", 27719 => x"00000000",
    27720 => x"00000000", 27721 => x"00000000", 27722 => x"00000000",
    27723 => x"00000000", 27724 => x"00000000", 27725 => x"00000000",
    27726 => x"00000000", 27727 => x"00000000", 27728 => x"00000000",
    27729 => x"00000000", 27730 => x"00000000", 27731 => x"00000000",
    27732 => x"00000000", 27733 => x"00000000", 27734 => x"00000000",
    27735 => x"00000000", 27736 => x"00000000", 27737 => x"00000000",
    27738 => x"00000000", 27739 => x"00000000", 27740 => x"00000000",
    27741 => x"00000000", 27742 => x"00000000", 27743 => x"00000000",
    27744 => x"00000000", 27745 => x"00000000", 27746 => x"00000000",
    27747 => x"00000000", 27748 => x"00000000", 27749 => x"00000000",
    27750 => x"00000000", 27751 => x"00000000", 27752 => x"00000000",
    27753 => x"00000000", 27754 => x"00000000", 27755 => x"00000000",
    27756 => x"00000000", 27757 => x"00000000", 27758 => x"00000000",
    27759 => x"00000000", 27760 => x"00000000", 27761 => x"00000000",
    27762 => x"00000000", 27763 => x"00000000", 27764 => x"00000000",
    27765 => x"00000000", 27766 => x"00000000", 27767 => x"00000000",
    27768 => x"00000000", 27769 => x"00000000", 27770 => x"00000000",
    27771 => x"00000000", 27772 => x"00000000", 27773 => x"00000000",
    27774 => x"00000000", 27775 => x"00000000", 27776 => x"00000000",
    27777 => x"00000000", 27778 => x"00000000", 27779 => x"00000000",
    27780 => x"00000000", 27781 => x"00000000", 27782 => x"00000000",
    27783 => x"00000000", 27784 => x"00000000", 27785 => x"00000000",
    27786 => x"00000000", 27787 => x"00000000", 27788 => x"00000000",
    27789 => x"00000000", 27790 => x"00000000", 27791 => x"00000000",
    27792 => x"00000000", 27793 => x"00000000", 27794 => x"00000000",
    27795 => x"00000000", 27796 => x"00000000", 27797 => x"00000000",
    27798 => x"00000000", 27799 => x"00000000", 27800 => x"00000000",
    27801 => x"00000000", 27802 => x"00000000", 27803 => x"00000000",
    27804 => x"00000000", 27805 => x"00000000", 27806 => x"00000000",
    27807 => x"00000000", 27808 => x"00000000", 27809 => x"00000000",
    27810 => x"00000000", 27811 => x"00000000", 27812 => x"00000000",
    27813 => x"00000000", 27814 => x"00000000", 27815 => x"00000000",
    27816 => x"00000000", 27817 => x"00000000", 27818 => x"00000000",
    27819 => x"00000000", 27820 => x"00000000", 27821 => x"00000000",
    27822 => x"00000000", 27823 => x"00000000", 27824 => x"00000000",
    27825 => x"00000000", 27826 => x"00000000", 27827 => x"00000000",
    27828 => x"00000000", 27829 => x"00000000", 27830 => x"00000000",
    27831 => x"00000000", 27832 => x"00000000", 27833 => x"00000000",
    27834 => x"00000000", 27835 => x"00000000", 27836 => x"00000000",
    27837 => x"00000000", 27838 => x"00000000", 27839 => x"00000000",
    27840 => x"00000000", 27841 => x"00000000", 27842 => x"00000000",
    27843 => x"00000000", 27844 => x"00000000", 27845 => x"00000000",
    27846 => x"00000000", 27847 => x"00000000", 27848 => x"00000000",
    27849 => x"00000000", 27850 => x"00000000", 27851 => x"00000000",
    27852 => x"00000000", 27853 => x"00000000", 27854 => x"00000000",
    27855 => x"00000000", 27856 => x"00000000", 27857 => x"00000000",
    27858 => x"00000000", 27859 => x"00000000", 27860 => x"00000000",
    27861 => x"00000000", 27862 => x"00000000", 27863 => x"00000000",
    27864 => x"00000000", 27865 => x"00000000", 27866 => x"00000000",
    27867 => x"00000000", 27868 => x"00000000", 27869 => x"00000000",
    27870 => x"00000000", 27871 => x"00000000", 27872 => x"00000000",
    27873 => x"00000000", 27874 => x"00000000", 27875 => x"00000000",
    27876 => x"00000000", 27877 => x"00000000", 27878 => x"00000000",
    27879 => x"00000000", 27880 => x"00000000", 27881 => x"00000000",
    27882 => x"00000000", 27883 => x"00000000", 27884 => x"00000000",
    27885 => x"00000000", 27886 => x"00000000", 27887 => x"00000000",
    27888 => x"00000000", 27889 => x"00000000", 27890 => x"00000000",
    27891 => x"00000000", 27892 => x"00000000", 27893 => x"00000000",
    27894 => x"00000000", 27895 => x"00000000", 27896 => x"00000000",
    27897 => x"00000000", 27898 => x"00000000", 27899 => x"00000000",
    27900 => x"00000000", 27901 => x"00000000", 27902 => x"00000000",
    27903 => x"00000000", 27904 => x"00000000", 27905 => x"00000000",
    27906 => x"00000000", 27907 => x"00000000", 27908 => x"00000000",
    27909 => x"00000000", 27910 => x"00000000", 27911 => x"00000000",
    27912 => x"00000000", 27913 => x"00000000", 27914 => x"00000000",
    27915 => x"00000000", 27916 => x"00000000", 27917 => x"00000000",
    27918 => x"00000000", 27919 => x"00000000", 27920 => x"00000000",
    27921 => x"00000000", 27922 => x"00000000", 27923 => x"00000000",
    27924 => x"00000000", 27925 => x"00000000", 27926 => x"00000000",
    27927 => x"00000000", 27928 => x"00000000", 27929 => x"00000000",
    27930 => x"00000000", 27931 => x"00000000", 27932 => x"00000000",
    27933 => x"00000000", 27934 => x"00000000", 27935 => x"00000000",
    27936 => x"00000000", 27937 => x"00000000", 27938 => x"00000000",
    27939 => x"00000000", 27940 => x"00000000", 27941 => x"00000000",
    27942 => x"00000000", 27943 => x"00000000", 27944 => x"00000000",
    27945 => x"00000000", 27946 => x"00000000", 27947 => x"00000000",
    27948 => x"00000000", 27949 => x"00000000", 27950 => x"00000000",
    27951 => x"00000000", 27952 => x"00000000", 27953 => x"00000000",
    27954 => x"00000000", 27955 => x"00000000", 27956 => x"00000000",
    27957 => x"00000000", 27958 => x"00000000", 27959 => x"00000000",
    27960 => x"00000000", 27961 => x"00000000", 27962 => x"00000000",
    27963 => x"00000000", 27964 => x"00000000", 27965 => x"00000000",
    27966 => x"00000000", 27967 => x"00000000", 27968 => x"00000000",
    27969 => x"00000000", 27970 => x"00000000", 27971 => x"00000000",
    27972 => x"00000000", 27973 => x"00000000", 27974 => x"00000000",
    27975 => x"00000000", 27976 => x"00000000", 27977 => x"00000000",
    27978 => x"00000000", 27979 => x"00000000", 27980 => x"00000000",
    27981 => x"00000000", 27982 => x"00000000", 27983 => x"00000000",
    27984 => x"00000000", 27985 => x"00000000", 27986 => x"00000000",
    27987 => x"00000000", 27988 => x"00000000", 27989 => x"00000000",
    27990 => x"00000000", 27991 => x"00000000", 27992 => x"00000000",
    27993 => x"00000000", 27994 => x"00000000", 27995 => x"00000000",
    27996 => x"00000000", 27997 => x"00000000", 27998 => x"00000000",
    27999 => x"00000000", 28000 => x"00000000", 28001 => x"00000000",
    28002 => x"00000000", 28003 => x"00000000", 28004 => x"00000000",
    28005 => x"00000000", 28006 => x"00000000", 28007 => x"00000000",
    28008 => x"00000000", 28009 => x"00000000", 28010 => x"00000000",
    28011 => x"00000000", 28012 => x"00000000", 28013 => x"00000000",
    28014 => x"00000000", 28015 => x"00000000", 28016 => x"00000000",
    28017 => x"00000000", 28018 => x"00000000", 28019 => x"00000000",
    28020 => x"00000000", 28021 => x"00000000", 28022 => x"00000000",
    28023 => x"00000000", 28024 => x"00000000", 28025 => x"00000000",
    28026 => x"00000000", 28027 => x"00000000", 28028 => x"00000000",
    28029 => x"00000000", 28030 => x"00000000", 28031 => x"00000000",
    28032 => x"00000000", 28033 => x"00000000", 28034 => x"00000000",
    28035 => x"00000000", 28036 => x"00000000", 28037 => x"00000000",
    28038 => x"00000000", 28039 => x"00000000", 28040 => x"00000000",
    28041 => x"00000000", 28042 => x"00000000", 28043 => x"00000000",
    28044 => x"00000000", 28045 => x"00000000", 28046 => x"00000000",
    28047 => x"00000000", 28048 => x"00000000", 28049 => x"00000000",
    28050 => x"00000000", 28051 => x"00000000", 28052 => x"00000000",
    28053 => x"00000000", 28054 => x"00000000", 28055 => x"00000000",
    28056 => x"00000000", 28057 => x"00000000", 28058 => x"00000000",
    28059 => x"00000000", 28060 => x"00000000", 28061 => x"00000000",
    28062 => x"00000000", 28063 => x"00000000", 28064 => x"00000000",
    28065 => x"00000000", 28066 => x"00000000", 28067 => x"00000000",
    28068 => x"00000000", 28069 => x"00000000", 28070 => x"00000000",
    28071 => x"00000000", 28072 => x"00000000", 28073 => x"00000000",
    28074 => x"00000000", 28075 => x"00000000", 28076 => x"00000000",
    28077 => x"00000000", 28078 => x"00000000", 28079 => x"00000000",
    28080 => x"00000000", 28081 => x"00000000", 28082 => x"00000000",
    28083 => x"00000000", 28084 => x"00000000", 28085 => x"00000000",
    28086 => x"00000000", 28087 => x"00000000", 28088 => x"00000000",
    28089 => x"00000000", 28090 => x"00000000", 28091 => x"00000000",
    28092 => x"00000000", 28093 => x"00000000", 28094 => x"00000000",
    28095 => x"00000000", 28096 => x"00000000", 28097 => x"00000000",
    28098 => x"00000000", 28099 => x"00000000", 28100 => x"00000000",
    28101 => x"00000000", 28102 => x"00000000", 28103 => x"00000000",
    28104 => x"00000000", 28105 => x"00000000", 28106 => x"00000000",
    28107 => x"00000000", 28108 => x"00000000", 28109 => x"00000000",
    28110 => x"00000000", 28111 => x"00000000", 28112 => x"00000000",
    28113 => x"00000000", 28114 => x"00000000", 28115 => x"00000000",
    28116 => x"00000000", 28117 => x"00000000", 28118 => x"00000000",
    28119 => x"00000000", 28120 => x"00000000", 28121 => x"00000000",
    28122 => x"00000000", 28123 => x"00000000", 28124 => x"00000000",
    28125 => x"00000000", 28126 => x"00000000", 28127 => x"00000000",
    28128 => x"00000000", 28129 => x"00000000", 28130 => x"00000000",
    28131 => x"00000000", 28132 => x"00000000", 28133 => x"00000000",
    28134 => x"00000000", 28135 => x"00000000", 28136 => x"00000000",
    28137 => x"00000000", 28138 => x"00000000", 28139 => x"00000000",
    28140 => x"00000000", 28141 => x"00000000", 28142 => x"00000000",
    28143 => x"00000000", 28144 => x"00000000", 28145 => x"00000000",
    28146 => x"00000000", 28147 => x"00000000", 28148 => x"00000000",
    28149 => x"00000000", 28150 => x"00000000", 28151 => x"00000000",
    28152 => x"00000000", 28153 => x"00000000", 28154 => x"00000000",
    28155 => x"00000000", 28156 => x"00000000", 28157 => x"00000000",
    28158 => x"00000000", 28159 => x"00000000", 28160 => x"00000000",
    28161 => x"00000000", 28162 => x"00000000", 28163 => x"00000000",
    28164 => x"00000000", 28165 => x"00000000", 28166 => x"00000000",
    28167 => x"00000000", 28168 => x"00000000", 28169 => x"00000000",
    28170 => x"00000000", 28171 => x"00000000", 28172 => x"00000000",
    28173 => x"00000000", 28174 => x"00000000", 28175 => x"00000000",
    28176 => x"00000000", 28177 => x"00000000", 28178 => x"00000000",
    28179 => x"00000000", 28180 => x"00000000", 28181 => x"00000000",
    28182 => x"00000000", 28183 => x"00000000", 28184 => x"00000000",
    28185 => x"00000000", 28186 => x"00000000", 28187 => x"00000000",
    28188 => x"00000000", 28189 => x"00000000", 28190 => x"00000000",
    28191 => x"00000000", 28192 => x"00000000", 28193 => x"00000000",
    28194 => x"00000000", 28195 => x"00000000", 28196 => x"00000000",
    28197 => x"00000000", 28198 => x"00000000", 28199 => x"00000000",
    28200 => x"00000000", 28201 => x"00000000", 28202 => x"00000000",
    28203 => x"00000000", 28204 => x"00000000", 28205 => x"00000000",
    28206 => x"00000000", 28207 => x"00000000", 28208 => x"00000000",
    28209 => x"00000000", 28210 => x"00000000", 28211 => x"00000000",
    28212 => x"00000000", 28213 => x"00000000", 28214 => x"00000000",
    28215 => x"00000000", 28216 => x"00000000", 28217 => x"00000000",
    28218 => x"00000000", 28219 => x"00000000", 28220 => x"00000000",
    28221 => x"00000000", 28222 => x"00000000", 28223 => x"00000000",
    28224 => x"00000000", 28225 => x"00000000", 28226 => x"00000000",
    28227 => x"00000000", 28228 => x"00000000", 28229 => x"00000000",
    28230 => x"00000000", 28231 => x"00000000", 28232 => x"00000000",
    28233 => x"00000000", 28234 => x"00000000", 28235 => x"00000000",
    28236 => x"00000000", 28237 => x"00000000", 28238 => x"00000000",
    28239 => x"00000000", 28240 => x"00000000", 28241 => x"00000000",
    28242 => x"00000000", 28243 => x"00000000", 28244 => x"00000000",
    28245 => x"00000000", 28246 => x"00000000", 28247 => x"00000000",
    28248 => x"00000000", 28249 => x"00000000", 28250 => x"00000000",
    28251 => x"00000000", 28252 => x"00000000", 28253 => x"00000000",
    28254 => x"00000000", 28255 => x"00000000", 28256 => x"00000000",
    28257 => x"00000000", 28258 => x"00000000", 28259 => x"00000000",
    28260 => x"00000000", 28261 => x"00000000", 28262 => x"00000000",
    28263 => x"00000000", 28264 => x"00000000", 28265 => x"00000000",
    28266 => x"00000000", 28267 => x"00000000", 28268 => x"00000000",
    28269 => x"00000000", 28270 => x"00000000", 28271 => x"00000000",
    28272 => x"00000000", 28273 => x"00000000", 28274 => x"00000000",
    28275 => x"00000000", 28276 => x"00000000", 28277 => x"00000000",
    28278 => x"00000000", 28279 => x"00000000", 28280 => x"00000000",
    28281 => x"00000000", 28282 => x"00000000", 28283 => x"00000000",
    28284 => x"00000000", 28285 => x"00000000", 28286 => x"00000000",
    28287 => x"00000000", 28288 => x"00000000", 28289 => x"00000000",
    28290 => x"00000000", 28291 => x"00000000", 28292 => x"00000000",
    28293 => x"00000000", 28294 => x"00000000", 28295 => x"00000000",
    28296 => x"00000000", 28297 => x"00000000", 28298 => x"00000000",
    28299 => x"00000000", 28300 => x"00000000", 28301 => x"00000000",
    28302 => x"00000000", 28303 => x"00000000", 28304 => x"00000000",
    28305 => x"00000000", 28306 => x"00000000", 28307 => x"00000000",
    28308 => x"00000000", 28309 => x"00000000", 28310 => x"00000000",
    28311 => x"00000000", 28312 => x"00000000", 28313 => x"00000000",
    28314 => x"00000000", 28315 => x"00000000", 28316 => x"00000000",
    28317 => x"00000000", 28318 => x"00000000", 28319 => x"00000000",
    28320 => x"00000000", 28321 => x"00000000", 28322 => x"00000000",
    28323 => x"00000000", 28324 => x"00000000", 28325 => x"00000000",
    28326 => x"00000000", 28327 => x"00000000", 28328 => x"00000000",
    28329 => x"00000000", 28330 => x"00000000", 28331 => x"00000000",
    28332 => x"00000000", 28333 => x"00000000", 28334 => x"00000000",
    28335 => x"00000000", 28336 => x"00000000", 28337 => x"00000000",
    28338 => x"00000000", 28339 => x"00000000", 28340 => x"00000000",
    28341 => x"00000000", 28342 => x"00000000", 28343 => x"00000000",
    28344 => x"00000000", 28345 => x"00000000", 28346 => x"00000000",
    28347 => x"00000000", 28348 => x"00000000", 28349 => x"00000000",
    28350 => x"00000000", 28351 => x"00000000", 28352 => x"00000000",
    28353 => x"00000000", 28354 => x"00000000", 28355 => x"00000000",
    28356 => x"00000000", 28357 => x"00000000", 28358 => x"00000000",
    28359 => x"00000000", 28360 => x"00000000", 28361 => x"00000000",
    28362 => x"00000000", 28363 => x"00000000", 28364 => x"00000000",
    28365 => x"00000000", 28366 => x"00000000", 28367 => x"00000000",
    28368 => x"00000000", 28369 => x"00000000", 28370 => x"00000000",
    28371 => x"00000000", 28372 => x"00000000", 28373 => x"00000000",
    28374 => x"00000000", 28375 => x"00000000", 28376 => x"00000000",
    28377 => x"00000000", 28378 => x"00000000", 28379 => x"00000000",
    28380 => x"00000000", 28381 => x"00000000", 28382 => x"00000000",
    28383 => x"00000000", 28384 => x"00000000", 28385 => x"00000000",
    28386 => x"00000000", 28387 => x"00000000", 28388 => x"00000000",
    28389 => x"00000000", 28390 => x"00000000", 28391 => x"00000000",
    28392 => x"00000000", 28393 => x"00000000", 28394 => x"00000000",
    28395 => x"00000000", 28396 => x"00000000", 28397 => x"00000000",
    28398 => x"00000000", 28399 => x"00000000", 28400 => x"00000000",
    28401 => x"00000000", 28402 => x"00000000", 28403 => x"00000000",
    28404 => x"00000000", 28405 => x"00000000", 28406 => x"00000000",
    28407 => x"00000000", 28408 => x"00000000", 28409 => x"00000000",
    28410 => x"00000000", 28411 => x"00000000", 28412 => x"00000000",
    28413 => x"00000000", 28414 => x"00000000", 28415 => x"00000000",
    28416 => x"00000000", 28417 => x"00000000", 28418 => x"00000000",
    28419 => x"00000000", 28420 => x"00000000", 28421 => x"00000000",
    28422 => x"00000000", 28423 => x"00000000", 28424 => x"00000000",
    28425 => x"00000000", 28426 => x"00000000", 28427 => x"00000000",
    28428 => x"00000000", 28429 => x"00000000", 28430 => x"00000000",
    28431 => x"00000000", 28432 => x"00000000", 28433 => x"00000000",
    28434 => x"00000000", 28435 => x"00000000", 28436 => x"00000000",
    28437 => x"00000000", 28438 => x"00000000", 28439 => x"00000000",
    28440 => x"00000000", 28441 => x"00000000", 28442 => x"00000000",
    28443 => x"00000000", 28444 => x"00000000", 28445 => x"00000000",
    28446 => x"00000000", 28447 => x"00000000", 28448 => x"00000000",
    28449 => x"00000000", 28450 => x"00000000", 28451 => x"00000000",
    28452 => x"00000000", 28453 => x"00000000", 28454 => x"00000000",
    28455 => x"00000000", 28456 => x"00000000", 28457 => x"00000000",
    28458 => x"00000000", 28459 => x"00000000", 28460 => x"00000000",
    28461 => x"00000000", 28462 => x"00000000", 28463 => x"00000000",
    28464 => x"00000000", 28465 => x"00000000", 28466 => x"00000000",
    28467 => x"00000000", 28468 => x"00000000", 28469 => x"00000000",
    28470 => x"00000000", 28471 => x"00000000", 28472 => x"00000000",
    28473 => x"00000000", 28474 => x"00000000", 28475 => x"00000000",
    28476 => x"00000000", 28477 => x"00000000", 28478 => x"00000000",
    28479 => x"00000000", 28480 => x"00000000", 28481 => x"00000000",
    28482 => x"00000000", 28483 => x"00000000", 28484 => x"00000000",
    28485 => x"00000000", 28486 => x"00000000", 28487 => x"00000000",
    28488 => x"00000000", 28489 => x"00000000", 28490 => x"00000000",
    28491 => x"00000000", 28492 => x"00000000", 28493 => x"00000000",
    28494 => x"00000000", 28495 => x"00000000", 28496 => x"00000000",
    28497 => x"00000000", 28498 => x"00000000", 28499 => x"00000000",
    28500 => x"00000000", 28501 => x"00000000", 28502 => x"00000000",
    28503 => x"00000000", 28504 => x"00000000", 28505 => x"00000000",
    28506 => x"00000000", 28507 => x"00000000", 28508 => x"00000000",
    28509 => x"00000000", 28510 => x"00000000", 28511 => x"00000000",
    28512 => x"00000000", 28513 => x"00000000", 28514 => x"00000000",
    28515 => x"00000000", 28516 => x"00000000", 28517 => x"00000000",
    28518 => x"00000000", 28519 => x"00000000", 28520 => x"00000000",
    28521 => x"00000000", 28522 => x"00000000", 28523 => x"00000000",
    28524 => x"00000000", 28525 => x"00000000", 28526 => x"00000000",
    28527 => x"00000000", 28528 => x"00000000", 28529 => x"00000000",
    28530 => x"00000000", 28531 => x"00000000", 28532 => x"00000000",
    28533 => x"00000000", 28534 => x"00000000", 28535 => x"00000000",
    28536 => x"00000000", 28537 => x"00000000", 28538 => x"00000000",
    28539 => x"00000000", 28540 => x"00000000", 28541 => x"00000000",
    28542 => x"00000000", 28543 => x"00000000", 28544 => x"00000000",
    28545 => x"00000000", 28546 => x"00000000", 28547 => x"00000000",
    28548 => x"00000000", 28549 => x"00000000", 28550 => x"00000000",
    28551 => x"00000000", 28552 => x"00000000", 28553 => x"00000000",
    28554 => x"00000000", 28555 => x"00000000", 28556 => x"00000000",
    28557 => x"00000000", 28558 => x"00000000", 28559 => x"00000000",
    28560 => x"00000000", 28561 => x"00000000", 28562 => x"00000000",
    28563 => x"00000000", 28564 => x"00000000", 28565 => x"00000000",
    28566 => x"00000000", 28567 => x"00000000", 28568 => x"00000000",
    28569 => x"00000000", 28570 => x"00000000", 28571 => x"00000000",
    28572 => x"00000000", 28573 => x"00000000", 28574 => x"00000000",
    28575 => x"00000000", 28576 => x"00000000", 28577 => x"00000000",
    28578 => x"00000000", 28579 => x"00000000", 28580 => x"00000000",
    28581 => x"00000000", 28582 => x"00000000", 28583 => x"00000000",
    28584 => x"00000000", 28585 => x"00000000", 28586 => x"00000000",
    28587 => x"00000000", 28588 => x"00000000", 28589 => x"00000000",
    28590 => x"00000000", 28591 => x"00000000", 28592 => x"00000000",
    28593 => x"00000000", 28594 => x"00000000", 28595 => x"00000000",
    28596 => x"00000000", 28597 => x"00000000", 28598 => x"00000000",
    28599 => x"00000000", 28600 => x"00000000", 28601 => x"00000000",
    28602 => x"00000000", 28603 => x"00000000", 28604 => x"00000000",
    28605 => x"00000000", 28606 => x"00000000", 28607 => x"00000000",
    28608 => x"00000000", 28609 => x"00000000", 28610 => x"00000000",
    28611 => x"00000000", 28612 => x"00000000", 28613 => x"00000000",
    28614 => x"00000000", 28615 => x"00000000", 28616 => x"00000000",
    28617 => x"00000000", 28618 => x"00000000", 28619 => x"00000000",
    28620 => x"00000000", 28621 => x"00000000", 28622 => x"00000000",
    28623 => x"00000000", 28624 => x"00000000", 28625 => x"00000000",
    28626 => x"00000000", 28627 => x"00000000", 28628 => x"00000000",
    28629 => x"00000000", 28630 => x"00000000", 28631 => x"00000000",
    28632 => x"00000000", 28633 => x"00000000", 28634 => x"00000000",
    28635 => x"00000000", 28636 => x"00000000", 28637 => x"00000000",
    28638 => x"00000000", 28639 => x"00000000", 28640 => x"00000000",
    28641 => x"00000000", 28642 => x"00000000", 28643 => x"00000000",
    28644 => x"00000000", 28645 => x"00000000", 28646 => x"00000000",
    28647 => x"00000000", 28648 => x"00000000", 28649 => x"00000000",
    28650 => x"00000000", 28651 => x"00000000", 28652 => x"00000000",
    28653 => x"00000000", 28654 => x"00000000", 28655 => x"00000000",
    28656 => x"00000000", 28657 => x"00000000", 28658 => x"00000000",
    28659 => x"00000000", 28660 => x"00000000", 28661 => x"00000000",
    28662 => x"00000000", 28663 => x"00000000", 28664 => x"00000000",
    28665 => x"00000000", 28666 => x"00000000", 28667 => x"00000000",
    28668 => x"00000000", 28669 => x"00000000", 28670 => x"00000000",
    28671 => x"00000000", 28672 => x"00000000", 28673 => x"00000000",
    28674 => x"00000000", 28675 => x"00000000", 28676 => x"00000000",
    28677 => x"00000000", 28678 => x"00000000", 28679 => x"00000000",
    28680 => x"00000000", 28681 => x"00000000", 28682 => x"00000000",
    28683 => x"00000000", 28684 => x"00000000", 28685 => x"00000000",
    28686 => x"00000000", 28687 => x"00000000", 28688 => x"00000000",
    28689 => x"00000000", 28690 => x"00000000", 28691 => x"00000000",
    28692 => x"00000000", 28693 => x"00000000", 28694 => x"00000000",
    28695 => x"00000000", 28696 => x"00000000", 28697 => x"00000000",
    28698 => x"00000000", 28699 => x"00000000", 28700 => x"00000000",
    28701 => x"00000000", 28702 => x"00000000", 28703 => x"00000000",
    28704 => x"00000000", 28705 => x"00000000", 28706 => x"00000000",
    28707 => x"00000000", 28708 => x"00000000", 28709 => x"00000000",
    28710 => x"00000000", 28711 => x"00000000", 28712 => x"00000000",
    28713 => x"00000000", 28714 => x"00000000", 28715 => x"00000000",
    28716 => x"00000000", 28717 => x"00000000", 28718 => x"00000000",
    28719 => x"00000000", 28720 => x"00000000", 28721 => x"00000000",
    28722 => x"00000000", 28723 => x"00000000", 28724 => x"00000000",
    28725 => x"00000000", 28726 => x"00000000", 28727 => x"00000000",
    28728 => x"00000000", 28729 => x"00000000", 28730 => x"00000000",
    28731 => x"00000000", 28732 => x"00000000", 28733 => x"00000000",
    28734 => x"00000000", 28735 => x"00000000", 28736 => x"00000000",
    28737 => x"00000000", 28738 => x"00000000", 28739 => x"00000000",
    28740 => x"00000000", 28741 => x"00000000", 28742 => x"00000000",
    28743 => x"00000000", 28744 => x"00000000", 28745 => x"00000000",
    28746 => x"00000000", 28747 => x"00000000", 28748 => x"00000000",
    28749 => x"00000000", 28750 => x"00000000", 28751 => x"00000000",
    28752 => x"00000000", 28753 => x"00000000", 28754 => x"00000000",
    28755 => x"00000000", 28756 => x"00000000", 28757 => x"00000000",
    28758 => x"00000000", 28759 => x"00000000", 28760 => x"00000000",
    28761 => x"00000000", 28762 => x"00000000", 28763 => x"00000000",
    28764 => x"00000000", 28765 => x"00000000", 28766 => x"00000000",
    28767 => x"00000000", 28768 => x"00000000", 28769 => x"00000000",
    28770 => x"00000000", 28771 => x"00000000", 28772 => x"00000000",
    28773 => x"00000000", 28774 => x"00000000", 28775 => x"00000000",
    28776 => x"00000000", 28777 => x"00000000", 28778 => x"00000000",
    28779 => x"00000000", 28780 => x"00000000", 28781 => x"00000000",
    28782 => x"00000000", 28783 => x"00000000", 28784 => x"00000000",
    28785 => x"00000000", 28786 => x"00000000", 28787 => x"00000000",
    28788 => x"00000000", 28789 => x"00000000", 28790 => x"00000000",
    28791 => x"00000000", 28792 => x"00000000", 28793 => x"00000000",
    28794 => x"00000000", 28795 => x"00000000", 28796 => x"00000000",
    28797 => x"00000000", 28798 => x"00000000", 28799 => x"00000000",
    28800 => x"00000000", 28801 => x"00000000", 28802 => x"00000000",
    28803 => x"00000000", 28804 => x"00000000", 28805 => x"00000000",
    28806 => x"00000000", 28807 => x"00000000", 28808 => x"00000000",
    28809 => x"00000000", 28810 => x"00000000", 28811 => x"00000000",
    28812 => x"00000000", 28813 => x"00000000", 28814 => x"00000000",
    28815 => x"00000000", 28816 => x"00000000", 28817 => x"00000000",
    28818 => x"00000000", 28819 => x"00000000", 28820 => x"00000000",
    28821 => x"00000000", 28822 => x"00000000", 28823 => x"00000000",
    28824 => x"00000000", 28825 => x"00000000", 28826 => x"00000000",
    28827 => x"00000000", 28828 => x"00000000", 28829 => x"00000000",
    28830 => x"00000000", 28831 => x"00000000", 28832 => x"00000000",
    28833 => x"00000000", 28834 => x"00000000", 28835 => x"00000000",
    28836 => x"00000000", 28837 => x"00000000", 28838 => x"00000000",
    28839 => x"00000000", 28840 => x"00000000", 28841 => x"00000000",
    28842 => x"00000000", 28843 => x"00000000", 28844 => x"00000000",
    28845 => x"00000000", 28846 => x"00000000", 28847 => x"00000000",
    28848 => x"00000000", 28849 => x"00000000", 28850 => x"00000000",
    28851 => x"00000000", 28852 => x"00000000", 28853 => x"00000000",
    28854 => x"00000000", 28855 => x"00000000", 28856 => x"00000000",
    28857 => x"00000000", 28858 => x"00000000", 28859 => x"00000000",
    28860 => x"00000000", 28861 => x"00000000", 28862 => x"00000000",
    28863 => x"00000000", 28864 => x"00000000", 28865 => x"00000000",
    28866 => x"00000000", 28867 => x"00000000", 28868 => x"00000000",
    28869 => x"00000000", 28870 => x"00000000", 28871 => x"00000000",
    28872 => x"00000000", 28873 => x"00000000", 28874 => x"00000000",
    28875 => x"00000000", 28876 => x"00000000", 28877 => x"00000000",
    28878 => x"00000000", 28879 => x"00000000", 28880 => x"00000000",
    28881 => x"00000000", 28882 => x"00000000", 28883 => x"00000000",
    28884 => x"00000000", 28885 => x"00000000", 28886 => x"00000000",
    28887 => x"00000000", 28888 => x"00000000", 28889 => x"00000000",
    28890 => x"00000000", 28891 => x"00000000", 28892 => x"00000000",
    28893 => x"00000000", 28894 => x"00000000", 28895 => x"00000000",
    28896 => x"00000000", 28897 => x"00000000", 28898 => x"00000000",
    28899 => x"00000000", 28900 => x"00000000", 28901 => x"00000000",
    28902 => x"00000000", 28903 => x"00000000", 28904 => x"00000000",
    28905 => x"00000000", 28906 => x"00000000", 28907 => x"00000000",
    28908 => x"00000000", 28909 => x"00000000", 28910 => x"00000000",
    28911 => x"00000000", 28912 => x"00000000", 28913 => x"00000000",
    28914 => x"00000000", 28915 => x"00000000", 28916 => x"00000000",
    28917 => x"00000000", 28918 => x"00000000", 28919 => x"00000000",
    28920 => x"00000000", 28921 => x"00000000", 28922 => x"00000000",
    28923 => x"00000000", 28924 => x"00000000", 28925 => x"00000000",
    28926 => x"00000000", 28927 => x"00000000", 28928 => x"00000000",
    28929 => x"00000000", 28930 => x"00000000", 28931 => x"00000000",
    28932 => x"00000000", 28933 => x"00000000", 28934 => x"00000000",
    28935 => x"00000000", 28936 => x"00000000", 28937 => x"00000000",
    28938 => x"00000000", 28939 => x"00000000", 28940 => x"00000000",
    28941 => x"00000000", 28942 => x"00000000", 28943 => x"00000000",
    28944 => x"00000000", 28945 => x"00000000", 28946 => x"00000000",
    28947 => x"00000000", 28948 => x"00000000", 28949 => x"00000000",
    28950 => x"00000000", 28951 => x"00000000", 28952 => x"00000000",
    28953 => x"00000000", 28954 => x"00000000", 28955 => x"00000000",
    28956 => x"00000000", 28957 => x"00000000", 28958 => x"00000000",
    28959 => x"00000000", 28960 => x"00000000", 28961 => x"00000000",
    28962 => x"00000000", 28963 => x"00000000", 28964 => x"00000000",
    28965 => x"00000000", 28966 => x"00000000", 28967 => x"00000000",
    28968 => x"00000000", 28969 => x"00000000", 28970 => x"00000000",
    28971 => x"00000000", 28972 => x"00000000", 28973 => x"00000000",
    28974 => x"00000000", 28975 => x"00000000", 28976 => x"00000000",
    28977 => x"00000000", 28978 => x"00000000", 28979 => x"00000000",
    28980 => x"00000000", 28981 => x"00000000", 28982 => x"00000000",
    28983 => x"00000000", 28984 => x"00000000", 28985 => x"00000000",
    28986 => x"00000000", 28987 => x"00000000", 28988 => x"00000000",
    28989 => x"00000000", 28990 => x"00000000", 28991 => x"00000000",
    28992 => x"00000000", 28993 => x"00000000", 28994 => x"00000000",
    28995 => x"00000000", 28996 => x"00000000", 28997 => x"00000000",
    28998 => x"00000000", 28999 => x"00000000", 29000 => x"00000000",
    29001 => x"00000000", 29002 => x"00000000", 29003 => x"00000000",
    29004 => x"00000000", 29005 => x"00000000", 29006 => x"00000000",
    29007 => x"00000000", 29008 => x"00000000", 29009 => x"00000000",
    29010 => x"00000000", 29011 => x"00000000", 29012 => x"00000000",
    29013 => x"00000000", 29014 => x"00000000", 29015 => x"00000000",
    29016 => x"00000000", 29017 => x"00000000", 29018 => x"00000000",
    29019 => x"00000000", 29020 => x"00000000", 29021 => x"00000000",
    29022 => x"00000000", 29023 => x"00000000", 29024 => x"00000000",
    29025 => x"00000000", 29026 => x"00000000", 29027 => x"00000000",
    29028 => x"00000000", 29029 => x"00000000", 29030 => x"00000000",
    29031 => x"00000000", 29032 => x"00000000", 29033 => x"00000000",
    29034 => x"00000000", 29035 => x"00000000", 29036 => x"00000000",
    29037 => x"00000000", 29038 => x"00000000", 29039 => x"00000000",
    29040 => x"00000000", 29041 => x"00000000", 29042 => x"00000000",
    29043 => x"00000000", 29044 => x"00000000", 29045 => x"00000000",
    29046 => x"00000000", 29047 => x"00000000", 29048 => x"00000000",
    29049 => x"00000000", 29050 => x"00000000", 29051 => x"00000000",
    29052 => x"00000000", 29053 => x"00000000", 29054 => x"00000000",
    29055 => x"00000000", 29056 => x"00000000", 29057 => x"00000000",
    29058 => x"00000000", 29059 => x"00000000", 29060 => x"00000000",
    29061 => x"00000000", 29062 => x"00000000", 29063 => x"00000000",
    29064 => x"00000000", 29065 => x"00000000", 29066 => x"00000000",
    29067 => x"00000000", 29068 => x"00000000", 29069 => x"00000000",
    29070 => x"00000000", 29071 => x"00000000", 29072 => x"00000000",
    29073 => x"00000000", 29074 => x"00000000", 29075 => x"00000000",
    29076 => x"00000000", 29077 => x"00000000", 29078 => x"00000000",
    29079 => x"00000000", 29080 => x"00000000", 29081 => x"00000000",
    29082 => x"00000000", 29083 => x"00000000", 29084 => x"00000000",
    29085 => x"00000000", 29086 => x"00000000", 29087 => x"00000000",
    29088 => x"00000000", 29089 => x"00000000", 29090 => x"00000000",
    29091 => x"00000000", 29092 => x"00000000", 29093 => x"00000000",
    29094 => x"00000000", 29095 => x"00000000", 29096 => x"00000000",
    29097 => x"00000000", 29098 => x"00000000", 29099 => x"00000000",
    29100 => x"00000000", 29101 => x"00000000", 29102 => x"00000000",
    29103 => x"00000000", 29104 => x"00000000", 29105 => x"00000000",
    29106 => x"00000000", 29107 => x"00000000", 29108 => x"00000000",
    29109 => x"00000000", 29110 => x"00000000", 29111 => x"00000000",
    29112 => x"00000000", 29113 => x"00000000", 29114 => x"00000000",
    29115 => x"00000000", 29116 => x"00000000", 29117 => x"00000000",
    29118 => x"00000000", 29119 => x"00000000", 29120 => x"00000000",
    29121 => x"00000000", 29122 => x"00000000", 29123 => x"00000000",
    29124 => x"00000000", 29125 => x"00000000", 29126 => x"00000000",
    29127 => x"00000000", 29128 => x"00000000", 29129 => x"00000000",
    29130 => x"00000000", 29131 => x"00000000", 29132 => x"00000000",
    29133 => x"00000000", 29134 => x"00000000", 29135 => x"00000000",
    29136 => x"00000000", 29137 => x"00000000", 29138 => x"00000000",
    29139 => x"00000000", 29140 => x"00000000", 29141 => x"00000000",
    29142 => x"00000000", 29143 => x"00000000", 29144 => x"00000000",
    29145 => x"00000000", 29146 => x"00000000", 29147 => x"00000000",
    29148 => x"00000000", 29149 => x"00000000", 29150 => x"00000000",
    29151 => x"00000000", 29152 => x"00000000", 29153 => x"00000000",
    29154 => x"00000000", 29155 => x"00000000", 29156 => x"00000000",
    29157 => x"00000000", 29158 => x"00000000", 29159 => x"00000000",
    29160 => x"00000000", 29161 => x"00000000", 29162 => x"00000000",
    29163 => x"00000000", 29164 => x"00000000", 29165 => x"00000000",
    29166 => x"00000000", 29167 => x"00000000", 29168 => x"00000000",
    29169 => x"00000000", 29170 => x"00000000", 29171 => x"00000000",
    29172 => x"00000000", 29173 => x"00000000", 29174 => x"00000000",
    29175 => x"00000000", 29176 => x"00000000", 29177 => x"00000000",
    29178 => x"00000000", 29179 => x"00000000", 29180 => x"00000000",
    29181 => x"00000000", 29182 => x"00000000", 29183 => x"00000000",
    29184 => x"00000000", 29185 => x"00000000", 29186 => x"00000000",
    29187 => x"00000000", 29188 => x"00000000", 29189 => x"00000000",
    29190 => x"00000000", 29191 => x"00000000", 29192 => x"00000000",
    29193 => x"00000000", 29194 => x"00000000", 29195 => x"00000000",
    29196 => x"00000000", 29197 => x"00000000", 29198 => x"00000000",
    29199 => x"00000000", 29200 => x"00000000", 29201 => x"00000000",
    29202 => x"00000000", 29203 => x"00000000", 29204 => x"00000000",
    29205 => x"00000000", 29206 => x"00000000", 29207 => x"00000000",
    29208 => x"00000000", 29209 => x"00000000", 29210 => x"00000000",
    29211 => x"00000000", 29212 => x"00000000", 29213 => x"00000000",
    29214 => x"00000000", 29215 => x"00000000", 29216 => x"00000000",
    29217 => x"00000000", 29218 => x"00000000", 29219 => x"00000000",
    29220 => x"00000000", 29221 => x"00000000", 29222 => x"00000000",
    29223 => x"00000000", 29224 => x"00000000", 29225 => x"00000000",
    29226 => x"00000000", 29227 => x"00000000", 29228 => x"00000000",
    29229 => x"00000000", 29230 => x"00000000", 29231 => x"00000000",
    29232 => x"00000000", 29233 => x"00000000", 29234 => x"00000000",
    29235 => x"00000000", 29236 => x"00000000", 29237 => x"00000000",
    29238 => x"00000000", 29239 => x"00000000", 29240 => x"00000000",
    29241 => x"00000000", 29242 => x"00000000", 29243 => x"00000000",
    29244 => x"00000000", 29245 => x"00000000", 29246 => x"00000000",
    29247 => x"00000000", 29248 => x"00000000", 29249 => x"00000000",
    29250 => x"00000000", 29251 => x"00000000", 29252 => x"00000000",
    29253 => x"00000000", 29254 => x"00000000", 29255 => x"00000000",
    29256 => x"00000000", 29257 => x"00000000", 29258 => x"00000000",
    29259 => x"00000000", 29260 => x"00000000", 29261 => x"00000000",
    29262 => x"00000000", 29263 => x"00000000", 29264 => x"00000000",
    29265 => x"00000000", 29266 => x"00000000", 29267 => x"00000000",
    29268 => x"00000000", 29269 => x"00000000", 29270 => x"00000000",
    29271 => x"00000000", 29272 => x"00000000", 29273 => x"00000000",
    29274 => x"00000000", 29275 => x"00000000", 29276 => x"00000000",
    29277 => x"00000000", 29278 => x"00000000", 29279 => x"00000000",
    29280 => x"00000000", 29281 => x"00000000", 29282 => x"00000000",
    29283 => x"00000000", 29284 => x"00000000", 29285 => x"00000000",
    29286 => x"00000000", 29287 => x"00000000", 29288 => x"00000000",
    29289 => x"00000000", 29290 => x"00000000", 29291 => x"00000000",
    29292 => x"00000000", 29293 => x"00000000", 29294 => x"00000000",
    29295 => x"00000000", 29296 => x"00000000", 29297 => x"00000000",
    29298 => x"00000000", 29299 => x"00000000", 29300 => x"00000000",
    29301 => x"00000000", 29302 => x"00000000", 29303 => x"00000000",
    29304 => x"00000000", 29305 => x"00000000", 29306 => x"00000000",
    29307 => x"00000000", 29308 => x"00000000", 29309 => x"00000000",
    29310 => x"00000000", 29311 => x"00000000", 29312 => x"00000000",
    29313 => x"00000000", 29314 => x"00000000", 29315 => x"00000000",
    29316 => x"00000000", 29317 => x"00000000", 29318 => x"00000000",
    29319 => x"00000000", 29320 => x"00000000", 29321 => x"00000000",
    29322 => x"00000000", 29323 => x"00000000", 29324 => x"00000000",
    29325 => x"00000000", 29326 => x"00000000", 29327 => x"00000000",
    29328 => x"00000000", 29329 => x"00000000", 29330 => x"00000000",
    29331 => x"00000000", 29332 => x"00000000", 29333 => x"00000000",
    29334 => x"00000000", 29335 => x"00000000", 29336 => x"00000000",
    29337 => x"00000000", 29338 => x"00000000", 29339 => x"00000000",
    29340 => x"00000000", 29341 => x"00000000", 29342 => x"00000000",
    29343 => x"00000000", 29344 => x"00000000", 29345 => x"00000000",
    29346 => x"00000000", 29347 => x"00000000", 29348 => x"00000000",
    29349 => x"00000000", 29350 => x"00000000", 29351 => x"00000000",
    29352 => x"00000000", 29353 => x"00000000", 29354 => x"00000000",
    29355 => x"00000000", 29356 => x"00000000", 29357 => x"00000000",
    29358 => x"00000000", 29359 => x"00000000", 29360 => x"00000000",
    29361 => x"00000000", 29362 => x"00000000", 29363 => x"00000000",
    29364 => x"00000000", 29365 => x"00000000", 29366 => x"00000000",
    29367 => x"00000000", 29368 => x"00000000", 29369 => x"00000000",
    29370 => x"00000000", 29371 => x"00000000", 29372 => x"00000000",
    29373 => x"00000000", 29374 => x"00000000", 29375 => x"00000000",
    29376 => x"00000000", 29377 => x"00000000", 29378 => x"00000000",
    29379 => x"00000000", 29380 => x"00000000", 29381 => x"00000000",
    29382 => x"00000000", 29383 => x"00000000", 29384 => x"00000000",
    29385 => x"00000000", 29386 => x"00000000", 29387 => x"00000000",
    29388 => x"00000000", 29389 => x"00000000", 29390 => x"00000000",
    29391 => x"00000000", 29392 => x"00000000", 29393 => x"00000000",
    29394 => x"00000000", 29395 => x"00000000", 29396 => x"00000000",
    29397 => x"00000000", 29398 => x"00000000", 29399 => x"00000000",
    29400 => x"00000000", 29401 => x"00000000", 29402 => x"00000000",
    29403 => x"00000000", 29404 => x"00000000", 29405 => x"00000000",
    29406 => x"00000000", 29407 => x"00000000", 29408 => x"00000000",
    29409 => x"00000000", 29410 => x"00000000", 29411 => x"00000000",
    29412 => x"00000000", 29413 => x"00000000", 29414 => x"00000000",
    29415 => x"00000000", 29416 => x"00000000", 29417 => x"00000000",
    29418 => x"00000000", 29419 => x"00000000", 29420 => x"00000000",
    29421 => x"00000000", 29422 => x"00000000", 29423 => x"00000000",
    29424 => x"00000000", 29425 => x"00000000", 29426 => x"00000000",
    29427 => x"00000000", 29428 => x"00000000", 29429 => x"00000000",
    29430 => x"00000000", 29431 => x"00000000", 29432 => x"00000000",
    29433 => x"00000000", 29434 => x"00000000", 29435 => x"00000000",
    29436 => x"00000000", 29437 => x"00000000", 29438 => x"00000000",
    29439 => x"00000000", 29440 => x"00000000", 29441 => x"00000000",
    29442 => x"00000000", 29443 => x"00000000", 29444 => x"00000000",
    29445 => x"00000000", 29446 => x"00000000", 29447 => x"00000000",
    29448 => x"00000000", 29449 => x"00000000", 29450 => x"00000000",
    29451 => x"00000000", 29452 => x"00000000", 29453 => x"00000000",
    29454 => x"00000000", 29455 => x"00000000", 29456 => x"00000000",
    29457 => x"00000000", 29458 => x"00000000", 29459 => x"00000000",
    29460 => x"00000000", 29461 => x"00000000", 29462 => x"00000000",
    29463 => x"00000000", 29464 => x"00000000", 29465 => x"00000000",
    29466 => x"00000000", 29467 => x"00000000", 29468 => x"00000000",
    29469 => x"00000000", 29470 => x"00000000", 29471 => x"00000000",
    29472 => x"00000000", 29473 => x"00000000", 29474 => x"00000000",
    29475 => x"00000000", 29476 => x"00000000", 29477 => x"00000000",
    29478 => x"00000000", 29479 => x"00000000", 29480 => x"00000000",
    29481 => x"00000000", 29482 => x"00000000", 29483 => x"00000000",
    29484 => x"00000000", 29485 => x"00000000", 29486 => x"00000000",
    29487 => x"00000000", 29488 => x"00000000", 29489 => x"00000000",
    29490 => x"00000000", 29491 => x"00000000", 29492 => x"00000000",
    29493 => x"00000000", 29494 => x"00000000", 29495 => x"00000000",
    29496 => x"00000000", 29497 => x"00000000", 29498 => x"00000000",
    29499 => x"00000000", 29500 => x"00000000", 29501 => x"00000000",
    29502 => x"00000000", 29503 => x"00000000", 29504 => x"00000000",
    29505 => x"00000000", 29506 => x"00000000", 29507 => x"00000000",
    29508 => x"00000000", 29509 => x"00000000", 29510 => x"00000000",
    29511 => x"00000000", 29512 => x"00000000", 29513 => x"00000000",
    29514 => x"00000000", 29515 => x"00000000", 29516 => x"00000000",
    29517 => x"00000000", 29518 => x"00000000", 29519 => x"00000000",
    29520 => x"00000000", 29521 => x"00000000", 29522 => x"00000000",
    29523 => x"00000000", 29524 => x"00000000", 29525 => x"00000000",
    29526 => x"00000000", 29527 => x"00000000", 29528 => x"00000000",
    29529 => x"00000000", 29530 => x"00000000", 29531 => x"00000000",
    29532 => x"00000000", 29533 => x"00000000", 29534 => x"00000000",
    29535 => x"00000000", 29536 => x"00000000", 29537 => x"00000000",
    29538 => x"00000000", 29539 => x"00000000", 29540 => x"00000000",
    29541 => x"00000000", 29542 => x"00000000", 29543 => x"00000000",
    29544 => x"00000000", 29545 => x"00000000", 29546 => x"00000000",
    29547 => x"00000000", 29548 => x"00000000", 29549 => x"00000000",
    29550 => x"00000000", 29551 => x"00000000", 29552 => x"00000000",
    29553 => x"00000000", 29554 => x"00000000", 29555 => x"00000000",
    29556 => x"00000000", 29557 => x"00000000", 29558 => x"00000000",
    29559 => x"00000000", 29560 => x"00000000", 29561 => x"00000000",
    29562 => x"00000000", 29563 => x"00000000", 29564 => x"00000000",
    29565 => x"00000000", 29566 => x"00000000", 29567 => x"00000000",
    29568 => x"00000000", 29569 => x"00000000", 29570 => x"00000000",
    29571 => x"00000000", 29572 => x"00000000", 29573 => x"00000000",
    29574 => x"00000000", 29575 => x"00000000", 29576 => x"00000000",
    29577 => x"00000000", 29578 => x"00000000", 29579 => x"00000000",
    29580 => x"00000000", 29581 => x"00000000", 29582 => x"00000000",
    29583 => x"00000000", 29584 => x"00000000", 29585 => x"00000000",
    29586 => x"00000000", 29587 => x"00000000", 29588 => x"00000000",
    29589 => x"00000000", 29590 => x"00000000", 29591 => x"00000000",
    29592 => x"00000000", 29593 => x"00000000", 29594 => x"00000000",
    29595 => x"00000000", 29596 => x"00000000", 29597 => x"00000000",
    29598 => x"00000000", 29599 => x"00000000", 29600 => x"00000000",
    29601 => x"00000000", 29602 => x"00000000", 29603 => x"00000000",
    29604 => x"00000000", 29605 => x"00000000", 29606 => x"00000000",
    29607 => x"00000000", 29608 => x"00000000", 29609 => x"00000000",
    29610 => x"00000000", 29611 => x"00000000", 29612 => x"00000000",
    29613 => x"00000000", 29614 => x"00000000", 29615 => x"00000000",
    29616 => x"00000000", 29617 => x"00000000", 29618 => x"00000000",
    29619 => x"00000000", 29620 => x"00000000", 29621 => x"00000000",
    29622 => x"00000000", 29623 => x"00000000", 29624 => x"00000000",
    29625 => x"00000000", 29626 => x"00000000", 29627 => x"00000000",
    29628 => x"00000000", 29629 => x"00000000", 29630 => x"00000000",
    29631 => x"00000000", 29632 => x"00000000", 29633 => x"00000000",
    29634 => x"00000000", 29635 => x"00000000", 29636 => x"00000000",
    29637 => x"00000000", 29638 => x"00000000", 29639 => x"00000000",
    29640 => x"00000000", 29641 => x"00000000", 29642 => x"00000000",
    29643 => x"00000000", 29644 => x"00000000", 29645 => x"00000000",
    29646 => x"00000000", 29647 => x"00000000", 29648 => x"00000000",
    29649 => x"00000000", 29650 => x"00000000", 29651 => x"00000000",
    29652 => x"00000000", 29653 => x"00000000", 29654 => x"00000000",
    29655 => x"00000000", 29656 => x"00000000", 29657 => x"00000000",
    29658 => x"00000000", 29659 => x"00000000", 29660 => x"00000000",
    29661 => x"00000000", 29662 => x"00000000", 29663 => x"00000000",
    29664 => x"00000000", 29665 => x"00000000", 29666 => x"00000000",
    29667 => x"00000000", 29668 => x"00000000", 29669 => x"00000000",
    29670 => x"00000000", 29671 => x"00000000", 29672 => x"00000000",
    29673 => x"00000000", 29674 => x"00000000", 29675 => x"00000000",
    29676 => x"00000000", 29677 => x"00000000", 29678 => x"00000000",
    29679 => x"00000000", 29680 => x"00000000", 29681 => x"00000000",
    29682 => x"00000000", 29683 => x"00000000", 29684 => x"00000000",
    29685 => x"00000000", 29686 => x"00000000", 29687 => x"00000000",
    29688 => x"00000000", 29689 => x"00000000", 29690 => x"00000000",
    29691 => x"00000000", 29692 => x"00000000", 29693 => x"00000000",
    29694 => x"00000000", 29695 => x"00000000", 29696 => x"00000000",
    29697 => x"00000000", 29698 => x"00000000", 29699 => x"00000000",
    29700 => x"00000000", 29701 => x"00000000", 29702 => x"00000000",
    29703 => x"00000000", 29704 => x"00000000", 29705 => x"00000000",
    29706 => x"00000000", 29707 => x"00000000", 29708 => x"00000000",
    29709 => x"00000000", 29710 => x"00000000", 29711 => x"00000000",
    29712 => x"00000000", 29713 => x"00000000", 29714 => x"00000000",
    29715 => x"00000000", 29716 => x"00000000", 29717 => x"00000000",
    29718 => x"00000000", 29719 => x"00000000", 29720 => x"00000000",
    29721 => x"00000000", 29722 => x"00000000", 29723 => x"00000000",
    29724 => x"00000000", 29725 => x"00000000", 29726 => x"00000000",
    29727 => x"00000000", 29728 => x"00000000", 29729 => x"00000000",
    29730 => x"00000000", 29731 => x"00000000", 29732 => x"00000000",
    29733 => x"00000000", 29734 => x"00000000", 29735 => x"00000000",
    29736 => x"00000000", 29737 => x"00000000", 29738 => x"00000000",
    29739 => x"00000000", 29740 => x"00000000", 29741 => x"00000000",
    29742 => x"00000000", 29743 => x"00000000", 29744 => x"00000000",
    29745 => x"00000000", 29746 => x"00000000", 29747 => x"00000000",
    29748 => x"00000000", 29749 => x"00000000", 29750 => x"00000000",
    29751 => x"00000000", 29752 => x"00000000", 29753 => x"00000000",
    29754 => x"00000000", 29755 => x"00000000", 29756 => x"00000000",
    29757 => x"00000000", 29758 => x"00000000", 29759 => x"00000000",
    29760 => x"00000000", 29761 => x"00000000", 29762 => x"00000000",
    29763 => x"00000000", 29764 => x"00000000", 29765 => x"00000000",
    29766 => x"00000000", 29767 => x"00000000", 29768 => x"00000000",
    29769 => x"00000000", 29770 => x"00000000", 29771 => x"00000000",
    29772 => x"00000000", 29773 => x"00000000", 29774 => x"00000000",
    29775 => x"00000000", 29776 => x"00000000", 29777 => x"00000000",
    29778 => x"00000000", 29779 => x"00000000", 29780 => x"00000000",
    29781 => x"00000000", 29782 => x"00000000", 29783 => x"00000000",
    29784 => x"00000000", 29785 => x"00000000", 29786 => x"00000000",
    29787 => x"00000000", 29788 => x"00000000", 29789 => x"00000000",
    29790 => x"00000000", 29791 => x"00000000", 29792 => x"00000000",
    29793 => x"00000000", 29794 => x"00000000", 29795 => x"00000000",
    29796 => x"00000000", 29797 => x"00000000", 29798 => x"00000000",
    29799 => x"00000000", 29800 => x"00000000", 29801 => x"00000000",
    29802 => x"00000000", 29803 => x"00000000", 29804 => x"00000000",
    29805 => x"00000000", 29806 => x"00000000", 29807 => x"00000000",
    29808 => x"00000000", 29809 => x"00000000", 29810 => x"00000000",
    29811 => x"00000000", 29812 => x"00000000", 29813 => x"00000000",
    29814 => x"00000000", 29815 => x"00000000", 29816 => x"00000000",
    29817 => x"00000000", 29818 => x"00000000", 29819 => x"00000000",
    29820 => x"00000000", 29821 => x"00000000", 29822 => x"00000000",
    29823 => x"00000000", 29824 => x"00000000", 29825 => x"00000000",
    29826 => x"00000000", 29827 => x"00000000", 29828 => x"00000000",
    29829 => x"00000000", 29830 => x"00000000", 29831 => x"00000000",
    29832 => x"00000000", 29833 => x"00000000", 29834 => x"00000000",
    29835 => x"00000000", 29836 => x"00000000", 29837 => x"00000000",
    29838 => x"00000000", 29839 => x"00000000", 29840 => x"00000000",
    29841 => x"00000000", 29842 => x"00000000", 29843 => x"00000000",
    29844 => x"00000000", 29845 => x"00000000", 29846 => x"00000000",
    29847 => x"00000000", 29848 => x"00000000", 29849 => x"00000000",
    29850 => x"00000000", 29851 => x"00000000", 29852 => x"00000000",
    29853 => x"00000000", 29854 => x"00000000", 29855 => x"00000000",
    29856 => x"00000000", 29857 => x"00000000", 29858 => x"00000000",
    29859 => x"00000000", 29860 => x"00000000", 29861 => x"00000000",
    29862 => x"00000000", 29863 => x"00000000", 29864 => x"00000000",
    29865 => x"00000000", 29866 => x"00000000", 29867 => x"00000000",
    29868 => x"00000000", 29869 => x"00000000", 29870 => x"00000000",
    29871 => x"00000000", 29872 => x"00000000", 29873 => x"00000000",
    29874 => x"00000000", 29875 => x"00000000", 29876 => x"00000000",
    29877 => x"00000000", 29878 => x"00000000", 29879 => x"00000000",
    29880 => x"00000000", 29881 => x"00000000", 29882 => x"00000000",
    29883 => x"00000000", 29884 => x"00000000", 29885 => x"00000000",
    29886 => x"00000000", 29887 => x"00000000", 29888 => x"00000000",
    29889 => x"00000000", 29890 => x"00000000", 29891 => x"00000000",
    29892 => x"00000000", 29893 => x"00000000", 29894 => x"00000000",
    29895 => x"00000000", 29896 => x"00000000", 29897 => x"00000000",
    29898 => x"00000000", 29899 => x"00000000", 29900 => x"00000000",
    29901 => x"00000000", 29902 => x"00000000", 29903 => x"00000000",
    29904 => x"00000000", 29905 => x"00000000", 29906 => x"00000000",
    29907 => x"00000000", 29908 => x"00000000", 29909 => x"00000000",
    29910 => x"00000000", 29911 => x"00000000", 29912 => x"00000000",
    29913 => x"00000000", 29914 => x"00000000", 29915 => x"00000000",
    29916 => x"00000000", 29917 => x"00000000", 29918 => x"00000000",
    29919 => x"00000000", 29920 => x"00000000", 29921 => x"00000000",
    29922 => x"00000000", 29923 => x"00000000", 29924 => x"00000000",
    29925 => x"00000000", 29926 => x"00000000", 29927 => x"00000000",
    29928 => x"00000000", 29929 => x"00000000", 29930 => x"00000000",
    29931 => x"00000000", 29932 => x"00000000", 29933 => x"00000000",
    29934 => x"00000000", 29935 => x"00000000", 29936 => x"00000000",
    29937 => x"00000000", 29938 => x"00000000", 29939 => x"00000000",
    29940 => x"00000000", 29941 => x"00000000", 29942 => x"00000000",
    29943 => x"00000000", 29944 => x"00000000", 29945 => x"00000000",
    29946 => x"00000000", 29947 => x"00000000", 29948 => x"00000000",
    29949 => x"00000000", 29950 => x"00000000", 29951 => x"00000000",
    29952 => x"00000000", 29953 => x"00000000", 29954 => x"00000000",
    29955 => x"00000000", 29956 => x"00000000", 29957 => x"00000000",
    29958 => x"00000000", 29959 => x"00000000", 29960 => x"00000000",
    29961 => x"00000000", 29962 => x"00000000", 29963 => x"00000000",
    29964 => x"00000000", 29965 => x"00000000", 29966 => x"00000000",
    29967 => x"00000000", 29968 => x"00000000", 29969 => x"00000000",
    29970 => x"00000000", 29971 => x"00000000", 29972 => x"00000000",
    29973 => x"00000000", 29974 => x"00000000", 29975 => x"00000000",
    29976 => x"00000000", 29977 => x"00000000", 29978 => x"00000000",
    29979 => x"00000000", 29980 => x"00000000", 29981 => x"00000000",
    29982 => x"00000000", 29983 => x"00000000", 29984 => x"00000000",
    29985 => x"00000000", 29986 => x"00000000", 29987 => x"00000000",
    29988 => x"00000000", 29989 => x"00000000", 29990 => x"00000000",
    29991 => x"00000000", 29992 => x"00000000", 29993 => x"00000000",
    29994 => x"00000000", 29995 => x"00000000", 29996 => x"00000000",
    29997 => x"00000000", 29998 => x"00000000", 29999 => x"00000000",
    30000 => x"00000000", 30001 => x"00000000", 30002 => x"00000000",
    30003 => x"00000000", 30004 => x"00000000", 30005 => x"00000000",
    30006 => x"00000000", 30007 => x"00000000", 30008 => x"00000000",
    30009 => x"00000000", 30010 => x"00000000", 30011 => x"00000000",
    30012 => x"00000000", 30013 => x"00000000", 30014 => x"00000000",
    30015 => x"00000000", 30016 => x"00000000", 30017 => x"00000000",
    30018 => x"00000000", 30019 => x"00000000", 30020 => x"00000000",
    30021 => x"00000000", 30022 => x"00000000", 30023 => x"00000000",
    30024 => x"00000000", 30025 => x"00000000", 30026 => x"00000000",
    30027 => x"00000000", 30028 => x"00000000", 30029 => x"00000000",
    30030 => x"00000000", 30031 => x"00000000", 30032 => x"00000000",
    30033 => x"00000000", 30034 => x"00000000", 30035 => x"00000000",
    30036 => x"00000000", 30037 => x"00000000", 30038 => x"00000000",
    30039 => x"00000000", 30040 => x"00000000", 30041 => x"00000000",
    30042 => x"00000000", 30043 => x"00000000", 30044 => x"00000000",
    30045 => x"00000000", 30046 => x"00000000", 30047 => x"00000000",
    30048 => x"00000000", 30049 => x"00000000", 30050 => x"00000000",
    30051 => x"00000000", 30052 => x"00000000", 30053 => x"00000000",
    30054 => x"00000000", 30055 => x"00000000", 30056 => x"00000000",
    30057 => x"00000000", 30058 => x"00000000", 30059 => x"00000000",
    30060 => x"00000000", 30061 => x"00000000", 30062 => x"00000000",
    30063 => x"00000000", 30064 => x"00000000", 30065 => x"00000000",
    30066 => x"00000000", 30067 => x"00000000", 30068 => x"00000000",
    30069 => x"00000000", 30070 => x"00000000", 30071 => x"00000000",
    30072 => x"00000000", 30073 => x"00000000", 30074 => x"00000000",
    30075 => x"00000000", 30076 => x"00000000", 30077 => x"00000000",
    30078 => x"00000000", 30079 => x"00000000", 30080 => x"00000000",
    30081 => x"00000000", 30082 => x"00000000", 30083 => x"00000000",
    30084 => x"00000000", 30085 => x"00000000", 30086 => x"00000000",
    30087 => x"00000000", 30088 => x"00000000", 30089 => x"00000000",
    30090 => x"00000000", 30091 => x"00000000", 30092 => x"00000000",
    30093 => x"00000000", 30094 => x"00000000", 30095 => x"00000000",
    30096 => x"00000000", 30097 => x"00000000", 30098 => x"00000000",
    30099 => x"00000000", 30100 => x"00000000", 30101 => x"00000000",
    30102 => x"00000000", 30103 => x"00000000", 30104 => x"00000000",
    30105 => x"00000000", 30106 => x"00000000", 30107 => x"00000000",
    30108 => x"00000000", 30109 => x"00000000", 30110 => x"00000000",
    30111 => x"00000000", 30112 => x"00000000", 30113 => x"00000000",
    30114 => x"00000000", 30115 => x"00000000", 30116 => x"00000000",
    30117 => x"00000000", 30118 => x"00000000", 30119 => x"00000000",
    30120 => x"00000000", 30121 => x"00000000", 30122 => x"00000000",
    30123 => x"00000000", 30124 => x"00000000", 30125 => x"00000000",
    30126 => x"00000000", 30127 => x"00000000", 30128 => x"00000000",
    30129 => x"00000000", 30130 => x"00000000", 30131 => x"00000000",
    30132 => x"00000000", 30133 => x"00000000", 30134 => x"00000000",
    30135 => x"00000000", 30136 => x"00000000", 30137 => x"00000000",
    30138 => x"00000000", 30139 => x"00000000", 30140 => x"00000000",
    30141 => x"00000000", 30142 => x"00000000", 30143 => x"00000000",
    30144 => x"00000000", 30145 => x"00000000", 30146 => x"00000000",
    30147 => x"00000000", 30148 => x"00000000", 30149 => x"00000000",
    30150 => x"00000000", 30151 => x"00000000", 30152 => x"00000000",
    30153 => x"00000000", 30154 => x"00000000", 30155 => x"00000000",
    30156 => x"00000000", 30157 => x"00000000", 30158 => x"00000000",
    30159 => x"00000000", 30160 => x"00000000", 30161 => x"00000000",
    30162 => x"00000000", 30163 => x"00000000", 30164 => x"00000000",
    30165 => x"00000000", 30166 => x"00000000", 30167 => x"00000000",
    30168 => x"00000000", 30169 => x"00000000", 30170 => x"00000000",
    30171 => x"00000000", 30172 => x"00000000", 30173 => x"00000000",
    30174 => x"00000000", 30175 => x"00000000", 30176 => x"00000000",
    30177 => x"00000000", 30178 => x"00000000", 30179 => x"00000000",
    30180 => x"00000000", 30181 => x"00000000", 30182 => x"00000000",
    30183 => x"00000000", 30184 => x"00000000", 30185 => x"00000000",
    30186 => x"00000000", 30187 => x"00000000", 30188 => x"00000000",
    30189 => x"00000000", 30190 => x"00000000", 30191 => x"00000000",
    30192 => x"00000000", 30193 => x"00000000", 30194 => x"00000000",
    30195 => x"00000000", 30196 => x"00000000", 30197 => x"00000000",
    30198 => x"00000000", 30199 => x"00000000", 30200 => x"00000000",
    30201 => x"00000000", 30202 => x"00000000", 30203 => x"00000000",
    30204 => x"00000000", 30205 => x"00000000", 30206 => x"00000000",
    30207 => x"00000000", 30208 => x"00000000", 30209 => x"00000000",
    30210 => x"00000000", 30211 => x"00000000", 30212 => x"00000000",
    30213 => x"00000000", 30214 => x"00000000", 30215 => x"00000000",
    30216 => x"00000000", 30217 => x"00000000", 30218 => x"00000000",
    30219 => x"00000000", 30220 => x"00000000", 30221 => x"00000000",
    30222 => x"00000000", 30223 => x"00000000", 30224 => x"00000000",
    30225 => x"00000000", 30226 => x"00000000", 30227 => x"00000000",
    30228 => x"00000000", 30229 => x"00000000", 30230 => x"00000000",
    30231 => x"00000000", 30232 => x"00000000", 30233 => x"00000000",
    30234 => x"00000000", 30235 => x"00000000", 30236 => x"00000000",
    30237 => x"00000000", 30238 => x"00000000", 30239 => x"00000000",
    30240 => x"00000000", 30241 => x"00000000", 30242 => x"00000000",
    30243 => x"00000000", 30244 => x"00000000", 30245 => x"00000000",
    30246 => x"00000000", 30247 => x"00000000", 30248 => x"00000000",
    30249 => x"00000000", 30250 => x"00000000", 30251 => x"00000000",
    30252 => x"00000000", 30253 => x"00000000", 30254 => x"00000000",
    30255 => x"00000000", 30256 => x"00000000", 30257 => x"00000000",
    30258 => x"00000000", 30259 => x"00000000", 30260 => x"00000000",
    30261 => x"00000000", 30262 => x"00000000", 30263 => x"00000000",
    30264 => x"00000000", 30265 => x"00000000", 30266 => x"00000000",
    30267 => x"00000000", 30268 => x"00000000", 30269 => x"00000000",
    30270 => x"00000000", 30271 => x"00000000", 30272 => x"00000000",
    30273 => x"00000000", 30274 => x"00000000", 30275 => x"00000000",
    30276 => x"00000000", 30277 => x"00000000", 30278 => x"00000000",
    30279 => x"00000000", 30280 => x"00000000", 30281 => x"00000000",
    30282 => x"00000000", 30283 => x"00000000", 30284 => x"00000000",
    30285 => x"00000000", 30286 => x"00000000", 30287 => x"00000000",
    30288 => x"00000000", 30289 => x"00000000", 30290 => x"00000000",
    30291 => x"00000000", 30292 => x"00000000", 30293 => x"00000000",
    30294 => x"00000000", 30295 => x"00000000", 30296 => x"00000000",
    30297 => x"00000000", 30298 => x"00000000", 30299 => x"00000000",
    30300 => x"00000000", 30301 => x"00000000", 30302 => x"00000000",
    30303 => x"00000000", 30304 => x"00000000", 30305 => x"00000000",
    30306 => x"00000000", 30307 => x"00000000", 30308 => x"00000000",
    30309 => x"00000000", 30310 => x"00000000", 30311 => x"00000000",
    30312 => x"00000000", 30313 => x"00000000", 30314 => x"00000000",
    30315 => x"00000000", 30316 => x"00000000", 30317 => x"00000000",
    30318 => x"00000000", 30319 => x"00000000", 30320 => x"00000000",
    30321 => x"00000000", 30322 => x"00000000", 30323 => x"00000000",
    30324 => x"00000000", 30325 => x"00000000", 30326 => x"00000000",
    30327 => x"00000000", 30328 => x"00000000", 30329 => x"00000000",
    30330 => x"00000000", 30331 => x"00000000", 30332 => x"00000000",
    30333 => x"00000000", 30334 => x"00000000", 30335 => x"00000000",
    30336 => x"00000000", 30337 => x"00000000", 30338 => x"00000000",
    30339 => x"00000000", 30340 => x"00000000", 30341 => x"00000000",
    30342 => x"00000000", 30343 => x"00000000", 30344 => x"00000000",
    30345 => x"00000000", 30346 => x"00000000", 30347 => x"00000000",
    30348 => x"00000000", 30349 => x"00000000", 30350 => x"00000000",
    30351 => x"00000000", 30352 => x"00000000", 30353 => x"00000000",
    30354 => x"00000000", 30355 => x"00000000", 30356 => x"00000000",
    30357 => x"00000000", 30358 => x"00000000", 30359 => x"00000000",
    30360 => x"00000000", 30361 => x"00000000", 30362 => x"00000000",
    30363 => x"00000000", 30364 => x"00000000", 30365 => x"00000000",
    30366 => x"00000000", 30367 => x"00000000", 30368 => x"00000000",
    30369 => x"00000000", 30370 => x"00000000", 30371 => x"00000000",
    30372 => x"00000000", 30373 => x"00000000", 30374 => x"00000000",
    30375 => x"00000000", 30376 => x"00000000", 30377 => x"00000000",
    30378 => x"00000000", 30379 => x"00000000", 30380 => x"00000000",
    30381 => x"00000000", 30382 => x"00000000", 30383 => x"00000000",
    30384 => x"00000000", 30385 => x"00000000", 30386 => x"00000000",
    30387 => x"00000000", 30388 => x"00000000", 30389 => x"00000000",
    30390 => x"00000000", 30391 => x"00000000", 30392 => x"00000000",
    30393 => x"00000000", 30394 => x"00000000", 30395 => x"00000000",
    30396 => x"00000000", 30397 => x"00000000", 30398 => x"00000000",
    30399 => x"00000000", 30400 => x"00000000", 30401 => x"00000000",
    30402 => x"00000000", 30403 => x"00000000", 30404 => x"00000000",
    30405 => x"00000000", 30406 => x"00000000", 30407 => x"00000000",
    30408 => x"00000000", 30409 => x"00000000", 30410 => x"00000000",
    30411 => x"00000000", 30412 => x"00000000", 30413 => x"00000000",
    30414 => x"00000000", 30415 => x"00000000", 30416 => x"00000000",
    30417 => x"00000000", 30418 => x"00000000", 30419 => x"00000000",
    30420 => x"00000000", 30421 => x"00000000", 30422 => x"00000000",
    30423 => x"00000000", 30424 => x"00000000", 30425 => x"00000000",
    30426 => x"00000000", 30427 => x"00000000", 30428 => x"00000000",
    30429 => x"00000000", 30430 => x"00000000", 30431 => x"00000000",
    30432 => x"00000000", 30433 => x"00000000", 30434 => x"00000000",
    30435 => x"00000000", 30436 => x"00000000", 30437 => x"00000000",
    30438 => x"00000000", 30439 => x"00000000", 30440 => x"00000000",
    30441 => x"00000000", 30442 => x"00000000", 30443 => x"00000000",
    30444 => x"00000000", 30445 => x"00000000", 30446 => x"00000000",
    30447 => x"00000000", 30448 => x"00000000", 30449 => x"00000000",
    30450 => x"00000000", 30451 => x"00000000", 30452 => x"00000000",
    30453 => x"00000000", 30454 => x"00000000", 30455 => x"00000000",
    30456 => x"00000000", 30457 => x"00000000", 30458 => x"00000000",
    30459 => x"00000000", 30460 => x"00000000", 30461 => x"00000000",
    30462 => x"00000000", 30463 => x"00000000", 30464 => x"00000000",
    30465 => x"00000000", 30466 => x"00000000", 30467 => x"00000000",
    30468 => x"00000000", 30469 => x"00000000", 30470 => x"00000000",
    30471 => x"00000000", 30472 => x"00000000", 30473 => x"00000000",
    30474 => x"00000000", 30475 => x"00000000", 30476 => x"00000000",
    30477 => x"00000000", 30478 => x"00000000", 30479 => x"00000000",
    30480 => x"00000000", 30481 => x"00000000", 30482 => x"00000000",
    30483 => x"00000000", 30484 => x"00000000", 30485 => x"00000000",
    30486 => x"00000000", 30487 => x"00000000", 30488 => x"00000000",
    30489 => x"00000000", 30490 => x"00000000", 30491 => x"00000000",
    30492 => x"00000000", 30493 => x"00000000", 30494 => x"00000000",
    30495 => x"00000000", 30496 => x"00000000", 30497 => x"00000000",
    30498 => x"00000000", 30499 => x"00000000", 30500 => x"00000000",
    30501 => x"00000000", 30502 => x"00000000", 30503 => x"00000000",
    30504 => x"00000000", 30505 => x"00000000", 30506 => x"00000000",
    30507 => x"00000000", 30508 => x"00000000", 30509 => x"00000000",
    30510 => x"00000000", 30511 => x"00000000", 30512 => x"00000000",
    30513 => x"00000000", 30514 => x"00000000", 30515 => x"00000000",
    30516 => x"00000000", 30517 => x"00000000", 30518 => x"00000000",
    30519 => x"00000000", 30520 => x"00000000", 30521 => x"00000000",
    30522 => x"00000000", 30523 => x"00000000", 30524 => x"00000000",
    30525 => x"00000000", 30526 => x"00000000", 30527 => x"00000000",
    30528 => x"00000000", 30529 => x"00000000", 30530 => x"00000000",
    30531 => x"00000000", 30532 => x"00000000", 30533 => x"00000000",
    30534 => x"00000000", 30535 => x"00000000", 30536 => x"00000000",
    30537 => x"00000000", 30538 => x"00000000", 30539 => x"00000000",
    30540 => x"00000000", 30541 => x"00000000", 30542 => x"00000000",
    30543 => x"00000000", 30544 => x"00000000", 30545 => x"00000000",
    30546 => x"00000000", 30547 => x"00000000", 30548 => x"00000000",
    30549 => x"00000000", 30550 => x"00000000", 30551 => x"00000000",
    30552 => x"00000000", 30553 => x"00000000", 30554 => x"00000000",
    30555 => x"00000000", 30556 => x"00000000", 30557 => x"00000000",
    30558 => x"00000000", 30559 => x"00000000", 30560 => x"00000000",
    30561 => x"00000000", 30562 => x"00000000", 30563 => x"00000000",
    30564 => x"00000000", 30565 => x"00000000", 30566 => x"00000000",
    30567 => x"00000000", 30568 => x"00000000", 30569 => x"00000000",
    30570 => x"00000000", 30571 => x"00000000", 30572 => x"00000000",
    30573 => x"00000000", 30574 => x"00000000", 30575 => x"00000000",
    30576 => x"00000000", 30577 => x"00000000", 30578 => x"00000000",
    30579 => x"00000000", 30580 => x"00000000", 30581 => x"00000000",
    30582 => x"00000000", 30583 => x"00000000", 30584 => x"00000000",
    30585 => x"00000000", 30586 => x"00000000", 30587 => x"00000000",
    30588 => x"00000000", 30589 => x"00000000", 30590 => x"00000000",
    30591 => x"00000000", 30592 => x"00000000", 30593 => x"00000000",
    30594 => x"00000000", 30595 => x"00000000", 30596 => x"00000000",
    30597 => x"00000000", 30598 => x"00000000", 30599 => x"00000000",
    30600 => x"00000000", 30601 => x"00000000", 30602 => x"00000000",
    30603 => x"00000000", 30604 => x"00000000", 30605 => x"00000000",
    30606 => x"00000000", 30607 => x"00000000", 30608 => x"00000000",
    30609 => x"00000000", 30610 => x"00000000", 30611 => x"00000000",
    30612 => x"00000000", 30613 => x"00000000", 30614 => x"00000000",
    30615 => x"00000000", 30616 => x"00000000", 30617 => x"00000000",
    30618 => x"00000000", 30619 => x"00000000", 30620 => x"00000000",
    30621 => x"00000000", 30622 => x"00000000", 30623 => x"00000000",
    30624 => x"00000000", 30625 => x"00000000", 30626 => x"00000000",
    30627 => x"00000000", 30628 => x"00000000", 30629 => x"00000000",
    30630 => x"00000000", 30631 => x"00000000", 30632 => x"00000000",
    30633 => x"00000000", 30634 => x"00000000", 30635 => x"00000000",
    30636 => x"00000000", 30637 => x"00000000", 30638 => x"00000000",
    30639 => x"00000000", 30640 => x"00000000", 30641 => x"00000000",
    30642 => x"00000000", 30643 => x"00000000", 30644 => x"00000000",
    30645 => x"00000000", 30646 => x"00000000", 30647 => x"00000000",
    30648 => x"00000000", 30649 => x"00000000", 30650 => x"00000000",
    30651 => x"00000000", 30652 => x"00000000", 30653 => x"00000000",
    30654 => x"00000000", 30655 => x"00000000", 30656 => x"00000000",
    30657 => x"00000000", 30658 => x"00000000", 30659 => x"00000000",
    30660 => x"00000000", 30661 => x"00000000", 30662 => x"00000000",
    30663 => x"00000000", 30664 => x"00000000", 30665 => x"00000000",
    30666 => x"00000000", 30667 => x"00000000", 30668 => x"00000000",
    30669 => x"00000000", 30670 => x"00000000", 30671 => x"00000000",
    30672 => x"00000000", 30673 => x"00000000", 30674 => x"00000000",
    30675 => x"00000000", 30676 => x"00000000", 30677 => x"00000000",
    30678 => x"00000000", 30679 => x"00000000", 30680 => x"00000000",
    30681 => x"00000000", 30682 => x"00000000", 30683 => x"00000000",
    30684 => x"00000000", 30685 => x"00000000", 30686 => x"00000000",
    30687 => x"00000000", 30688 => x"00000000", 30689 => x"00000000",
    30690 => x"00000000", 30691 => x"00000000", 30692 => x"00000000",
    30693 => x"00000000", 30694 => x"00000000", 30695 => x"00000000",
    30696 => x"00000000", 30697 => x"00000000", 30698 => x"00000000",
    30699 => x"00000000", 30700 => x"00000000", 30701 => x"00000000",
    30702 => x"00000000", 30703 => x"00000000", 30704 => x"00000000",
    30705 => x"00000000", 30706 => x"00000000", 30707 => x"00000000",
    30708 => x"00000000", 30709 => x"00000000", 30710 => x"00000000",
    30711 => x"00000000", 30712 => x"00000000", 30713 => x"00000000",
    30714 => x"00000000", 30715 => x"00000000", 30716 => x"00000000",
    30717 => x"00000000", 30718 => x"00000000", 30719 => x"00000000",
    30720 => x"00000000", 30721 => x"00000000", 30722 => x"00000000",
    30723 => x"00000000", 30724 => x"00000000", 30725 => x"00000000",
    30726 => x"00000000", 30727 => x"00000000", 30728 => x"00000000",
    30729 => x"00000000", 30730 => x"00000000", 30731 => x"00000000",
    30732 => x"00000000", 30733 => x"00000000", 30734 => x"00000000",
    30735 => x"00000000", 30736 => x"00000000", 30737 => x"00000000",
    30738 => x"00000000", 30739 => x"00000000", 30740 => x"00000000",
    30741 => x"00000000", 30742 => x"00000000", 30743 => x"00000000",
    30744 => x"00000000", 30745 => x"00000000", 30746 => x"00000000",
    30747 => x"00000000", 30748 => x"00000000", 30749 => x"00000000",
    30750 => x"00000000", 30751 => x"00000000", 30752 => x"00000000",
    30753 => x"00000000", 30754 => x"00000000", 30755 => x"00000000",
    30756 => x"00000000", 30757 => x"00000000", 30758 => x"00000000",
    30759 => x"00000000", 30760 => x"00000000", 30761 => x"00000000",
    30762 => x"00000000", 30763 => x"00000000", 30764 => x"00000000",
    30765 => x"00000000", 30766 => x"00000000", 30767 => x"00000000",
    30768 => x"00000000", 30769 => x"00000000", 30770 => x"00000000",
    30771 => x"00000000", 30772 => x"00000000", 30773 => x"00000000",
    30774 => x"00000000", 30775 => x"00000000", 30776 => x"00000000",
    30777 => x"00000000", 30778 => x"00000000", 30779 => x"00000000",
    30780 => x"00000000", 30781 => x"00000000", 30782 => x"00000000",
    30783 => x"00000000", 30784 => x"00000000", 30785 => x"00000000",
    30786 => x"00000000", 30787 => x"00000000", 30788 => x"00000000",
    30789 => x"00000000", 30790 => x"00000000", 30791 => x"00000000",
    30792 => x"00000000", 30793 => x"00000000", 30794 => x"00000000",
    30795 => x"00000000", 30796 => x"00000000", 30797 => x"00000000",
    30798 => x"00000000", 30799 => x"00000000", 30800 => x"00000000",
    30801 => x"00000000", 30802 => x"00000000", 30803 => x"00000000",
    30804 => x"00000000", 30805 => x"00000000", 30806 => x"00000000",
    30807 => x"00000000", 30808 => x"00000000", 30809 => x"00000000",
    30810 => x"00000000", 30811 => x"00000000", 30812 => x"00000000",
    30813 => x"00000000", 30814 => x"00000000", 30815 => x"00000000",
    30816 => x"00000000", 30817 => x"00000000", 30818 => x"00000000",
    30819 => x"00000000", 30820 => x"00000000", 30821 => x"00000000",
    30822 => x"00000000", 30823 => x"00000000", 30824 => x"00000000",
    30825 => x"00000000", 30826 => x"00000000", 30827 => x"00000000",
    30828 => x"00000000", 30829 => x"00000000", 30830 => x"00000000",
    30831 => x"00000000", 30832 => x"00000000", 30833 => x"00000000",
    30834 => x"00000000", 30835 => x"00000000", 30836 => x"00000000",
    30837 => x"00000000", 30838 => x"00000000", 30839 => x"00000000",
    30840 => x"00000000", 30841 => x"00000000", 30842 => x"00000000",
    30843 => x"00000000", 30844 => x"00000000", 30845 => x"00000000",
    30846 => x"00000000", 30847 => x"00000000", 30848 => x"00000000",
    30849 => x"00000000", 30850 => x"00000000", 30851 => x"00000000",
    30852 => x"00000000", 30853 => x"00000000", 30854 => x"00000000",
    30855 => x"00000000", 30856 => x"00000000", 30857 => x"00000000",
    30858 => x"00000000", 30859 => x"00000000", 30860 => x"00000000",
    30861 => x"00000000", 30862 => x"00000000", 30863 => x"00000000",
    30864 => x"00000000", 30865 => x"00000000", 30866 => x"00000000",
    30867 => x"00000000", 30868 => x"00000000", 30869 => x"00000000",
    30870 => x"00000000", 30871 => x"00000000", 30872 => x"00000000",
    30873 => x"00000000", 30874 => x"00000000", 30875 => x"00000000",
    30876 => x"00000000", 30877 => x"00000000", 30878 => x"00000000",
    30879 => x"00000000", 30880 => x"00000000", 30881 => x"00000000",
    30882 => x"00000000", 30883 => x"00000000", 30884 => x"00000000",
    30885 => x"00000000", 30886 => x"00000000", 30887 => x"00000000",
    30888 => x"00000000", 30889 => x"00000000", 30890 => x"00000000",
    30891 => x"00000000", 30892 => x"00000000", 30893 => x"00000000",
    30894 => x"00000000", 30895 => x"00000000", 30896 => x"00000000",
    30897 => x"00000000", 30898 => x"00000000", 30899 => x"00000000",
    30900 => x"00000000", 30901 => x"00000000", 30902 => x"00000000",
    30903 => x"00000000", 30904 => x"00000000", 30905 => x"00000000",
    30906 => x"00000000", 30907 => x"00000000", 30908 => x"00000000",
    30909 => x"00000000", 30910 => x"00000000", 30911 => x"00000000",
    30912 => x"00000000", 30913 => x"00000000", 30914 => x"00000000",
    30915 => x"00000000", 30916 => x"00000000", 30917 => x"00000000",
    30918 => x"00000000", 30919 => x"00000000", 30920 => x"00000000",
    30921 => x"00000000", 30922 => x"00000000", 30923 => x"00000000",
    30924 => x"00000000", 30925 => x"00000000", 30926 => x"00000000",
    30927 => x"00000000", 30928 => x"00000000", 30929 => x"00000000",
    30930 => x"00000000", 30931 => x"00000000", 30932 => x"00000000",
    30933 => x"00000000", 30934 => x"00000000", 30935 => x"00000000",
    30936 => x"00000000", 30937 => x"00000000", 30938 => x"00000000",
    30939 => x"00000000", 30940 => x"00000000", 30941 => x"00000000",
    30942 => x"00000000", 30943 => x"00000000", 30944 => x"00000000",
    30945 => x"00000000", 30946 => x"00000000", 30947 => x"00000000",
    30948 => x"00000000", 30949 => x"00000000", 30950 => x"00000000",
    30951 => x"00000000", 30952 => x"00000000", 30953 => x"00000000",
    30954 => x"00000000", 30955 => x"00000000", 30956 => x"00000000",
    30957 => x"00000000", 30958 => x"00000000", 30959 => x"00000000",
    30960 => x"00000000", 30961 => x"00000000", 30962 => x"00000000",
    30963 => x"00000000", 30964 => x"00000000", 30965 => x"00000000",
    30966 => x"00000000", 30967 => x"00000000", 30968 => x"00000000",
    30969 => x"00000000", 30970 => x"00000000", 30971 => x"00000000",
    30972 => x"00000000", 30973 => x"00000000", 30974 => x"00000000",
    30975 => x"00000000", 30976 => x"00000000", 30977 => x"00000000",
    30978 => x"00000000", 30979 => x"00000000", 30980 => x"00000000",
    30981 => x"00000000", 30982 => x"00000000", 30983 => x"00000000",
    30984 => x"00000000", 30985 => x"00000000", 30986 => x"00000000",
    30987 => x"00000000", 30988 => x"00000000", 30989 => x"00000000",
    30990 => x"00000000", 30991 => x"00000000", 30992 => x"00000000",
    30993 => x"00000000", 30994 => x"00000000", 30995 => x"00000000",
    30996 => x"00000000", 30997 => x"00000000", 30998 => x"00000000",
    30999 => x"00000000", 31000 => x"00000000", 31001 => x"00000000",
    31002 => x"00000000", 31003 => x"00000000", 31004 => x"00000000",
    31005 => x"00000000", 31006 => x"00000000", 31007 => x"00000000",
    31008 => x"00000000", 31009 => x"00000000", 31010 => x"00000000",
    31011 => x"00000000", 31012 => x"00000000", 31013 => x"00000000",
    31014 => x"00000000", 31015 => x"00000000", 31016 => x"00000000",
    31017 => x"00000000", 31018 => x"00000000", 31019 => x"00000000",
    31020 => x"00000000", 31021 => x"00000000", 31022 => x"00000000",
    31023 => x"00000000", 31024 => x"00000000", 31025 => x"00000000",
    31026 => x"00000000", 31027 => x"00000000", 31028 => x"00000000",
    31029 => x"00000000", 31030 => x"00000000", 31031 => x"00000000",
    31032 => x"00000000", 31033 => x"00000000", 31034 => x"00000000",
    31035 => x"00000000", 31036 => x"00000000", 31037 => x"00000000",
    31038 => x"00000000", 31039 => x"00000000", 31040 => x"00000000",
    31041 => x"00000000", 31042 => x"00000000", 31043 => x"00000000",
    31044 => x"00000000", 31045 => x"00000000", 31046 => x"00000000",
    31047 => x"00000000", 31048 => x"00000000", 31049 => x"00000000",
    31050 => x"00000000", 31051 => x"00000000", 31052 => x"00000000",
    31053 => x"00000000", 31054 => x"00000000", 31055 => x"00000000",
    31056 => x"00000000", 31057 => x"00000000", 31058 => x"00000000",
    31059 => x"00000000", 31060 => x"00000000", 31061 => x"00000000",
    31062 => x"00000000", 31063 => x"00000000", 31064 => x"00000000",
    31065 => x"00000000", 31066 => x"00000000", 31067 => x"00000000",
    31068 => x"00000000", 31069 => x"00000000", 31070 => x"00000000",
    31071 => x"00000000", 31072 => x"00000000", 31073 => x"00000000",
    31074 => x"00000000", 31075 => x"00000000", 31076 => x"00000000",
    31077 => x"00000000", 31078 => x"00000000", 31079 => x"00000000",
    31080 => x"00000000", 31081 => x"00000000", 31082 => x"00000000",
    31083 => x"00000000", 31084 => x"00000000", 31085 => x"00000000",
    31086 => x"00000000", 31087 => x"00000000", 31088 => x"00000000",
    31089 => x"00000000", 31090 => x"00000000", 31091 => x"00000000",
    31092 => x"00000000", 31093 => x"00000000", 31094 => x"00000000",
    31095 => x"00000000", 31096 => x"00000000", 31097 => x"00000000",
    31098 => x"00000000", 31099 => x"00000000", 31100 => x"00000000",
    31101 => x"00000000", 31102 => x"00000000", 31103 => x"00000000",
    31104 => x"00000000", 31105 => x"00000000", 31106 => x"00000000",
    31107 => x"00000000", 31108 => x"00000000", 31109 => x"00000000",
    31110 => x"00000000", 31111 => x"00000000", 31112 => x"00000000",
    31113 => x"00000000", 31114 => x"00000000", 31115 => x"00000000",
    31116 => x"00000000", 31117 => x"00000000", 31118 => x"00000000",
    31119 => x"00000000", 31120 => x"00000000", 31121 => x"00000000",
    31122 => x"00000000", 31123 => x"00000000", 31124 => x"00000000",
    31125 => x"00000000", 31126 => x"00000000", 31127 => x"00000000",
    31128 => x"00000000", 31129 => x"00000000", 31130 => x"00000000",
    31131 => x"00000000", 31132 => x"00000000", 31133 => x"00000000",
    31134 => x"00000000", 31135 => x"00000000", 31136 => x"00000000",
    31137 => x"00000000", 31138 => x"00000000", 31139 => x"00000000",
    31140 => x"00000000", 31141 => x"00000000", 31142 => x"00000000",
    31143 => x"00000000", 31144 => x"00000000", 31145 => x"00000000",
    31146 => x"00000000", 31147 => x"00000000", 31148 => x"00000000",
    31149 => x"00000000", 31150 => x"00000000", 31151 => x"00000000",
    31152 => x"00000000", 31153 => x"00000000", 31154 => x"00000000",
    31155 => x"00000000", 31156 => x"00000000", 31157 => x"00000000",
    31158 => x"00000000", 31159 => x"00000000", 31160 => x"00000000",
    31161 => x"00000000", 31162 => x"00000000", 31163 => x"00000000",
    31164 => x"00000000", 31165 => x"00000000", 31166 => x"00000000",
    31167 => x"00000000", 31168 => x"00000000", 31169 => x"00000000",
    31170 => x"00000000", 31171 => x"00000000", 31172 => x"00000000",
    31173 => x"00000000", 31174 => x"00000000", 31175 => x"00000000",
    31176 => x"00000000", 31177 => x"00000000", 31178 => x"00000000",
    31179 => x"00000000", 31180 => x"00000000", 31181 => x"00000000",
    31182 => x"00000000", 31183 => x"00000000", 31184 => x"00000000",
    31185 => x"00000000", 31186 => x"00000000", 31187 => x"00000000",
    31188 => x"00000000", 31189 => x"00000000", 31190 => x"00000000",
    31191 => x"00000000", 31192 => x"00000000", 31193 => x"00000000",
    31194 => x"00000000", 31195 => x"00000000", 31196 => x"00000000",
    31197 => x"00000000", 31198 => x"00000000", 31199 => x"00000000",
    31200 => x"00000000", 31201 => x"00000000", 31202 => x"00000000",
    31203 => x"00000000", 31204 => x"00000000", 31205 => x"00000000",
    31206 => x"00000000", 31207 => x"00000000", 31208 => x"00000000",
    31209 => x"00000000", 31210 => x"00000000", 31211 => x"00000000",
    31212 => x"00000000", 31213 => x"00000000", 31214 => x"00000000",
    31215 => x"00000000", 31216 => x"00000000", 31217 => x"00000000",
    31218 => x"00000000", 31219 => x"00000000", 31220 => x"00000000",
    31221 => x"00000000", 31222 => x"00000000", 31223 => x"00000000",
    31224 => x"00000000", 31225 => x"00000000", 31226 => x"00000000",
    31227 => x"00000000", 31228 => x"00000000", 31229 => x"00000000",
    31230 => x"00000000", 31231 => x"00000000", 31232 => x"00000000",
    31233 => x"00000000", 31234 => x"00000000", 31235 => x"00000000",
    31236 => x"00000000", 31237 => x"00000000", 31238 => x"00000000",
    31239 => x"00000000", 31240 => x"00000000", 31241 => x"00000000",
    31242 => x"00000000", 31243 => x"00000000", 31244 => x"00000000",
    31245 => x"00000000", 31246 => x"00000000", 31247 => x"00000000",
    31248 => x"00000000", 31249 => x"00000000", 31250 => x"00000000",
    31251 => x"00000000", 31252 => x"00000000", 31253 => x"00000000",
    31254 => x"00000000", 31255 => x"00000000", 31256 => x"00000000",
    31257 => x"00000000", 31258 => x"00000000", 31259 => x"00000000",
    31260 => x"00000000", 31261 => x"00000000", 31262 => x"00000000",
    31263 => x"00000000", 31264 => x"00000000", 31265 => x"00000000",
    31266 => x"00000000", 31267 => x"00000000", 31268 => x"00000000",
    31269 => x"00000000", 31270 => x"00000000", 31271 => x"00000000",
    31272 => x"00000000", 31273 => x"00000000", 31274 => x"00000000",
    31275 => x"00000000", 31276 => x"00000000", 31277 => x"00000000",
    31278 => x"00000000", 31279 => x"00000000", 31280 => x"00000000",
    31281 => x"00000000", 31282 => x"00000000", 31283 => x"00000000",
    31284 => x"00000000", 31285 => x"00000000", 31286 => x"00000000",
    31287 => x"00000000", 31288 => x"00000000", 31289 => x"00000000",
    31290 => x"00000000", 31291 => x"00000000", 31292 => x"00000000",
    31293 => x"00000000", 31294 => x"00000000", 31295 => x"00000000",
    31296 => x"00000000", 31297 => x"00000000", 31298 => x"00000000",
    31299 => x"00000000", 31300 => x"00000000", 31301 => x"00000000",
    31302 => x"00000000", 31303 => x"00000000", 31304 => x"00000000",
    31305 => x"00000000", 31306 => x"00000000", 31307 => x"00000000",
    31308 => x"00000000", 31309 => x"00000000", 31310 => x"00000000",
    31311 => x"00000000", 31312 => x"00000000", 31313 => x"00000000",
    31314 => x"00000000", 31315 => x"00000000", 31316 => x"00000000",
    31317 => x"00000000", 31318 => x"00000000", 31319 => x"00000000",
    31320 => x"00000000", 31321 => x"00000000", 31322 => x"00000000",
    31323 => x"00000000", 31324 => x"00000000", 31325 => x"00000000",
    31326 => x"00000000", 31327 => x"00000000", 31328 => x"00000000",
    31329 => x"00000000", 31330 => x"00000000", 31331 => x"00000000",
    31332 => x"00000000", 31333 => x"00000000", 31334 => x"00000000",
    31335 => x"00000000", 31336 => x"00000000", 31337 => x"00000000",
    31338 => x"00000000", 31339 => x"00000000", 31340 => x"00000000",
    31341 => x"00000000", 31342 => x"00000000", 31343 => x"00000000",
    31344 => x"00000000", 31345 => x"00000000", 31346 => x"00000000",
    31347 => x"00000000", 31348 => x"00000000", 31349 => x"00000000",
    31350 => x"00000000", 31351 => x"00000000", 31352 => x"00000000",
    31353 => x"00000000", 31354 => x"00000000", 31355 => x"00000000",
    31356 => x"00000000", 31357 => x"00000000", 31358 => x"00000000",
    31359 => x"00000000", 31360 => x"00000000", 31361 => x"00000000",
    31362 => x"00000000", 31363 => x"00000000", 31364 => x"00000000",
    31365 => x"00000000", 31366 => x"00000000", 31367 => x"00000000",
    31368 => x"00000000", 31369 => x"00000000", 31370 => x"00000000",
    31371 => x"00000000", 31372 => x"00000000", 31373 => x"00000000",
    31374 => x"00000000", 31375 => x"00000000", 31376 => x"00000000",
    31377 => x"00000000", 31378 => x"00000000", 31379 => x"00000000",
    31380 => x"00000000", 31381 => x"00000000", 31382 => x"00000000",
    31383 => x"00000000", 31384 => x"00000000", 31385 => x"00000000",
    31386 => x"00000000", 31387 => x"00000000", 31388 => x"00000000",
    31389 => x"00000000", 31390 => x"00000000", 31391 => x"00000000",
    31392 => x"00000000", 31393 => x"00000000", 31394 => x"00000000",
    31395 => x"00000000", 31396 => x"00000000", 31397 => x"00000000",
    31398 => x"00000000", 31399 => x"00000000", 31400 => x"00000000",
    31401 => x"00000000", 31402 => x"00000000", 31403 => x"00000000",
    31404 => x"00000000", 31405 => x"00000000", 31406 => x"00000000",
    31407 => x"00000000", 31408 => x"00000000", 31409 => x"00000000",
    31410 => x"00000000", 31411 => x"00000000", 31412 => x"00000000",
    31413 => x"00000000", 31414 => x"00000000", 31415 => x"00000000",
    31416 => x"00000000", 31417 => x"00000000", 31418 => x"00000000",
    31419 => x"00000000", 31420 => x"00000000", 31421 => x"00000000",
    31422 => x"00000000", 31423 => x"00000000", 31424 => x"00000000",
    31425 => x"00000000", 31426 => x"00000000", 31427 => x"00000000",
    31428 => x"00000000", 31429 => x"00000000", 31430 => x"00000000",
    31431 => x"00000000", 31432 => x"00000000", 31433 => x"00000000",
    31434 => x"00000000", 31435 => x"00000000", 31436 => x"00000000",
    31437 => x"00000000", 31438 => x"00000000", 31439 => x"00000000",
    31440 => x"00000000", 31441 => x"00000000", 31442 => x"00000000",
    31443 => x"00000000", 31444 => x"00000000", 31445 => x"00000000",
    31446 => x"00000000", 31447 => x"00000000", 31448 => x"00000000",
    31449 => x"00000000", 31450 => x"00000000", 31451 => x"00000000",
    31452 => x"00000000", 31453 => x"00000000", 31454 => x"00000000",
    31455 => x"00000000", 31456 => x"00000000", 31457 => x"00000000",
    31458 => x"00000000", 31459 => x"00000000", 31460 => x"00000000",
    31461 => x"00000000", 31462 => x"00000000", 31463 => x"00000000",
    31464 => x"00000000", 31465 => x"00000000", 31466 => x"00000000",
    31467 => x"00000000", 31468 => x"00000000", 31469 => x"00000000",
    31470 => x"00000000", 31471 => x"00000000", 31472 => x"00000000",
    31473 => x"00000000", 31474 => x"00000000", 31475 => x"00000000",
    31476 => x"00000000", 31477 => x"00000000", 31478 => x"00000000",
    31479 => x"00000000", 31480 => x"00000000", 31481 => x"00000000",
    31482 => x"00000000", 31483 => x"00000000", 31484 => x"00000000",
    31485 => x"00000000", 31486 => x"00000000", 31487 => x"00000000",
    31488 => x"00000000", 31489 => x"00000000", 31490 => x"00000000",
    31491 => x"00000000", 31492 => x"00000000", 31493 => x"00000000",
    31494 => x"00000000", 31495 => x"00000000", 31496 => x"00000000",
    31497 => x"00000000", 31498 => x"00000000", 31499 => x"00000000",
    31500 => x"00000000", 31501 => x"00000000", 31502 => x"00000000",
    31503 => x"00000000", 31504 => x"00000000", 31505 => x"00000000",
    31506 => x"00000000", 31507 => x"00000000", 31508 => x"00000000",
    31509 => x"00000000", 31510 => x"00000000", 31511 => x"00000000",
    31512 => x"00000000", 31513 => x"00000000", 31514 => x"00000000",
    31515 => x"00000000", 31516 => x"00000000", 31517 => x"00000000",
    31518 => x"00000000", 31519 => x"00000000", 31520 => x"00000000",
    31521 => x"00000000", 31522 => x"00000000", 31523 => x"00000000",
    31524 => x"00000000", 31525 => x"00000000", 31526 => x"00000000",
    31527 => x"00000000", 31528 => x"00000000", 31529 => x"00000000",
    31530 => x"00000000", 31531 => x"00000000", 31532 => x"00000000",
    31533 => x"00000000", 31534 => x"00000000", 31535 => x"00000000",
    31536 => x"00000000", 31537 => x"00000000", 31538 => x"00000000",
    31539 => x"00000000", 31540 => x"00000000", 31541 => x"00000000",
    31542 => x"00000000", 31543 => x"00000000", 31544 => x"00000000",
    31545 => x"00000000", 31546 => x"00000000", 31547 => x"00000000",
    31548 => x"00000000", 31549 => x"00000000", 31550 => x"00000000",
    31551 => x"00000000", 31552 => x"00000000", 31553 => x"00000000",
    31554 => x"00000000", 31555 => x"00000000", 31556 => x"00000000",
    31557 => x"00000000", 31558 => x"00000000", 31559 => x"00000000",
    31560 => x"00000000", 31561 => x"00000000", 31562 => x"00000000",
    31563 => x"00000000", 31564 => x"00000000", 31565 => x"00000000",
    31566 => x"00000000", 31567 => x"00000000", 31568 => x"00000000",
    31569 => x"00000000", 31570 => x"00000000", 31571 => x"00000000",
    31572 => x"00000000", 31573 => x"00000000", 31574 => x"00000000",
    31575 => x"00000000", 31576 => x"00000000", 31577 => x"00000000",
    31578 => x"00000000", 31579 => x"00000000", 31580 => x"00000000",
    31581 => x"00000000", 31582 => x"00000000", 31583 => x"00000000",
    31584 => x"00000000", 31585 => x"00000000", 31586 => x"00000000",
    31587 => x"00000000", 31588 => x"00000000", 31589 => x"00000000",
    31590 => x"00000000", 31591 => x"00000000", 31592 => x"00000000",
    31593 => x"00000000", 31594 => x"00000000", 31595 => x"00000000",
    31596 => x"00000000", 31597 => x"00000000", 31598 => x"00000000",
    31599 => x"00000000", 31600 => x"00000000", 31601 => x"00000000",
    31602 => x"00000000", 31603 => x"00000000", 31604 => x"00000000",
    31605 => x"00000000", 31606 => x"00000000", 31607 => x"00000000",
    31608 => x"00000000", 31609 => x"00000000", 31610 => x"00000000",
    31611 => x"00000000", 31612 => x"00000000", 31613 => x"00000000",
    31614 => x"00000000", 31615 => x"00000000", 31616 => x"00000000",
    31617 => x"00000000", 31618 => x"00000000", 31619 => x"00000000",
    31620 => x"00000000", 31621 => x"00000000", 31622 => x"00000000",
    31623 => x"00000000", 31624 => x"00000000", 31625 => x"00000000",
    31626 => x"00000000", 31627 => x"00000000", 31628 => x"00000000",
    31629 => x"00000000", 31630 => x"00000000", 31631 => x"00000000",
    31632 => x"00000000", 31633 => x"00000000", 31634 => x"00000000",
    31635 => x"00000000", 31636 => x"00000000", 31637 => x"00000000",
    31638 => x"00000000", 31639 => x"00000000", 31640 => x"00000000",
    31641 => x"00000000", 31642 => x"00000000", 31643 => x"00000000",
    31644 => x"00000000", 31645 => x"00000000", 31646 => x"00000000",
    31647 => x"00000000", 31648 => x"00000000", 31649 => x"00000000",
    31650 => x"00000000", 31651 => x"00000000", 31652 => x"00000000",
    31653 => x"00000000", 31654 => x"00000000", 31655 => x"00000000",
    31656 => x"00000000", 31657 => x"00000000", 31658 => x"00000000",
    31659 => x"00000000", 31660 => x"00000000", 31661 => x"00000000",
    31662 => x"00000000", 31663 => x"00000000", 31664 => x"00000000",
    31665 => x"00000000", 31666 => x"00000000", 31667 => x"00000000",
    31668 => x"00000000", 31669 => x"00000000", 31670 => x"00000000",
    31671 => x"00000000", 31672 => x"00000000", 31673 => x"00000000",
    31674 => x"00000000", 31675 => x"00000000", 31676 => x"00000000",
    31677 => x"00000000", 31678 => x"00000000", 31679 => x"00000000",
    31680 => x"00000000", 31681 => x"00000000", 31682 => x"00000000",
    31683 => x"00000000", 31684 => x"00000000", 31685 => x"00000000",
    31686 => x"00000000", 31687 => x"00000000", 31688 => x"00000000",
    31689 => x"00000000", 31690 => x"00000000", 31691 => x"00000000",
    31692 => x"00000000", 31693 => x"00000000", 31694 => x"00000000",
    31695 => x"00000000", 31696 => x"00000000", 31697 => x"00000000",
    31698 => x"00000000", 31699 => x"00000000", 31700 => x"00000000",
    31701 => x"00000000", 31702 => x"00000000", 31703 => x"00000000",
    31704 => x"00000000", 31705 => x"00000000", 31706 => x"00000000",
    31707 => x"00000000", 31708 => x"00000000", 31709 => x"00000000",
    31710 => x"00000000", 31711 => x"00000000", 31712 => x"00000000",
    31713 => x"00000000", 31714 => x"00000000", 31715 => x"00000000",
    31716 => x"00000000", 31717 => x"00000000", 31718 => x"00000000",
    31719 => x"00000000", 31720 => x"00000000", 31721 => x"00000000",
    31722 => x"00000000", 31723 => x"00000000", 31724 => x"00000000",
    31725 => x"00000000", 31726 => x"00000000", 31727 => x"00000000",
    31728 => x"00000000", 31729 => x"00000000", 31730 => x"00000000",
    31731 => x"00000000", 31732 => x"00000000", 31733 => x"00000000",
    31734 => x"00000000", 31735 => x"00000000", 31736 => x"00000000",
    31737 => x"00000000", 31738 => x"00000000", 31739 => x"00000000",
    31740 => x"00000000", 31741 => x"00000000", 31742 => x"00000000",
    31743 => x"00000000", 31744 => x"00000000", 31745 => x"00000000",
    31746 => x"00000000", 31747 => x"00000000", 31748 => x"00000000",
    31749 => x"00000000", 31750 => x"00000000", 31751 => x"00000000",
    31752 => x"00000000", 31753 => x"00000000", 31754 => x"00000000",
    31755 => x"00000000", 31756 => x"00000000", 31757 => x"00000000",
    31758 => x"00000000", 31759 => x"00000000", 31760 => x"00000000",
    31761 => x"00000000", 31762 => x"00000000", 31763 => x"00000000",
    31764 => x"00000000", 31765 => x"00000000", 31766 => x"00000000",
    31767 => x"00000000", 31768 => x"00000000", 31769 => x"00000000",
    31770 => x"00000000", 31771 => x"00000000", 31772 => x"00000000",
    31773 => x"00000000", 31774 => x"00000000", 31775 => x"00000000",
    31776 => x"00000000", 31777 => x"00000000", 31778 => x"00000000",
    31779 => x"00000000", 31780 => x"00000000", 31781 => x"00000000",
    31782 => x"00000000", 31783 => x"00000000", 31784 => x"00000000",
    31785 => x"00000000", 31786 => x"00000000", 31787 => x"00000000",
    31788 => x"00000000", 31789 => x"00000000", 31790 => x"00000000",
    31791 => x"00000000", 31792 => x"00000000", 31793 => x"00000000",
    31794 => x"00000000", 31795 => x"00000000", 31796 => x"00000000",
    31797 => x"00000000", 31798 => x"00000000", 31799 => x"00000000",
    31800 => x"00000000", 31801 => x"00000000", 31802 => x"00000000",
    31803 => x"00000000", 31804 => x"00000000", 31805 => x"00000000",
    31806 => x"00000000", 31807 => x"00000000", 31808 => x"00000000",
    31809 => x"00000000", 31810 => x"00000000", 31811 => x"00000000",
    31812 => x"00000000", 31813 => x"00000000", 31814 => x"00000000",
    31815 => x"00000000", 31816 => x"00000000", 31817 => x"00000000",
    31818 => x"00000000", 31819 => x"00000000", 31820 => x"00000000",
    31821 => x"00000000", 31822 => x"00000000", 31823 => x"00000000",
    31824 => x"00000000", 31825 => x"00000000", 31826 => x"00000000",
    31827 => x"00000000", 31828 => x"00000000", 31829 => x"00000000",
    31830 => x"00000000", 31831 => x"00000000", 31832 => x"00000000",
    31833 => x"00000000", 31834 => x"00000000", 31835 => x"00000000",
    31836 => x"00000000", 31837 => x"00000000", 31838 => x"00000000",
    31839 => x"00000000", 31840 => x"00000000", 31841 => x"00000000",
    31842 => x"00000000", 31843 => x"00000000", 31844 => x"00000000",
    31845 => x"00000000", 31846 => x"00000000", 31847 => x"00000000",
    31848 => x"00000000", 31849 => x"00000000", 31850 => x"00000000",
    31851 => x"00000000", 31852 => x"00000000", 31853 => x"00000000",
    31854 => x"00000000", 31855 => x"00000000", 31856 => x"00000000",
    31857 => x"00000000", 31858 => x"00000000", 31859 => x"00000000",
    31860 => x"00000000", 31861 => x"00000000", 31862 => x"00000000",
    31863 => x"00000000", 31864 => x"00000000", 31865 => x"00000000",
    31866 => x"00000000", 31867 => x"00000000", 31868 => x"00000000",
    31869 => x"00000000", 31870 => x"00000000", 31871 => x"00000000",
    31872 => x"00000000", 31873 => x"00000000", 31874 => x"00000000",
    31875 => x"00000000", 31876 => x"00000000", 31877 => x"00000000",
    31878 => x"00000000", 31879 => x"00000000", 31880 => x"00000000",
    31881 => x"00000000", 31882 => x"00000000", 31883 => x"00000000",
    31884 => x"00000000", 31885 => x"00000000", 31886 => x"00000000",
    31887 => x"00000000", 31888 => x"00000000", 31889 => x"00000000",
    31890 => x"00000000", 31891 => x"00000000", 31892 => x"00000000",
    31893 => x"00000000", 31894 => x"00000000", 31895 => x"00000000",
    31896 => x"00000000", 31897 => x"00000000", 31898 => x"00000000",
    31899 => x"00000000", 31900 => x"00000000", 31901 => x"00000000",
    31902 => x"00000000", 31903 => x"00000000", 31904 => x"00000000",
    31905 => x"00000000", 31906 => x"00000000", 31907 => x"00000000",
    31908 => x"00000000", 31909 => x"00000000", 31910 => x"00000000",
    31911 => x"00000000", 31912 => x"00000000", 31913 => x"00000000",
    31914 => x"00000000", 31915 => x"00000000", 31916 => x"00000000",
    31917 => x"00000000", 31918 => x"00000000", 31919 => x"00000000",
    31920 => x"00000000", 31921 => x"00000000", 31922 => x"00000000",
    31923 => x"00000000", 31924 => x"00000000", 31925 => x"00000000",
    31926 => x"00000000", 31927 => x"00000000", 31928 => x"00000000",
    31929 => x"00000000", 31930 => x"00000000", 31931 => x"00000000",
    31932 => x"00000000", 31933 => x"00000000", 31934 => x"00000000",
    31935 => x"00000000", 31936 => x"00000000", 31937 => x"00000000",
    31938 => x"00000000", 31939 => x"00000000", 31940 => x"00000000",
    31941 => x"00000000", 31942 => x"00000000", 31943 => x"00000000",
    31944 => x"00000000", 31945 => x"00000000", 31946 => x"00000000",
    31947 => x"00000000", 31948 => x"00000000", 31949 => x"00000000",
    31950 => x"00000000", 31951 => x"00000000", 31952 => x"00000000",
    31953 => x"00000000", 31954 => x"00000000", 31955 => x"00000000",
    31956 => x"00000000", 31957 => x"00000000", 31958 => x"00000000",
    31959 => x"00000000", 31960 => x"00000000", 31961 => x"00000000",
    31962 => x"00000000", 31963 => x"00000000", 31964 => x"00000000",
    31965 => x"00000000", 31966 => x"00000000", 31967 => x"00000000",
    31968 => x"00000000", 31969 => x"00000000", 31970 => x"00000000",
    31971 => x"00000000", 31972 => x"00000000", 31973 => x"00000000",
    31974 => x"00000000", 31975 => x"00000000", 31976 => x"00000000",
    31977 => x"00000000", 31978 => x"00000000", 31979 => x"00000000",
    31980 => x"00000000", 31981 => x"00000000", 31982 => x"00000000",
    31983 => x"00000000", 31984 => x"00000000", 31985 => x"00000000",
    31986 => x"00000000", 31987 => x"00000000", 31988 => x"00000000",
    31989 => x"00000000", 31990 => x"00000000", 31991 => x"00000000",
    31992 => x"00000000", 31993 => x"00000000", 31994 => x"00000000",
    31995 => x"00000000", 31996 => x"00000000", 31997 => x"00000000",
    31998 => x"00000000", 31999 => x"00000000", 32000 => x"00000000",
    32001 => x"00000000", 32002 => x"00000000", 32003 => x"00000000",
    32004 => x"00000000", 32005 => x"00000000", 32006 => x"00000000",
    32007 => x"00000000", 32008 => x"00000000", 32009 => x"00000000",
    32010 => x"00000000", 32011 => x"00000000", 32012 => x"00000000",
    32013 => x"00000000", 32014 => x"00000000", 32015 => x"00000000",
    32016 => x"00000000", 32017 => x"00000000", 32018 => x"00000000",
    32019 => x"00000000", 32020 => x"00000000", 32021 => x"00000000",
    32022 => x"00000000", 32023 => x"00000000", 32024 => x"00000000",
    32025 => x"00000000", 32026 => x"00000000", 32027 => x"00000000",
    32028 => x"00000000", 32029 => x"00000000", 32030 => x"00000000",
    32031 => x"00000000", 32032 => x"00000000", 32033 => x"00000000",
    32034 => x"00000000", 32035 => x"00000000", 32036 => x"00000000",
    32037 => x"00000000", 32038 => x"00000000", 32039 => x"00000000",
    32040 => x"00000000", 32041 => x"00000000", 32042 => x"00000000",
    32043 => x"00000000", 32044 => x"00000000", 32045 => x"00000000",
    32046 => x"00000000", 32047 => x"00000000", 32048 => x"00000000",
    32049 => x"00000000", 32050 => x"00000000", 32051 => x"00000000",
    32052 => x"00000000", 32053 => x"00000000", 32054 => x"00000000",
    32055 => x"00000000", 32056 => x"00000000", 32057 => x"00000000",
    32058 => x"00000000", 32059 => x"00000000", 32060 => x"00000000",
    32061 => x"00000000", 32062 => x"00000000", 32063 => x"00000000",
    32064 => x"00000000", 32065 => x"00000000", 32066 => x"00000000",
    32067 => x"00000000", 32068 => x"00000000", 32069 => x"00000000",
    32070 => x"00000000", 32071 => x"00000000", 32072 => x"00000000",
    32073 => x"00000000", 32074 => x"00000000", 32075 => x"00000000",
    32076 => x"00000000", 32077 => x"00000000", 32078 => x"00000000",
    32079 => x"00000000", 32080 => x"00000000", 32081 => x"00000000",
    32082 => x"00000000", 32083 => x"00000000", 32084 => x"00000000",
    32085 => x"00000000", 32086 => x"00000000", 32087 => x"00000000",
    32088 => x"00000000", 32089 => x"00000000", 32090 => x"00000000",
    32091 => x"00000000", 32092 => x"00000000", 32093 => x"00000000",
    32094 => x"00000000", 32095 => x"00000000", 32096 => x"00000000",
    32097 => x"00000000", 32098 => x"00000000", 32099 => x"00000000",
    32100 => x"00000000", 32101 => x"00000000", 32102 => x"00000000",
    32103 => x"00000000", 32104 => x"00000000", 32105 => x"00000000",
    32106 => x"00000000", 32107 => x"00000000", 32108 => x"00000000",
    32109 => x"00000000", 32110 => x"00000000", 32111 => x"00000000",
    32112 => x"00000000", 32113 => x"00000000", 32114 => x"00000000",
    32115 => x"00000000", 32116 => x"00000000", 32117 => x"00000000",
    32118 => x"00000000", 32119 => x"00000000", 32120 => x"00000000",
    32121 => x"00000000", 32122 => x"00000000", 32123 => x"00000000",
    32124 => x"00000000", 32125 => x"00000000", 32126 => x"00000000",
    32127 => x"00000000", 32128 => x"00000000", 32129 => x"00000000",
    32130 => x"00000000", 32131 => x"00000000", 32132 => x"00000000",
    32133 => x"00000000", 32134 => x"00000000", 32135 => x"00000000",
    32136 => x"00000000", 32137 => x"00000000", 32138 => x"00000000",
    32139 => x"00000000", 32140 => x"00000000", 32141 => x"00000000",
    32142 => x"00000000", 32143 => x"00000000", 32144 => x"00000000",
    32145 => x"00000000", 32146 => x"00000000", 32147 => x"00000000",
    32148 => x"00000000", 32149 => x"00000000", 32150 => x"00000000",
    32151 => x"00000000", 32152 => x"00000000", 32153 => x"00000000",
    32154 => x"00000000", 32155 => x"00000000", 32156 => x"00000000",
    32157 => x"00000000", 32158 => x"00000000", 32159 => x"00000000",
    32160 => x"00000000", 32161 => x"00000000", 32162 => x"00000000",
    32163 => x"00000000", 32164 => x"00000000", 32165 => x"00000000",
    32166 => x"00000000", 32167 => x"00000000", 32168 => x"00000000",
    32169 => x"00000000", 32170 => x"00000000", 32171 => x"00000000",
    32172 => x"00000000", 32173 => x"00000000", 32174 => x"00000000",
    32175 => x"00000000", 32176 => x"00000000", 32177 => x"00000000",
    32178 => x"00000000", 32179 => x"00000000", 32180 => x"00000000",
    32181 => x"00000000", 32182 => x"00000000", 32183 => x"00000000",
    32184 => x"00000000", 32185 => x"00000000", 32186 => x"00000000",
    32187 => x"00000000", 32188 => x"00000000", 32189 => x"00000000",
    32190 => x"00000000", 32191 => x"00000000", 32192 => x"00000000",
    32193 => x"00000000", 32194 => x"00000000", 32195 => x"00000000",
    32196 => x"00000000", 32197 => x"00000000", 32198 => x"00000000",
    32199 => x"00000000", 32200 => x"00000000", 32201 => x"00000000",
    32202 => x"00000000", 32203 => x"00000000", 32204 => x"00000000",
    32205 => x"00000000", 32206 => x"00000000", 32207 => x"00000000",
    32208 => x"00000000", 32209 => x"00000000", 32210 => x"00000000",
    32211 => x"00000000", 32212 => x"00000000", 32213 => x"00000000",
    32214 => x"00000000", 32215 => x"00000000", 32216 => x"00000000",
    32217 => x"00000000", 32218 => x"00000000", 32219 => x"00000000",
    32220 => x"00000000", 32221 => x"00000000", 32222 => x"00000000",
    32223 => x"00000000", 32224 => x"00000000", 32225 => x"00000000",
    32226 => x"00000000", 32227 => x"00000000", 32228 => x"00000000",
    32229 => x"00000000", 32230 => x"00000000", 32231 => x"00000000",
    32232 => x"00000000", 32233 => x"00000000", 32234 => x"00000000",
    32235 => x"00000000", 32236 => x"00000000", 32237 => x"00000000",
    32238 => x"00000000", 32239 => x"00000000", 32240 => x"00000000",
    32241 => x"00000000", 32242 => x"00000000", 32243 => x"00000000",
    32244 => x"00000000", 32245 => x"00000000", 32246 => x"00000000",
    32247 => x"00000000", 32248 => x"00000000", 32249 => x"00000000",
    32250 => x"00000000", 32251 => x"00000000", 32252 => x"00000000",
    32253 => x"00000000", 32254 => x"00000000", 32255 => x"00000000",
    32256 => x"00000000", 32257 => x"00000000", 32258 => x"00000000",
    32259 => x"00000000", 32260 => x"00000000", 32261 => x"00000000",
    32262 => x"00000000", 32263 => x"00000000", 32264 => x"00000000",
    32265 => x"00000000", 32266 => x"00000000", 32267 => x"00000000",
    32268 => x"00000000", 32269 => x"00000000", 32270 => x"00000000",
    32271 => x"00000000", 32272 => x"00000000", 32273 => x"00000000",
    32274 => x"00000000", 32275 => x"00000000", 32276 => x"00000000",
    32277 => x"00000000", 32278 => x"00000000", 32279 => x"00000000",
    32280 => x"00000000", 32281 => x"00000000", 32282 => x"00000000",
    32283 => x"00000000", 32284 => x"00000000", 32285 => x"00000000",
    32286 => x"00000000", 32287 => x"00000000", 32288 => x"00000000",
    32289 => x"00000000", 32290 => x"00000000", 32291 => x"00000000",
    32292 => x"00000000", 32293 => x"00000000", 32294 => x"00000000",
    32295 => x"00000000", 32296 => x"00000000", 32297 => x"00000000",
    32298 => x"00000000", 32299 => x"00000000", 32300 => x"00000000",
    32301 => x"00000000", 32302 => x"00000000", 32303 => x"00000000",
    32304 => x"00000000", 32305 => x"00000000", 32306 => x"00000000",
    32307 => x"00000000", 32308 => x"00000000", 32309 => x"00000000",
    32310 => x"00000000", 32311 => x"00000000", 32312 => x"00000000",
    32313 => x"00000000", 32314 => x"00000000", 32315 => x"00000000",
    32316 => x"00000000", 32317 => x"00000000", 32318 => x"00000000",
    32319 => x"00000000", 32320 => x"00000000", 32321 => x"00000000",
    32322 => x"00000000", 32323 => x"00000000", 32324 => x"00000000",
    32325 => x"00000000", 32326 => x"00000000", 32327 => x"00000000",
    32328 => x"00000000", 32329 => x"00000000", 32330 => x"00000000",
    32331 => x"00000000", 32332 => x"00000000", 32333 => x"00000000",
    32334 => x"00000000", 32335 => x"00000000", 32336 => x"00000000",
    32337 => x"00000000", 32338 => x"00000000", 32339 => x"00000000",
    32340 => x"00000000", 32341 => x"00000000", 32342 => x"00000000",
    32343 => x"00000000", 32344 => x"00000000", 32345 => x"00000000",
    32346 => x"00000000", 32347 => x"00000000", 32348 => x"00000000",
    32349 => x"00000000", 32350 => x"00000000", 32351 => x"00000000",
    32352 => x"00000000", 32353 => x"00000000", 32354 => x"00000000",
    32355 => x"00000000", 32356 => x"00000000", 32357 => x"00000000",
    32358 => x"00000000", 32359 => x"00000000", 32360 => x"00000000",
    32361 => x"00000000", 32362 => x"00000000", 32363 => x"00000000",
    32364 => x"00000000", 32365 => x"00000000", 32366 => x"00000000",
    32367 => x"00000000", 32368 => x"00000000", 32369 => x"00000000",
    32370 => x"00000000", 32371 => x"00000000", 32372 => x"00000000",
    32373 => x"00000000", 32374 => x"00000000", 32375 => x"00000000",
    32376 => x"00000000", 32377 => x"00000000", 32378 => x"00000000",
    32379 => x"00000000", 32380 => x"00000000", 32381 => x"00000000",
    32382 => x"00000000", 32383 => x"00000000", 32384 => x"00000000",
    32385 => x"00000000", 32386 => x"00000000", 32387 => x"00000000",
    32388 => x"00000000", 32389 => x"00000000", 32390 => x"00000000",
    32391 => x"00000000", 32392 => x"00000000", 32393 => x"00000000",
    32394 => x"00000000", 32395 => x"00000000", 32396 => x"00000000",
    32397 => x"00000000", 32398 => x"00000000", 32399 => x"00000000",
    32400 => x"00000000", 32401 => x"00000000", 32402 => x"00000000",
    32403 => x"00000000", 32404 => x"00000000", 32405 => x"00000000",
    32406 => x"00000000", 32407 => x"00000000", 32408 => x"00000000",
    32409 => x"00000000", 32410 => x"00000000", 32411 => x"00000000",
    32412 => x"00000000", 32413 => x"00000000", 32414 => x"00000000",
    32415 => x"00000000", 32416 => x"00000000", 32417 => x"00000000",
    32418 => x"00000000", 32419 => x"00000000", 32420 => x"00000000",
    32421 => x"00000000", 32422 => x"00000000", 32423 => x"00000000",
    32424 => x"00000000", 32425 => x"00000000", 32426 => x"00000000",
    32427 => x"00000000", 32428 => x"00000000", 32429 => x"00000000",
    32430 => x"00000000", 32431 => x"00000000", 32432 => x"00000000",
    32433 => x"00000000", 32434 => x"00000000", 32435 => x"00000000",
    32436 => x"00000000", 32437 => x"00000000", 32438 => x"00000000",
    32439 => x"00000000", 32440 => x"00000000", 32441 => x"00000000",
    32442 => x"00000000", 32443 => x"00000000", 32444 => x"00000000",
    32445 => x"00000000", 32446 => x"00000000", 32447 => x"00000000",
    32448 => x"00000000", 32449 => x"00000000", 32450 => x"00000000",
    32451 => x"00000000", 32452 => x"00000000", 32453 => x"00000000",
    32454 => x"00000000", 32455 => x"00000000", 32456 => x"00000000",
    32457 => x"00000000", 32458 => x"00000000", 32459 => x"00000000",
    32460 => x"00000000", 32461 => x"00000000", 32462 => x"00000000",
    32463 => x"00000000", 32464 => x"00000000", 32465 => x"00000000",
    32466 => x"00000000", 32467 => x"00000000", 32468 => x"00000000",
    32469 => x"00000000", 32470 => x"00000000", 32471 => x"00000000",
    32472 => x"00000000", 32473 => x"00000000", 32474 => x"00000000",
    32475 => x"00000000", 32476 => x"00000000", 32477 => x"00000000",
    32478 => x"00000000", 32479 => x"00000000", 32480 => x"00000000",
    32481 => x"00000000", 32482 => x"00000000", 32483 => x"00000000",
    32484 => x"00000000", 32485 => x"00000000", 32486 => x"00000000",
    32487 => x"00000000", 32488 => x"00000000", 32489 => x"00000000",
    32490 => x"00000000", 32491 => x"00000000", 32492 => x"00000000",
    32493 => x"00000000", 32494 => x"00000000", 32495 => x"00000000",
    32496 => x"00000000", 32497 => x"00000000", 32498 => x"00000000",
    32499 => x"00000000", 32500 => x"00000000", 32501 => x"00000000",
    32502 => x"00000000", 32503 => x"00000000", 32504 => x"00000000",
    32505 => x"00000000", 32506 => x"00000000", 32507 => x"00000000",
    32508 => x"00000000", 32509 => x"00000000", 32510 => x"00000000",
    32511 => x"00000000", 32512 => x"00000000", 32513 => x"00000000",
    32514 => x"00000000", 32515 => x"00000000", 32516 => x"00000000",
    32517 => x"00000000", 32518 => x"00000000", 32519 => x"00000000",
    32520 => x"00000000", 32521 => x"00000000", 32522 => x"00000000",
    32523 => x"00000000", 32524 => x"00000000", 32525 => x"00000000",
    32526 => x"00000000", 32527 => x"00000000", 32528 => x"00000000",
    32529 => x"00000000", 32530 => x"00000000", 32531 => x"00000000",
    32532 => x"00000000", 32533 => x"00000000", 32534 => x"00000000",
    32535 => x"00000000", 32536 => x"00000000", 32537 => x"00000000",
    32538 => x"00000000", 32539 => x"00000000", 32540 => x"00000000",
    32541 => x"00000000", 32542 => x"00000000", 32543 => x"00000000",
    32544 => x"00000000", 32545 => x"00000000", 32546 => x"00000000",
    32547 => x"00000000", 32548 => x"00000000", 32549 => x"00000000",
    32550 => x"00000000", 32551 => x"00000000", 32552 => x"00000000",
    32553 => x"00000000", 32554 => x"00000000", 32555 => x"00000000",
    32556 => x"00000000", 32557 => x"00000000", 32558 => x"00000000",
    32559 => x"00000000", 32560 => x"00000000", 32561 => x"00000000",
    32562 => x"00000000", 32563 => x"00000000", 32564 => x"00000000",
    32565 => x"00000000", 32566 => x"00000000", 32567 => x"00000000",
    32568 => x"00000000", 32569 => x"00000000", 32570 => x"00000000",
    32571 => x"00000000", 32572 => x"00000000", 32573 => x"00000000",
    32574 => x"00000000", 32575 => x"00000000", 32576 => x"00000000",
    32577 => x"00000000", 32578 => x"00000000", 32579 => x"00000000",
    32580 => x"00000000", 32581 => x"00000000", 32582 => x"00000000",
    32583 => x"00000000", 32584 => x"00000000", 32585 => x"00000000",
    32586 => x"00000000", 32587 => x"00000000", 32588 => x"00000000",
    32589 => x"00000000", 32590 => x"00000000", 32591 => x"00000000",
    32592 => x"00000000", 32593 => x"00000000", 32594 => x"00000000",
    32595 => x"00000000", 32596 => x"00000000", 32597 => x"00000000",
    32598 => x"00000000", 32599 => x"00000000", 32600 => x"00000000",
    32601 => x"00000000", 32602 => x"00000000", 32603 => x"00000000",
    32604 => x"00000000", 32605 => x"00000000", 32606 => x"00000000",
    32607 => x"00000000", 32608 => x"00000000", 32609 => x"00000000",
    32610 => x"00000000", 32611 => x"00000000", 32612 => x"00000000",
    32613 => x"00000000", 32614 => x"00000000", 32615 => x"00000000",
    32616 => x"00000000", 32617 => x"00000000", 32618 => x"00000000",
    32619 => x"00000000", 32620 => x"00000000", 32621 => x"00000000",
    32622 => x"00000000", 32623 => x"00000000", 32624 => x"00000000",
    32625 => x"00000000", 32626 => x"00000000", 32627 => x"00000000",
    32628 => x"00000000", 32629 => x"00000000", 32630 => x"00000000",
    32631 => x"00000000", 32632 => x"00000000", 32633 => x"00000000",
    32634 => x"00000000", 32635 => x"00000000", 32636 => x"00000000",
    32637 => x"00000000", 32638 => x"00000000", 32639 => x"00000000",
    32640 => x"00000000", 32641 => x"00000000", 32642 => x"00000000",
    32643 => x"00000000", 32644 => x"00000000", 32645 => x"00000000",
    32646 => x"00000000", 32647 => x"00000000", 32648 => x"00000000",
    32649 => x"00000000", 32650 => x"00000000", 32651 => x"00000000",
    32652 => x"00000000", 32653 => x"00000000", 32654 => x"00000000",
    32655 => x"00000000", 32656 => x"00000000", 32657 => x"00000000",
    32658 => x"00000000", 32659 => x"00000000", 32660 => x"00000000",
    32661 => x"00000000", 32662 => x"00000000", 32663 => x"00000000",
    32664 => x"00000000", 32665 => x"00000000", 32666 => x"00000000",
    32667 => x"00000000", 32668 => x"00000000", 32669 => x"00000000",
    32670 => x"00000000", 32671 => x"00000000", 32672 => x"00000000",
    32673 => x"00000000", 32674 => x"00000000", 32675 => x"00000000",
    32676 => x"00000000", 32677 => x"00000000", 32678 => x"00000000",
    32679 => x"00000000", 32680 => x"00000000", 32681 => x"00000000",
    32682 => x"00000000", 32683 => x"00000000", 32684 => x"00000000",
    32685 => x"00000000", 32686 => x"00000000", 32687 => x"00000000",
    32688 => x"00000000", 32689 => x"00000000", 32690 => x"00000000",
    32691 => x"00000000", 32692 => x"00000000", 32693 => x"00000000",
    32694 => x"00000000", 32695 => x"00000000", 32696 => x"00000000",
    32697 => x"00000000", 32698 => x"00000000", 32699 => x"00000000",
    32700 => x"00000000", 32701 => x"00000000", 32702 => x"00000000",
    32703 => x"00000000", 32704 => x"00000000", 32705 => x"00000000",
    32706 => x"00000000", 32707 => x"00000000", 32708 => x"00000000",
    32709 => x"00000000", 32710 => x"00000000", 32711 => x"00000000",
    32712 => x"00000000", 32713 => x"00000000", 32714 => x"00000000",
    32715 => x"00000000", 32716 => x"00000000", 32717 => x"00000000",
    32718 => x"00000000", 32719 => x"00000000", 32720 => x"00000000",
    32721 => x"00000000", 32722 => x"00000000", 32723 => x"00000000",
    32724 => x"00000000", 32725 => x"00000000", 32726 => x"00000000",
    32727 => x"00000000", 32728 => x"00000000", 32729 => x"00000000",
    32730 => x"00000000", 32731 => x"00000000", 32732 => x"00000000",
    32733 => x"00000000", 32734 => x"00000000", 32735 => x"00000000",
    32736 => x"00000000", 32737 => x"00000000", 32738 => x"00000000",
    32739 => x"00000000", 32740 => x"00000000", 32741 => x"00000000",
    32742 => x"00000000", 32743 => x"00000000", 32744 => x"00000000",
    32745 => x"00000000", 32746 => x"00000000", 32747 => x"00000000",
    32748 => x"00000000", 32749 => x"00000000", 32750 => x"00000000",
    32751 => x"00000000", 32752 => x"00000000", 32753 => x"00000000",
    32754 => x"00000000", 32755 => x"00000000", 32756 => x"00000000",
    32757 => x"00000000", 32758 => x"00000000", 32759 => x"00000000",
    32760 => x"00000000", 32761 => x"00000000", 32762 => x"00000000",
    32763 => x"00000000", 32764 => x"00000000", 32765 => x"00000000",
    32766 => x"00000000", 32767 => x"00000000");
end wrc_bin_pkg;

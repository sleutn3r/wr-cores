// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GYfyPCsTIevWVcG/9uvLesBOJFW2+Z93BCflHuzDPi7pqPDZNP8vBrcG8sst3cYg
CY8IztIQPRfos+uMTwUjoE+rydwFHmdXvhp4Nu3KYWsWn+VVgcOcJw2FAvG6qniL
IDxKbEMndDw4GShlFBwAczCQngc3p7vUwsX4QsWXRJk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12176)
ftBW5ztfskNqEBHnoxOCYC8neoQC6rQMb7wzGvxtjh5uhQouaMqcgbDA5R+OcpuZ
moC7btfZ23k/MKIJYhN/3jQxtey9kRyCCi2rORhYEeXisUWY57uiJVs4wzvuhG9t
FjkDRw+CNKPwqooIaOxSEue14bC7x7XqDxjJ4hF7I8ivvFA1pKiWA6IU+PQlgr87
or9ALqn8T+9RmsEVpog+DD3y+8a+EmMVveaaeaBXvLjZMyIFS9Sj2ur232zQWFcq
ie8YGi1Zm5en1yRl8yC6XqeYYNmAFasZBf+6c3dRwBR9pD8ZeT8/M73MuHOfl2/5
EHGHft5+npce6nCAEKjOCKQ6Ev4mIBi+3ECGAVEZoXxrAacshPxJsFhwb9I7RUe7
I75KHamvygd16EpfOpydcS2KSgOWGJl5yohZCtgfgQ5kd26zj0LCaIxj7KbzmOSB
OGZ/cMtmzb7PeOglWUKer7FU4jr3vmIwUFFzE3ALhG/udbV5k3teyeFVmRMe6ajf
RXse2m2ogy1cjdoiamteIrlbhWP5apFTjdYUOEk92lygksm8M0As4Bqh27P9gyh8
rqens3YKNDBNmLZknqgnq0Q4L0xl7kItPce1H81lh58ERTjtCOl1vRphhuet8klD
dGKutF70aNlLq2Cwr7FQDqvRvJD/wMQQikjhLvBW6xqecZYywFNnpKe9awgYM6Fl
IUcbaAMmHzUMaZ+mgmw+dG6qALAJj5so1/w26YHkuHU0/oNoTLEWijCpPEfgXoAg
L93+HWDeyEWZ6J+S2N0kaR7Lne/cOIIhqjDqufG/gxVfHQ8iN8fBLNN11VkPSxbQ
crHtB881F6xSg0hVYNCFE/cBB6ZkC1W5fLo/oO7uhIT08M8YbVIqbG/1+UveVn5J
2G1ZRmLgN6OXgHC1scvrWflw5VAfYStLrdVo0776uW82wY7cVvHb6sqSQS8JTXAU
dCHw7tthfkc5zaMXt5ScPbKszmXoNvKfTFivBET6VzWPN+DXVJBNo1wLeyf821wB
VqcfwgATCB0IQp1pnbS4bd/5Y/ZtHOoTjDnRM/wzpjK7Bh3ZP9CC/fRS1hu0E22V
67XubZ02BqBKJLWNdOZ+G7NsqN6rlSDMAThj/75nkrpOmPeBsetcIfPbOt7V360E
C2i34xeyMAA8HMSL1W7RPxqjM89Sm480UEVBRgDrUXFf5+gYGIO6TnS2oJn1alp7
Xyg0TeAPhAylWMTtQiRcMyeYy80opIDL0zRpMyo2VBhvvImdhD9a3mK9ZCFFlk2d
Vbpxfnbf4DZXIVLIdmcNL009/eA6bbCcvte+DypmDG74YeeLWZ0lrdAoUxMzUf5u
BO7de9nK90UTFj5tc7HXIEaQkOUNIEJopDjDTZNs3STDlJaS+/EOiw+P+F2lp0+P
SBaGCTQRYtT58g26nectTTg8FItNreXOhklblZMn2wat3eeTJq43vv2s/opADm7N
p3DH6SCNuGtSdyrycetF68aGY1nwvopzmWLi6EbXyT22IobaxqPhHXQc234jqA0L
eN7GtCkJOPpEvs+proS9z/DaY4mqMXINgwzCZt+HP6Tp6xcZXyhI2+SZliAnlDAV
aBoBlIJkEPeNUGlkYp4L0r8zRHnrWHahWfdTb9qzI5iskGPc3FwCiZchVbfkorc+
vxNehGQDEkKpY4/BNP4sKc3M9VjuMYilkHB4iJdzb3sz0qCAbVn18jwyIySnc+j6
YhZA5wXpGuqc3v1FdGk4zSpIbm2BaRMqKyPjUcM5FJ/lKGFmepfU/Qqe6MBp+tq+
3rATN489mgZ6ZIMLkMkFYbMrjuLuXcIr6vickrqw2ZQXQJ34/KiMejnNJclTdB/s
pa5/Y8z+cE3FhMSCnvzkCn5NTNO11gHncJgRV5fyzACk9eIvw4ToZ66uGfQXh3gS
aZq1BZzKkeK3ZHmvaKrScg6pwblt6TjhxUqwG4lwXXPWvL/25zlNiJ3iUBJDvQHp
/zneQ7Ri0Mfimqv8w19HqVT2YFi+54HlrJJf6L3KdngLg4084EWW6iM+5ud7lvZM
+mgsxbFAWqtMv0+CBx9+sVJh7N8TGBPC/bumPXwWATBQjZxh8og9vfSu0P5hH6SQ
byxKZyJy8062A5LPoEDon8xEkTWEG/MlM0W2bvgDYOfBQbd3ev7DtjnsdjzTTotv
2rqTgw7aJZoLiFk6VTHMHLXVuiipiVlsWroHjfuqqo7fT+yEBSck/3piRVYpbo7m
L2MTkBsMCi+M8zcS3AraLcqmsGJLifH8ki55/K3vP1+M9Gn97D0JWVAH3l2B/Pip
MfoDUjfRx3ahDc6QPBQN7IpdKtGUJDNKi3k0Nof+Wd7XtFDx80hUne5CknsnSvgU
zdWURmptHxL1Rg/3fjtEgEttcji3lzPvgKJebZLKhMh/POAaCcjoUPOLMF+StQDc
3Xjbvefnr9EecZhoASTexQPFVaneEoIRxfBku9IYYPcChQPaevt9eJlMcZGv7hvf
6cv9ZURyevMIMw0bbpreEyknVrmBnOuJu2vZHeig99Y79+1skI/E99USU3U1KNWB
S4NXQusV+dbkJmPsK6sHjUKU7XSMj0aY5ekh4ctSVDkQDk4EnbVhhIXyh7gxVKAG
rUeWyXNi2kYQ70lEqo2ZZdOJuezsGNkijvtJIWmZZZcZMrooVMXfRLdNf2r7Yvb9
4rlBx+UEEnzGFGiGH79OPQ6g3RWvs/j7P9kY3pyq8x2AmbzLZvi3PZbZdlO8T7ZM
/pbJkHB+keXAm+aGaJOoJM757OSfAhgwVx13UebcmkTA4z87t43zMhElo1lrwNl+
CSp7gxJm/41mXXWnfotLl7qs80xxpKnCbpzMS7R67zhrXSwiT+PdubYHx4qir1mo
MzGuFmRJC/anU3wyRW82JFKWRErNN0MThLunlV16m+i3LH5Y0CyoYdt69fuaqAbS
A331wLGWLQ+9c+k1jtAMy5y/2WFgtbNnw0jBDIH8wDqcnL59xpqU58rvCQSTqyl2
s0hVDJfcZWTdn1doiCK2Wku2RbDFt4lux6oo2vYwmZPyBiXlDkq07SZ9kM6aOoG5
1zDm1ZYxQoJHN4Xorc6APW/zcYwOGx13+ufHfHfgyetqCqbx1bzzoDyH8OfkyB+6
WjJHREgl87xv8piEPg0M2v3lWosNx6hQ4Hhnd7f0GO6+hbF0/mvMyq0bSNtxc+Hl
aG5AdfIbPKoq+QCQj2y3ogbKWdS/JSSa1ufOlhDaovd/TSKWNoI9ZTFuSexBKc2k
DOuBOXr9nKD7NIeuj1IpCebYbunQ4vJZ2i3rPz1BOJ4Y1ZhqGrZxWQKFjUz0wfpB
aSSh+G4tNj2KgRj6TuoNBoXrWtfKYMrykPqYyA1V7q5nm+1F9EcReKeOmUuL6tih
UIGHsv+Imv7cNiPpsYCbya7gLT5H15o6wbi5dVvBn9gYnrdmQyKEb0/ZQUGdEvbb
RpQ1Xw7sRfcIXVPeAKVxbwaSvPwQUONnSwtnYoUJOYerQQAMg5lWpvtUMN6JhiY9
ZQMhi8/jBJv7bOHOeaARcPj/2atcF94RPEgcEhfG3PXKxFY8FxaUvzeLQS4etOVg
bawWP4JZDWOPrYKU1tjg1Cbu/nfGSgshKMFfuHHNca92+e6B7OuiNWXW1kqKXlhU
zMTn+TVFTQkruvB4nS7P+XPK1wVmobj0lLFRLnwLq6uPVBnpfGy8gSb0Uu3cgiFp
VBqXJqTAo29Q+ZR4UctvM50IIOXdjh4/rGfpbDBLkoBpuYYb2eViQPoxViEbGHRn
S1rqBCs2c2b08kIlEHwR++FrljjkOsgsi4rxrtBPFeDK92RURiyp+ZDFrKclEi7y
yfIuhsZ1TrdbdgTBAo+b0xiWVhH6pFFHVAhsoHfxS4QSTLz0x5RsNKG4yTRRrM6H
5elyjwifmO29s0AvH7Pf8I3Cq/qt/vchZT5gUKS31gDk2FjMX52Gdghuq5HYlIyE
9O2BFPhiaQudQzyMoKpEnCedwJ0WppCL47lqGw1mo7eMVKq/yEiP+MEPv+rspikb
MsuP8RFnP9fuodtT+mHkicXjKBIATyLBiH1qYEUdeSZWNt3zWfOc6ZpJSv81hdSz
oY1DtVQvDoZLk1YYLgVTFZs9GAByIAGSEldbM9ThTBiNPdL6CBXE4kRZpMjjxfgb
nxTUEZdvDNuZ5cRK1ZDFAtSkdzBtoaolC7BQRnz9yhoEybXpcjOTNFEx60gDq/Cr
3uVXiOCzUO/tHN4qmjEAcXL3tA0q9ooAmsQfCcX1ZYBY2nvE5/2O91kjFeit+c2U
LHlCBnXe6fFAhSi4w9/o2YdHXz/N6jN0DTY2T12qmOS4C1+dVeRrDJI7L6ATbqJa
BrRr8ZJfcj1aHpTlrLLMfkmHOtu/Cfe0dfN5IlxuEaYvH8Y6M9GIiNlvbcHHpkyU
jAcT9ezn1paF3gMn+XXEIbv73nf+qWjKoouLz15hGTmtD6sDcCsl0USGyG90LLO4
0wici/FkvfsmPybZxeBaS2W7kAHJPkEiDf4BRkJsmL9AJ6B5S8e853kAJ8oN9UxS
+WhQ7zKPvD5bQXck+UrHUgLV/rYXnvO4zTGKp6AdOmg+xse0PbwZfODa2gRkJHHy
LErgSs/VaZzS5R+uRDxqPpa7Jkt/JaV0c8SBYOwRZ8fYySz2V/M4h0+u+Gplxl0Q
5Trs3i39YnNCNefE91kfBy28fi3GDvAb9StwrZdaPCqoTTVqn+x6mxilthmzeSwD
yA2o0DUPJtpS5yBf7hQ0OajACotwCKEqiuQrTp7sHYmJPl8Cmd+4OdztduuRtsiu
UzaKH86VEQy4hlroixmKLk+aHXa9iiH57CFdMvuR7HQ5hbsmyH9yCuY723eNBXU2
olr1FqN6m5Tl0tFJ0t6EeFQf0txlEOW9hfaPJRPjXkGrivVAWjQuhBWabBoB28pz
PJf42MmBb42RkhMnbc0Qrgq+Dq6lbGZNBV9gWic9MgF6eKe/26tmsa6lOvEC1hWL
N/1LziaX4foTJnD6ke8aA0q+Uwlm6eZhBODZ1uipMp/19QmlIeUyjj6m6ASGyq9j
QZYcctLKQgg8PkjMpHYIX7zxmKRRBQzPAZawXXbsvGm+dVg4Hd+tefjel3ffQKB0
GSCUpI3uKafi+9CNpedAOSZ0iHJkFNf1CokQBlvBJHVVI+Ey5AWrj38nbjAyaj6l
iCsjmkkK2quUl+ZBQ46eAE4sK3KMhZvkbAJHoP83VKfRWo4uRAPOI3dTO4721Jww
Owb8yXajBn5bzVQ6QBOWX16my49IDhKrMfYkG3spJ7rbB4gCvbPRsITYHKnwPr0T
KhpRMQmOiISbzoE4VsNC51frxjTsGcimD2mCC6+mT8IS2OgVFCjl3WYQWp9/v6SD
CqZE3/M34qRV6VxtyQrORb7Lg9V1My92GBDzgiv1qIh2t3CdLshgHdcdJRLUNrdL
/q8cwmV8efKNKvCHomND8uOLNKa5yfYd7rHV0LQnwj05ALKb/4C+qj2XM6P6mZhO
oEJPeGNtBnx4PcXS9qmb0H6oNWAyeKAyQKWfN0CVXoaFUsdxDpvqagknIwp5VHNt
zQT/nEXxn5+1vx6Q3mSDQBHdAstVvkN8FoKiPDVFG3D3VWQhL/cjtDWVwjGWcXRq
jINcbITS3/DuUgq3NMxNVqvOyFGH+jxSd2oePXNwaFjOjcI/GypihpSM9ZA5y/ug
0cKNVoLa1/wNKxdT7YQ3lhA74J86dcg0mwjwxjV1ZnK383vB7Ktd7Bx+fA4RsAX2
ig5otVnIXJ+5ieBZyeNwRV+5sl7rFpU7GrlW1E+sVCsTXMNNghcfSU+xOigxoi6s
GoePAvTF1ltgDDC74r2ZJG6WS5qywY03zImNHnW+G7LdkezEGys2oK2FyC3Ln/9s
Mpj5KJI8RU6jIPNLJRBBcorxXu6jW5NBEnxhRZadzmOY0AQCIGH2C0y+SiY5nvdd
kvsaI7d/S7VyVZwez/CjPNAVu/x/nznzUpblBR0r8V5tzw211BoE/S2NiICpVZG2
OKrk7LMSKjPz7MuR0DcoAai7xyG0u4ueAdKFb5Pe4iey+KSKmAMve6zEAjc8Ugvq
z8GrI7hvZ6KoXw3VgMSoBSdEsyqL/2deomLrCMd/2MoN/CfaV3S4qd3iz4bjt8qq
NSDUD/D+WTcQbUMdzQra4esAJcFKezfrvOsvb6RXntCheyEgC+70+Xxtf+0PXWAv
b0FD93WpZwNZZ6Mp04cIH/tgXqaq0G3+qbm5zgqrKjWs3xpI86tZVohoQ+quAx7+
SPq2zTOHUlrvLUK9VBT4LBFTmJgVVKzDyqH+5A4/YDoHe+nXGVlJFaSSLWzK6kLh
PlZs0SC36rf8h132MvS8JE9/Byqxauljs8uBYF/v9+A79LnjfBWuYFD00FS9Nemy
Ucrs61sXjUPU1MMSJBMizelfqmVy7voKStcBaihruaghyDM3xBB6+yF8h+tyeNwu
zDv3Xaw70OGU083y0uBjEfTFTS9OgBFJKrm3nWft3qAed9nGuB5FxHzbdoaIGVF0
lZB2LfUtBxdEqzTSSovwUR6gZp+c3+w5qwxnwtBXr4z+/HiTmBdytz6DufF6NAQw
QTwOiyNKdHYneTXmTPgKtYG6gRPsVk/tMwQU2+oT9wNmI6dlCkWu+78KzovgkjVO
/sM+bImfWwlwpQu1LC8Q6Yx+9SPzh9jVkukrWrXybP/waRpJPDgfHNvE+258LF+U
8v7ljtpsacuQjRjAVGnlUVlwUHf63qEduPN10C1J7gKznU5BfwWWu00MO4+Ix3ZA
X9RHFlwjWycwYzWhqK8OzJNjqWmvOxo+4PqQtEZ9TlWvNNDrOxOVW/qEHv/xduoV
cRYv4An6Nmm9UcVdh2u7tOx5uTTZSWpXPqv+YfT8qSW2ZqA8kWei0cKdSF8v3yVB
MU6yEnQ1I90MTQ6huqIE2dYKe5qqL9Yd8csqgCey1/EoJSLpj8kKzKtuinRy00RE
TWwYTHs1hy7SX4NUMhxzZ+jOQ93lcft79tPuEGemyvbZUKbf9wPieAHdLUPzwGIC
F7Qqfusiq5j4Aw/R0s0viUb2gHStwOT4RdLnm7nnQ6NhLsA9cLPM+zCC1niktHqu
PVYsnRPRVXiHHbgnMcc/2q/yCLrk4nfuVqSzBlqQqOF/ANVRtV4ItvljEdNNlBZk
ckGBthIGJmv8aKg0AZleMm5rMFAN87WKDCJEKnyN4JZsKyCxjDbUy97Dd7jn/QY0
62/zSKkoYm6ChTKDO1Ff5NhiIK/R7+fnVtI4QYVFLGsERFg8ZZFua+r4s6PJYYHd
9Kuh0EAaEqSCHQnw53vQsnISfzyXT7QNkHfYJWyLO9yJa98VmeClaVDvNE46HC3s
XV8ZevUYJQY8/2jiCL0fBxeyUkAsf4L5zOYOgPPCSnSWciHO/o2/Iz0CVfz3X3d6
nkIo/DdK1FaiZOpfhOaf8xGI/41mYrSQ0raQZxfZE+vVWNlLm6B9TNh8LVYKsGMK
ACCvogN+fM/Wp/4zjL1XwMIPwRBwdOey8cSeo4AwwO6bnJXsSlDf4CJHY3FiZo2Z
DZ083IQ9JgiPOshBaCMqKQFG8HZYObKvorbHdzaMHbwc+SC0A6YNd2qznGKwIcIK
DFp7j/Atq+eSN0lrhKz5suGcdwg/7/FoatsQL+xLMz7PpJqkYWOn2PHdz33Dqifo
UvXdT8AJ0dEI4+v0QdFdsz9yvtUEFhJuksTNT6+INJkw3j+Rub8hI1X7uAwjnLt9
ktuR670KuGmMJ6JUT/+uFhoqXnpk863r3nRHs9/1jjD14HagDERyEtC0+8NZykUJ
dJg0xwjxFQYpc8yuBT78VuMn2Ze8inZGLzzRu8+heQ/eXLZmMPPfIens8sLhc9Au
N/hyXlh+8magjmwiQXbxY1wD4C/Iev62T8aLt7xMymVT2uVH+5hmLfoV19jcOPeM
2bP3lF4ava0qRUZM6v7cw21vhXfo6l/nbAsvPD+mo2SkpYzu1qVUaUphpMVGHnqj
1zK5GGIfBtk8vgXBIEnf0DXJddU009O7W6iEWiSCfYzgxz48odwHxHfyCpSi2UHb
E29hP2/styho0ePcUFOdoDyJsyX28KGh2UDzm9br4URXQ1JaKKRTGADZLixvSnFt
pyJ+ly48rpLQhz3ArFWwduZfe7Eu65odjpeDsNfptoccasl2FHm2a4J/3Tu4rjIe
MtE4dPCjYJ4++b7/f7sQ8RBkTjvJ7SHABYHpsPyTKmCkewS9rc6xCKDFZqjgg0fX
IBxke5Wx+tImL/+OWxsbpYr2nbF3ZO1cm6Yi1Di2jFsv3TCF+xjCTfwI0T1OQWmw
85o7x+E8RWBY+YiWx6RbmCfz43xfSsgE14iesjWdOy8YG6Oc46dbKraOBGdtaBLS
45TTE8Cqp6oPcJ4xZdeoDoK4Bx7vx06XzsfVvjq8AbUlzP7IKHxbSGZZ5j6z8DGC
trJf9tiGOX/xKSH0rZA7mWpdGE2VwOOKsRebG3o8ViL4X0g6+43wdjLf9/xzkCdi
d62cfdatPn2eEWfMO0AmZHy7bvgALGVpPi0H6487I2QmILNvXs+cVirv8p0lR7RT
9KOIHwBVODFOkYMUmBtCK+aQxZY5yqdgAI2mjoslKdDJTqiIbEe65FsA5p39HHbx
edsxiyo3m0ck85qKndto2z5KbOSztDYYeZSfxdExQgvcMs7cIO6LDRfXePEKan0M
LAUnwVAwkmuuRW9/huJWQAXQsJZvsF544DLyEhJEexqEJzkPMcM7CzdQkLkXCBf2
J7sbmtZCBT/Wd0VTrSy4xgKR9rJ7ydShjXX4iGF6yVg8TUXcGriS6+ein5p2RATp
vUPMVDJ7WKTe7/YBm2fJtJ5z1o0WvJREMd86oYOLEK9Q8PXHWtV/y6Kcgb67Unmt
wnbLbuSrTfo9wNRtr+Rrj3nP1UA+jGtCTEslp4z15CS2gmFnrqJyipiJRCHH1iRr
xjezFkxGU043icDWTCuf1M5+BMPfVwAkYIkL1EhgVw30TRgxCaiiEzO2OdY8Rtku
iAJq3QJQNv9MspGJGGOCJOyH23gzBoEOVCXGZqpl2AaAKIVbtK9B5eFTa9hBbXSg
p8EtwvRFeJcSXzuW1QbBRUhHMEjBaqRzW0hucZHONiJDkcaNtFtpGtU9fQywvdA4
JguAgvRQHPgqzveYzQUJnDH05MDaf51d4KvXOTQ19f2x/YRPhEunn+0LUJdZJVY1
0lNkwuDQO4bR3HBH7MGroxDg0Cq3qvB6gTXUVTFrsvLgiyTOk6RfgpvEvTL49wK9
kigs1bUyTOb1T67hu5Wsi+iJhavKP88oFZWUY638L5PoVpRcW4uSBMvi3EYBd5lk
WzmZpBJ/B8ghauYPGxGuC6Gf48s86BYKKJVheamZ1JPnhf+b83b4FB19qImWJcsR
UuErBmHNu+FWpPCrw/gWPAFBb/SdVygeRFoPfnCsoUQghN2vrZYyMwbv0wXBWWCi
w4p3yLrGw0lTGLiCKNZ5GBEqdc2V05g1GMh9xVpVEH8MUQ2Se9OCgIhEfx/N3gJl
y/7l8npkD0JhxDOHs/RckjpcMdPhdWrDSqdya1031JBQD4g00bkBEjbSaaOf/NyE
HKCti4JCRXsEM4dgGeSQ5iBq7P+ppNg+kaQVSvrH6iIrxNnj4rPdWxg8bdmNAWSs
NBo0ERFenrIeOyYFD+8Za2SLQqcEIicK2yFQEgU8vxswBBU3575C3DFI1PcplQZ0
lvhnTLMV8oXJ1LsxRFyFlW3RGp49Jfy8K5dsQ6lcD+LKm1cGvQSgLXhZFnZb+Qdu
j8sftOJPDv6JyI3nMfWgnHANfn0YQqkWYwF+UBrZqZ2Q58tEpUG6FxNUHNhnFMtf
9eIzm135MNMboSot+Ow53rbTOMCw9rTAj4Dtw1ZluUFgI1cqqH5S3N3qfwVgJK5W
AJ7j/0qv/QZrD8J2ILn87T8EloDq/oP7fz0vNxLS/HjJ1QliXPY2cYID5ZNPsIn6
bYkm/NAp0lcb0X1kuCnJf3G0GbvKryKuZHZHfUN0Hu7AAeKD8YeEbai4EyOsvGxj
hgoVtzrngzwHI92M9HRX3qRww9Lc9KfgBFlDmvOg0Evl+1JKxAspnXGOFbLU/Vav
8iSY0VRHvBgHCtfChjZSIBJ0WrnXEIzUjEGVvIDTCxMI2vHbo9P5zuV+U+oOZ7RE
OG1DMTBzlZ3+fBvbr3NcjmxnY55WhwSCv+EKciK6uJq43VvMOS4xvfeMoweDh3gg
ueZkWZUagZxxnvJ4aMmx1UrXHd1unR2n7cuuOK71IEeutulkPc3Td+BF7Gy2XTbp
u6cb+So/StVPj8GebFpQnvE8ABRhQXUMYa8PzNOH9KVYjFNdQb8XVKpQAoxhIqQD
DxZHfHbju0MdHTIyLAyWr8KrVUfJhGLHjBaDC3H/h6NOpktGRofx/dxJN6n5e624
giHATrxFhnMNgLbt/auu433iW0pi/WBsl3T5oKIYP2bQ9B8A92lZl5QuTwGpo0+H
wpypN/5bq+lAY7jau5KML6F2LqzFlwsWikRFkWU00VrcBTohGVwJFcBdZyZedsY4
928SBgME07K631jG2utzRsErDIVnB2eLOZCsxOq1BaZ8Rf4hWv+4PJ8RbghBSBfs
fKjD3FLkNQhnjFh/V6YjXvvs0+T/Nmcah65E0olSRxcA3SUBnjQN+QwNFgccncPQ
HXCrtpqszYWA8at0zTW4Ht5BitBNre4SmuPDTX3K0OLlgW5W6R8F9t8v69wrbbOP
PXa4DxJQwaPkMyeL7OzfZMiJeyvFn9CbqpBJmIS80lpq5hep2N6k3slszJby81an
H1XOWZ3prrjEHIwRlfpZQtY3+P3w+SDBkuv1D20BktioQ1kXBCCOBs0idvEYAbAL
KRJAcxQDRD0eWN8GH1cwEMTbwMPZ0JIhCPj1/2yfrNQSfhikth1xTJFAk2Eyv1uG
P2mFtdgHkzSz5nPMvTh71dz1/d1wc5idNhBn/6NhhUrtMedKrgef1PmRgbLOXjWh
1EG+5yTafbKrP3fzO5nzZEjwlSD4rakQu2HSv33AEIZf96BJeJcEydB4C4EskyLq
pOyRdS1OK67Fb2OmJ/cL0cNCIW9251FeEVWfjRKu3ay3AheXM9s/jWqSGiUbg3N8
MPHjyVJC2huybuaA+L7wmX0E9up3NgPaFwrjwJ6hswLrsnzfYKJBmWgeBZGK2iVX
I5X+oGJgVAAXjQXOeDPHJKigYokmgEtLARzEm6Bos0RBI+T7MI0GN9Ns2l4C5En+
4EUI7zR4PKk+Afj3udYeY2FxoZ109lSI1w5NmtajN3OGiv2wS/CMmLEqRbvAdUry
XPtu2qsaDKPNSPYBCjryx4aej6+GLMz1spdTxJzpSFZvkZYd/kKTG3N2cYECNV0U
wN2JbfRJ86Ly/sjjSMYn8QG389HQxBIG4NbXm+91FAAdUFxqP7wusFP7f6BbXkcr
qXYXa23xsc05YscOAT6suXxXJgefBf1Tt0EhpElL+iuBzufmCa9viD7uop+52kyU
VJbmba5m2BEHQpGTwJk4Axh1pIfYUehINhJqJpEZkoDr9w0N/X/YJWV4RB/7UTfd
U8aWqtmvhBFP7swRIjEuCVzhtn3HadqFr8bpkIBowJZXz12dkmBsBnLmQHs0N5Z/
c9lADMI7GwXIjcUhZf6sBLyED5OA4wo3Yl/HlVxcq13JfNOTuOV6S5RP6YgzRDZ1
2NrSGQDBs5qytqI+XOrpkjPoCyYKpLUsE4Wul6sCyqRBFLN0f0EeKjUJss8tKOLo
i87DDgSYxO/1n70X42goIxgfWewsquB9kesZ634hkJH2X3LIWod/FWf1iOqcQIvl
vBUZHaVPuoHcLoeSpNDeg49TKqC4V64txvAWdX3W9cTk1ETMgk/C54+e0x+3Rd2K
jrxAbC/xlH+qpTulaEwHeTWrSA11W/1y5F6LujvtvU5KnCmJacl8GHOXTesVqN8x
vi8dgc2Y2XvQ5utqTxzeAzCvHYkYKEQy906W549UK48dNeeKacFzp8YFeVWJ2uhb
7SQDH38Gd5EXwyO1j6AG1MXeeDNFfhYSNoPtMkLDyhoXiL16u8EPrkjFZ7Etpn5f
nSullBvfgDLM2UL8jJk9/LMnuyZtE5/Irb44BjxypSgvFrpEHszVY6did+vScx/1
PYgFzLDyPRHQB/0QsT1Sprn1/UxTMVUlJfXhXVgBz1NIYkx1JJKoybuCqHnVA1+A
dQHzem/sl8cNfUivKrPdKiZTO8/EJ81xfdNgPfMYj+nk7Lov2JBSO6V1y30ks+fL
utmbok12iIr7RxPM11/+9hRYxDpfXgjznlzg30ng9J+zTCHIjOu2NaZ+SDltRVK/
wymqySm/iuwkF1Bcx+eVeqeZL5rbeQaVpnxWn062RuiGYBlHYaA/674+ddAupfi3
et3n7PTQYxajHt6HLPYT0KEB8g/zbo80loJHypApGbFmHYum7sNi1ri+/h805Nxp
LI4tdyghpnwNHFoY6IRXBo9Ueee0LsKB5b40SA8SLq/GA3VAhvKMWD9+9fcwctRY
hB5nRyOaHnMId4u0Pb4X7uhrzXM01c98SLC013MHLTJY1XyXo6OJMnqO1bs3j1fb
LFVEjon7Uj6jJJ3tnOJTYtk6a5qYyblDfdR8kRz5VoXdvPuiNep1TjGa4GiCqxjX
qHDwBj3j1aJEo2J6fJ4J9i0QFgELjd3PICw9y3Vjesw9Zc8RXjH8+3Qf59lU3CwO
/19AVv9TO48i2XT8/eS+EMpjCDG2h0WhCQtjCR9y1DGsHwJ+J6rTsh8GD4AuAb1U
iTJACFP3LI43wkqs376+lRxoKNnEaMwyuq24ZFK81vVtJLUaZcXAbeypNk9oNm7t
Z9Uj/Q6CL0a/3gLr2fi3edEtwz/pTbR3p/JBHfVtOnvLvf9cJ9zJMHgAiOx+zy+M
m+r+5vizQhGFxwJlEGASi7XmWhw0QESZK40xb6cNzAXBRnqoUDxSx65BurZXcpaA
6cgW8PrAs5zvMutokjs1mg/Ak0WFhpRBPzEx2zxN6OaF6wEHdw9r94NwC/XkK0jc
hI73v7hJZ2Kj1WkRq3QZJOe/db5Xsi8zq3yEe8EBM0IcjTmdagwmr5hQyRuY/Wa1
D7PwOnQu6Nq5VQ81tIS92cHsIxTWetI2F9rU9onSR/1H/jcwHjRs9dxkZOKNNm9l
tNM83bwai+nT+VrqDFeXXKvLu9esHjbuVFaATexAATj+v3IcM4jxSza0z05BkU/5
OcnGhPKxug2D/ZJcGSKKVrMxEnvBOxrafFCu0KjiqOT/w0fUqO1/dIiRP94nJZs1
BhPibBNUAP+AKFi/D4GqGNPoodBSGcng58hDXHpU3n+aeoieBHZrr8C0PMnfdkCt
zXwr/7n7XTAIW+Pp/4kULTSC/NoQtg2p/QD20xw59zofqFhHwXxU7YHE7ZgHYjN5
E6DCw1neIty1SU+Uh4uc0HFdj3lBiV8JPpTu6oAQj2CMYPw4vMZYMax3pCpZBGsJ
sQLDVMNRr+0qyD9Gr/8US13d7us45c/cE1tubjP8PqhO+Mzz0D4XoC9QHre0buZ/
zMO/HDLbiIiJ+JzQQeBe2u3KNnc132Jba278REwYXxOzgTguNg1pGfL8QrnAEYVa
PoPtBeJoXDObEtj3XX7expDANrEiusm/hY1KGaOG/WrIQEdT0iTFKJH1eSBDKiBq
DAno9kxgB0pOidQKQEsW9jI85z7ZdVynHhZzILuARRZ6+olohoKDI+zGEf5/Rmwf
1k9YvHCyPqqukWk1ZDjPiEfBgGgxYAwu2f1O0HzLHEafRB1b01//qxVdPIB4Z5Vh
5B2ljIZbMdvnPS7ocxKKTeu08bmbYkl1bRMT9Q4ieaqIEAaESnwcMJsm98Rjcuxi
1vj5t5A4AHhGGQOlsDU3yYXiOQD82968W+olRQO00VL9DITBJuRgTv2E7Y8YbWYZ
wBbcg2z4khK3JvRLneofXxY18WD2UGT257HVHgxgA9wM5YSeV7mOmEdweoEfPyqw
uiAsFbMkhoIDBLR4n/D0XHtalOLW1KRW10+DzTRDDSIjHof7uLSfMRz7eokye16z
u5gdI1CZPGYV0lu+Jpi9E6jBXW666TV0Yt46TWXCAqJGbqcLbt1ndA5cBy3jM1k2
rWLmxy2vnr2gr7uqewWTg2mTn7HjKEeSM7Wq/cUfn2JM5xQUOL/zIfmBPfQU/3D5
8Dqet/CkFSzYQpEq08wzzs1go3YqBqH4f+FNqy6TilWm+VC2XumRqT8hhgdGNYti
EtKsZCoEh/PrG5g8LvVmToWxa9dPMUU/jZDvLVCN3h1BTZywzwlJOHD8qqZdqgKF
DlmB3oS+oa910EXwqccIbRGV3Nf7v+YPDbCmqd+wy0nIvY5uh8x5jcdNtWdmaBeM
OWzD92hhJBUfrM4atoFANgbm2yPBjyfsCI/gELRc4CHv01/3MHdAeFEIbS6gymm4
Stznarp6djl1ZCiBR1KQSUSOk3NLeDdVGi5edAX9jG2HZsQQzaN54i2sm3WZtxb4
hKvNY9SjWxYsb27FiDVTkjO8o29zQJ6FZOJFJ5dWO/JcfDSPvZ/aM7bAjMKLp26Q
Siq89hmeoqNKIsKWg7n3wG8tC0RZV2ZAG3TQE8Kt+NtONEn+kbQ/YkZkFr7vqdcS
h8ZfYBB695AGS7rkQyuGZnONrBSybXFzdR64UdJH3nN2aCHpO7yyCTA9Vaa1Ka1w
tDtTnqd6ZDnykmotKiBVIlAsh0nsfHddL+KM7UdpwNSQwlWdwcpPONxIWCsYAvJc
B36UZiacGO+7tzxU+78CHq570t6VhDT2Aqv8LYi+nb1Z9i8XDiPnteKk/xFiZMn7
tE7dJjJxe29Vf7Qwbwa+qd/HivG1tSd8r44Wy2k5rQPJFDTYTM7WJwrx0c65mLU/
06Iq2ZsOreU4DB7mRQEjdxMslmzHhvIvU+z4C7R8y/VN6uSer6lk/aV7mwW2H+3o
ELuZgJ0ockhOSmTDNpxaRWzeFMVb0KSeU+FNtKyIlyD5XSEL5sb4E+N/ZL9p06oF
NKBbratkL3tLQaL9NjL2GLd5Ai0L4f6EvTV6dE6EjA9Pf7H0pNoF9pJFEHvdo54f
1Oz3MEsd39rAUe9h4SXgXr9miQGo8YtV2Sp3UxqGEkk5Oekkhtxjec87bb9vCokD
d/X0Da1qfFS1Ffj4DpS+a+LRaZMtPf+aLa+Rx7UpNaqLfjJuKsLpPxYwBYPGr/1b
6IECRCparGSefDI669vUPn3YVMzd6FwPqxyGD3oengy18+cMJbvQcWm+E9+A73bi
osvnqL3DsTU2GswJyem214z1rC5lwQCtTh2AUrmMXKenmloFsUNrD3ZWKcadS1+1
2vu5e0ViWq9QDXZKwYfk0R5C3cK1zf9jzkn2XIy6VNSXIlcI0wHAnmMw/B1O5pAt
jmfhXlXUZZ8wofQ2dJwuD6/pvD0wLzCw/lETPQqit5x/ImBpDvnREgUENVrE+QMx
E4FHSWExV1GhUrxX8cU1IoIe3213slGnSLf3EqLKQZTlSAdcJtim+U879jW1RRGI
MDluIhbCDrJuonx8429BHl2ljGYldSd0dRIDoDZ8lF2z54wckhMicB5/oVbHBd1l
1/glmBR+ltmuqgvwfhnQsp8F0/OzFcX30vubhBK3iLh6hCVJctL95lyFj69bE8tp
iUsyKZ5GexdRCl/1TwMogpGRlXvD2HtG9492RUg//Cq5u8bB6zA4ShnXglGrExM/
LBOe4uCGIdL3NfRRymcrKLd7EYR73QMz3dV8vnh2x7RfKpwNjAxpkppahrlETo0i
545buzQtA1sGcIqTHpvkS9hAd0nxN3hGsHp4yixAsV0z4wcUvlqeY8YmT6ttsLdG
7t3kr3k4lDz9TQv/+xgAjFG0g0JnCaKszXwReFHoum5PaGroQaQFgj59FVY318ki
Imr62LayDVFfazzIyzUmJQtYdk/5f49d94dXnZbMY8eeiivdg2zDv52ZwIE7TPau
pBqsSBtUI+xLsysxpgh/0kvihkUSML8q8M+8WYVAeFxiY+E2Q29LmeL57XXzc/ho
RinR5Kr+z8HT30Y67Ke+Vhd+VCo5AAWaiNvhXIHZlmzn0nBh7HtxZD7nRBM3MJxG
oXsfQ5kJ4mhXcozaX2d61O0bNKL8MFRvRuNdvZHaEJeoy/mJQHbaZLxUqC8EJBJ7
AqOtHHKtdk2Tn0rBg2UWHLrDm9MOQH8H657ZONWfW84=
`pragma protect end_protected

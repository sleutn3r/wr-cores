// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N2Kco5xayZak692V8FvINTAanYL87lz0bbvuUS0ZDnl5SAZiMGzW+Rh+HbYusm4s
inu2KLzOAHSTnunQBqK7ZmaiioX4s4Al34ET1mo90UW8UQDoZFLbWRsF5yeQ9RDT
yLK7PC4RF55WFerlt5509zdqrti7x9fF4woNcoEwFXQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2976)
71vy+CKybfQgrRE8ly2NGpGZArXsorCcuxH/fq3dYSnVfBqT2zt5jPdkHmZ/mSnv
roBFtauEa8zucyjJyKOI0PkS2J0XswrWPuTZQGgtwaeiDiv6cxEpN9apA8tQC3AL
ol/CUNbm62s/r7jF60JS+1+XKw102EKgf+MH6StP0yMcIq5c/6eqhFvAEjWtKzUd
Ih0f7eVI/lH8whJkBv/DO9h3L+ZCOlDYhmuh0RnqCqK1KH4pFulZ1is1flX12zZp
HlEQlCaBBeQ56ow9j+C+OdIN5gyGBCs5A1ceEXXNdYasCa3XjgByfqJqEAA8/5yd
fzrMfWum5yW71T1a5C8WAbXEH+8BCrkB3/fI6sDEGyeFJK7oXtFSRs1SCI8nnGji
yQ40K+m/rBzvv+f8BOKqbwBiHAnyeTOp4QHkAz750Y07WiYvypaM2OJ5kzLX/aR/
DoXsV1vPzNS7lUMqmPLSOl+dyw+EMsWwSSRefvjRF6mPdwle9ipGg/gQzNYgFBG5
1nPK8DYjly0r0RcaGsECByCe88Sz2XbjsKUFK/coB/YID6oacGjGctCkdwUOtKWV
TYkXkkOEmlDpoJU530pL68bYnQAKoP391WglNI+PuPjkERlREniqR9MiPMpR5mMD
vbZjYNJIhJpL1+AQigfrVKWpjiZuj+hivsuVC4NXTDNaVDjme7OdI1OlgoyTXZaG
LeuadIresXsDBsdDhwwK88W5w5PLTPrFJd7wRf7qXJxR7/TTz3gkE2PjG4RF+fQV
3ZmBwa6sfRk4LPm8QdBLm4xeusBbWxdByQ2Om+U2kKTQgfPVKElVE7/dVCWnZ5LW
t8JXn/X9TeOEZ2AuX72UI/Zq72itCFeNLl7CSoPPvrobo0b7f3fdBWWTFdwmvdTT
PqbEh38uNXHVXoV0O/xIfNZqW3cVzTqUAOcW/mV8ZkXgxCGZZjhTxkH+DhnTdPfz
vvTaFFKe8ZOHHnDA8tUKjJJwpz2xo8s25Ydea4xPnVQBKwDyXbsNUJUP0lJqR3ua
LOE2dMSCG8vHQSgTaiDb/474ukx9E6D0fEx/VQ/w/vcODfr2oQsahVNnW5Nh85M2
YO99qhBjKLmfkfihcWtxURU8C0ez5Yms6mLKDftG5nGnfC+CRVHQFb2ajjBvDHoc
8Q2/cDx8c7V83n5AES9vjwp9zNEKlJOVsScAAKpXgJRgP+3BSeKoMrukzvSINMfA
KhIx+9NjsN/DGJ0RIXjSdxS70J/Tz7pMf6pOqBIYw3fTKmpTmx88rNsG4GQwfCSF
XMoRVLQwtsvvH2GgfTA9jgx1y8WjdxOwERLXKQsfMMePC1SwqElwVClqwYHOs2yH
PFHvLL8V8WzXFX4xMQ+CwgSY5eU8qLlbXWjIwZ+FID8JGubh7EVeMLHpKAv8GPvb
6qZ26NHHdjFKODsdLM9Zk4yDoh+Xxul1COP4YmrH4Qfaa2bAjr8f9h2X1hNcuAXx
/ZaysrbOk0hb1rikOgBvYWODhmHIFqqf7pYgAHKtvBhdTaNXRwzDutH2giyYMYQU
erHdYMU03XMRCyjNlCC6gREE4kMQcCcD4o7SahAWV/AIO1GalTQCCWonMbfpMrzu
08kDavYD1s7iAe0FYE0kDF5/obguTNvXxoL3OhyZQWCV5Pf7GvvabEYosLk547QD
KTLe+UcPZBxK+19jNlQBPECeaF9cAuf9F1DjjF3D6yiOwIkNugoZUk9XCUZxzoCN
yTyH8hgIjaDJ3/EcTGTWjnlN9whMuOv4afFqkxAdFYNlFBigGc7mLBYuG4oKsr97
ybCYl3kQNqkSu7pOcqiLZulgE+XxUAchSBR/dgodpodtz5tnCH4CfKijqsr0vuup
1fPxgehI4eAsetZl6T5bQJz6OrsRXA85BpoRjA8zpto973d186LNfX+uDp8hnlRx
RcpA8m5LlvsTkZ0uU+ej67t0cZtwV73N4azhPDuXHg5mfUMFcsckadwWT/YGyMWH
TVNy/zAl013ub/RykPRo2rAgsFz6SRye8dLpk1a7nRzfz268SSx858BLKSWgwdeA
dQ1UTW/XRVy3OmGvO6wCj9TEl/f128ez/1TM7eLmImubl34bYhedv9DSsFA+YMKi
c0MWWevCPlympIdcqwqR2M3LG2U8RHIu1ifI//6UIxcTCsyKk1qX8dVPalURpgx5
zliK4rf8EYGICmfa1yzGLoMusCfghOQGKWmPIg6niPUBdngDAUO+f6bnCOJrD1bt
t3Kf88kX3gAWNX05RbT+3c1zKwY4sYfONBAlvoU5KU8HMFC/yTntj6F3re1oC1wG
V7mHlJkVH/uPIwujnbUoQBrU/0wY7OfCIoNV9sJY0iA+7W+FBp6kywL7bu/29vHN
KlOKs1MGmygPw9OCmQ0I2QdO0p0tjv6Lkof5toxRR9DTi+/a4Pxo/O565tTJ+POS
Cmkziw1Nh2vrOreBfGgTbGtUrmMlRoQA4G+cU2ZnwK8h36M7NmsBt8ZbLE86atYm
fMfEpjQC4XrD07AjbTwpqbcYiGLgduQCqXt6UTmTvsaWJck2+0P+p/O3lDIZzi4z
j0HPvrdiFRHLOH59d/wWHn/TD1SBxbmvcuMN7q8JmCA5dTzttJCFvzyHOaiYvAZt
wWqTTo6mNJjW2ggZjvSyD6TJa1mX7qsEbdFQ+xoaRnBPkeqvMxDVUvnwnsZDf0+w
YyUautmoa/kwwU5J3jC5YPKjOEwkwgwKvIib4Zdcb1u1HvSJSbLqvu1MRMCzhoGX
02/vMOv8YwGfBfXVXk5cdRyww243UwozFDRomqhrYchrxwd/fnsQKePadX3SDHdz
9BImm1fn3s0bT14AWB+NqPUdEtIzGMP7olRC+nFXzJhOtcwckKtlRF7KMfXsiF1h
e02jtWYnSPXVFFET7X4hB2NDIYNmk3DP4+qHarisF9QDLLO73myANijwjlpNCUu3
n/f7Fx9vz6MGvO9WxaG12yeG9tP3qDZBNjydrNHkey5a2FDGY4mhwN4Op7LMs9ww
25cREYynnkJE2Ehpk3+6gLfdZmBPEf1jIhpXIUiHroyuHKirJVXyjdM4LNgqEgYd
uZmF9FKsw+57R+zreSgLf4P06hjsO5D81eFCjC1FtQGhaQ0wWz+YZz2W0NhUKcPW
JGbEXwii2L3h+byAyALXI3mDXw85LsRXVX0nLcPjNZWIeMhrUhE7Bym6RgjECjP2
s5bub+Xj7FaVI92W3vol3enaCEmPQ6mXX0aDNCX2fJ56d5/bLn6mIncx74cFVQBW
YZs2BPjyvnMG9nLAPsZqFzGYH4rywhrjIVYGUf3pRpWxshHs7akBFI00hcGzc8Mi
jvg6EJKmjj81XjoFiEcBi59QBXdDpRZXZtg0PZwZR2puSDfTVJWraNal02yVfZ8L
jLJ/gMKq+BglExAEyBMKGyeoki9dcKSb4PGEdGtuBMumMAsyp2R9ThkW7XO/7iS7
AWM7svh/S+yEluLLOkeIQTjVhUg0uJnJ1EyQF592Ig3KUOnT4JqABbJO9RgGsbZm
c97xpBKf1QFkR23rcEpHiKLur2yijSyPAdaq6GrJkqUGoR2EyxeaUMTioHDgvRxf
XCYT/R/SK6nHeCph9uoS9eFRjYSBkMilHKnxr0d8/pYY/KFK5cDPUco/9p+SPlhk
QicCpjlRA5UET6GI1pyxOuMFyRUbJfg+UCCJMav4RI1qN1k5qiYKFULdWk7V+HMe
YkUi7VAbN9qZBSfvmi7fBYCs2+p9jbNvOfWVP+XrUVt2oE6fzPbln54k2VNoUxdw
AQWCsmWoLA5bcuVqbFlywt/G5aqaTSfj8GFi5Yd3jtTa0J06iYANC6WSC2DsaUU1
raBz41hAU3T3J/Irg9Pf5HJiVMTDuWUnTfT1VFrAFQa0S/l+5Kp92+dAeB2CGdRv
KE4jcKl7el8L7kPJP7eOuQFhNhJ1D68JJKwX5/FCha7fP4OTFJnZ7boRZHGzGcu8
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oRPt6OdIrBBs4hnAoL0kl5DN/2L7zJWA/G0l4lMXXFpqwtQaSwmu3FTwsU/K2mYe
RSSySLPVS7RGEQAQieewwhAyLZIxdnbtbiZmCgusfXRpAxWiNlOJEMSAVaFpwizW
GKnoKM5LgPAQA8eNl/+9iTkyc4hY1D+OrCkn/5wmlU4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57024)
tQQYGWZMM4N0Z0rjmgPhSpbDuBC1TafDL6w07o8ERWNscjlDgl+vJfY6D5vjekx1
dYpzr/x0S+HFthsusoZkOK4x5TJSCIpQtB3FQFJIiFEcoVUmbQomN0hL7j2pwJ5+
r/pteEEIrwnP9RuGiuW73j5j63T+cM3Cag9PjHfaPMIUcYGk2VIgZZq0/GqGF8Xd
liaq1iHFpK8YloadxRn2jtMKOZAxPQUQdUfUBrfpAdIlnQ4OzWUty4MvCY2vEyRX
XY5ya6ujw1iwObMBnqAtzyQotgy3K2Szqtl6DmiRMrHbC4evUjfxyT+sTYFbaRBi
7n5TBS8MnNbUoa2LLYci1MB2eIoAF7SfldsGq46URoOVg5/gNVb4dHk1/41tRyha
6bGm/tyF0AgGa1K0I9MdBNOc0lYuuuELKwG+H0lqfKP+6iLGErEB2OSf75S3GYrq
CDkH8VDHv3MZvCUKxINRor9WbmhS6L9rQGHbwMXglpr6CJeWzP5qalNsBl+PExRz
dbBCPbinTugTeRQ4Dk7SY+BjPKPhNcs9LJ+i7stW+1joo8wIcyr5FjLR1dgh1VNC
hYFe2JqK3Y4xK6YTEC3MAiFLDTEAtKV5q7jv36MAViLfb1xukvyaEjaDWjXNQgCT
TsSlrNUmPSFSZbwFHHTRx6g0P+x6nnWrkN5EJ9P2JogC+qH2HpTLrkCMWwJNOJgO
pkjSoLTIZgor9cwqGnHT9ka4UYa75ZDMwrgDY6y8wBnB7AIzWoXmRfFyX7nOYN8j
+kG0lscGVEi/ZMNym5XPrHv6M5oI8YVhz/NAPjSnEjiz9vDQf3isEOjyW8uqfrfb
oAb34T0Gcm/Ho5tEsfW6zADiKf/mGYiU43oohIPJ8+nPugaO1JgGVecSxtzs16dU
2dmYralBU4KTVA12knu28EMxxMO742/1ccJDe6s9AURzVQ+GcnryDZYsW7DU8G5P
V1vuVc4QYd9Uw6RR+wl0B7c34uWu4aGAQle2o0LghnBoKYCtwSYvCY8iBz51JX2H
sS45wFQG/fJkYvsqXi0c9qUkS5frkGd+808EV19ZtREj7ga6JqYVOW0xPHYlZhIO
nlwzgyzQxBmfppcIrB/3pRAgqfu5x+2hwnWyo8Q37TLi1KWttk3pAtgCBFWZ6Bea
hhVMFhyRrcvjB6T4Z0ztkhcXD5s5rIG9KsYP+KFvz92ceWk2Sj3gFhN//2bjIJsh
9Cakm1k2FlrZttFdLjsNzYdQ3xG1C9uw8eqpxzNw3kLQX1T++4v9qTRIeoC9DnwA
KfnWR+szFcU7YCTUFwmGnvZcq9n9AE3dX7irAGlxxzZKSoxVkEnlB5vYYHaipdWo
AHj59QRCuueEdREU3i8nrtposAiSBKPlHZlb/14X3Z2jkHeSoe3eOs93Zem8rQk2
2chXJf38hvN4TOEm5L42Py7voSYINP8reT55wcFXmVHz1Ugo2ahw6tbkk/wluMFi
gNRWAScbgEOzoCgCJaTPnEU4GbjUc1Hdr2wl57x2JH5C1NRERipUAn2Kern3Zs4J
wkEf+NLho1c5tkO/8SpsjF6uqvXWEcSbkg09yhmAZo/TS79Z+Tzr9sp1+57EWu6m
Iv6axVlpPzBkK/WMGc/XY91880AUnJGkTJrgqvyRTpBmR2+jOroZs5HU3x6FYwKt
4+ToKzXiIfDPI2LpsIk8QZN2x1c4nVd4CIzM2Vo6w2jL3zWsa+F2ODkcU5bvK1eF
LBCpqti/SuY6tcUygSBvZAwls6gqObbg3x1j3kMryuBpPY9n2EYHTuAylvoh73Db
OORmBjrzCrbo70LM2qeKpPT1lnufvA37C/szeIevS1cbYZ7Trx4ByWGNmSz3NE/8
UNSUR/5X/XuRakXFDxk5zOvbv318aH2zvEnnz8BKoAKJIn8pBn8EC88MpbqrCfey
e6vopfXOHqqkNQbjMmLx75Ql6GjZ0uiuLVH8kIf+WmcLjcjUZ+Gnt9waQqw+G26p
OUj1MaH94eyyz06MPsizZHqf0YpCiqelqBLaCvyD5CjsXe/cM1OS0rEOJ/8vlFVt
S3wFubAqqpxi8iV1kY3AzdNxPSSEtltJASPOI8Wtj5pEhhiZTrkNS+m+zCb95x2I
7ymFej8HJ5hSaMB2FJ9tsIfYwdhK8mesqeNdyeQOPJ/BVLxU4lfFNJGxG+rKABj6
MUcVUb7g6i0UMRYVwu818sFLjpxvCisJtN0bG3iHXIXnyINaOxKDm0GA2FaBZycc
LfGi1P3W4FoMo2jM2+n1W132p8SrglQf6eENH9B+o8j267cIEOSQUm1zUefof3wj
3RS3NkBoBKZ8UDa+T+7xq/3ANsNyWP+DgeD+U364QRKf9wyW3mlbewJIKA33fBb5
CKh55aRGAbc4ihWhib1XA6PUIKdfzt1WyrgZNxV/CExWFVYBkOO8WopZM9jW+SQC
G07roC6Y3pOy+6rQZ++TpvXItTx6wHVrxef1fOPKvzBhenO0wG2aIcBSo30PeCT1
qB4OS5ZOTO+cc6gqyIC1k+a7uwvOajQIuLKHmxr0To7XiKl2Ou5p6k7ZN4fgV3Xd
uPnyXDz916orJhxbuf1T54UTxaCqKgCvg3G/pITK1KLVPmReY8e99uBVdK1yPhLe
Ifnrsc+hm5zzMRqG5qQH9Jfe3szxqJ/huXKpAfSfqz6OuZUuBsXCEdcpBNEADAjg
AefFZA8/Qjq4RFXl+H5r0txPAt3R7gSVnfPZVubR1nYApRXc509Zl3varUHaQJtU
HC4DfFMsC2D+djT18oAxg9yaucFx8VnhVigGT772q5ohqdIabzWzUecPZl/EWBUP
1NaqcRkeYEDrQ3jZjtxoE3q2w3oS3fCAUZd6liTLq89PCGTDrbkATZp1G9p0wEhs
wVOJ7JEJ++bF6K0VDCMBsLAe+4NVcLbIbYAxN2FAkypTIFRgyahgTasFmZ/ofCUH
x+jWj2qqcsLk2bQ7a+vIAgU8dZIKg/2ttP8+908j+wsih4jvzwTZORbMDjFFSLnv
q+qcluU5kRrokHJYxPZEC+90kXgiDLRyxC/pDzY6q+lClFIgLYN0mHmqklybNwqO
fMcx7mL6w9w5VfuVjQG2s+fig/stBgJfv8u3TAvgrkv9vBHMzLII8y4HFfeYHJvg
gNPDhyR+Mj29uHJNlgysqi+aWB377X/0Q7vakOfJsujdLZjWTttCAhBWEv8ReA5i
CgOlKh+xkJESz9eNHcDTFNMkBJpH4PCsTKhuoXYsK9qwATg1uHeDmlxs3LkVk6X8
aVbfYHvRBNfPDzJzwUi8TozQdznnHX9u9TsT7xhZAW/L2r0QRogrslc95D0sr4Cc
3kiCFxPRnGJLcrYyBur6OnwqtfmOySKpQBm9W3UWQFNf6Y6dBBez4C/VCrWDaliG
CvIgKRGku4TDscE47KJed/WZmtcYPip6KOWg0uj9jq0+kV8XnNy9wDHYcLi5khcE
S4ZjN8BvtH/FB9MEmt1mMoGjs9YcRyF39WJVzrO3PD+ALFl1fXHudUmlcGBOI3W6
AhqwhEY4KJJ9TiZZ73S1V2llKLi6NFA2RMqzbsw9JYG9WJaTI4Si4M1WBzEaxmdJ
xeP4Nyii9LgAA/zmq3vLPk9D9vxo3yQX/wLKTZXnvHeNvjqKgoEFoTxtMTe+dCth
9U30hA57+A3x4RMjwp7b4CjEYdAw87IJcB12qBnDKoHNDlLbUOBm6fF4ww8ojKzB
07UCJFBjEsZGlZk7QEQE8HACzTdLvJ282GsfRRJWj6uY3MdW7jGO1e/Gb+IJdKDM
n5HDIIk7kBDlMWvblFG0GUJUBa0pRssAsTucAUh8petLkjjUg37EkXtqgOPabS+6
z4j77eE1mKJtm1J1ecrrytPf5GUzrPhU6hboMbDVjC2GhPFCGUBavwcC8pNK1oqc
x6KIwm3ajP5R5704U0ojUx4F16xzMeah4/p6kanv+kuHuwVlzSfnuD//4llKbFPz
xkdZ9ICEjrXHACIquH7NAQ7Py9TiS62YVUvyTYYAzng7uYicezGvf1QnVRUYbOvC
BRKH1IBgRnQkWSRe4sRFAJj7rbTE1HIqi2RZ1r2vZNCBN7ETvj+dyE7jx9VxcAOM
fOULe4lOyhfhv8hVidKd+1SNOcpvcA1ED62AZ5m+7vLLtOtQqQIKRWV8zFIGdgzx
1UEW5roA4QJ22mWQyg4iYJYdhUQTObiYPP1OEqNthjNQQAjykxIJC0oDjAyj0Snz
/P/iupu3yVQk802KRkiAXZSjnvXpQ+pd+ZPcHpPzz2hRyPNFhaMFz7EwKyRh09Vd
xk1G5Pn8D3L0obn323dkORXL8k+/qiU14vS/CQRZUFuHy7GNoLfxYlj8ToQowFrq
0KxKrMrNrNdZaHzViSCBbMdoAuf/3sE9Cw0gjDrihNDHMiXtko9l48M4Fg09Wckl
EJTb3FOOq5cK2lx3KQhM1tnZbhQrDw67CLUmYp56SaikJ3VHhcqYuqGu5uzAIMmO
eaWBoVpe+BbphLxtnC89QPMh7lE00RhIsyGdSlTEzmLCANJu7gm4PmDNnDfty+D7
fgBJQwkKtQZiKrdMxc/j9NoIKiIKxOInLB5CSNzc8JYghQ9qcB2W0oEpeU/GilJh
B0XVnwI3Ha64R0Ue7iig5J5Y7Y3sdAa8A3Q3jmko6EiE8zxVJ41y9ynDvXNoCcSg
WSPShZxDzTW2tTUbQtzTtcBSRTxlyDaXzZqJDhAjCNQocB2F1BvRyixPutlOgBV8
NAJuuD97JRdm3kO8rGz6RwcZVLj8b1GyFJ5i06m3QUhHbOi19VP921+4sbe7UJMZ
aZkkfqWPDASIReTuRxKESqEXRVEROtklm7oNQM79K9GPg4sQ6bbeYgJpmpWouNsL
JnosO4GV4umg7Lysh1eK7EU8xtZ72sS9e2c05aG0wiHoiODujQoOqQLSf+gbwKFd
Dblnnhgc6c4kd30S/Qqe/gOERPY0xzTpVe7tjgmSrTvQP5Ry8ndngtfYY9y9j/6t
WFab71V/NdW+Fw2zhVBDXgmTdxOOgw5cRKi3evjVM1ago4R5GWlD88jQzZx7brzD
+ICC52Kc380I9/tds2AB2nvj/sovreVLUI1M3suKoweFfoT1e1vBe1TZ6Vunr5bP
mGRITj1E2UZd3ywxqPqhT2Ij4um57A3eLjiwBM+nsRvSOgaGPd82AvbnUDWndULu
mVWncMQrN7DnWbUUhFnkRVL4CPmHMc/6iHW8s648GOuWXGhKwnkrvB/P35l+cP6E
cSBbM6X3Y/CvJroiUr+9nmEFbtF5belwFHabb5C8BC4uk+Ow6Xon4cbVb2d4pflW
rOX4S+uaAW0hdAZShcgf3xH5/vmbJz5sf143Hd6r6EE4x46/nyZLjoLcuPC6HRCQ
NmN3e1DyQRB5jaZdu+L5Dt8mGz0YHcRMx1WVp2lZDRBu41ZPscumTA/yZXfmLFyf
JUK3kSlaeCUDhgn+eX3zlYL84Ve8gN8PYcludZ22+LNj13mx5ILNp3GfYRGEpcq4
fAcGG1Jivm+E9KUC3IahZEEO68OIaMzpyarUzIHGqxw676fo2E5z3UsuWSQjBGiZ
xraNO2eqS6ODqAJkzZLBDKYqsdHTdyrVMnuceUcck1HuJDk89yRC8SNJ9wzZlcD1
P0s+L/uEBEBloxIosDE1R1oU6iqrdOMPDwmm6VnRCffubmJtw2Qro3D61Ht5jiRf
GV1oOos1Te9U4zM5aTg61vbkk0PgJEdM9WPzhxsqdYJ+fggx/mzYz2oJ5jKe30oR
CsNp5ffJYcdelZe4g5ZkRzLjPHGkMjRS8LtqrgfSUBDfxJ/7AzH8vih7JDvOaGN9
sr3GuaM85HZe7/ytwDA34R0h7ICn81a7i7GOElYmh358CUrfiaSc0OBQK3BpMMcE
O5y2y7W1N3SVgA+wcmc/iN5tabsEwOvX0HQHqddT1t/3/ONKpDJUIFVr5e0T5SVi
xSg8trrQuqW8nzDi1FxRoBwblal2A81b8xkY6tQKo654F51pn+MYHc3GX/lMM9/R
SvJPa3Siw1sgsjovM3mUaV+nHNvYHnu8wtTlxWP5H/iaqk2BlbPF54MR7P0PsUm2
95NXFkA4pF0hutjow6cJcRmpna/X7IbmiX891+3mp7Aur1Nt83nKI3JwI+F9LDfg
E0PWOMVFtOOn52+j9iGKZckuFrFM3uPqUGswBVdFYydusS8FalsoYFU7zwNTPy4h
QHHcW8JMxwWT8FXq04L+6927sCRl9EYhsF6Y2bIe1Dbltx75lIOpjbiy9nAaJLVB
qQl7f4CMwoWUpAItbaULoMk5G1/bdT8vm+gRgLGvBF48qvJP1q/PCo6zcOxdB1OX
aCRWI9QYB+u2zzMLagiSJtvp5UOtWK5hFhTl/ipJJIo50cQIKkQcDC6B2+cbUieH
ZPjGqg8cMi5tHAW6lsSB3RRfZlo6NWNzNURB0bsL+MxGso2ztrvPuqHnw7hGbY0t
ZM8f50Cbo0K7Jjhvo4+4SEJdOdFC/skPKtLhxPnlcgkVG1Za3ae/nFeYjm8fWSSg
cS+yNMi9vl7+irpOsqrR2VAkNvYhR/vTfDjWVF7DIJ0KaTRFoF6oVmFIakjwRsI0
urxD8oycQlBX+EwDG6B1pio1CGNWozxfITtDu0jCDtJX7nCldl1HhtV4ziYsy8rx
S0yzQsm4RNGVpNZQCn4Vj9OclEOFnTzy99AoS9pheuA/qGMR+wKpt4W31dR17bQN
5OkWMBnodQdpUA/2vIcs4RgqU2nIcC6CxgXacwfbPAXfaqjdTnQN7CES9i9OLVEZ
2pSO1fzEZ3jYFHydia4U53PG43582XEj5YqONXZUQKY2HBA0IDmTpKeqB9wZNag+
0jT924uQWgWD58zufXAzOrISVLT4GlPWsty75oBepbaz6Aebr7eRVjjRIv51+7GS
I6aKva+qASTdfr7uhBeGaefx36SqUV/+jxw+1dZhxnCifD/wrG9CyJL7ois3MY8P
rzTE2+webOaVHLmBHyBe0RatoWCf+3CwIoYMpq/P9RlaQZjNON6qAH05hPT8UA/r
xeTjIBA+2dMrjIr7pxIxb7JM2o0vOqKCfWn8VVPJ5O/cAC+VrDT0iCqFqxGnIB6Y
fUr62FcMdjSTBA2vrFo2ZP4NM/zo8dJAZj41h8FrRihkJ8dGioiV5CT/b9YDwDOd
nM6+lW72UDhFQzXyCfCO8SIZpBA0CT0HRWIL62yx/MkxgVcDztbA9YvWyhoNiHDj
Bqp6VeylAZZAKGcsgzRSEJL6RirF0AYBM4fgadm4tln58LPVHLv5ht+HhuxOS+4R
DqO8d6DX67fPWHIBgrE2/5UewdfCQ8i+P3Qbx4I/X7TaFoYH7uoeIto42ve4Kyiu
KpVfryc/BrVlvCf8f7crkz55k56YpAOQ3AmgAga2v+RtkLVLhUfgIYqvKj0fS3eA
6zeVf3PN3g3GSStbfqlQjqGKdqv7E4KoFMLrgdH0a/skaD5MF3aD4g6tYKNlZG/o
OeGsFsUDxiwPbo8YZPaD0nRzDeXXe1jnX9tBUYCqMbKX3nR1rkSNPjrgXFIVHDhe
NIDRkmfVCON5XD5kU22HXmknwY0589OplfWduASaS5G0u4AxJ9q9hWoyZckCf/Mc
lB0tdFC3i4PWDxPDqk1Xmsee7RMccsB8mVfewsF26hT7VN3/dQ2nJnI9H84e807X
yHC0qKX1I364cAdxP81KLiS+X8QPOcvcGea5J3LrcP0oKPXiKe9z8BZ7Z6JsKIWW
A1TOLN7SdkcYvXXOQIJM1PClLKg6MFh/ggMxxIPrtpV+SMNLwUEONR7YFnCbw/Ui
+8XaRu1D6zPRyz9xiI4us53IUHC/lRc5d/m09KM17hbQm6VCNwK/t/hKE/YK0Io/
y1lYwL6x1ZT0qtt48hQ5duqTTg4NIE87L+k78ofXBnG/bdKJcHQigH8awmu/Pkmu
U0wfVRfSwPpG7GPiN7+QfVqSedUnDc2jzvHwA9wZIAKiS9eP85trdPpNExgCKNxQ
ARHHHgrdD1DOHBxOPbFfkxlKdOAA59yz7UC5N5/jmNhueU7VPOFVNnVtMnBwCO8F
kCWNO6KcnwCg0hayoSkXyQPEPSRXBoXcpbi/mr8/XYOlx6vzfSxfaul/PgGnxLKc
/uXL8CFoqW5vJGpXWi1yP++WsArAeBqCETXEj6bBTpswOM6AwIzWIGYqTe/GXq4M
Vj3J5ge3wdzE0bMAUQ4YtJtbZjFNq5UuimnxmgypeBzur1v+Da07cC6JIL0WRmBF
c/YXJRFhGyvyC+dqI3VwGTIfqrtLyXl97T5MTwjtcSXjq/Kb9hhAThNzfshH53us
pcMYBA1SA7EjVsLypdfsaE+PC1cjiKm6AK3vClAqr1sytm8yXP0IeHF82+nnqKq1
HghK+4lCSeVXfE9DxN8w8vIBLm35kF8zwegN+jhemt1op/yqXdsZ/uy8z8ufoJPx
/ACzkJ5i4DWXHNQsSA21iPb90URAV4KnJE9+km4C21S+7kgSQy8oPeG6G2wxwvmg
6wTkBIhsV2Gdm57yCigvk9ApyGyWNx4BVIGzY3nBJpLhII56NQyo7ohSA6+H/mhD
uTxgkKhtrKSyvhSxJfoHJUeZFPpnjiqcIgkAW7qR9mXQSDHYuWWN6UNEG4fVrxNu
FSGXPpTnz/dIOu/egTiDg7Ql8zAyeWS4N0FhWp7JbhHCnP/FW6Zj+4nz9HxanMqK
vkUi6HjOWHl2AQ5cD8dClzSDbP7+knxiH9z2+kWf+U+ChsJkcrf4ms3Q76v959Kx
aVMQmKe3NCVmG6RP/LEe4ffDIZMiEHW93l7bt0WAERScOkA4iK1oB46QFYjPtQ6F
JYn7TRnhkgV62OvrAi8HO00Sg3/Cbahu8XAi2urUIIDIxKF7NRlzpqCPp6B6fOwK
lWrZkhFpjb++CprAp0VVlPrTtCLi9HWnyxktRxbunsEDq9Djr2NgRYkRevNTUFBy
0wSQF0JhgJxwbnE6YO6WHdbbLIOjAovz0nVFlqvxOHoS2dyBLxayAej7wTMVvotJ
nI9wsmH/Fp1nZV4jkAnmEa0ld9zqGu8rrqrFQqVQLEP7A47NmXEKr5L+WWz/fbWW
wuiL0LQf5KlzaDAyj66+xFPUgiLtJga0VBmikrmE7Lc7aUtTpAHdoWkyzhw496YS
lXF3cnES0QUHCIln2jpx50RklAMBt+HZOpgWShVd1Wfc77D43jWnOywemB2d/bw5
H/lZSOjC+8kFmANp3t5fUprI8Oc4zthlsE3Oemsn+smj9uh05ubAl9QQchO8OQo/
p+OEQjZXHo3fpIi2xnQ6xz1Sei6+5iqG1HxW3QlUwYUM1HtT+ntoRuFHbTLfx7FU
mceqptqNUwTtt9pFuE1/r7M683ZG7Xiikab13INJcknnyLrkW40n/Ol/zEkv7Ukg
q0IsQBmZH3nncaIk9O8n5Z5ZzTLsfRNpue+cHnWXtZfUBzIZuP2YqVWt/sC9eZVX
0sCrEYhyS/vvMXObAmk28n7B4bojqfH3PZupl3TVnNayIt0Qy8Xnczleeeaa4YLQ
q4FxyqWHrUaAvuKAC0ijmUUxb/RXJnhvUi6wBNn5/ahyrjv0WcC8nf8p+mwSGyXm
vnNqC5q/Y7wNk9uHjyJq5mVaRCrxbrum0XeiSPEtkZ3Cne5qEf4jSbK2WfKKTqf5
uJ9eRZz6fW7PHrD/nPIjNU8IbaXkwRcLcMPdgQEjFsRMAzfqcKXQndJ3WxVRm4HP
06LmW9lQfOKsRcc1JqwKVK0IayUQTf2CEldkPfacVy/sICrUcUeFP5FdstmEtmvH
Ge9mQnUtHV9NubgD6Oq81/Zh16O3C7SgE7t7l+Yrk4oef8Y570u874Nchd8zfs/L
h6MD6Mug0iA9TsSNKuS2k1ppyyRVv4qxrikiudLUgNON2rT2Gk2j1KxyRpk8Iqsu
UXnFIw/GbrYLmbrfq6zii1RyUaC8Fll7xsW+sd4/MLZpebk72Jb0lXBhzTxYsLly
7YW5CHhHZQkQ03zl8MZmEnlRIgdXMqpyAROoeIj8hqO3rIioE4yzlNMrZ7AL0Lrd
0rtrw5n1eiVRqtsRwAH557f7rL9/34qFvgNaOqinBSFZ1bJFV2bh4IrS15LRF1h5
Szk+NcdCGY8MT2EnwU3W3cAtr6uTcQxIkTbAFVMmtjPT7osKgf3LSaRPDEWfvRgU
YSK3MgJWVHB5SC4YvS+wmBo4qVIKS9yYMp+ZUaDDrDnRbHvJlDOGmn92Fbrg9JwO
/cys8NRWNcCsN6ZPcPn8dEoGRF9VYsX+bJBxMwI1z8kfC53UgGYwaxn626dd6ur+
PtEx49usE/zHp4b/d9SP+J+NQLkRklzI5Q2ha+NxaiDgE6/dS/7m1oDrx+qvKxW2
ztuPTeaC/tjiVrLoOib9mNqDSfpPGD/P+IuZZCbYYTwN7tqSh6wCo2ZmN5nB6URc
JxxjOTdlGPo0tiILrDx9i5WgxLdF9iXhh5Y/j42ReZRLPcMAUJYvU7Q09FB+q9ni
DhmOGnfEyodaI3OYuBtGLVMCPaTsJtOwcygfqCHryCf2j3paW30kb7qOuHUy65Ie
S2GLfT9QN2/793+tSHeTkgrIIW51UgyG4OfeLfPkzjNlmOqe1ptFbx+La/53yEyW
gre+noe8/fzC0x33gQabNIF6pQlzPrUWB5GqZqJJpeXUNxRtAwaKbsb0Er8y3krD
Lg99YzGnLj+TXfwt245x0OWKzc5nxsHKIu/fOGE/UFqmQP2fplRBXlJ1DbLFDofs
OQRLBxeZaaeCopPcKOx3xYKKxoZQ6uU9lVPXkH9EFy6y+JTRMDRh0IgNKvhCvsWX
6zvuXdeuPQM0qUA1utmyDjvp8/K72Pxs5P9f3kyoJ8Q69HwolFMUFYyZYoEcVTjF
3+dEzErTeCluXPWXAMNu6CwQYYc/1wkvk7lcd9XTkZeSLv/nNKNMFi2JNM6c2YEj
BLFJgsrMYyiJIqfyqj+rPTlXmK1eFd30MSvqDk4sxxfV+oBn3N/lnED20VBbAjH5
clT+Xyd1i7mvTDSk1L1rMpo7zANTCpdIPr183yextfANTy4znLwVGUNxEzF/chAY
TP/CTRpzPhsihB2qbkaBcb7V86s1Wridgcc3eHjo7zPAzF9Dh9BRWLydpi3/mZy2
DITmyZxDEpD5Mo4iL6Rhy4XGao1+QrTFZCYkepp+dOCCeuWZoPuGiZQi7EuB1V43
/HgDG1gPMdEhyvjz0LckMldYzDGdGxkVDF7ZrQsT6zaY2HfFEJcj4FEXdnft8f90
0Hxnjd2+riPEb/KJv1MuqWnU2fRWn9EBOlU+ilgUvb2q0/6XI5EykR2llLFFsfwH
2eosvZhQpR1A2wF49dgny4S7bXPzkYmzv6aL9kMYwvVfCfBLz46FCO2mkSCxZB0y
MlS5qohmWX+84UOkemE+pnOi8nKG14LhI3ZfR2nkm1cK+8ctWY+6ZPFbJa6S5T/F
B0Y0ucfRW9uvn/e1nO4j01Aa/uqti70ZQyMTnxuWbyZhrg27ELJ76+g1Z0prBYXM
vvGVsO6hAdus5nLRrTsK2kX/WmIy+gOu0VWfs4eSo/QDA7tsfHEjxjzGitMdUexT
FXGCd25wRRNkrJR4YpOqWmeLjW2bwWT5maEsR/J5tethhY0EP0HZO6tZc4C0ZXgP
qe+sU8WF/c8Db7qmg3elpttIDZe7+L89tAr2adfvz2pe/Jm6LJq8wevpa1nyZs+q
rapzYFq1E9tDkPUX4T+hUguJ233/wxzzfecYncPvP4831kwqjjkhB1lKXA4HUTgu
1Da7p8SFjulsfmzQERXJ8zviHxA1t0hLsLJh/GvAVHseq/YcaPCaUvhoUho/ZzvH
y55TnCctrKIaYG/82Quf+DEcwoeZGa6Pz+j1cq6Bev0C/eKkUav+wWZB6tFi7E4O
MwqBvYz3YV1VMbzUt1nMZWSiuP9eoi7LyNEf1fJ6agqaGVFm/SgE8IIOzA+bFX/7
vLkE0US2j77/pwXTGwrdPo8/515uOxUykmx1pJU8aV8I1vPwrEi/WmpoxS85qn4l
Y6N5dDGVR8Hz9kd+rt2xSNnv5fzjYqkw6+teD5MOzkSEB6dNDes2UrmQebvTiWwQ
Ly1AGHxa5O1cEznNELnjy6tP5yPmv9sX3cy9dIS7bJLMF8jTHuN2xAUh+mFxXtzi
Ji1rzPm0R4V+tHN46YReaaB7shsvlHBUbJY+UZRKYIQENmCn2E2IZSwdSEspFVM2
T2KR4TZIWxwomLFSXc2Vocv91sfVECMsk7GEMmCLRDTY6CK/oMftxwk/Q65HKi8r
wBvO9wtOGSofiutsUuzVa7O4jw2vUE6pXkDxwsxzq6xe3pj/4DoZshuoVi3ahkP8
0DBEMKlUvui9L5gQfmKjlOrhJILmouw3nSzxHpcXkkDVb+S4haH/kgaru6meYLvU
/fxB1Jo1jfetF2qRnZn5RRAuYTLEB2dYd2TYpCxkm4gsWbzDyaZsE8n/0EB+nvrY
Cs6lmYNYIS0awIDovGgG8y5K9Z3ULGOmXmABPfF4rMmtQcwLmWY6GNvq/bmoAyb3
Orhg2mdc5X4o1N9xu7GwR6J9bNZNrZyDDuRRuk7CXICvlLkO8k939PdjG+5xLxE/
+XL24X9Fi6uju5QXWd4z3TvtGHqxyZEhvOg3o5wRMT7T5xqgxNh5DhO0qKjsFTpR
3YIXphU2PAUcsT/uF+ptOLES1EU+inZg9+Py4IkeKJ165lFKiu6KroQBQQs6+fOC
dLDA+2Tdrq0PtKR0HHwMsrYrNK1XBV5QMo2Hj0rb//hhfv0hKAIYpD5EM5b1TKW0
QQoPpmnher3XDLEu3rb+d0lRvrCdhL9wj55AeulM6JwOj0iQ5JGVMdWqVmM+VjVT
GMYYBO7sZR5BTMUOduQObuIeFOekWIaeAKwarZcACb9KCwFsp5LRF3AvxToEgmuG
/98Bql3OYsmieGRwc2qsQYSrHsiSZ2EJFYr4iKN9YtnWmJI22r2nXiok0luGwSj5
CAlGA6WzUW0aAYktguKZYC5L1NBLsMolHtQKppEUDooNNcf0z2qKSn6Ia9aF1RQ1
FVNMTZJqcAZWFT4qxRaejlEQbhkPHZhDD2YHdDLccfLYcW4KTMP3rg8KA4/JQA+N
KkO+6xc2Llybko1rP0w1Prlo5PuZNAy2WPuERNm2IeBVLQLad34VdGCvHHSqWWzS
AdTGeoo7hyNHsyybndpe4EYsGo0ltZ1x+BX6ue0UeFQ5OVLm4yNPfCO3pz7cJeb5
pT0MJfQ++n9hJkC0ZK0/GAqwhesYfwO69WiUW3wHqCn8YL1QIv9AzPDKhuUxErH8
BbjLesqdaKr3XPK6zucn7Yk4IT/JWEniFTh7zROE+goMJEY6DSQJGcSQ3pxeoz2j
zZrcwOXBQ1eciLAG13/83hsl16kVcbnNCPBmxJ3o/+/xVgIGXhYphzv7WizkVN24
RjKx9CtJa0IWt3V4xIAZSKg45tAj40yLVcJhbf0oUJ5+NNc9NIPDgPlckMwCtGWe
m8buSjdvpu7Xi/agIT3PRkHEs9j9+rDfVwbNS2LfnhH15afEhYQOCy8PPfVUX4QW
Q9yPhWdn5hScC4TheCGdJDKDeeSnxz7C7k9K7qw0dPXRmIu0D8bIvnezA6rGjARy
zOYSEFGNNnzevjvd4eSjWQZwfH65rGfoG8QO1veGswoKXNsLbu7s4lLAqfhJdPCm
/khlols0SdGofYgiL+vwQ5W5YHxl4q2k75Trl1MTY6NBUOEUserL99eTLKcLs0yp
OoP93vIR/lSp1qua2FZ81/w2qitvHudITRklNPGCQC0R/OnKAA9aAigeGRtmcREg
Mn6q2T12X3naeXNk8ciCb1HQpTNRazrdrNpoKXhpWS0XBg/MEkorR6hOBSzwHGUE
zxR9J3aAA5JsbsYRZBPwUwfWS1pK19l6oMvZdDaJXkTeYYkWTpxSPFnf1dduFLLn
Gao+hTKUQEu45hefxIKZEqUQG2MTzWa8yTWukbiOVZeZA8mEM+2h1eUsK1hZ8K9C
ogvvceJWzSaR4B6NOrEO8UwmS1c62jVx4VMcPxcLPrPYSNkEwuKuqUfpNFW/dWn6
urA6MWNJcV8Y+7NiDguoJlUlonYQpx0G83N2CyjHb9xcbw1yUKLxpU8KazQOa5qg
1ylI1QqQsdX+Mw4m7STm/TjwoJj0JxnEv0F9wLD3ae7kv0GLRFRwOntnnp636oif
NKFvSKGawdu4IAFpkx0cnFGWukBIdVx48qqS1+Nd5fxsyY48LCetZDA8BaSY/bUN
HDOR7FOWHGXd0F25bzUYFSd/4Oek5HkpTgBONkAq5WR49dfNsMzLf7oJ4Va4LaEa
Hu7ZmPxXErZysHQ/azT/1qNYOwjwQ+/fPW9o+fQIQaP4L48X4SzszyFUQtTSUaLp
Sqc3eEVNs3w1wdLPXNRTUBFoSzO2U8v4kmtBuQ27Dun3pPvrVP3yV5ybajZM0W6z
AjWtjWJaOI0SUcThYwVnJbAsUtVURCcrq8GTXiXji5Ni4f7yIzMp4QgapSLyxvd2
+JS+I5dOmR87tzoVp9WPH4hZFDy25V3jI7uEOeypuXlgMx1zl1/apHBmVaJ1f4yE
TWWqXrzdDppsmXOPTWzMsc90j4GUPR+kz7JGc41Ny3bMJHWYEiJ9nExKvN20nbz8
77CCArZKTrQmTl/2mJOmuBRcGyTjMddRCMpxXGmfTV95UzYzhVjtyIlE87svcLCY
v0wPgnDcaAm4wVt718Ph3gjrTIrQzlZqDBxreAepcg3j6Fv70GWz8LVcKzYQNa7r
+n/Py3u0URCHQuXfeL8qh7E44ZXggffxeoMgjhIFp+oVyJmtLLRoZ/ZS3jNd+70j
IrUphI9tHcv7Koccjn1KPapG2iOIuRoHstuVLwQxVZumUogUoQ8PbJyWzRKNcwTV
TNqAUVP6YJjca6pSQYXhkma5OyCuIDoMKLaGZD0c5wMSWRg5wD2ATR/+JuuYxpWd
c7OCiZ52nsXfI/oXvFWrFjPd9PbExyZ15sL0fiM7Dv3Nl+dQhklZ6RR0k0PkbW5C
m+j14dxPdMJ5DOkisYVr9887/gmcEQbX3ylXGny6jAZ0En0lG5M0Bqe+xL3bdC3n
+hwcOGd/5/NsMHEWLYnXqtHecZ6Y1+m2B1gfWCf2y7t/IGoCg6s2RkNmReiz63mn
oyPzDLTcaxCPv75O+Bc2hiTwTae9PEidsJW30OUW04GLIQtl0s+4bo6JC0i7+gVT
8Ng9zVCZW1UNXtOPonSbwEjLI0tcpoRrpC5+Q8O5/zHYNucy3WMi6y5Dn+L1ppuO
/q+5V3R3CfRmXojfY1c1b2SCHVk6GU3p1yyP8Hx+HsEKZF60o2gOCqHvSek2IU93
5KuioTrtblqa0MIO5b7/3czNulCgv0Z6ZQVVmi1UPwJsIkZpJ5P99dURQe3mxgx8
QUMx+7mjMm1wIBVDOYAuZcqskKbBP2eSHuYD4W0PsUg7+bx68ir2wEmiya96LCT3
i6kaLZgGwJixEGtWMBPcRWL42qYEj/ddqZV8+jVdU7aKXEbW20EonSu5SzoV0rym
MLtKPPXdDjzI4yQCU/Bnn8A2e2etGRM+wkjr1McTOYUVjAKrmDILRoLkMSesynoJ
U3F/YapWHnza4P9f4vJKlKZ3Qlg4VhDy+ZhLoNa3ZFdqbkFUW1cGWW4hbM0et27A
imRtN8VxCHc412xkLLZffCpLu4Fp5CP/vGOnHKY2CoExTotZm3nj+JZdxezPrDWm
xkgUDoLzg/Kp7ydN4YF7UfXady3uOT+CUB9vr+tqVluwbDkB9Gkpe7QCmvJExFTF
x0apMAhHJsh4RmpZkUQb27Pd1FJN/nRd6KX+pL3J+71h7jZ/Z5BfJ9eCnLQhpwmj
X7mNbrBo2KmtLgV4Twqrie/RlaRXZ6VilOn6rR/4hQ0EeQ78V79bKJpEJM1SZyIv
d06YrY2U1gzNz5S86DGmeYYHirkFey7b5akWS5C/XedxJLY+alhsLWu1dyD/bYYo
YJBVFqCujRPu5eQMXs85qcoULdIH8tS4/ZcVu+SQ2rOVMLsWp7BR9gstu5Rkpdql
2IE7XYfAw7qrxNv6f3STNIhQK0pSyWSvi1VSyZNtmV0EzB1PZA/nzo3zdCOuCKNj
VM0E7EtZE44kNz6IpOjYeWWExqNS0eAj4knexvzDBhGTlUrvcWkRnmTIOTT4bASv
XfcYT20LgXlezz2wsb4CO2Yu7quRnxKo2/CRq0O+MczUS8Frr4tzjVwvWsGNgCiP
LdYwVoJsqV/Xkv2vME2PCXSwQeEXklxdBSVCDXYTyYV+bcAu+LxmPdBYnpEYJ8uS
HxhKHdCUdiawmFEYPQsX0U7hjc9Lchusd3/1N0R4sEuulcJeFRobnaZbHTReEke2
TYP+SBIsyTB0FS2gXNJt7O/1265yl10Yeb/VaBIicB290sabK2aow9dVQ6YLZXem
aEOWaBsoglwWtV4gRQ8MdmDnKR9+h4Vq6Ltj3ctJYrRESaOCm+7dHC9l4/2Vv6z6
c3WprPrd9aA3Wa+8z4OwhfbrWHzjf2RBkQUMfe3KIeJgzZxPytlgGmhY2aSKUnKt
bN8pCwHu0hPMRLNe4qzMLvVsHqg9Oa4Ncg7TOkI4SwkDYSxdQ0ztlPGaY8Q/Bg5K
qaaG0ZK0vsigs9CcA9rDQlfTs+MwKxZIRFI2U5W8caMuohzx38kh0FRHllOce47u
wBT9eDan+l/UjM/bXilgW2Lt37ADQxz7z9Z/UYwX7E5xipv+1fliVpU32B5T6kqq
qIioo07xPqMuWLOJFijsDg30R7/n3ej14Krxi/Sj3nxHb69NjbLut3JwEqqPFn5k
AJ3v4dUpGkud/bL9PkjtGjEgd8ZpWPlGdrpi5xSHyUcvgCSIryzjTmkpezOUYNX1
KSLifdSNygZWJmn6E/WM1BLma7NXvrFohRiUsRNEkWHC1FiQw4SFAFarX/xXVo5G
nWssB6tE6+D7wg0/qKo3q2tZou0MYR9A81sKhs1/QVAf4ji7LCKQbPh/FwG4NfnD
kuFzq6JSZpgeFxcZvYUiAjSUaDVBTdD+rmiD1n13qHz4K8i8R45gMyVGB2dYaxYn
hBH7sU4h/oqi019C0EOOt9IHjF3PQXdLdiIMJwrHJCBNoUEJ2VuS2D1wc5k5UQK3
BeTZA4otCJYIlf9xu2+giZkSCM2RUjWmve/LriP05NU6shXev4QAZoTH9gmZLlfD
vb6d39JMWFFOwyr4RMdRLZ5/3hTAyCZUAawy8vAB6KCoI63aEqzbSw/7Iah0zb2c
Nh6PMfQnykxIZ4Isgj10LZat+ewR49PWWsoNE6zNL670Sd5bYysYYeU3uyHK6Att
lywFGC72Qo70sTUrxjBBjJoBtIwk/+k3dRHVf9zkAJEUwFfPbjF90BTzFdBlXtwY
ppYIp6KdfSV47BYY2Ba4AW+2vQyTdkXRtPd7m7P01KDiwPJPd3215Mw0lVdsCI19
Lwi8cvjIPOhn81ST/jcPvTWHxTrlT2fRUUpN8oj/u9DJyqgR8hA9peZKiJx6Hncn
KiRxarU/33AXdwwpwnLlol0TKKam182bhEmmnRCwxI1E9Cop2yKKohfn47/spVPI
zxXg74bqN75UbpI0Q5KzcanC4APovPuZeeRxmmup7Dj7hvfN2k1Lq3yeSHOUtwtq
+AwFTrHDCU3MnuUhtduJfb4z4LqlqA71MP3SPsz8troMUOAp8AI4CdPPbfuPix84
W53rh2kVhwH9Enl3XCRkzdDDdeTIcM9XgnhRoncuYFCj/DUeFXQaDoFTxGsXRN98
C7xODwphvXemdh6grkqPs1HY6liphIg4zmY4Q3+o9K7smamkXzIniRHqhBHhLBYt
1zIcp4Z18xFNMnIcgVnRwmNd+UANs6I0geqo6mA1PKP0MNU/U+xm/z4UbMiIffe7
t/llvS1nj1PyRkRSJfBlkNVbsdauoLHokKwxajAEu8MlNu178mnMF1139LINSW9E
hQBzXR7eaG1BYIL66foFDxVEdNzIwJa2/SwcWU6pbwTfH/z/sIZlfeZNgNJKslyh
IChPqTTmS5VM3/YaXOiaktbfn0EfsSiLq1UTwkwwv8yATjYvZTtvR8w2gqp2GmTs
yvLq2ptmblcs+ZTqNx7RPGWKT7R5WI+SaqxmnmBJYfX35MsUJK9gJTcOuSdqoZnu
cKY86ZJgbLQhLmKI306Yz9wObI8+cOo8EPp9rDmOilvQ9gnTVCJ98TrchWOREpB8
okn8StppCoHRMhS3DfmMypAIPzVmO07K7JSroSGExgn2yQKBYy2jjIA04D1FyFk6
qGNwBkHTdAB0hodIwOPZ4e7tcRq3tyA0KYJQuDI4mpKmHcwM7889MFGx7TzDhbRr
PHn234TFXVaUdB5e5Sov5pdAjnVUanZdhDgTDLh/LbU5pjJAfIPeXLgKGL5cpQrZ
GY5yujz5lnvVaLDtDQSBbEVUf7U5+YTJdnL14omUkH3fxGQoyLwKfNrDnHNhb9oZ
XvIQbIk5UlUiA7Dl00vuPadDmVr6tHA0nmAcXoL8/Xt0WGHOl9pyYd4a2psCm5C6
iuzXWq2xF/vQIVy6+iXlJD07MF5BxrRLZwvTRGtDr7NsdVh4e9FH6RHe3pfbCuVi
s1/uGF/1LJD4SpYyDXTlngXiWtHOzKhPb3Rioosu8eR19fESdoMVEP/8gJ98J3xS
+tyPint08YRHY26lQeoEGH9d1KoLrGxKI6PaOyLrR6J92BYDm/sZ30lbEXqFKPYG
oAKogGgB/h8p72XfGYBLf/DSWicQe/odJffvfYyXnpJvaaSsBZvCIsiOlquXKHdU
oxzkgF6p5PcRs0J71sKjdDFhynad+VTW0wdC3XBdrI0CjNzi8jRDdhSqOHMCsyZs
QmdgARxKHyGTUcDcpqdz7PhPqbU913WRGwNf+O4i7CnOC0xFOKxXa+BN+UwtHd5g
fUCKsDDD9ZUP4zavzgFVSj7AcTJCgkO1kfGzMoab0N+kDiwmUd0inC7W4f9klk3y
roeXYumUa7N/DCEA2jUoUwPrtGeLBtD7W4UhoihTxi99kaqKrLjTGMjiQVmr/XOw
ai4b+r2WXvCN24zTafAh0SsgZE/P/p1tA8X69XpHu3SZqfDlkrRW2M9q5pc8kBfQ
RPyZNlZ3CNC7kfW6hYzvszQzejlZRQODV2au6JW9AtoeFtFsky+s46MXTtsY1htW
uyxE2buIDWe3//g5neYyUbr5G4Nd6hNwiHx6KsC6MJbwCn9rIaspsVw7W0Ga4DWj
2HvEOp4WpJ5cUtSh3wvz1gI2VDbHiK5rSubCiSaHHsaCoXCyPf7pIrHtCvriPZya
9vFAvc6CrDXAe8A5v8MEUlCdDtp6cS9fN3AGBREjERVE/IzGv+C0E9JcQFW4kKM2
yjQhTGXaHQg9l3kOfxFBM8kpDfW6aygsXtzq+Pil8j7r/C2vEJe1gYoO8PN/DLwu
mPl9xgK2fTPQcbhZqjDL8SDfPgQrBvkokMWdsYKQPSB0DcWgfEBErd/Iru+6grGF
PpxuBexLLj3VfzJvRq41OlETrqux2UBx8FtrFEwz1+Ebg5sttLmGSOQZwh5WBs2C
410ppATQN1WTLtYExfNa69fzsVl/yoqjYufKTZ8k+R6oerl2J6RVpNCnl/E4wFzP
aEZ7kaIDHhM3J+6tOEnQE/EjkjFNQXFkab3ljRz9dmhpl00tfhw/dy9LHoAm7wB/
NcyzVec7JTxkIdAJjGhFKC7nQPNVL2HoUgf3ZnEAXf05+r+opYArPao/mObyxFO8
MNdSJzYxHA9Hr7LX3XE+/FMLeM4mdq9RVfkp/9Xfv1t+620RuxIDaZ8bd9gJfFOX
uLQmXd2GpPlL7/dRRy1f43vHAxbT9IqKQUmuAplNqVKXoa8raOY9gv/zWb2ZRZ3o
fa/MtQvvJg1CklI5/W5uNJQlSLRZRFGuarf3DkmWGN/VuZW9x08iPSAY1mccordS
y7fsuS2JuGQTbygT6kqQb/lF1vex4hqOM1FyQ3VsKGuEGQxJBYpQRag2oOMfo9eH
2mx1rvAUys7rukhapcqjgUMKcu08ZEkVjUqVVd+RlWmyKu+kwfi726GWvXlZApLF
vtGGy9Du9ttgwiafc60bE5bgaBeoLN8Yx1npBRU/V/qRrGXcDfHHBM+vE8X6b+V5
In7M+Sn1tPpKZRrarFG/ovHFP/WsW1u1b1cB+UHveHV9xWk7bu3wjgQnwybBp3tA
w/IoBMNepSeGZv5cgbtSAAfA7mdI0nQmzkqmiCx6ctwIyn/hzUx9wAjMd2r6AQLQ
OT3egFZJDqvLQcskVv844nuIhDLejGtCg/NjrHRRfDZ6+AzjPDt4hJ6QmFzY6ji6
oJMLA58Bba9Z0bIE6BlZKg0YQcYMYwmYiA5RM02I9qQhVKj+DH1AzZLtP0gpojh0
ezNekBGf7SVVlfGivVwqMXvn/dfjCWtPk2pXm01H3yCKlMsDyMxOJK4ksT28niLi
VJSa3QB9A0hfM0jAee30NedpzQPgiUCYC/ZEs2eJMzhe9tRa4MRKdQVl1jZQmlIi
2voxGmvottJtw7dIUNRwjmL+46RVP7Ku40qcV6T0fq0WifW9F1rcL5171wEH0fYo
+RTvqhuFo9Nbk5Gyh/lNki7CE+LIuHImnrpEYEllu0tJiUHBq48N1r96KQelcNjB
G6ZCIxFSG7DwYFEe4TXwCF2Qp6ghg4JN8AVnNhrRn2Y+lbt1KoeqizOQpZ0Zsdyi
o/ESHfuUPuLZh74mKp9w6ozJh07ntF4FWnqmki1R0cdhxgFeBaa2DsXwSun9uvhT
AnabHVEUMRzgbW6JweGlPyRR9GLeAqwnCH0ChTZl9ASvqMH3edQKtuKkUDrA79ZP
F/s5GIkKynhO2qz5I7Wy3+X/jOwzvWdZiutKHNE2i99ScMWSwS4tAXqFM8BjrYxp
GzAPgTKDgJjtaP8kQkYVaF654iPwgQrTLS5OvMK7u8GqQplmyCNkec5mt67VhHGf
xufMjHwDZBroFnKrkxIlOExgMUwukllI1FnOje7FyIV5kUNnvBdAvkPo1X3NYTbJ
fSldy9R+lZkwwjqZJ4hmTMvTXGPKxWYTKlGBC0PqFpXfAYSjAUxae2YUbMbP7JvL
qrp+v4uHNN0fQSsmW8n6/FVGb9rYjopG7PwgViwIeUViRfj+s/uyA0rVLUQ4OnDh
nI1Kz4bwlflId8TGKnQ7fVrr0XughgjQR/IQ7fwF0SnpCmA4zK0bBNPg55SNgOPo
eDYHARNKPWQakftEIlij1CDOk72Ion82+W+j/GY843fv8p/ceSy3eyIU/Fmn0Amh
fD/8l5fbeLiluNW91MZZyqOY3glHVDM0Zqv+yDXi250RpEjHh+5OiT99XHi0Dhld
CLQj68dXoDsw7UKVzEG1oD+mcXh2ZLjAolHGwCvB0k3JE4roJRJN1Ib/yZhd/l1v
g6CGX7U6LwUzSq6fkgxVnY3+2WaT/0pmYqSoDNoOKHz9pfnvEed2hMwr6D4hl0H3
65AFe0JXLtU3f77x25OyQ1k+ZzgDiYh+CP0qjSy2x4EyadX0+YIRpu7VZpP1wNQr
dcYr38sLB0RBbicwevgr/ZBvC6jlT/pdLFv7Ifjb+XStX9gpT8tRxD99PFKmZz9Y
odrdAtJkKqGScuWapeffU+Q0ehEstBIG7Dpxo4xT+4BrgnlJfiOTtWdq5uAnQfX5
qOe/wAWtVo/hBKM8TmZYxqosTv2cRQ2nRe8ecl01jQGYE42D28dBsmiCuxZ59eQ6
SHJ4P5cBZNqSqL6AoQbqO5fbJI+BnIc1PFPMbDP/gDLTbpTxfrEm3Zx4zuZv1fAQ
AqDF593XkfEukIQCwM6UBfSEOnWdp3y+kSppR5d9w9UvMbbbYAJ9H+VM5v8cpcGW
Z5YGKEz1Yr2dy8SRU/ZnyPxMiXQsnNeNnidAnZvVhLziZ+GnddtUK2JQWhAbCp77
J1uy4n7/VByVpCzVGZg6aNaXUc2dLwGVePdM3jNMcT0B3IxPnbEEVTEsaRvTgOWS
T2IiOEIq9ioWDK4VT89DZKFXn+GCxSxdhHEuYZFk5eckLeYCy9s3JqbR/v7X3/lB
1ntojEp7QiIMUHF22MToDXQiV8366C6E7A3jH5ct/D2LhGGVxWLDi0dxvXAklRo6
VEcRvAbZsqI7zvX4p7QDfmt/IHQWtDFZMSgNJai92IY2gMqGtKVQSklcrgYVZJWH
uXVQWzFMrF3wMlks53U9/SZRnThE5l5ubNITuObBhT6VnEOa80OBdqNLjmu6sTh7
tYvO2SfoD1maf3kueIMswTeNIHLjT4gyrNVxGRuHCV+T3ARFOC5m+JTlGyNw8BiW
IrB/vgLU/Qrehob4MzTiVYFMfc7YGmqlJpwd6c9rvKNMy3YFFDJHT7fSzGxaMCFZ
+TKzXNbHe9Uh6N5sCmRkApwUzaAfuHXiYLOgPZli1bs2LpiYYhK/cnLAKKrwG8zc
/v8rmgld8X7NHweNcOa2F5mtQkkqftGBX59EsTrM4vWxUHJPTxojWOH2oCEDAdWY
gB1OORtUN/RiAAhqoWPr7lz6y/e67GQ4/FWD0J6VA5l+ERC+0bzmMTJLz0ipANER
GNeBG5vD68phn/cEd84nCEPBzfoqYC2UYt6blayMX2xMx4FU1xqMRBmcKIPXcIof
1fDYphNI0pYlXhU84K8RHXkchQdpUII6zpreKoeS/bVlX8XOBWQKs+3MQ0xemTVB
wxZ68gtm0dfdTsjVWLwyoji06LOLYpYy/iGTmiu0YDsABLWsVD0evUesHvko77YH
FyX85x9LeKofJmDKhlx4Ubi1Bxf2Wy0DYGoq8mzs1IYl22s4ubwsTDiEN+yPts6r
tipVJi5UJzr+Nwef6efwhx6ih6NczipMcoKf5VpY0x9DEtYs18l+RyJpBYgTzeTo
f6WnCI3VMXGTnktT8HFZtCq+ecXZk4wHwQuLRnjMJTkBSuidT4SMjklGetjONl1I
fEn6vc4Ish9PWF8tzpeSz3FTrkV7UoqLuWWxY3zEBnASsvoaheqoHwQwf08NIFJ9
LkeCdUYMaMB2H3YiWkOiM5NaWQuRkFiJylcZB97tmiv4PfTF8AXgUi5fP/VModQO
baNQjDywuUKkwHWGhej/xelAIY1UYNCby7+wzzPU9i0PaYBkBXZY6x0P/NBRr6UM
o5U7AWxiLV9CnTq4ehpML2ysvu5zLlwdEq5nS4793jXWS9eJXYEaJw3uoJvw6Bua
WkbNTwExX5UItCV1FaT/cyaYeQGfYv9xg+LqqWxvwzchdCI8cgmIdAxe5tK9cgu4
0FBh7j8tNJqD9Pi8jZE0e3M3RoAjmWyRFXTWFve8IT5Zf+Vpa5trK8JPG0XIoWOP
M8qwX99CKCcdK1J2yBGwOxCWXQEK2zRx44pa0bdZP9E1n+mXmpk4Mw12AwIsNYY2
RxRky36LSjk/D2UNhktw5HQHlrBn9stnpLBrDSTWY3ajEPSWH1WcVxHzHLgEpPDK
qZbqRmt4lzEpAQOgc2x+iliuVKPEdC7vVoiBi4M+3YlLAxn/cKPb1+dA2R4CN8hl
J9rBLQjzMjldbsesvCOsdFcU8xWJsUbxDDGzkWCm9fcxdvO7zCrRW5b88b8DMZFJ
+iHzxniue//zIJ0xD/d76XfNBJs+gF7jXfIeE0OeawGgisjCO6rDK8pkA5G5ks7P
jizFBZZcHkV8VoHVY81+RF3XS1GW9V6cQYoX0x4V67azpf0UQdLBctJsRAw8DNEa
jHXHb1TWbFdEcJdlqy3yAU2rYxpN+ZS2IWpulSwLiJPTT0Qr+tQ1wzWaygfIjhIZ
lCG0+Fid4b/eD4jC7p+VkR32Uv9hDnPtjMA7MOuX5Y8Kk5z9c66+m57Z3QeuznV0
lkPli9w4uD8IG2RQpSxxvvZ6m6+bFkXSpEhgQyI6MIED/+7G5lAEoHJAtgsHQNiF
MOvYvTL49YdHUkx4iwuOAlbF0PGDQvHgzcF9lXfc/7Wdj/xk51ZYLAITi5oCr6wW
MCRfEf6N3TBbCQ8elokTbPurFBN+gg9PrsudqJO0Opcte6hgL+jeE3T8d0nbw3bJ
onn0cIJ4nMEAXKsgIG5LwH4w1FA0lCl6ZbxNiQSntVvYlt398drGn9eUXOQ19TQJ
yiTEfBk2qiXi6uFu2b3vxQbNfde4CZT7o6SoduvRqj30k9oAH6mtHdd0+GRf8DZX
5Dw5126MHMLdn9KV49VNlSV/W8G/9fRFazKN4LfMuOBCCCoDDt5yBw3fJ2L3x6Ar
TzeukKTVC5RWz2vBDMkVSlz94jZ6lv+uKfQ+Z3VjKv8zUsADCMvY+pxVHTDT3ju+
J6OjvSkniUQ08XrcHmo9IXLygxcu+bNh5naTJSirdjjSBzccRjr7J5hZiZJ+hxRs
UoTjeI9OnrRyO5upgxnevX93g6u0/hSM8TEadVOoVLQOB4/qBUb3DFxZ5xBtOo9f
de3Il5552pKUEf2gXXuAoOxPPsMBPjiA/13D7fXnZSBR6fWx09xjfCXezz09EL5S
IL/bhPJlxacB4RXBC14HerqATPEIhh92CRZf/JLCi9oveVfA7je5wvM34QRsNk85
khOCP7n+XbHLmRM2lLaIlTvJIo5fFJbAQNRwKzLvWpP8PoM8Tc38LzWUcwb9XpRQ
Qq1a2fkv+cObe+tAVowrnO1KDQMvq1sncc4oAlLt4vdqhOkUlSkKyVl6ghz0DDZm
uHZjAuocWkzedhT4sfNmuny12YxVA9Jf3KhtKrcqPBE3ZcFTYkTejBMa3ZXZVDPw
HKZxmT0yFXuF55Qs5Mahq31xcOV0zWYlZRSdAXlSMeaHUIfNvABPUDJmzp+ayGG0
ydDFU6vB7O/+ix2t6gnQ6ekeSX7aCGtUiMh90vWDFaWex5E9cw/9swGq3Cga6WCr
AsEBNogux4sPXP1rhBI4ZV72LZ2ssQfSJhGrrEhBfG6N7EXJ+edPtYfDjimjSDqp
WdAWKZfN42K2Qp5ASQ7lmrqbuN7l/YY4xU4RfcFUeqcx3SkClU3tLJdZnPn37lPR
FHYjoY3vaG2Nr5gkNfdbhX3owD5E8YsNGnTW5EaOu0X59U1hrBG1RV6Tqu6w34gW
XSZtrAboSGQ5vFonlJ17O82GFhViXVkdX7StbrbJt4unI8aze+JX+1XhrHelfpP0
HzwJX0wUgaTStn1a5t51n5YtTOtLmoU6Cwu394z8MA8h0NjfA5Dld+MX1ExPDXyc
OfWmSFspcmhaM1Lbpa9ZWM58YK6GI/MRYGAgZTxmNsaCl14Mtyw7tpoFWokvPL2/
GEl2IIcucQIjBSNW6IMb0g7P+QXxv05tBgbfKhlRAD2TnWJpSJySLsc3tUX7x3g3
MD8bHiCHR/Cc4tjiQwwaQ3L+MzjgOklBiySzxnIoD54Memhwu9ONNRNvby8iVRJg
UEETCMH6XPhrvr16y/dCEkISCaGLxckW28VGenkDCp5VR1SfjzKWLXC3rsKke0zI
mSGDr8K48YENCXzBLey/jXykpiQjs+hyZUzcqKoJvmmIFYCvdFtvFSBLe3a9wKtc
jfV30tRADYP/WYuo/G5OSDXqsB9U1nCWB4lwN2nV7fsUfYtNO5y0HXLJYkRTo6P+
HrW9mVLNnSlfc8COZZsWoyJtYiab2+bOzjcYIl5KInPT3Wma8ri6tK5K/llml053
ut57JJLN7PdWuObE6L2Q9m9sqfHMepIN+0Ssea4aMMkBm0qjalJdO5PSRYDmTYah
fYsiKctkq6hn0rULgqaR1wdYp1WMxqLYSSg6dGURAFqXy20wkaC8CcRt6sfbqZUy
6kyL1h27IvN0Isu2Up6xchNQhBZSiYqfku1NqeHvhwKtssxMSxE5kjEY45Qz79Tg
ztLf4cIMtX8/Oo766fzp8YHAg0acDB0W9/H0hnqUfNPgLO+h3ZjNRJaw9wwUgfnm
ymWQg/qn8aXrx1CxBxvjGfR/+FY8v56jbbXbt42fXlsKb+UfoGvVO7IVAKGyyEej
vkPR0p3gW92ZkHYbhvTZdO7+ga63bcy299DispMBWDSVZah87n9wFrwBkJ3s2m4C
30OchWmicQx0/BfQHvJ7bxOIFCNdSl0E397RVowxe7JTuTTP5hBc6G0RZjWYsYML
3vSsE4uU7gl87h/uLDUYeJ77BcB3Xm7OymoUmsICZzvyHNyvhot/vBnJYiZL4PE8
c39xrUHIVz5YZA8SjKFMuMeIyw1YdAZk6JqGH04vZbnQDTAUDz/To0FtAl++WTd3
EtJ/cK8cI3uAbRf0SPU1c/RPa7kBh/w/Rl2BKDyJ7HEkoKVqGIoG4Ejoqj53W5BT
a4ouL5OaIHWtij9+X6UT2nM9i/R7Gw+ImL33mjCrfEqPr2V/T6UjpDVCCF3FdkuG
9JI0kUVsTHG7b1NdlRi/tANMJzSwzBbQTl9e3BOeJYYzy/TvRUYZx+1nmhLer6j9
QtymRyOPh4ss/er8F9GQexqUIQDlSaXiXVsHSpeZfHirYtMPqYgTAB4+F15ep+3z
dkQdMfv++VOg8ew0hJanOZLVi2HDMMmQeLuUzLYenZLkpW5q0uWECFrslJbUbMqV
BrDBoZ6BMvlXHFXCynasZHmAwXdcxwfAg7jx7FnQVmiHLw66Sjs8SUaNFWVLJULT
dBTt6kgBOlhZ3gSu5I8GstaLNnNopSSMtLWgDEPt1IaIA6zr8FS7pWG1Et1xgewO
K/TBNmnIi/W196/YLPNLzMPIXpy2Bqig+w9GWi6B8I0wDnj126kG6iDlGirRkbNk
49rC7Mq7MvrVDpOx4tfeEZROZ54IjKg3gLyLgVnFTYsYJY6B4wKkepX9tKD8Dgk8
nFf1CCiRvX3QVs+hOUrPUCPZdi7ar/2WcjBb5vR0MihCAfgHk98nBFUa6r8rQrVC
DH6A+v9y1Cz7N0faLI+vk0OxVASCSQWX4YE0u34s/I748I8gatjQ5gfcBVwxCFnO
HPAahY/aRiPk0C/MBdEXc2lZ9RzjFv0ZRUT+y9YcDr97G4vf3WRma2FsxtObvD67
5We6ax5i4Dn1XjRpdkXwh1P5y0TKsKPDodr7WPJd12EjpnChEmkwIOyDKZHt3mBo
lLX3W+9VotDHXTm/34ViaZ9xaePOcbfZatF1ElE7evKxsn47hpki+WyuCKWjETmC
LsNyEg3P8XRqCLrsdprthxO8UpTPmx2p8sn+42KLC8Oe6oLwJ9AuH1KQVQC1ZsEt
2kf3rBsPfCXzfro+HjIy8q5dljwFdrYEhmTyeuvbZ5DVo3snIf+c3n+TYiBQwMxt
3JgbThd5MKVnBKgV90rYT8S2EVj8JgBRpcwpd/cSe9Lb6Oy5gRFJ6j+3adGP9AaK
1G+dNd7TmQ/+lmgwQri1wDfuEjfDMs/Gym+03AcKBTFBXmB1rqoAm7XW1lKD1mvS
QhaIPr+yyIXQfCxuJ0Lf719HaM43dKOnTGDGdU7vY/Gyjm/frdKG/Ghq7Nnopw3C
cEMjM5mszdo091zupYIivK+soXqlJ3N3ULu0IEQRBNF9DSu/rcRhFgxRyLYZjn3Z
M0I78NCa1qWwvR15Lg3LxJa8JupDlCXNo9GtsVYLgKgcdlV28/muqWXQENKi/RMK
3+X0KcuDH97f83KpG0j+8p9VM0ohhoci/3+Jsisr5KbqfZgOtd2nMjRKkf6w4i4l
FInfapK61/cuSY8+nzii9Icbax3O9Qp2kmLoUbpDONmjr6c5ON62cWqVjtlvs9x0
fqvxxWRCqrjg0RmZaiyYwgIQ/BgbfN6dErzCNCXDvU0Bh2sSAa6CR/j1Ivmscwun
oQ7UGBNbUq3sC82cEbwHFevpqsZDFp7JUpMfdY28IOAGl27OQ8kqbEwtasejiMLd
Bk/qWujEBXCJ4Led03cFmDjXCHwht4YjdmHHwsca6MU3cJO9HXz+SyqwBtar4M+P
9Mz5ecJuZ25XmqK9pYijML85xAC6frzP2HfIiAsqak+Thy2ADurRF86mbNqwf2sM
zgEt+CwN/rJpUfk5Y3WoldmTcriJN6+UY482NXknbNRCFcPOr3G/p/OwFc/1GaTm
kdVr5ROmj6DlsvGcAJwIhmSWA4fb1Uu5Bnt5zpJVLlywXZTXouorAiEcFAUoLgo1
JHy2T6CK0R/DKFIkS2GLo7oWdpnhFyAMtOy4szvotkTkcBqaVe+b98jjoJV9GeBC
jay7l55L7FbDoixK3TOHYf0nXZz/jO0cS0PbaaSyN78N8Z0uMu+HmLZFX65Ugz6u
73radf3R7/IpaDO0rUvk4mka4vS5MQZLSjHJ/uw5yOCS8uKe98Qcjl/xw9HsiaK5
fHPCPGlYHlSkteQL1Kx1kr0UtbSekLYYCY2qOpRVvY1rym2r/0c/p+EagF2nG+1W
RzGcVV1VCaTzjt/13/cELUfYa/nejbjwMdgYleFN0m/cktx8F6Gp4Dkk6oVvfBlu
WL1AJ7FWqQo8eQ1tskA1de/WBjabUQirkySL1X8IFfFLOmZjvrSksWRBGW56nxX7
NRF/Xhcrps6VV83KnYUtMaC1czTVsUmA2aORFUod+XlOyW0xX3rE7Tfps3JlwJ85
tFjJVrgE8SjhNhkjY+1XTAh3HNW7L1p77c8CO+RXgwTFeQ+TLhQz86CWDxs/DMU/
nqszsJj43TXrIun3/Gh7WCCHkXQYvdorH+NY8HFYFh1EadEPI/koDisoZQVgrq3+
p8+gI1GbBl/P5kB3c/Vszy4TAXyXdCgNMABnTL/K+//9pawaHu288MW/N0sPpCYS
tebaoA9si31rVQ+IUaopI4yaObPM5xCOy46FaqvN58kJow50slW9VNJ1tFsBKS18
J+zLl+1/dyJWcWjSUHpM0NfEyXOJ7oYwaRwZk3Yuv3DYBJzdK6jo+wwbXqP79Kgr
4RkbV3HKklVDnGRWrwVdVq0H7o30bXRnRaVWIcCwL4flWhKWA6CEoGdJ7tOUa/oo
BerdG9SKGuA7uHz0yDpXN5nU3MGQndt+3ant91t+g6l8KGXsgI01xAE8fBq3WpyR
3s2Bf7+skG1PpsXb1wn6XZDYxn0UHWwyEAC3RfYaHEMMTi8dXKIU4u9ma1IDPFcR
Jgv0iwTRnr9doWJq0wIEIrvwEGGFz6V52D00wWicvJzhfGjE2SD7E8655qWbgO0v
HcO4Zol2HaX9n+3N/dTUWiF/k91X+LAFCf8oYRKK4/EcCVxWyhunb09RyEi9PeVO
hPkCEVnndK5eVDXnObbS0onAkLIR6GbPgTuf6O+AcpgWe5AvVTAXrukK/a5Wk/Jc
x2ByhoxFcOIphWOpr69nYrG+2OwM22fiHz93dbt61I9cjChXVKdsArMRb3n2MOfh
ytXwVPkO0pQQSiArOXUAk3Cr3i4S+xG6PbkRfQ0aQNmJSUxwu2aO5SaXPQHtute1
kZVUIkVBh2j1cy6ProY8cVEq3+V9d5RmthPIT8dTSPmrwaoqSZoQpp5yFzZAeLAT
u8SnZMyNI29ZExw/AuGGLQ0Fm6OXzx80KvO9npJJnyNxPG13skD8OmBP457fsqfr
oKJWMXwxp2e6KMajE74YipvaShgaUeMXAuZtjp1dWCA0UrpVHm0V1urvSGmTUUaD
HljNRCaUm8SXC7NJfLS+9f1fHLfQ96FT8j26QZIKuG6di737XpGd/YLqEsgVFzoV
0jOPT3vhH/N+0KJmZXGXz1QX4IhXH1+haWwGs8FxLlyiHaqW2mxEhJi+KTD6StWZ
sOYhw8DCxueutlxmiObLWobH+HUMn+Kl+HjNO+iuw2Hh8S/i+xZZuiZEKqzPR5/h
1WOo92UHQOCj7I7la2MODFsSIKvqofQLVbycAQimbPzRCdzd9NeHUw0tR9xyaz3f
gnqe0Tut3Bfx/W5k+oBPqqc89IAXxvA4TKC6470biQFiYha7gYVuWC9eoouQ3tBI
MoMiFjjuI+AD+LNQhF9x/AwyOQaXRoTZt1A9/Qz9Av2kzGxgrD69AV2EOgmSgfJS
DICB5zQq8k9eOwBRcOUzKI6i2bnUApmvvLTtP+abn89ZyL4RAdnTesZ9ogfzc6lg
2+TaQC9kkZOPsWxHy8bzSVTOFxw4qJzTb1+OCUW/x3YzcxhT0Dwqv8b6h/kWCYqv
CoMIF6NGSBH5rZ0Jlf8B29psB/pELqB3v67UvZPM5/7C4kn5R68P7eDnNxxiB8z4
/P2p6AkbSOy/h/mejYE8x8iYz3V9J83qX7Kq56FBZF4wfNuEhGbS9HYN1KrLEQb8
iyzSiBpUw5IqCAaz6iOmpXdkjPqKt2KqkGhEyt7w8zCanS+LAJSQ1tz5/qQorpWQ
oGsapO5fpHG5vroKphkhzlg8n2vOIlVWiCEdI8MjFv3vn/yX6FXVgwIln1KGKyVj
9G1TK0c0vYo/Zp5dYOQZvL8tTiLuytlFg5nWqduVcho6sdujFgdb4fdchrgwoHDX
BEAFfJXQtKsdNrM07gfp7gxq/3helZOuK+kfcPdqMNWZuM3UPXNQHGGrXHb6KV0p
Fh/5AoQLDf94t+gce6iq/hGh2oRjF1/i/P5bc2Ogu9ucKpgaU6tIT34K01kPCWZa
ki8wYtSTTNpI2suAqzpc0CpzwVUYho2Ko7d7f7zS9PuQ1HKMkugxWfdC/69WqjmE
kRPe21fyxP18pxj9DJjRTjErj/ejtau88H+NGD3RIekNRCcaL3yn+Sh7GA24CNxE
c1RiH78RFSvxjsUPk5PAl+1LcOQ41d5s5J1A7ZeKxYri3ckwswPLwODdStBt4f7h
lSFulEF3t3ci0L2GykHL3zcvAbVHJNa4wjGFLd4ATafE8F1oJdJvOcp5Rpo2nlVv
mFrJGF6u4k0OJvj4l6t6EwKiNMZdbevbtyEMiLjFLM/hxdl4+4UHLNGiVCum+s1o
tUX004OmIr5G8eEZHRvmf+skcft2AOXaesKx39L+GnMO8u8w88YIChH5Q9XW+KGH
jOsqwMaFkZfJ9V0lj4ETMGXLwzHxpB5VZtDsrkAvswqKQOkmu/HcedWRPYynyVlu
R7JrBMNx5kYbHH55N9iFwfNwOLz4E/T8InF4kTBtJSXZtb5830e6q/IWSYwITI+R
tdpiSArMgbaMO6ehruzheAqjSXpWsw68or6bqArKB+OIODuTp4EtGSDh8sWpRy5I
4Mp9lxnLarh1wFOlYFh4NqUHOYyFx7lpgNyCb7i0gkG9dG8WUKXjH2I9HA6AqWeG
v1M17IACBIZqE3vmBNu1BHqEBflZ4/Jq/h2i4MWU1yI9fm/BvTysQOfRV22tEFbP
xQ5pKMjIQlxxqtRVwkZb2ArhrbdpcqCTWuSvpTN8xbNJ6OJPWE7i6kgo01fkOpFa
pnFK3j8RViATYQHnwpM+nGDAySusg48EDzdSGaN323suRPq+yZzTjXZc6SOqmEjX
Sh2bVs1aPVpTnaHedoCzarBmsRDn576FKCeX7OkxnvTKmzDnQt4Nc9km6jkQjnon
hRZdMv7YT181tyo4OJzDOL6s0cGpgEjOHuJixRQNyZXeKCPB3qKKGKKaPzFFj/TJ
PWwRBgR6PgXtKndTIbcSNOrh6Eq8ctOqCNGMqpwBvCXuhkCYm6iSJH1y6laZJYPL
T0kjM4wLC/+9l0FOb0vfEtzSfwfjB6Mh5vfVnpTiSPyqTN7ccDgYgGS4AmSEImjH
IzluF9McPunoTBhSo2lyRkqiW5zk1942980t4k1xDzFdlHfdEFbvQbx2e6JZfgDR
IomBHLysRk8QSLwUydB+iUk0OslykR58bNLP5CpblYtMz5erxZ6b57hDRqLDjSqr
6SNMgax56T/kIivGmvNkViRvKFIQXrQuPzA+ASKdB/oB9t8pwRIYvuwhrT5qXTDO
4MwFOeTge9/RXfUMqCm83IF6zomgMEkTAPTEW06IyzGus9ZsTCYJdLeAjmZpdW/3
WVtbTTRb0RTR4gTIK8JHEtL8xXetGgG45cZITPw/qd2sUmLkxYO1PtK+0rE/nVGj
Xu/46RyCVYNbYcBsDhQNaKHkGvhS2QTK1UF1fbSJnENuk1GeJbU6QsAGIWZ5Tc3d
skM9e5eQIp3SSFceqLVmPLNT4W2iGSzJ01OnThFyBJuzwvF3n1XFeTUJr0bLjsef
cSMg0qXjBeflhGvj2/819SpPv0YrIx5amEXWXStdZd0ft4yzSVNr+BLPgMAHPwZl
6nIe+p8bub0XgOeR4BTkNAe3dvwRO8Z4NOqA+TiCq9l0LNyBh4sMXeH+d1CrMX9J
DQvat3ZlRZwHxLl6Mg7YcVI5m67GRbAVjtvX5Hy+eRZPruljwwhyo3xpnA1JwVBv
7sjG0VU4tX4f84PqBYMtfFkXpSp1EnGau2dk0Cdmp1GGrHXT3KuhHOnC5MKq083C
3N+uqPU+eoTOPKOGhEknZUUAWDDEwZ2IU39A3pNINULT5MEUqpkKRyzToSKfWDN3
kpBWRar6jDV0KgxPuKSITE0HBd6moMOz2Zvqp5OFuI9SxjN+BsCZq7Y5zKCsyvlf
rh+X76qcqiUKK2SJhl5tu0LP1wolKPLVwi36bfdIPGzKszIkbo0XLaUnAJb6KtoC
V+3mcX9n/XhJ4wdvq9dhJF0+ba3+2jMUEeslua4/wwcgfWwMuhwx/qOEL0thdbb3
GCqrH4d47u/7RfCvBJGohk7F5lQkmEBhLSwxkKodOClW4eSlOUd/ykrzzxM6zytS
uamqdYSe9ALTOJqAH6zqW+wvf9hEJnKSDehb/elNONRVdMXoUx11aM20gFWoJjjX
t91EXofpM6Q9JOLjmT73+6zZ+H0OZlUgBdW1vXqlU9WS/A1FNliq3kkiWmsb/Onz
eGktN1Az1JGy2Y2klW7CNgdUpezkcdhjuSaAH2DzitKtePVRCOXSOiOTGLLHdgzA
tZzaw305CddTfNOi4g7s/6tRBJzOjXgNDRcry1uzQMwd5UCo9KXkRpIInWCwsBQV
7tYUTmio9NeOBt7C8xYcV0qIbd5wkoVsEo9uyxLFmTFhjfNEUUHQuqbg3PYZz9mf
vV8m9q7FZ09aQayTEfuS9ed7y/1iGVz9awQ/VBiPPojTe99wilGm2FlqobIK1pc9
P8y2+E7FknfxbAiq83DpNcOfQ7ChGhQFIK+6sJLb+fvp0TzL0eJQLBAlLKIfLHYR
WMS7VfLgk8CjmJBs38tWovPNneyR9gNAhHSy+jySJ0TqX0IOugPOHh4npNKc3vpo
hZqCVnBVkPlYS4/pF1AJjyny256rRDMQlBqRqTtVVbUAedRRQTkDh0U/iHMt1wMH
Ngrguyl2bQ55pA+9DxbB+QMB/QKvu+UhEg69t8Bzh4cOlbX/9eJBErmLyq0jGJio
E0h3ARwqeN5i2wqPOXHdPIjctR5KQskiBktGLg39EIxJBgU5sBtaD0WWPaoArob4
BbHS6c+HKQ126IUnEpquBadoxzLAWlZ5o4Ok9XBWK2YbBhE8v4FmtVGdKmTf8MpO
uRlsMh03KyZzSW7AswC/Z5PnfYuZR0T7DRjcEvPuWIk8tmZE5SpDGuS5nWHLut/z
hi07hlnOnHxoowZiSKErfi5WdYxLzlE1bih7qtdMhqm01R+FnwS67PSfA/SVfydt
l5//92xvFvTqTkWD+9yOYg8ojcKk6WrhtmqXG/x9aduHcJA4II2zhmaxZCU9HyZY
iAhzM6LPKjtAPdoGDbHrqjsRo0XmetlBV9ZgtJaLVDQjsQawysAqJieMprd8jhPQ
EEuD62gjyrBqUV/YYpidxirJPm9tKG13VPk3iugnh0/wpuuqo7/Zt6S2gfGZdlLr
wYgSEpC/fOhcd8bUo3uym0TKD70Q8dueR2wvopyIlcR8TeZxzZbHkbWeZfTyki9C
VwsozVSV/PvqoU/nUVPyHzvg9xNFVm5NSVrY0h6eWJHkzUHUa703dSSMfMJKa/cc
Lr8BohtHfVb/7jxlqrjyEWK73ml6UYJthNGEOQoEGqQFGqunBl1ERxJyrF7m5Tz1
1v7Nfi6nv+mRU3/jAVLeIk2/GSb5wtNzz/NAJiAQGLk/jcXZ5YqXvT/Yc+F9f+e0
zQV0iq2ZWrwB/8ibMsaPkZxwKowSWvBY3NSg4P6Azwl9a0Ls48nVZHqioo0rWO3u
G3Y0q6FoHC98nNr7184sUkYIg3WlB4s4pl/pD78QBCdAu5ZDMHsZXgD7cZcfmxhY
2gzLejdjq55J6O6gSgXfuA+qe5kfFP3/VPA7aF1IOPtjFkYWjYH2r+fPQk1/QqLL
oBkdKx6fgoDzhqPucpXl2n/jhITwMKQHxeylY59rF0bB9OnQv4GOJusGU0cpNpa9
GnSo2z0RY3X8x3VCv19P+2cPuQJf2BmzjQoYkpA6u3G0BSx6S4lwhVskaLHOi9qA
LywGYX7tewrfYVKsbjueE4izrUPzRx67SK8R4W9K7Ta/c5DpQo33xf7KI5N8gYKL
KWUhoCOodQLxQTE1OL9h7fDDf6/92jtrmpli1Ix3uC6HXQtCIzSmtMwz+VM/H3zk
DbQYS18TMYh/6/C85ndlfZzmSGU9sQkj9nQIwQ8YD31Ng0kb2JPCxVvKtgiApdt7
/YfKDrdFVVhiT0xrthQgmT8DrM3N6oDWsIaHH3t3dBOsLoRhndseYf6aAL30xdzR
o9sZJsXkDrO6ZJkaXL/2XgZQQCP2DnKbwhlgDYwq9HIAb2tyuKftpIE8abIVxI9z
d+lsahHUF6wGzi+2PT3PSSfjQgRDD4h8o5BCE+CbwJVIPCLTIK0J3A17TElkMNSm
FxaEisCVqrG7+ZWtGRpwW3lw88yEritGZXnIwpG8RS+7vwQKU8Ixy24ef8R60D/o
8Q8ghUrENH3S9iYt8bFBilDkBtPZvFDZ/jgjeBaRzkSOPxYlZPWboDc2n8Ej01MD
SnYq3GLJPY1wrl8Xh2xkUDvMhJ7Riimgll2Och5hNsUOdLMp5BfqdgnU68b0Rw3n
wmDHkeR8tV+z/y6xpCzk3UGykVz2oteAgywA5JNsJklYKmiGul+G4St3smfnBxxg
BPk1cTS3oVp6ZDrbkUIfdGNog14EKEkaVMklsUbfQHHL9hZEl+SJn3wnfpaylAbq
oHj2l0JjrofIT5e/Y8MZzTKmG6rcP+BGAip9oItQYvuX3l+bw5f3/7OfVtOIDYdD
hq35V7u01t09gybzegngxaGlUgWDpsXgyxZbQyRo/wDsoda83CGHoaP9S5BH7TvM
3UtOeInz4naRjbzK142y09TyiHJAuCAuf3iN0vaknb73v0xgBi0bPA+3OGvFNnqA
VNvxkQZRoq77PxG2V0H52RG1fbLs6KHq4vZHbEj7cOXtV5fYC/HcN+KavXWfyyi2
BEp6Oefq5HWQCAP7bWwxjbrEJ/ca63tCeXnR/RSGApqrlZI6h+efW8g0B4VYcoPI
HVyMtiQeYsoBvmYaYHpeVkQ5WifSnLVyStParb0r3vcAubIKmnw6M3v0xYzq1Q1R
IOki7MRU6yWr/9h02sQ+Fy5BtVMdVNYQCAz2PXB/9rURHNzcPQohzT8Xe1ptb4Kw
lWVeizg9Mq8H37PKRn9e0ZwWbwVmh2blRwJLl1yR27nSQahDlA7gneK7c9TPtfqE
DyNNqAYqeLqQtAlHnyS+ExgN74s6DfqYKm4BTq8J/KSNSdSTqWwMFaQ6LufsqFxB
8INY1sSHNgVNizj2q9qN+eV+8SZ0VTlqGrDz9GwDegxK0zdKdZ/JAH2I8WQ/JeJh
X8vKhblfUxLobZG6XWOPMbA37IX8LXyuGud+XCTAYVdmwtN432Z8XXYfhy3Nobpx
Xj3q0b/++3ODkCKu3alUcreE0kpPPGmL6NY7uyKfuOQ0sf/WPVt93A5uWBvHo6N1
A+1LDSTaax8L+E/dfTfuoiwviQp9XIhGI55trttnUWbTxDPWfwE7hoSqv5MfqFGZ
dmZ1k+0jYrd5edh+JWyqUvxElqQnrG7Ll8W+TfsctdtVe2F9kvMSPMmD7zF0juqQ
46KMtGKRYv0AAFjHnlUM+DWby72sMq0/Ci8GDEwYuQnnp0p5S5PaoH3DJO80mkhs
Z87EzhwVdoRiP/xgxjQzZmMsPx2SJTFfTdtDYqKXZcfZrHwDCIJWOLuemj2snaJ8
qFHT9L0y/4ZnCc6n+3RYrkO8p/49zf7U30LNYs4MaXmJy3ilG8d5Q2oGZKotROhr
QXt/OaZZoIRfjhqEkRJGRYCbjhhokilhUVYfmqoaFW5itmOoHcM1gEI22/Ew5gbG
cchKkcly41JvVWKHKP0/BtAtKzlV7c4bO6I2ueUFdHgf9tBbkWaLqzngUApJVQwZ
Fgwk3pDZN9zNWM/9YhHwPljoc8YR6CcztywC5aMKd34WLstoSsk7wysIOqbZPhVJ
hQyBybp6apZy8kInqHZSxlAgpuM65hZKb/LZlqQKCZFpAQe93dus0h3O0Yo4XGtA
vhHfSyx9W4ADKY8wLe0oHO0uL9DL/OTbSkEBU6SahLqckXHuWBNZSpkMrCUgl8M6
L1/Bn8oHwpnazRyqSDgMDakH8QbDeheS5+/0cwOSx4xlu2hg1uzKKgPhAl1AN0uD
TlaVTJrlBuG2h1B66aBR/m3H0unFQpEaPY9mBxWw5f+tHjT85iLwBCTaHqPp7gaU
ct5nl03LvQdWxCwRTgsGlEP98MlR7c21qnbHscXrhfF1/E7217qOZMgMoJeoiDaD
6FC+mIh3GYo4h6726N1DUO+WmWZdYSIdg5lo+4U+DBQ3wrM8jDgZBUXkm6Okuz75
p0gkSJUvSiG3xND9bsJ3yP671dO4wdTajeuoqlaO1PHqe++rEZgrMQap88MJtaSb
zyB48Ycw7i4PMDX3cFhAPsCS0LMLospZSDCeVEP6ZguhKxOIWz80ZLccgXa/7Q1A
bT9dH9g1eBRCcB3ijVHWG/cbCt7GChS1z5/WHab3e1RkP2PikPCdF9p15mRSVsrI
oGX7iHwx7vodHJUgzCNn+oANEkif5p2WxdrwpCiObFaCGz6xT3HsI91sajgyi+n6
CGRpJ2vai2xJeNmg32DC7c+RWfeAO4taN1/x+lKq3jGcH9v7eJH7oEWBsT/LA+EK
tA4OV4XWBXWudd9R+6Aek2r4LOVVUw5QBdvSvLJ/a0EaenZqdmD79gq24B8SS7Jf
1ZwBd8x4N9ZE/sUOoU4TLnz8IEVcQEXhjKQLKzsYPiBmxgNXjkMObnekJ49c6Yjm
ArrvQr57Ru/zcMKF/QFgG8BBWr3y5VGueANS0vlaV3o4mfcHVtT1zBy419u6fVAE
fr7047/eWwZfofzLACPY9uBeb2F4tHokNQzFOVjukzDXaLWkYHBMsjXkEhKc8Ycm
MPC7mniOvyd8EqmqsCmQUJlLJwC1gq6Nv8hBhOfY6hNCazqPp+PaWSb+R40wwmR1
+E9a5yCKQv39rL2a6BxW5aEgLcQ0ewA9KCjOaEDu35P6Wd7k6w9Y+RSpfnRcypi9
T5eGvBVZaUCf3Mvd/UGlvzhiMxzAqdHkBjIIGdAHsGzYa9NTrlDQq6SNnW4b8Hiy
UjqYCBYwn1NbFSytdEPUK+tGB3fSv8+4sP5qpVEEpQE86lbJq7nkMw0DjbHgNDjP
hlhNPSKBI1iGyIewOq9ATFVuyo4YxdGSHrH6H5SAKEOwst/DnNhXLm2hjK3iu525
QvZU7pC8TMENnvBBdAbH+g5VKNt5dskkxfRi8P4ci5I3kWUFM556od0cvp4K/A3r
CaGXJ3CDuxLfs4pxl4FfSuHnZiYWuJjMheDx2UDurBKyqKU/RWs2fBY9s7sfjNpU
p13u+RSkhk0oUyNDpl6TRJ36ssbrXPMMmaVWMCPaO3iX+Luvb6Zhv+USndyW9lQ+
vpxgdA3VBIltyfxtSAwER1D+WMY59PKw4+vO4+nxkugAVPGgGDwPcnM1mPCaI0e/
t25VU3dK0aK5T3/KQX+s22lzCO9hDDU4takYXEPaBrmooNTIH129DOBE4qqBfB0f
7qzlHEGnfzdWsgSuT0fhZEeZuJpy7lwz0od2znZNy+nUGHbAU20udcioHWRNPPkY
DZgXYGvS3GhMzUh2xqj3tKF2MVa76UAjEv5e4WLol4k/X5deGZHXBClOBEr2MZvN
fp2dqSXw7faDneuPx+WRQ8t5cIhP29/asFa+aOhcED2/BfuLAFd6Um+hEOiiVCB+
ehIz2pPoXnfmIPQ9mH/gcW2EGrI0XhiDMrJWcVxVljY6oDZ2AnFgnmMwZkDRvmmo
5Cw7/gmYrlqYWki+sQsMvmBOsY/eFbT+nrOAxS6rAMrTVetjfSenwpNJ1mc7kTIH
8he6cSDMsHp+Kd+et0QqYYfKToeAYT2GwcHvUqxR9l+/kTmMKwOOIFJWxldGAZLG
F+zDIu294L875Hnfe5SA+bJR2wex5FurAdx+KUjCDtRK2uerCZ1f89/gC9PU7slN
2p7LebhH7P2cijUsKpi/en/FZRXlPCrWA64c/rRnjenC03v/Fv22tidGFJqPQ34Z
o1PFge+hBseA/VOLMSNz9dQpaf38NAA5wMrsZIYhrKo7bMgZCZKzbWUyL/eIndDd
0S4bJ8VAgCPpWJ5r/KIesfla69DLH+tcRhkZIP26wE/sOybRqwTOmK6LNBCvwSuV
D9XcNbfFiIBCcRVh77wY1nf4nFh/oFVvjAKfR7iQT85hJAIfOB2tZ5+7Ou604XX6
QDMuhclLCIGcU7tyEBMHP1uyZWy9RhNcaErxYToaQDdBlMA2jJbCQQsykVUMjFQK
+l237oOyK9v+kQJ+pcizEa3g+jPVffEsiXk4GiRmNucBxnlWQu45Se6bZzNYYp5b
9i6r3SklyTPgKdLAOtEwkEI80HAX+6AKR53E8fmTSPvaorsq8nTwTJUvBBwYf0PY
3slY5OaFGOMIEiP7kRF7FnVX9T3R1vVddzRanCS4cV0cvrzuBp4h+yAOv2NUVezf
GC4hzR6F0CO5lSLD4vdQ5Xgmr9MvTdu0a70PTKc9XpliXmPmS+4FCjjxrNqhA+MP
a2M6Yfq6AqIQGPPfEH8ByXHwcS5hHg1d9hbfh3xIfqglF3ANlN/G+UvFoo0pz+OK
9UyjfG1UGGt1e7FnnbAJfhBbKMoD2oDI/8oGZTXHsoNwxcnbCHZWh030onb7D+ss
7kFC9h2gyJQwAwgQJW/NF66PJkklOM22sCIIp1oET4T+jkLXtLqnRLv+QJAJfaZt
SjMBkyiGCI8By/jKuZ33l1HRGLy8/WZv3WdbLJi7tHgN4UBntodChhE4nsOKVApJ
u5qP90o3wASaAsl64Hig2h4HhsvfelDNmN20RDZtd2fyr/GGBGQE6lEVYp+nBQop
xK/KVOLw84JCDkX9dFz+mwRYpKpb1UISZwoFgFzummDbJuspJwP28PUBI0L1pooE
pik1i0+VLesE34/2XpMMvoNPTYWzvsxE6PmkvObKr0Z5cs5L8n2vq4N8R25wzf5e
vQCi0wAgmaiNojkIvulZ7IELJGfdP/aEcAQAmTaEFjRfD5Yn/G/TloO0erC1zW8e
caGF1/vZx+4xLteYtDKchBNyRzN0fzl4Yp+9P6ppvXsmKNoyz2eL8WQWoXIeb1bc
efrKx46pSkz4GNzHCi70p12K2JqhO7BmYwgDQbeJTf6YVq6QlyMcZUXBWvbERS6w
s+N5b8cjO4NijYTB0WQBgW2XILU8sQd3jGaSCsTkOcuo4faTI0Z/gFp4QTZ8cFaz
nRCpOiN71FfrORfnE2hQFapJ9cBsyCf3pJnWQtKldEucIyKtBNHj91vg9MhoGc8U
F3AbGtVpBcyDKROWhCeYIaVLHsA2Z8zoytMtsKNWg3E7fgzOdHywQbdZJ6lLJskO
ajc4dQBM7JiU7CE1ImuG5vAk2olHqoimL+xRbAYRtSLCSf/dDScJMnUrBhFWD2kU
6zOhpSciuOn1OLmWrJhmN+uarQfgzzbqrsk+KsaSoCHr1msuUucs9AY5LylMjeBd
6AP3mg+0KJ3c70qq90CfmX6hLgTGNy88qq7deXWyol+Yn0P0YNtLE1ZUgGoTkUm8
AIRpXLNP+s6dQA8z7agA5OV89STFEGd+r/783odeFNNa5xt4FaG8FmYGH5aJAZsC
jFUkF0C0DEWktG9oHFa52hCY3Y31ysD9ocYekSGt6XOXy8/xzOt9zfvf9xQhYvv7
4mzQw1Sh0HxlCzJVvNGPk8iPC3MZhCMQDfPGETwC9CNJbkMlGb4rPV0LFpahPDBJ
pkAkeiKeZnLcsriaKDCwrkJg3tGM7mDrJRIVjuyT9y2QbhPp1J3Wr6q9B0Xk+wpA
8p+uEZbTGyRpdu0ZylUwGF1hxQpNn6i57ZcufHmJko2itDNFjSvIViWubApbU4Vk
dLu+88wfzC63ePgV/KJ2TSsg16A7NYlul6R4gSi7+A39JoAlHFvoOLco/H1F8Aax
vDFOPVgbVLIxNYZIdnKGilztGnPsM9B1k/7bD6jkbu6tcuA8Wt8q9PvgNjNhD5A3
gKbH0P9n+BhvVk/DOJjLZTeprpsX3xlYLditrwgy1PVjC1KxvZ/Qo8kEYjkfRI3F
KWfBdMSj/nTfYfoXqrga10EJiOxAHUcya2oasgGlcL2REfPHTbR6vYWll9x5ABFf
Tl1cJlUNe2c1LiqQjxX8X1t81O9ry8EhtHnZcQYpQVGQl/UAnwgsysk1UCcZLzXx
/KpDvX39LQzazyt1JrZMdcS34kkhc/Ij+oROCVo03rpDrrjXjH1dnlt42v1g36b2
JWeD3ejLogfQI6KZvKUv3geID5GXnvBwVY1xFckufRF6mejToEW1fX2z8exBviYI
cSPQ2VvJK8g0KNFyzlVn2voDY2ZIbGkwPoY+wNuP4+vVtp/HPcvE2xrwfswhCv5o
swWip1Bk4a3DDvq9NfG4jjY9gcKNRJeBxGJuP0055ZE0G+Z5ttyLLlcPJFwWJ6LJ
psMDHa0uQrrzza7BfPVRGiVFv1j7+Yg5ft3g0iPoPwQgiVcysSr6tB35pUcnZAsz
H2RUOb8XHzx14/EcHQgnF+7FLheSA9526DdFUi5rhFlndUirfw4QkF02MxKQjAKu
zzrhpIXcZzgie0QxPe9pjdN2vHkcyaoeonnoXpdl5uh1yAMPZpXDy72CVKu7KZDO
jwSrl44/Hh4kt39ZFGX4QyFJoZZ7wOurEB7B7r3eddWLmcSbAaDO60g+6z4qSkuw
dPIZ8DSabc3Fm7eFup02RY6VbXmPYITvdVptxvVP/neQRPwbxXB+Gz3T+OYVal20
IucPrQgqcfRyTdMOikmv5P1d/B8ViPOS5lM9H1az6m1jkjFh9+OJq9H3uLSNPIoQ
Zu04XFRq1rpJyZ8+dbZ0VP89d9JPdL6SFdkM82MDBaaIYODdqB69JwqDRx+knYFm
FUTsmw28dkvUNVF9l9LI993gsKeM2QBdGKXzu2BppCniAxBr/y+blCldl9I5jxfZ
XpDyGaxw+Cclz0Us+KCWvr6cLGYiiGw/k2RE+za5V3hAGRSZfgCq84XBuCEm7fZX
5V+eE9K9H16KoeiUOErSxoP9e+M/prTbEByAWOi0xySd2t+eSmIokqDVsPNJRdxT
KlFEHBH/rY7YnU/JbOMpfF/3IuTZSk/DZaAddHd2RcL96OINsZ5XtFU1d5fQ7Rx/
r/+grhBBSlcXfhGPm4lx51mqUF2jzKz930rtKFM6M4887iqElO3mKQFWo9HpsOv7
wGWx+LElmATxBlPz+a3R5RtpnESTuyKiz/3ZfMRdzrxv9ifuAjavEl2cv/VNqwzh
k1vmIzIMANVnnLarPrVupos2KZOfk++Rg8f7EzvzLEtkcWGdlKCZhUKSGAGdun/Q
oYXCQNuQWXe9hkmFMuY5WBj7jgk6VvpQ4/hw1XNBYDpAhEBiUf+AlSzg5HW8RpH7
arHjkXK3byPhYP8+zVaD1Jpcr+bO5m5U4+9x1ucFtQ4CRyHhUmp+c1cedJcDuIbc
hl9RjcO6/PVENucF0ek7nVpmlhAGQxIdsYwCxFdCa2j8NvYrsFOZMOkAXGKQniRk
EQ15X+Oj5alafhKQ6QoqCC/FAsSloU+Ml4ySm4HQ+k4nAeVOsv5xHMv0On0u1oyL
+nJ0e/hBQm1iSnMufIm1W9Yuss/hHOH6OsAplzBenEHKWT+9h+c0JHjG+jAPDLRr
OfgGW1qGr6FhpHOxSexqGxG3luP9798ZNbhYXHeiAtsiYL8RQWzFEdxpT/TpPagp
KD+D8CCVFkvV+3WqXXtFTHSjbOM4toiVACr0olEvp//qgsPd5FnQJaB9ikqclA+L
via46HgDakayWWAXTfo/YXcOXTahy572ETHegqeZkAv/2CPRCmAMACXOxN9SGQu/
i7YRyKCaZqp866YMMKNbzFAr8912rM19uqX+dm+BXKtzazvQE/h5uPh302f2lofC
y/y+Sv6Vlq4AXWXkNhFob7aW1gHMU9uC6K9iXrvK2bneyjGTRuv34xMyx0i/GP+/
PZNaBB11jfkmtWavPIf9xWFb0l3kDBHsIkGA3hdeqo4grzqK/0lTZEWsuFCvziRL
ZMP/6sKMdcymE1lB81KcQbUC5NvRPDqcGz+XUMOCW7tjxoZgL3iyGTOGciK2se58
anmSb4XYoey/pQUymUpbznpo0SUlY2MjzDfYN8Do1+m54u3gqtUzuOGSzekBXAui
kf+tYtgMYSnMxdlT9drl96P/pYzd0r1euoDhdHMMtDINZSTaRioODgERK5zUcpqm
1PuNRy6JeVKGnIrwH5pNWLrhRhmz4WiLsGfPddnlxfgyZubw8np0KQKOVcyuhiOd
LV3kysYlJ78KM6BCXbsgRGdABVve5YVexnkc9R1fRrohhhlbOZMFI55XjnU72fKA
dCwSE448G3v6jY/91S1LzjAI6U90mEwghZc5NUVREQylP8ieg8T1lsMptwom//To
LIkKCHhxyhKiXrODuT7XMEpcMBcIkjPwE+YR+h7eojcyetu2NzbakbBcNvsKrnjW
eIzjGAHW/Hh5TRcbIxMmzbwZTnC8Ks8w+4tx7wpmOZv4JsQhoIq6VxowdN9V1Fdq
cPFKWkHtny0ZpCj36GF6LVuquY6LpA9HBBoS/AeTTryqVMpGvRg3u2mFAnI5F5e+
ISPKNLbdmT9suV8qtGcVA8sgeXdPBCNWi0fjSiUwpkk3DN0NWlXie65fTeeGJ8FY
dbW5TbsHr7H7VGkvMyqE7b3BcVg3LtzpS8bGJDXpCsv8WRRUN+Zhg6NvGUvtZNdf
GRqCvnEbcrlUlA46KS8KNQO1lO2cnsaqvyfC+9sWGdM3230UlUhRXuOXK447nS+r
1tSbN6zm7sSJlJxKkOHoDD8UO0EXR1m1u4E3MjYSd5GpEwJBaUSlMFA6Oe7IjhyL
6Q/5PXyxrWSxIzyFPej89uDdeCYaNF22X88L89YkYESg9xfIXKdxMTuSpisJx2Pq
BZqXg535uqSohterQvvcHDzqi8PqL2it7baqQD7+V4Zkqg7sjoiLu62YTO/YPbQS
zCtEkLDk6eajlLmYYC/bGULP4CctUpJB5VAXYY1ly0hGkwAP+y6t2v83AxrUIvJy
95yTvskCAfAbxOgsnCVg4hVO2PbyMCjVCkT8byfA8po1y0Rr3eiXZgDKQGghq+Vi
0vtMSDXZfuuwKJiTZym9CUCHWb2MKmoZmDxCXrKX5nwP8kM4X9yCi77uGXcwgSX9
G8mjL5JGyxKGK4dkRmmA8Q7So0yb+8/0f2EZDho3Bt9h3dRNcG8WftsN3qgvyzOo
lhDg1Lyum3PVOLkBuRnGewJjJCRX5GJDzo66+IfMMibyIt11a1LcFP+0FHSv+ve8
QMdlHm9VurmXgtFe6l/EyxqtjNPHONwFkqWCx1lgciGLOLwM36n3W/tBrF23hX7c
r2FjgvCVUhqOXNMFKt3iNA3Ru8c83gIpAU6MGxth7EeVY2sWKHNhZtweOus65wxu
s0N/eUHAacgBoNxC7N3A3gpZHNst6dsxsoqCWF/g+WG8rI49jPWDrdyGUtmLXl0Z
YAY5Z01YlvnGi7RysRdejPdHLlqkNQ7WdpTN/ZvxI1XgMsPaujYnUnHjq15klPfW
cuytth9dmbF4mgd1/ib4Lc9oVDkDaeIgB0kKnmB/zUTUPekS7eOhcooPk4aeSIpa
6YVwEo01Kf+p2A3aKBr25+XMUfjuvwln33co4rae208V7eMZ/sx0829hOFQcl9Ip
OKfzAlT0T6ZlTz8Wu/MpYYoxzoa4ocVRHFYzpR+74qnWrinQFtr47L881bnLy5yb
FjpVP96C9LwxtyoKTHc5tZ/SGigiLY88VECEyl0w1/4eMAwA72X/l849QcNX19KX
9TSsvjDGPw2sGbsZI2YTEeBKgrthXK6UhuyOabUF/pAAy1kOD3fHIj4BXhNSxJdd
xaJsyM+RC36+ag8mHOHOC4HgdPB5DqIAWqhrxE3H73sjhv1oGK6EAL4nyrL7vhxJ
62H2Y5qCY8xWKj6KEQ1q3J1AWOegnxhkkRH0HpkaXPDBnV8+5eCSOxuaSXPer1nd
lvibT169tcShGbWfytE7ZKyDeW4haDvXuo6L6C/Iff5oHSOb4dafm6hnSokk1ynb
zti9ceC4N51awVmDpBSjSp2sG53Hze4r7FXNtfHTEbGnf+oqciwoJ5AJCVz1jIV1
tM54sFOAE4Mc+mAc40x2TafcrUz3T61PJ8Vavq4JCEANr7BeFy0jobrnp0deZc2f
QutijYiLtv30KVuyAwFkRWM9YAVt95zlcOuWx61fsga8JjW0ZNV03972UhO0/QHw
hVUY9YsMPOSe4w4FXBYAEplvstdtGGwlFM0IiG88cTGR3jVh3YO1O1Hc9QPDeinY
jB+g191wWwfF+Ovj9ihe2mOirT3Fut+Ii2NRNm5+fvvu9e4qvLLqSftRnIaSJxmo
OL9xLn0u8aVb+GHgvGkWDNwp5XS1LIAFwmhnx8t9UD64nMepCUh4OQ7N1Spk7ETg
Vk9tANE4LU5ckSi2Fnw4a4x6lCXZmZF2b/FijUlOccWdkHTx6RkvOevb8F2nhsBY
2Dtdl4Py6+d41GHxABcHr11xu45Hl08aSqn/rTlL4iDMudADEsn9EPkbr23HCBB1
cSoqZp674NlVF0V+YyzupAkk8FPHtgFgdBRtuEwTN1aMkNfF8bUKfdcDwMPYM7KW
ll3ZeH5Of+b1cQ1NQeISwCxBXzOmD+KbPnw+yJLT2yzwNHYDsKOympr3V5cXTD3d
j6kKpZ2y+89GAuKHQzLyKfQImHuzuRImkrtuHZ7zGt/hMwv7dXZYFqT68gNhWnKS
9LsUsfDNvn6Z5GWbAW1gXgJ8AkLPE6x8NFf+cL1wteDjSM8RTDbdYOChEyJXUrvb
/7GauopgFT3G0oMDttTilNzU0eeZ+r/AOUOyLR8CXg55Xv32eEgjG44od9BYqB3h
JPx10Yuetlvbf+TrkKGV2XwoeHDI9Fj3X6j1Xmv02AeHT2wkyyNg/FI2s53j8+b6
kg6okRCoeWlIzvsmqpCDI6sXYOStS9dQeFqKof17bcV/enqWxu3uG6jxLBeRwkk7
1T9C3hyaf2us/Awjtf+G6ZEoaHlxH0LKnJihZvZo/udH5svbH2hP2YIpyMu7kqJa
USXqjxSeG/1z+ncENq7aTqydVzI2AB5Jj29fFsXM4ck5h2W6bqVHzmVvaIyn6lNk
bMCuBLWpq3hNuQrL7RabH7ei7GlT67jY6AsK1BaYdj6cQPWZd0vOBnA8idbE5TdN
O86cHcCrfDi36ff3BYMbBMd4ngwsFlW/zwiydja+s5sVO3MW/2GFOBpwIDaNxQVV
R26vnktINQPREdnoSVYJixHN3H/VCXHSj0T33grpkMQxVXgqCYC8CJ+akqgBuNSk
m461PO+sBqvQdSCCsJSBjAw2vhEd/Foe/aLvj6hN94wsuK9IeaO8aSuvmN1eLZsr
Tqz0h+j9rN29dw1G4/2G4dtj/3HvPBErpSLLV/X4VlSlPwQP9el9VkqCg/BIBVp9
55Z7SSyOA0O7BOiHN7HrSRSwXXXyNYXvbJpV559tvk/1ruSHSYPb3yEFqub7+Oyo
NwVQ8KWhxuxYD08xJ4mCWjJbhbO6KJBjQNotx8NBRnPHd4M6KvE9MBHJIIeLf4ui
HpKG75j1ght+T7YIYocLN66eMAhRm7KKgSmY6p5BJt1bI77cy3fzOElH9FCfTRKm
z2lweZeb+zXmFduSF/XArXbKt1kXe4aQWI0Awejd3oTqdSfFmFND98iZ7UMKQzwu
9Ud2LoB4n2n2efYVFowmKAZPJw1O2i6GtsUg78PpTs/FFjG4oh2doW2Oj9jvbcL9
baOccYJuPI0XSGqDvsVUpdu2suNXrCgAoJrWOvKG2XqP3ZIaCra2WYnnIiVvS56e
KLTbrjo6KZyXyVwqZok8WvwWGeU3dZiBYe5Mnh1toJU1dcRYHzf1VGS0Si9e1pFV
+bsi0brxskBcua+Gn33ZXcf+HNNJVBQkZq0zPIu7LAHw9iL4FDFZNbl7avxu4ffR
dR99p2dpHFJB8RPQw3w9ch6RlD0aTftwfh4FU/8TEIHz1u7xvOjpMdZ3ORQV7OEc
TuVTDES+Etzx8IuH9isFVBBy74rvqIbX1kcaQdCw+4L7Yb6s5wjeY98OIMo18WIL
6GgNq+RsnbtTL3wpsC2aqdgdTJMpS7VOXkPZyUbCMVUMej7QUXBXTZbwZ2R+l8GK
p9ZpSpgJisNl0dcX0sjzJo+02AonuMwdLUscs4bDulWkDbpIJdg+77RZ7ExyTtBo
nlrI3I9ziKBIj8raXMyGLglZ0bjgZDluJTHXIFNOCJwTYUsWKD15UzIpVtCvMaV8
vrmlp4Hn2qmkxnlCzsZTeifFuLO7dKlph4tY1NJJhVw7OueJnL3j9jlZzgmF59RU
ptXm8xGoorg/TQ1v0TyIYynODfTgW85YjSUw5ipEYpDXgnCREO6W5lfVqSLfiPDc
qZia6e/SuGTdgjWbqC5/RxIc1iT0KFNzEuq1yyG3k+XdFNriH34j0n3ZAZl1z+RO
LrHgmi6kAFGw0CpE8GeJFCu4X+yjmvgsoF9CwyWwIhpAfz8/3wX1b52D4Gp7HNkB
DjVfMbThF/vJLPR/hhVdHK4KEVsK0N2VwbuZWaPfwJ5sTQBI3882UDW5q4AWFVHJ
tJAdR6V59DteNPRmJMmr5O+BZ3c6mC0eKzJrsambXd6Zoxm+FaqFRbHon0wwuvXH
MK79cSdbxPYb5kwWg7U8g41aI1bMZ54NWBiSq2g5jaGQoAzwAIdWG/Nsb05pRZpP
LDIsvBHHVu+D3oRb/J8sMBlEM+GXkI/XrZ2k/a77QjB7/lJX9Jd1YAwM6iJu0d3Q
bLRC8IiITDZj9dxBOokmpxZJ3AymTHqiaxV2Qf4DOVN8by4wIbaI3Q5ktRjPbbPE
SndSBdqvjO8OrxHS3fK6rslwDi8ufNO6+BlJXLkpJlNjjX1VoF0flpJ3cDRSmCUM
QY1+M3/0/0uDPilqasPrSRiRHwD75lFxARoMsWKspN30ZUGhPUmjmKba+9DbYJ+z
eWN02QQvPzMZJewmx2Z+8RZwT1FwlLfO+//4a7CFkuIwC4te8f5C8pQGLR+8dj7/
PTTVxrcMf6BUNGvlqpfin0bkxsMdSpY7tN8JLfA1bKkrhBuyqCj1091AqxiraL5X
+uJUHY13fYMGIl3mSxNzXQnQ+1P4NLv/sWNLUy+sBaIdPdjlRS6GbWsRAsQvj19/
btrvOMY32juwXp+vFLjDObhod4Lu7WVgdxiRJL/DAonAIPo4mZp3sN6k6Wloxuex
6m2proAKJRLh4fC1SJl1XTa1RAxPNx75VE79ph8uxVrOU3NLuwCjjL3VTEtDjcbX
CQKqBLsupjIwqmtvcCm7vYzhjRfZvK385Bsiyd8lEtg+LYR68baR5YgVLvSO1NxF
PC+Zhl8hVfYBPGNTK9XjztcxLZlWqcqGLvmrmOeRudpO2x9FVVsZGLHX+cx1mvd8
lrdt2FxNaU+OSaRkNRPgOtV5cwySx6FUftQrv7TAQDITjikbHZwikwC0i2XNW5eI
850J8jMuFYIZqTtYsE7WetYLXpdgH82tmlBxlhESklUUZvUpGgF6z5RDPuZ3tNTm
uAwzRu+xSQCnRQbe/iftsIKLdj9RgSRCSjZFgsprVfT867rYcCIE7MHe3CowgRq/
5ovCbAPYAjJCR71b9GNS9occQkUlqjglOmWcNXBO8yHoodrGOqj0qg08R1U/p4ZB
dbi5aHG3jwwgG/3kNzfrnIdifKONb0Zft8++z3OfefOvu50t1aLId/z3ajI0l63A
RYOFNPIIL9qzG19mFLFcgdSjmkYhkz/l6fsusxh7V8THgyOmycimYuyegYn0WlHG
A6vv8GT+gR95fmmpXodQ8HCiSaBFLcpL2HbJqNHvia8Jrc/XHzc/uGr4T81cdQBT
D9nwvQ0m25JEb9nlgHZ9iSBOsooYqHjZmVQoAAfDniWF3wvoiyCKFXQhT6Cfjwc4
o1Q3b4AU0XYxstxGBhTFkjWUMg7rOK8d3IhBXHb9eNuTGfhVIBy3nbGyoFhLGB8W
HVJCdLnGrs9EFescz6gotWDx8J68xQEbaSDLqMopkguR/93597Q6FgGxsJ6FNvGa
o/W46SqZZLzh8os+pm8US7/hzvXtBnsB72eBhkcT57Mbb0tIY3rNJoulUrXbuQly
1WW08YFtJ8i36BRMR/+lHkbY8pmie2zJcvQb1yQLsu/XG4ZuvSreni0VzOqtkN8F
aEK4Q7ruve+pZkZocTY6/cxGjd2U8KzW/ExLRzAZmjFG5ZBUHs1ZQlwAu5akxJ8D
6v8JohUCsbXfaoqIe5EK/6U4+VGtHpvSieWCiWcEfOt2gJ3VYNrihfgcDkz+s9Nu
4JDQk3LRyH04TDm58usLVei66iJytKSdbspKQilop/uGHgbLsEqH5dhb6K4zUM8r
qs+jR11twl8klsI6OT9CMGs7nGx9mVLpbh9/iCd/YTplyIpcm6nCQdjC/YuFHEUs
f8FJln4W7d/R71rdQbpmObiAhjLB9GEglhu2xUrYY9t/4WGOYUBxgd6BBhS1/mHq
TSjfMN/VEhQp2iEz1MMEbLHvSt24Va7Li6zZ9kpIH9khuqI+yFoFazHJZDwJT9mz
6Ex4/1MaEEO8CNg3sxdC5L7RVf3kJw7uaMAcP4DYO3WC+QMg7EHFb7XsB627OHwM
JwgAVkKhEGbGXx1Ej3dODBoojkM6z/X5+4WmwwAsZ4J0bPMkYpXvJPsOEqsoykj1
gr/PazIx3o99KXxSF7ptmTFKVq8zta5WMV/G0r2dmi0aV6g91L+DOn+1UOtRfhVB
WSuSzbZ40M9h2OPF8eBEOri3DuBSNYZJNZDSKIhowyipryXb7P91xPBpFwXNcCJZ
RtKq2nCWN0c/VYR6d00Z8kDYcGzdsh8hwQdgq+Jrq87jEicwFh94xkfOqSnmHTUw
6USgAvVJQvWjVWxXtHGHRB9VWgWjZiq/Ai8Z8+7cXBfFqsMLdjiUGHOswmaLFPBH
ZZmbW58u44DRfjGb/6q97grAtOoxjnELcCWg6r6ztPC1YnY1WpUUCuTAUaFYZIMY
VQp9a5V1AleLlRVPrqDp+p4Grvc8QwOYdRhufLAuCUf8CDzc/viZaNOnRB2MdKpY
5+2a6ubyeaNzV0O6w/olB2+BS5aCe6atAubLwTf7bvUAjv1ckpb5zZzj/BWawp6A
dZdoRP9mAbYBI0YCc+9JRZFfcMRiYzG3+oaaEo6VZ/MlLMrIWXXscJhbwEDAbXgT
sKfYkFu8R/Ha1zcxjvC0+exOTQ9XQESeAig1GdnzFJbALWoSdXZGiYOBEJnVw5oz
LvdcepIRae1Zvs1PcFqkXbHZCN1kXTBVpj2WcQkV7ZDpo9qXiCu0DgmgWEkgepnu
qSMYO+1EQInx7vj2+x24zjPdoH5c02vmAJMRMg0So8OyBK8nRR/UeCDKyaMDT1DB
Wi7l5gd/ZsvZhfPGUxiL6i+iHO0VyRKrg/rGg4mLo84rNVdbF3a0T0zrvtxcqOnK
UB7XobGIGYHRhz+oeqq5L+mzDdkJY2/HTPPTiTOkUvPyvUX+WykuKmcXkHmqIkjE
+GNK5P8vi9EE2q0+Un10UefGrGmhbwFw9of8o/W06uGa13anDmwXr9fdHG+3HYcW
Ru3mtDp/VrDqTxOAPkunQGVUWA+UBcXWbG0Zvq36XOVLd7+CEBpxQ4PKapoB9Z1F
PyHHPclMVpRWtxVCFFZTnDyJNUVUFILlZm+0vk+FpBt5Hh5IwdxQkWjB0tPb73mF
h13x04AWoLaR4NCwgwG8ox1XMwwLmupl6sdihr0LPFN3XzhJFd8ho2LXJ6Ek22rh
pEmkg0uun08yvUR1N3ohkNW2LdP1tw+91/D0l53Zmnbra4rJF/Ew8r9gjv8TN7Kn
6ew9+G5AW5gfG7WaDZtlTcxKkxmVglNS0gP2dAbp3LfePNB5IXqkXfegR2/W2NJ4
klPEsYGJyaUqgW2qI09vmRjTIWdKualpquI3WVmqzd99KiEpFEEviVdlnX/9jXl8
U1oDL8kQeDUXrcYCa1BjlxLtKxdALZVBclVdUWaebYex4FARI7w6c0IFOMyVDgNX
PbO1kk8Hn9mw05IU/bowKEu/JGmfhfTOoPxzhj9I/8EfiVoRbyqiFD+GZKX3mfNv
7N13ER7/0JvHsOW52WsTNSfSqiYJe/MxdNJ7ItNvBHAl7OG/jpRWzL8x7Kyn78z/
XZD942Vcf5TlQqP7zO9NmZq7xMszl9togdL289g7+mMvdoukTb0QDEYBWOHVmQuL
0kJGTma+3Y8XVZbmayWXymYzu1VsRUfJf80J1RraJZm19r6ts+9xoX5VE9dfCQRz
KYFMQEX0sOAHejMkX3OGT7OPXnCwwRDkNcdIhWRAK4YQUZcloFiJUZz5kpOzoyxJ
EIkFwAn88vye9noR3rcD6DH5L8wD8JeyCX0o6xQ97C1AHk1PJsyriwhUVwyvTNGe
JEXXfOOurApr17TXwvBsIiIlIK7NvtjWY5xtFSFRjWvpC5xZp6iXQiI4I+HEKxDp
3dmliP+KwyLRI4OJxprPLvRpik/so44eQDpNFKEHgcRDbM8g1oEQWf93OMGUlRCS
bUPqpswsdDN0lELjgVMindFP0OdchGBOthSwrQZKYLXNDIm5iV6XRkXfXxbm20e9
IMUr53laIl7Xjnr2apuFagbz8mbcM1CEys/F/4xetcsMyAocHU+Y2VfecDkgX3CM
aZCJJQO7x6E9dhFmnIkopO9Nk4G+HtWh3bnWOtpRiw7SCkwCJ5OIlGkvKWvcPoIQ
SbQNvY653Vsfp6eQqRRK+eAPE/ZSvl+6o1/iJVWt9ZQv/a2g/ehu0VciP/g/Mbbo
RuZhHi+GlAnhn17U1m7yDkOA56LY/CclY5wVRVp86la8WT9r+LKUMkUSkCp8qeW6
UK4AYfuO+xjxhxuziMoFdXxH3xRZ/yRm0dZMeFdlwrvMa2rL+PHdjzCWYbIMxBpO
4ihEjpLc62yklL5Upj8mrDlD8dkya37gDdtokhdRiUEX5ZF4cnzxryCXLq6GPaYu
DKMSzOrX4LIP8GIFqbysEgbL4GXEPZUQT+4NalLuWZlm3XP/X5j3Hx66hDE8G1Hf
no2vcgX90ASrFNc0awDfAq0DQhQ43bs+A6A5RZSNIRG0jA2J4hFHdXQH+sYP+0/9
uNQ7MuC/psmdwXBlHayYWzYH+llaeVyz9Hgbb8A+JYLOVhkjADHwf2skj+kRPwhm
Xl6XPLOlefKP8zOBi2TlIOcAUit2sk/MBKHvpFLzxXCKkN70Hea6bVU37ookIvW0
KUi6sAdwBlp2aY1TyZ5vMcMteoNdKjJSMmwtdH3gu/UbpbDXKNqQZVwB9suHbsSu
MsDro0AXb5D3eGXGBEWBjmRNt+nsB3Ww9uOtJjBasANAJ5Yx0eytVabykTRwC3h8
0dKywK/qCgmHkWhNfTUbIxqeOIcGVXCX6k7TTYaDehg8C6MgnnfF8gDYePLC3PVj
yxLVYqVx11gGuABazEQYmlvKrSt8PlAxvdxz19dpL6Viz6/o4GCJ58NvsCqh9A2t
lP0vGWN51w/e4k7DwJ5U99NYcVQvQBLnmCjYktcvyXW3sOfkO1ghfCpGcnwCUa/M
WYMzMX7AUhUI4X+QES/bs61eSzTUFT9gViWyijt8NHbIyO60adst8kbgW01z6Sab
vr5hSJ/32fykWbI2jr82cR1u4iriKWgs+Encoueapyy/D/t+vVMpVTSmT96ZjsQx
KtcDg8o3zs7gE630pHDZbix4bSrInCng7oWPK556veAxlOTbrm8UEUze2EivnStn
9vP8u5TOALFrDYwMDEFm86m4xiWkpE2HKzhi9PZih86UxAaOlARpnFOKFbkCzfWk
wLcV8rU9SyTYSlz4ElW6q+imlSeBYQbnmHKSHD2xqe4uQtFlOiuNo7w5XVHkJvg7
AJO1uDjLDqxNAfa12HrTDkb/QPwYLTueKsOossq+wL/zs/l5Je7AylKAwQeBwl/Q
HzRL6B/DzLigDJam9quXTNdGuuae0dcIbI2avBCCtxiM1PjUfvqgloW6bSzGs/b/
Unz9Z9Hpd4r5D2+4qqk1UX7uPg0XAzN6mrgQqU0RBD8QSMsXMmJOYBEzVOqFOmlB
oQpvSAfwYHqtGbW8khXcRFyGVP9DOeri5ALfJG+WigN12JVgBprA5++PnJtjdwrB
fuhpD+yOncpoFWST3CfEBVHs0w3lHJrOjOrudJ3IE570bJpTO5n6SSAqaKP/+oXb
9Tz90l5YH2KspZN2LGgh4WX21EA4YFRq8ag7wivuaeq/+o+e9Vp7z/wimSJd5eJu
7Zkkyh36iIQAavCNTy+UCkLWcu0jI3ovg6DavKVBrMnQhozhitQW+xTAhbPhmzzU
qLayS1bk4P5dPNJgaWogsl0NR12nCT68oqCIhMSuh5QR0ok6cGonXDllsRy521Ig
ivhDAKA1qndqTAyrf4qDjZjeke7ktTlgGlSDV8h8BRREDo7Wg1O9CTTPDXjzgGhO
j06OpER/Vi2DlzZHlOsOw3XkyFC7jK1J7QfagX787Y7clTsW8pPKnTydxEVMHk33
M+qTrnK6Df30Y52EDjRwXphAtLx9O3oeZnZQhPcoft7ft+Iv1dXID1xOkOnX43Os
+B+SHpmo7DHWB7PW2P8a+M8u0mm+thepWOa4ewqEStuMAPsxEQmlVWRLHQ2/AXxv
wphGBapR4KKb3/HEnrJmJ1tnaug1BqhVlBkFIBvuG9eWI8jR8KyyEWu30cdLJrRt
kkTUT740TLHPuYlizP/rjVO/UQP8c1iMTGgKKgu1BRa4vtVoBvaByCgH+uCPD/jl
lr37FMD+CJK2UTeArIt7QGpZ1Dp+T9ySjKmKr1PVwrmw5wFKYOij1Yrb7QEW8hoT
QUJHQ90+Fhz312AYe7ksYDYbt5xH59qlzO6k98tjJPCYvszda0aMqyNLfCOFaA7K
poSWulNPfq1PcudTgAZ+LBhWVAKwZxvqCLDJeKmXD8oLwe5tKVFokI5Cv0U72Rbt
38lFNgejx3jL4bgkQ+nVVHo1aGRuBF4ORoaXSqLnxJuyxLDgD+54a5ghYcs8137M
y1wWcFfuXrnL4cA0wq/0tNMymFhhL7jza63/WR0rABYBGrHILgySamMjj1S9m87v
tkK/2EUJ6dN8PNouObJXuph1i7xL1xg5FBALSgxYxsb1bRprMYoXUQ73JcTbzhwN
XQjPZyXlcXNcPPllEXbXuZM1bpkFEWrlZz7NgdqmjHnDbQgZofBrjWlzywpil7v7
+1R4FklToJiozngbycEqVB1lKnzx2saGAFXej10Ew6lBvPocePdDj5Pne17TdrCD
lXr52tbL3wWLy6YILAaa4G/Gt+UIOVKA4rpm08ztOPad8SQP8CqKr9p1ZIYFO0jF
hkJnl06FrVA6O3TaX/N8K9CMZLhjk/QR8dp5JAN4QeHTLpmTdeQKJ8nnXXXCD8TU
14DWzTzaz69lwdhjOee7bbdTy/Ug21ZUt6p8JppKs8LjDKUxR6S3kJ0mhYeHwu5s
1G2xTdcvIgGOMG8H7Zw3dm03u5CGSiDTFaZMWqzoHeie8UgbC7oPHdDMPX9LfAF9
GP5KLnnmV6MhSi2gdRQ6KiccF+YNsG/CTRec2TcLVDin6Mu1K4rw4FThcepaiCjb
ioIuRSxsXTNxxriC6HJuLLocxUWkG3pxm6PY8uoAlc5jSKGpcvFK9SiqmfZEaThC
TG901s3ctvqRoTL6QPEeMMzf2DySyF/Tkimr84MEZyYLH9HTaf+ioh6FYfhB+i0Q
gjnd4cNc0DcSLw9MwNjtiSf9Me7buCnaMZMLUiDDOnQAc2FK6OprcQq67yyC07mz
c6iIvXAVoWfmHcKZ9eitOps32nwcRadULXZh8TNvREnhAr2DSgYRKk9yOr6a22AH
+FEB5rbLzTtEKjwgdAMcILTuiW/Feb8KocggvAOWV27rB8Ds+tq2rsjjS0voDBbr
lTemntbalKKHSjx8UMIOe+BbE2RIEU+8HMO6Ki+PM9Ju5URbX1auYgkGOe/fPDX/
1iF7iqMwAlYYX1OGS0u1i+olha5LLlnlOoBgTXVLn+Ktzj0bLn0AclivNHd3DP1o
xe80jX7t5s8sYYZnNYeRM29Ntf2KfC+aR8fJr7mDoTBRuYxksghECQIQTskXuaUr
ZWAHX9w0+Vke5jszkZm60hTMsX3GGd1kXYYBFwyC8SSV268bvIiae93fgFeKZBoJ
3eHCr2vEvxq5eCG11fq0xerdOG0W6wVmqQAg+HLUisKX9VExv03b/FBJCiiuEfhz
TGgYnjxeGDONx6S0jZWfiwAfXwFejnsJ8B5PDZwui9Whm+8oj0sbRHwjowmf55QS
E4Sjljhhu1DH6BjtxtKxrrV2VDqWlQSSvBv+f7n8Kf+1U/8lfMwCdMdsBwxpU4na
gR+SP4jGufeTCOeV3p65P8zvdHTQRwlWkkLM1p8hRMR+68jQrdX/sG9ecnpQbBJT
0H8n2Db9a4nthgqb2C8yCK350isV2jswvEW6knN6ahxK935jVXVPaIy25+c0AxCf
73/Y94JtcoFiVB9HlvQce5tCpbTk8HUIeVzJyZdq/JuiOTop9Ld8HuRL1cTM4HDR
GfcbT2KRbuoISjKWfdEzRT3NfWeH14yoy3QZ7jbfhSV7iEyRnL/JEMXdfRoX+yXN
50P0OHCdebPS0rTceSfYVsaMiSeULBa0FgsbAF/3fGDFFkFxGa5PhX4foeV424Ec
1t9GTbyFBr2HwiN7bIDzb+hm0uk+KhoBOoVgC98lwwPry2qZHtHyUOT62pi+ktZq
gYNmabbzmuAjeL7Aa5VpMfY98slZNutUnUAZGeLioWreI++QvBeras+FCBHX2gpf
QcyJbdzfAl9tP1BIA0iQeBC6xukq428GxXh8RvgWbxUa0hS/Zt1mhabOa8KhQ9FX
c66yqLpvQIpzy2r00QDZ9XFiyryjT3YZ/KSIbbEZdMNLORxzr6FxY23bWry1daeT
Bg8ryDtTkdRR5j93yi/fmGQ7cyPfh+c2UtqBi72kG6284cgeeWxt6nxpF8zmCese
tpYtToHzdOZZ8GwEXszvbINDCn7dezqbP24JtopAZTFVr2E5MW2DhsB0Ehk90n+P
cabkDJAM/sClPOFOXD56LJkF8QW/ROyk1VyHSny3hgsfssm4s0GclMXR8gLRFETH
y/9+j40T7Hf5ooiu6m4cYAHrlIZ7T1CrEN6PQ4J5rMKTw9+C09Dywc1NKwIsDxio
raO0dZq3zCcWPXQwq5mH7L2sMWx8+GWUY4xNs/X7rAmMJ6cNT2xxFJ2xo9Ck3Nzk
sDtbvpokR2Wtj9gyl9IiJmPdm/eKKOjizidv7eShYwAtlJVbmCli7Bsrwd5DKnUZ
kHeI5ep5EqqPuGih6a5gyIjz685q/bpv1EfylO205vwbzMeSgrPoBvxs2O2Y9Cwl
LqqUVcSjYXRMDyqPzFif/2PtpJZUT+pJAZN+gPKwZkhMbAZr2ZlzN7ruMn729B+e
MygOqM2SUJAvgXgZWpCkHCGPiFL6BIS8tD0KL/VS1Q0aRL4JcLTi+uNPiIbK7D2e
dWbzlk2BRpYzFscVWKyqhW53ZgE5tpfqPHyOtSJ0ulT7GjSYZq+6O8MQgGZ7Ja1O
4qoPE6MZS8zShujSBPxav9ywUTTreTMPtXnvuUgDcOpkOtluwbzSInX+o6ppRnf3
dZB7m4M9e0duEIpx1zi1/57wZJ4SX4IjQJSjWzf3xR8GFdbakORaUSJlYShz6RmE
wSlZV9ZmUwBEBhGixEYvlGDJfk8QZ4knvstNBebDmyQyoIuh5rKrCytpc9EFppUg
F1UsKWfn0xoLruWu9zR/7qlnj7p8ARrEcN1+QUhFhUPA96uLnQio8gT+/gNtBf7B
08ZC8DGwV1H3df2aAVG7iRrwL6nRXlgx1iBSdcE6vfRnSj059ZKE2FNAHVeTNEhu
wtQ9gLKGHhgaIqoW4OVr9cMVU4JJxwX18+PGim2nim19rF2eNawJ0KT1a7elMQ6w
xE1zMx9XKwk53mBEjddFMrNFiiwpOvj6Pw48delQgq6+WapGT1qCeHtjv6FPpd8h
Ltjkmt3ubIRaIP+IfalqUh96X7wBhWJlYkHW9EEP4plXnFKmRck/k63B6YeuuVA7
oVx4kEQO0ClZzKi4lVOchK4XvnrR+mUT6t473GNS2hwIww9PZNOYuXLzD1Pd1frI
f+D6GJ/ladF2TX/VNIkmSkEHsA6HK0AN3PaEMOs3DOYM9MGOHY1vOJVbLaY3AQKG
yYVBlPLQur/KYDiX2nEYmg8BRkD+TRil55BhrJ11VPhxVFZMbEc8OOhVtGl1HBjJ
/aWVUhCvaZoXy+Po/x3o0BbSvMwJG3v74J3kKRPRcGn0O564MuioCW3aHp0A7vBh
V5gRg0NG83aO34ONXLLc4K15lF7FjrdcqQWu5eo52JpzFQq2p1Y4TQrINLWXJs3J
B4wGYMhZ5LnfltcYEvQTTtn7HcYBjtAbFm/+PLVtYXESZkD2kIeCtaP9HtKdXVUK
kKqzoRmILWBpsSm4Gnp+z3lfbc+TK6zYuva1/YSIClTob7X/F6ySzy4erIL4CGzW
rGxJqFLdY0h+lj3+ZxI6rJY7tpldppycCZfQU3tiUqy5CZ/+6NjAKIkSUBivf4E8
BeP7J2+UXZqWLUH3bN6uvB3RCMu5Zyuw0p69COzu8NzQ/fxCZIv96Aw7kCp73T1Q
QhuUU7Xou9WyC7INPehOGq/SONHVPEuGD9tiGwQZdas5oiflFlr0nKg/7q56l73a
SHPoZviw0o30LV9WWU/A5S/LmuZl9YjABx+cMpycFAaqlMxy/k79BrTAm4EJsV8a
OUZU11aOPAKNQgC8uEIvzRt8fcUZ70TNNzOvgNnXXSu2QTuAklZxepoZO9KOGH00
bYwAGPg8zmS5D7OxDlYKsGTI79VGF+cbDpz/ILPiBlWm1X+rJRNk1i+VGV/1JY6t
s14g0WA+mBsMTgXAo0W17LN5bUdJ5CUgGqC31590iYNku7y3tPgxucEVOaIeHZ3f
fz7w7MZcG1RiecyS2CsqD8fxpITlBrgpd+hc/2JaLe0GE3SdS2YETTF8cP76m6pM
BUXsZaFruVDp2jmQCZwcpjOcN+K9/aOTUg2ssaZjiDU8wwy8Z87RXSxyfqbYGtSZ
LsJXVCS+1qL9tlPmT2LnRKFdGzt7fb35nsbbrb/ftbMN6qul4nm3WonYW6DzDm6Q
xhofgZ0Em0ht3nTbmAhTQZcsQD694LoOVPM9MkcVD+Hhq7L5o80Gw7Nspt5pCT5+
EclChXsCYdsPdsbrRpssHN3OLTwwz3+35F84cIpZ9iadcNe1VYGukgc0ZNj3gaiO
JrruocltQn+VMX3GbVlqJ+ON6p0IDGFW8/4Rr8YqC3yLAdQkqmbEh9VyWsgkosfd
NODeyUNspxqnGNkuahfHNL/lnNuKjmW6A2W9ZU2444qAq9pM/3jPBTLMJ7gZ6PNX
lBMAkyleHnPMF/z2BOtETv06A6wYyh0t8AC1CfpAYu1qcA72s/EhAbL9HKkCqxIp
uxFP7uUVmZcuSxDEDSrhxYLX3/v6MOxFYqGWXRQL5uLmIn8kAJLtAK/fEXZDmMEn
W9HZHMwRJTMqiwh7ehpvMhiZKhMEntddfum5jXxmz0OaXC2gfThzGN8/KrQ8onhf
nC1OlAuB7NzNFOqvvLybtfbYDmgWkGGP/WSa9OTzjqur8E7MHEL9VQU+qtvs5xiO
qctNg75R7fVdB0BL7vvo3YgWSqxQZVCFaasqtP0kFeqkiWWo6J/ejnHIGGBbU8Ez
tedri34Th+skBtqZoeotPqjcXlYjME0Ta1m4aydlOaex4KhKg346J4XLIfYesik/
U8QTAdSyyNF+1OBgPcWnZzjQXxSBIyTiDnPxAm6maFLbHi4MEkjgJaz/OVKkkVTy
m17adU7jP1OTw2jMnmv6ZP0wg4GwBDdUrXwUnKOkKM6rZKp1zVzf77/GAXgtoPic
9kHiQwtaNpiQuHfNG2PwlF26Wv8GKOqagX4AaxTy3uPPO0ADPMtuaY4MTD9tScwE
PUG/Wq1KF6HEGGe/OZKct0/AutizcwrcovIU5cNOyZV6r4FzGWf72v5wqtri99fZ
03mO7xM32XZwKIhvKTla/uyqORuK3WRbVhJAQJZio/bk3ybvnOWPBwXf6qcc+QBM
8EBJXscR3ZgRGQkEAPIUdpc/5WJ/mbUrpSaTAneOcG2oTt4gG+bJy75aVkIQQTkS
f6bitSNxivJMBVLx4kMCXTe+Z1c4eGrmNUHIzEtMIacRQtg/p5Z6djKd/AAJc3TK
PPKsvrIH1lKw4v/KX50DH51+ODA8MbnAVUG7AqWb3tWUDfu07Kjz6ESsOaFXAOME
+A0iS+cVERY7MhPT0xGHkw+/7klhfr1wRffH69OSLmatOm5FvkkLnZmLsW9MqxBR
HBRdUbsx8GNgikN/nV9CHfI692e3DB/Z/WTc4kFzqakXzMZh+Az4TEMHh3dMStCK
NtuaCu36inimTdbjBJf6Sdgl594zV5AubhmgXw4Uh9IUkOhVBGUshof0KX9Fop/p
Y3QY/f3y0twuuCXOw65OsY4J5oTwoK2Ra3JVKvgmKIUbU0LF6mpLdqAezl7ybN/m
SGIpBrQqzJvd90AcBy5Y8k5m7/hARrAJpHR6hQmwk4J/e/SCo+rjqFzH5uFjDHWV
jxULv3KlzNJpyHKbQLE1LmmGNVKfkM/3f9ukvAZCpY56ZyBD8H1gosBEgks4W/6l
gxFJiV3KcCRGVsKdczsTAWnv63I9GmSGhgLIDIaqDPAP7VSUVRFKQXhAjpAnDpVW
it3Z5hlsBCe5s6Hjysf4va+/4vabY0xv3KvcebvdIeGY2Comjf2feHXgbAOvsAyb
fig5XqD+iK8lJxbbUtyUYCOdnDNVyGv6AWidSjH/gbvgbb1kg1/AzEwjzdZcKXP5
4QFqPzidM+vvOO/+u0sL3S3zZKD743hzs1NRK8Leu3uuXWb9oTUZy9RQqua8Nyma
Xwe8Q9p3yR+g0G1agCMor09sl4Qzy/JRfoKJgFW1/BujA26IkHKyfYsxaymKJfoB
B6rWdtnvOTKAwnsWJ8HF+4oyGRBbCy3igpFw+fPYVy4TRf2ChejFVSMMMb3WTjyf
digMLO3dGu8VcCEtdOjxVW0ixnuVklpJATEwGjZJI/5tk03gNxf5ac9gNOj4gQy7
Zo+IOsvOsXgnhCp7rj1/HTq7bN452fGDc7c9J0pF9lgX/4n/w7o0WJe+9vZrCwG4
2nJoSwjUzhHrpJiOc7BZJN46td3F/uz95AYKT8c6EPMoQHuQ7LnFGWzL03MZCsrf
6EB6IoR9bBi1Ou4P/G2m/d1DqiFUoYtiaiww9oACoir0PpCwrA14ul7Tq9qZbRXG
0c/J2CvOkvrhRyihIU1+3AeEs+UmMrJpJJ6OAV34SfnlsZMbTA3rWWbHKzwojKZa
pvDkuN/BZGl5PRq14CdCDMKElK5L7X63OvHd5T+sHWQNmT5lXbA50cMYlBjJ5xf0
u9xWSJQMYUSnFDunpAtyDjRZiLHLCL+eJ9YXsrsz7saF8sA3x75hNUK/BRySE0xr
4CsepE1ARzdc2zP8SIcqTTejInzK4w8UOiMKw+q67QAu9TpOTOvIBlToqWrg9iZE
bEZMuOm35p2xF59O+vaJbZZXbhJIxOv9DV3hfc/00/uYHhPts56BskA5kQmcpF0G
NaVT9snuIMO9OhOhDrSxJfLFKTl0EH8ZBMT1yJPr+ixQ+qXYHkuaVtFbcjfcSVnn
bXcirIRYnxWNfv9KBwue1egEyj/o72J/YfdRy1/XJk1G94/OiKzQBsv/tqvGxdTU
HQzZfVej//z3SS7DktJRPWm1Hnc2wrnHQ74FmvaPaPXEQT9Dl5wy+v+sMLDic55l
f0yn82M9RAS5mW+tfASQjX/GKKivnb9kX5i7niTE5+ucZroXamlDM3FKanuN8Ywe
dvJDfPMc6SgcB4nI6kIdrW2uzwxd/TsSBTL7NHd5vlkwJQua4rfXaaO15FEi6DHi
HKrXTPFSC+7j89DJOq+xZxrGwxAGz2hqnyog4XuIj0ItqHbmZCjKVyA3hBynT40z
SvhVWDbU1CFD5rAK+rhqZrqRuGd4674ge+Vf2J4KtOGRuiKaSjORDqsLjhNl2rGu
NI96PiiwBpVueQZu23bRZ08n/qMSan4f3ZevVrfypsyM/v+Xehqol3VvAo70xt3O
cekZyZ4kQnB6rrCDa4ggg0AoAdIgqAfLKfXPscEgdQZ4lHp2/RXS7S45gL2BxXaM
mDaTcz/ori+qmVoX49H6eGd2ekXJSWrv/TIt3EsHcgyyjJhuBPrxWI+i83CUi0m2
jk6mjxyqytnJOaeEmUCVmcWl+pArpZgN+CGuQunTdMwePL1o4D16GM0bCOiK/FXe
U4/3iCykzp05+HyPU/wNu52iuA3ETRBr5SKmgNhXd8nsP0eegn3R5ZYUniFZ2RUi
nWsZhgJeE0m0BkJUVBJPE04ifVHyavVG5F4ycqd6mh2oIj68sqg+AroR2PyQG5ce
w6jrDU7NsvpnG4IfJR+dMBAEbGjXwZf1YSXiMbO2H1Wftw6VfhzSTrZEzFpMVVKP
TOGxjnY8DPbgZSSQw3VCCY2N719fvG6BQk5/gEsN45JTRocRShLTebCNbQOK434h
PIL61hjoDIeORHFUCs36suhQwtH8GqilTfop9fhvOmsfJ1gJQZhVdwDx/yTnB+sU
uhrL62rBrr6wpZxeX4Xkw9XgAWqLQekYi47Sz+RH1/qh3P44vkjhK4kTTNKYk8kH
aBAZBOzE+Eq+LnFsmDVsfmlZZk6GzdwdeBSValukRciO6EMbQ4v3Aaqb5mJlPxPG
bWwb5YTptbVVACV+ztBTKD79Uwu30rKJpK4SNc74Ee+o0Qxe7KHMoxiGpGp07yx1
EdmisA6rad9x4tCX3/JRR9vt8tirB7P2s2YTtvoY3Uas0pf0+vLKL9+9hjmH4Vq1
pL+8wSqesrjba2soyX/517s6rUyP58//H+s9MsyEg5Jk88P3cP6OyOgpBFgs3gnD
0ZRn2YnAI/60o/6oVbPzyDgFUSIloS+I9sEysLZnfOqsFKN20Xjz9SEzZx5LaTwp
zKZKz7d6Fgo/Tx3JzOovr3D8fhIhRMynM3CrnMggadlvarD/OLBPWTETa6C/1tBJ
G0gJEQ0TS07OVpYckWRX7wD8K63xXV9aMnNG6yk8NYId2kC6Z22T6nzWJpVdsdKb
nJ01a4tyrMU+AC1jy/zjgHl2oTcAhjORQb5d5+sBLO8QXmXrcyxvVKbtg/aDXnaV
AlCgK9ur7PKfFHGoS4R9QBVT9k4CnI5naWUeyGbCjHVoKWzbGlMKEjAiLPiyUbF2
W3nuiccH4Ej+gJ75CY7PcL7QYZSe3MA0hznEkF12o6l55fjl/PdwT637gSOYZs6h
zJwWUX8AenvHsw/VOtaz9kX+3uchCorPITslbpS0EkYs/F/7szqaE5Esap738rGQ
EgzOFMRNxiZ97LXirW9VU0mc2IqJZwIVRFOKIGUyRtI0vYs+PvjhsyRVkUur2Z6k
5nVInXL2i+AryCpBUMRSGFDwPr5Mynmrv85sWxJsFbwjNgEkVaF8ngw7mTWid6BX
rNcjdIIb0Km0qUE4uyevDMW/zNclimPCy4oiuuEuHTKXBXs5ncUmaiSwqcGlNKRh
wNNSrMxZeE7qZEo6FLv9CcjPerFxuqTfSr9hanuE9JgklmXUNYbXHXxW89vG3INv
AAHeQOs1KuD6s1StGTbb+3rRSKKyMa0Xz6OeB4eSlaXiCPmIUZ1UbV7xcwQZLuss
80/XwaB0XAA8Q1czXMk0L+JdrPZt3kfl3I1WGSuVM4ZMsZyPL2tWCZPBPvj8eg1l
M1YqjoPGaIzdolXBZpGwxCgMKiIDW8NrLyoRbNixoLf25gQXAQdc9N5Uw0a+7fd/
hMGg/imOmO7ijZ3DYWcTcWpqAido//QW1Jc4v4/gSTqiTkjqSXz7tKvJdr1DSgWd
YmC9sTR8xaWmY4HBu3/PyzExD/Wj9C1bHRU3+eXtovbqxDj3qBb63H3ElsBuUBhG
8ckUn0bvgTgD8yl0Axu0R81mZ3YXchoeJOqT7QbK2/DsjIRAcTD2nV0junH2YE9G
vjqffVgfkohSLrbHI+cNnDzLzPG12GcoFo8kT04CGzuPX0Oh93itVkDuwHtn5C9/
Oi7IYQBRd0SM2WTXnMN+TdozItzXIM0iRrop/A5yqLvYnIpbmhI2FGYfswxmeieo
ATTx53Dw2Q/zWmBJ2NFEBZ9EcDg+ciOa6kFqtGZ4d78qMCPZR643kwYe09AN57qn
8KM93+5gsUwpGxouZVfurUSJjRrynaBT1FQItW6xiysU3dh/X9bWyBm8K3iPXgDT
uVGfBsvgdrr2IfS9vkzWhtEG+kUXcfUNYZYTnvNPgDGTrLoDMCtRFbnKm6vWdwnn
etasjnDKEevGIHR3xdVfrL68jTFNZNpx/g8sL5JbnS1bJBVu5D12qqwy/ppDSN/P
gf5eDbCzJRNEfYrECue5VMWQl9zdRByZUAdMkovmYvaDFA4yka9QNmc4agNUUqHc
UXBVyupKiSea/lJvK3rqDmYBVJxA2YzIPbaatPRfZVCEQG6HrDsR+2UEdcoxI+fw
aEJvIRy2aN85vJitBIZzlIq2qo17JEfZ1vKxEA0xH+GBylszQa5mX+jVL0nzTx5l
nhq8KFT2HaOHOy/SYlm882exNnCjJL1ddJi/DgW2yEwOaytOMHPa5QDS3mAgOOWm
SP30sQ30mtrTqObT3iyJ/9auo5d6ZMgEl2WGqVARUQrqSi/kHDEr8XQXIa6pBt6n
Av5AlAHyrvj0uEgujMOWmjMil2/WQjZtw+vzdvnJ4ubWXg5HOQWjUQ3P6V7KVZma
IUYiw+Mk7DzBosfwhDD0qI9jUJtgpj/y0lHBsKnUWQdcfy/dQC51UqBWCGxr+aeE
xugGah0mT8q3XZWiJV19JGmj5DySXOHzRYqb0/d1Aga2IGz8/5kfQcXyyr4q9RbQ
nUA0Gm/wKN9UpvHQq7WBXQqOR+uyvcJbgS7uS3h0Xh8PFlDSdnjJJoc1xcyuzD++
YXltJKPo9Y1s15lEGfW4UZK/8EK3BLAY9UNwVYD06w3Gdxuqw9u2tevxHbTyMDg5
Tx/HOlQ/caTB9yPbxcpHqR8QVTIENnyyijy66cRPTAJFj5aYY1acSH3h9tjMomw/
3SmVXy++GTiJ5x6533IPbpLs4gVSkC4huMK6dQtABkBPsBj9Mi8izE3FmF3mObbG
4ic8XTha9Xh2tDOkXSkIVc3BXm+N17kd3DrW/q8BKn3v6CJtzHhsEShQjQNo5D+x
QQfMCnk2fb9jmExlV4dlgjewmYFgAKXS1+BaS/S8XFs9Ic/QWUfUTzflj4YgjRhq
UTYkHFG/K4aDB5vloWYMxmgv5Tt2YcKKCL5f3Kx8P+iWH4ugiMEiAB/rWURN7z/P
0WQzEghxnqF01ZWCRgP10BbkmRzZ4p/M8btxTNRyAWzXsrQMG0qwHVPHqOjdFTtq
9UmfOFH6otPMLHPGgm0y2kmQvh5WF6RT87idbg5iRhx5Pld8uQVE/cP5WY0ZwdMb
p5fBe+Dat1LNtoYZqNdUf/MaGnLEf4tFtAU+ipAUgGNKGHlzg6l09uzM0H/GouJA
9vNVYXHS0VQbFArv+ABsnHynJ7mezaCJeaQ1LU3BBSzGSRrZXPJckr+m5M5Vsx4s
1DZKisv/Wk5PHvJJbuOiymuZPXFf1AOlCRq++gfHzgOe0wxt2Ew/buf77mwH53Ld
l+ir+PB5hKoo1g91/zbg4uDknwlxV6mpjgwcPgeOHiw+za25aqXMywPj1K+zaNFn
kbEr6w3uB4KMaJwMvUNdZ1TrbWDswO9r+YOwKMCRQqwm51eNEmLJBI6ifnBK+e/V
H+cXpdh7I+EcbKGH/ZIygqhHZpHoqdmGXyWsZ4Ux5Jdfu3OEzkflLI6uEfy13COm
3C7U+ZRi2z6NB2a35WWuSTRxklSjp/JDwEhzqnr7DpxUE0y/ema4dyY9HBvtin1t
GFbe8mXQx01V6/0alJKNnzJgp/Us/AwTYHPd0SVv9jckyNP1gXHfkz/zAqYFMVl5
0nEpn0jW4myCkSRVcDcBeO0iTnfvF6n8xq8o37q+uva4rzMoa4LNiFYcaDSPJ0vp
1WlpKRI0aP7BuQlrjZFy9ZYH8yHkG1Es1xRTcn58N36tbeZcSNdakJeTNjL6P9jm
D+PshjjgZgMfXnh9R4v+h2wRVYzN8JPgIX60FiIzO5lE/WYIwOCbsvCvfceq23O2
V34akN4xtH1I4LhORd5djtBdSdUfrO3B2DNNXcvyHsB7Er6oLhmiF4EPuDLUWR5U
TVTdRhOnLPyfQQowN+D6gXhqQj2d4j2sU+HBuOsjBEjF+hpwWvYlkvnCIwCu5o5b
E3SIUSMJGRhbtGa0Ju45wznzTMkegyvZJyY4B9b+RXDkZfI7kcNq/hi/XwvdmoO3
HpROBzY7cYgeVT+8eQKVFGFCRS/EwE8c4sMewhBTnupeMWaI1D+YRFoz+Pol8n3d
+kw8lOaSKCQyHjlGi/nxUiKAPIhyvCFipCgFlh2fmQDte9mpW2TUKeYZrZrVmk/m
TYVP5lCpiUkam0HuAZlurNnsTdf6Ii89FY47mWp3nZEilHPjkZLJuHXq2cHnJbt+
wGMVHIaYo14UFrMonjUyAr3tyMOzWWMlUOnXZ8nxz3+Gh3waSutb/BEhVV6yJdus
MaFVrRfeAu78GUUKfm32IjVhe/UU6q8aTxzeDZxHJuNJli51yoKPbvu13F3NgER4
xj0UJqwRNXiyjMbaurfUj23lPiJZwKeDX4kiaexQT2WUhN5riCxL3RtvOQ7Q3jd9
l3mf+XoOfl+2Q4Zw82gPQKr8a6bmwHUU/PvvVzff+yE4IjGYukCqEaLSRoIWa9EM
foF3UaA2ZSX0BxaGF/v19Kqus1diYM7wCtkS3WGlCNhiwxNpoF9enYquLcKcCZwP
tSALclNf4rKKOaJt0rojjippswlp+IaEmBQuQ09strwzfc8hS1SnBh0iHHt8QZjJ
rz/7oTChdQZdJsy1jSoBNI7FeRkKc+BgyJlKWrjSbxshQWTEcfUzW7WUDcpXskKp
WNR1OyWm57MM6I5TMt5ZWAJdIMaaM5FOxojGfNrqi7Tb9clxkCgzcJyp+DdjYVab
S8N5+G0nJ+j1K0BdNjLEBaIqVWDUdF2Rd+U/ZpT0pR+CrS0ad4+mwGo8U45h94/h
L3n0tJOxtoiuoKq8vqv1Y/i/49eSTcREt13jvvEd22OPfEWYgyqhGFe/9CJjU2Qg
VgYWSp5U5yKlFSt5tBvhmpbV8VgWz8IMqyB09+cevfUQ75QLRwlMWTznLorDiDE4
HcXGwTVBLHaA9BkY2MhWS9YW++0VqNVzUhNfPg1hxE8h15DE6ZSAxrbvWGuGly7/
7RfaayY0NaYd9/L9P1VcT8OUKxkp8cFTnOfzYgsfN/9u1Qiph4ELwmwKgfL1NjUe
575rdG93GGiMJQYPDMphg5aLwKmtBenQAVo/LDrzrHvNeuJc7XbdoX9FylhB3e8S
fOSJRtPjVk3N/OeETI0USUzrLo5Q4EIbtBdplbPxeeEpa2vKaABicZBhQ5hAd+hz
RGDgB7LtYTMNVQPJbvNNSXizBGo1gqE1P4u2lcpdPYbbW1Qg7nQZciDYmgeypUv4
f1/UiJA1v1EioQYfk2IMS3Y49VDvPOqeqpbWtv6DKjj3gxegqJ5brfj/yOKJ9aE8
7hRJrERKXKEJgpJOKQCCE5u/o/PtF5CJCoxGgGnqscg4ZQ4O9dHwgoayO6InZsll
0sHwiHsPjVj2FEheMMnNWOeXsts8pI26jFXiRnHDiChEjh6rVXOeb/Fmi+IiBQMc
okhbMkn92rCbi9wnYviKQI4gjiKDuvweBgkaZfenib1Ig2vdCk4MQJ6/qvMwmS62
vwdnNc14BES3Dy5EoSfjKyXejvoNaVQyg4DvlUa8JRtRZ5+tWRZqEEbvvN3VG7u2
cZ+DN77PpVNHEwfCMeG15/SHHcjPZ5nkxnO568EgjDxx3SnD+xJwO1aSQiMEGWed
rncNdC74Pay8LuonnjK30/PMmKaJyCKWCzrCF8TxFKowoxRMRkrCQxNWaFEtk5lP
8ba2euGCEFg/9rrQYdO04GqbvjTMTu2QfSzeJTKw3fTKL+bZAVT4EAYz8GGTQAk0
bYL409VwIKC4O1qyeUSatWXwBznGkG5GxuN8VkvtvbIfwhc6nXHxF/jDDfN1C/LP
L7OTIirF+SoEUl4aMSDM38gPCdIw+sedxRxyfVBeTrFZ6/7QX0PVDeTogOvaGOmc
XW+B7y5r7z/rpQnOrbQbyxDUWR2qAl7e9PqMYLo3lQHv+A6ulEplKBSrX/uwzI9Q
sIc/BtPo8xg+M7Er6JpaQo+oVXb7UlybX7DGo0jKbguWLGK+vqxPDM7HLgIopSM/
JNc+Np4gvS7NL2geNGUds/TCbUbDj+zZExb4NB0ROQ04ouJ/1EP9mq02cf2k9nz7
XKrlsFVCMqpcshfsLTsyaMCeG9edT+HFidSqHN5kfTRtub5v0AXhTtF0dspQ+Orn
vNmxFQYXG9kqIf87z5Cn+ZfbCufbjyyBg/7aJbISFJNGjwkfGCsSJz4ilTYMMelh
22Gkg3j0NTLlBqo42a3y4ZmSWiG1+WA5kpA/NN3dhzaE0CP4A4DvzJKpOtvLsYF3
23y0PxNmfSuPcpCAVD87g2iwPyn59JyNZtUGS3ZiR6k0gx2roaFwsdro7B4Yi+iI
LyqmQycfA5XPxHglVqXut1+PTsxdg2EWH7GKeygdpmoDphrJIceizZtqscdpA0gk
x93mvb4V69SV5vonX4uGbMWJKVEUOUefnwReowDfwZTZ1DUGR+2j0dzOU0itLuzx
NQVSbVgMiX6zR5XRPnra4tPGINTkKzKSka8arOPWxoSY8KgM6ItgSWsfbvSqTlVu
XrsmZetHmAybgJhxnfqQqqCbggg+mJ033RuMzQNQ5z4Q6ZEveBDmRtsUG/9WlESL
O7YUIdlooXe2aMA51UbVW3lUsdbL0T7pcDTT9cYg9+bYSMudLgOmlR0Vw37t/k1r
pFFyhtMGZEEknBNlGL6T1D7SCKfD7qliqkhVcC5m51LxqT3VB9AHOf4bGG4tetuG
XJZ/u0XmLtf7F56Pyccalif7yThXuVGw0f0FyTe6ctJU4IRVxWmS6D6YUIAjQtrk
ix3HIYN2B81maTe4uqks1WWvmhS5SItY6FkC5oTlZDIXMWy9Z9AIah6WQN9tf8QN
CuvIjI2aAFB1uwNQpcyJ1Q4nhyP5GZC/gqtWWhCCY9uOzyvk1JJ/v/5ftdODfuYT
lOMAHAq2WeEmEEZ1S+KeStz9Dr9FXzZp9B7TfJ4LGMtdddi/8WB0a0J0C6wVMD9Y
lsVVht5Lvx19kCA8sv7JnSnQxlk0LKGqd86TvZpUfXcEBoeIM3tYAlyUC5HIYs1h
U7NKyOCvHbQalxuif8W/O1iRCR1H0dbV986uhjXodH8H72KMOX6ItyYxGrlmq3vx
rBUWPS2sb2u+b4TmbLbyNOr5mxnLeR2aoQgh0nD4t6bzIYFNh6RcM4tWEpP/IzuQ
HDE2Oo3lQfzTgr6Ga0DJJ29kiMYJ4sBJbsZyeKc90F96IXQv6LqosYtYqXrok832
g3fQbDyZn9QqOn4g4+qTsVWfG9oE597vHwXu+iyYPJG9wlUPEJoMKODPZq4xwZTG
pT/UsAqrHf5ykARZwQiENk39iB57rq5OHYo9B0nvK9pl+rgP2yo0NlJ7Uie5c1VP
hgi/AifyMSxjOG6f0bgZEe0pk6rUsxGb5Wce/R249/1GltRBXt4z26wsyILcftqN
HVUKVm3BAwBLZoIydxNNy8YpPZHQvXq1ca65gqLnaonyF5cft3ox/qPmKHeKZ67L
c5pXqLB6xgyVLo/DSYoUsHpTTwjRKidr61pfpBPJHzLYmbMvfGO2jX+ivOBtVGjG
iNdUZLacYUz/S9raeqmX8FwF5xF45a3sK6vnF8o7HLB1pnSKJeyaBV/6/gv9HOph
uOP8rNkPeYMQXguZBxs0grO0X7/4Pg1jRjZKDpC95iS4f0/DOTsVAcKaDkZoeIvN
otZVn4sygVlEYDzDiUtjSGVCVpRNN8z3Fk+1ZsEQF3g+UTqxbbSwoXVs3cp3gO0N
myVErNExMSNu/peqwHEAZiH7QSms7cIs+tvKi1BccpEq8kMv8TIH2HTROJM0nT0y
AlBrke33gvyGxDtulxC6vcN5CZ8db+cuzJWUikGAqQ7qvXbF8j8+MMzIHWjMatNI
HI6FR2XZdoyKw8oSoNKMEuvDTONtYjteWgHXdQ2QVAhvHVJgqh9By8Xkqe91umlP
2nnvvYgUGDXaV6IUZsGneUXOw3wimDf64hajxGfiWoKDMMOdzN6Zd59VgXNt228I
zPFqWXGE1IdxloLCajVgvriSATHN5DMSW+F19GGQC6S9InmK1UlOCw7gOq8KefYN
k42mrvILiJXT03NXnpjM2140cOmGQf09Xx+NaUwLBVJ2XLemda63vBHAXXAY2ol+
FWvSJKW4vJQTZ1PYzz97WQpixBUuB/K0EuwT3NCtEdoQ+bRNE3Hj/JNZOa07Ze/j
veJ7jn2Gemlv9TBazGnUS1xPR8EslLyLcdNLWOFHNHxyVWaDazTtg+Y464VT/PRl
OHBxVOlKYhzqB5TNdiwf2k8+TXt99XoEnq0UWa0TH1GP6aYlenQqLlCNyk8LOMly
StK/nfkSG0DBKSca+n19PBch80G3i4u/mSnpkR5Kx7XuAMpBgVef2N3sOYILfaLC
naOPLKPFhMuDGG+oR4gNQGkIQvMn7kqvzjOHyqsOsGcw5+vgOdcVRiefIYjmVHk5
jFDZo/6iHcpFvLwfo1MPimUl6MWBIIXUCDyiI9UcFIGbAlso1NK/qFwrNN8CgzNg
ccTLJD7feWnChCPy0IDSvdD50WiZew+X+RkJ21nUU20YxsVOApNrAG1w0n+42Ar1
D2IYBud2cY/vN6ectCHOKtsC3ylAgm94HGZ1ia8UfbzSjoJFkUg3cCePWMPdgA6A
J9UoVbu3aRUdjJzJH5cpce6vGanzVm0WURCSZSNdFccBP2PMpsnqdBK1Qp1f6ays
hdmp8mtn+u4y8Yn/ljds1u9BnTK6WHXJSyy8IuVe5OjyXoPvp+YB95rO43vg9k0h
lA8hH5sm2QvT12IRuTI7Cktn04qKDbgoJZTOxKWM7gA9+woTDQSaB38NbedtDjBR
2BZl9hfD3s5QeGo09A/uIvaa/fxw8ySq+/hSEtRezsq6ng+0FnRkfnew2kuvbQhN
UZ92MtX93cErcsT+SRhHHFkjzqXnhrYz53qRTXWy8X3Fs5b+s6iGzSNSjhiuhOz8
DBxZhwavK/YFzpc4bN9NFrjCx4tBzCBR02G+8zKbhT2NdCfhtS3204D6uinenOL2
AoECjvHGmnCYdir80pI02wG0UJgk+8mzL1h8zxAZCX6DHqSkERZe6WLS07dsD4tb
8ICCAHfIX3AltStRhcXNNzLzjFRDcITrS+gf2ial48gKoGhMplqPODDB4wE3G9eu
ALgmaFBgnRzT+t1dD8GBYzPwzZQhozRrVSpc94p047kyKV6dRrMLe8xXp9tH85YF
daYty4+TNeeH4SagKP5Nd1scejAklTP7t3/bgvv1AB4f7rD7Ob6R5/Whv2Otw1Cg
txaoesdxlIiuycaqHdAsUrKDqTkl8f+9HP3Og0YdC7k+ZoeUWPaIHwJiROA9dTxT
rMWsfOkV7TIoyDRmi1NuMwrPFQEv7N9kDCUpc+hyRYT71NDoQxxM0quibKw7G5WQ
CYmxNM9xwopKypz+rzj6Fu0MQKft6+rdKBNINrxDuE1ZkPqLUrfGbMyYEInUvkQy
hnNmlUnNJrkhRvY8z/XLuBWsnXisMQYl+5NzqVOwPSqFJmgjXEA7KDkG2Ki6NUKf
QRqXZQiA/FEICIlix+JwH7Vw1HXI7YwJeTX0kKxK0PGn8LI8tlOytMkBAxXuj2Eh
C0779luo6AGByS4Nc2H9XtMJ/CwSvff2Hi7wYnyEw5O+Lo6E1Y/yhPcUKKwV/ieh
tgfO7uCRnK5VRmNtiQIJjPGGAoJ4mIOVFVJ//3+xn+JEblXOQelgFnaSsQaH/ZnM
090EMVHaGcQZNf3rgzPjN22hfoek2pVFN2GpERovdId0rAIavR9sZb9F9Q1iIzaw
kzR7tmRmzC6HtvaRY/5pP6SxaXRUcemoRsvfSYq98d71rQTOyLovgNmv/ddJXSqL
cmWyXLaltOyttrOeAvB1trCO7AfujAgLaTTBNfXLdyj4azmVS9dTwSG8CEx/A/Eq
hMw1ssQOFwetE5z8mhZlKoz9iFb1nwuEtmLTcfU3ywKDEcaTGklXZeHOuIyi5GQT
qfOEKDYDp1Z7YNwVtquNu38cVfw2Cc67LKax39PWQQQ/66vr6YpLdQJ5sH2uW1/N
ccGcs5WSTymcGv3JIM+2TVjnUSj3ciLzPHk3/HEIpgsQMyXw2tdCVy5MZ2cyVS8H
bJEuk8MF8583avebCpqKGNX3YsqvaHCtr1AukqHb2rnrqMu6JM9F+/ec2VOoM6RQ
k23drZ6qNg+EqZdoShf1TCUM5R0UjMAZtoWZY4bSctVFaijTapIj3fJ9Tn+0XxJ3
a3jDfzN5ScHSydcG7Bj3tlSwKOpplsynpbxYxx2yKz/B3rUlr6hZ6Ml3kfNW9llz
aaV1dj4N8vasvvArxnVy0Vedg0X9/xO+RNQ+nHifxUHw6ICoezM1tn9Z+zUdddpM
S0ZRKwtDiBvSlq1KnavtiL037KkuR51Yf1Mb5AJgPCkFSvVkeWnCYVKHxaUhgl9d
8/bB4U58vQeGvlWq44Z+2x1fLpBhzNYMAa+GFaMoURkcJNQdWOEaYMayczsAYO9F
LRhpESz4xYmC6DDIMNl/shvunKcXseznDsL/CLyo0pnTziko18g4jr9eWcV5OkWA
fdyu3YR1plZw6eaQ+A1tZ8GQDoelONUCjEf1ufkhfSqCfw6QoaO4x+Uy79Sj1OVP
36hGOb88jYNsk/1LdVLSZm9jqM7ACV2R6oFG/I3QfCk3q/huwDr3AHVBM97VK55u
wLucnWcsoDIvmS/EyLhrojuZhrt67sSKGmotCSTzt4DYVPCT+PDbcsrODfza54hn
iC9BzbVNA3ZUcUbgGSrQJjD62yOqd2DciwOkfns3sFUNecjub/xmsjbWyjS5Z1gG
RXJ6/SLepPoXKu1sI0CT79+7/BO9EOtv2uHGxvt5LFZs5zxbC2F5gtAyDL0gzUjo
LwZ/2lPn2EVyRGEjrbWe4VUy29Nk9dQjgXk1H6Zq9ScgkMS8fi6mocXyhHjBv7cE
ffUumCoCly+AlD5rEIxiZORvug6N7ab+/e7l++hPKZIHm2C3CzogOnvvt6KGjZCn
XTIp9YrA4EkH3LDRoaIXW/5JofPW4OHVnG0Qi0tq6W/bC529T/WzEGgCcwtl1rUp
e7EZqWkom80lYEVa22mAZSLPPG3RTiQF5pXKCXblvITvqiZqlOFgUKWx1KUik4Jh
C64fr0SA4n6J4zyEI98uTF5ySEVd0ub71mMcKCpy1KKNnw1eUXRZbhu+sGb8sy1i
L0JXJ9JpJXQTNJdd6qlM0tQqVdiaK5gv+EbJs1b915vPB8uwmDm3kNdnmxE/QLHq
9kRIAWZkxarTfTbWOqF8SvYXKl8uzn9doBYMxbl31QUvqlGW6nFec6atqp+7LiTI
uX9LpRiaXbthW/l6cmrmvyhp8GHKWSP/70+uitzNUc2PxuX0Syr9d5ICVSru1Og3
/Hr5VCFsADiRCsLbVr9UchaO+HFZxcGBSL+9GQEXJhlTDTCDTYBt0b/9eyEigd6V
JiXk1WExJC05Lzfnan5SONERNti2Sju/1xboEihWN4pqhgX2Y7vTvvO3IAA6Zd8P
78jGNKZj4LkzBO3X7vRp28RJdr2MTzYTzx5H5Yl7M76q2lP/IMDp0Q4lS31DtK95
OIri5SiHLR+a0kPpcV/DYlpO/692OPpPhWheUC63bZOz63WsAIPnA1U1l+ddQOqk
VID99aUPqpgjjinYOsdMQi8S/cjHxjS6lE5EVwefNzaJ6xVj9A1SEpr+z0giC75w
kCD/rCRL4NIxw824/mKoNVh918BksII2Ykd/vpfOV9dWjV99iJAAAHev5khSExyz
xhrEd61yDDcbWKgHCMNkA7nqPAj68VQDNa8C3Tp/mAm0QCxjzJ4dyRR3iQloYenz
laqpRtwRHDzQeciqRij7XB7XTkBckQyE2VMVoCJ0ANGwJhJ0h0n7v1oR3VJSNP2U
XuRVylp022+oCjYxxptVw2qFiaepFq9oVxNcquFvPmKLK/RVjL2FJCb22x0o4GR/
mumES4ZZKN+t0kpNEK8uN3WBotJFUVu6wxa27F4Y/hCYFJpSiGzOvVIhkWvAn6j+
FThDH0kbu678o8sK/071nE2m0K9Klyis38RkzOW9o/tZHbLCILnwxShn/ofVxLea
LomrcIi1M46ctaInZZRCAqCt2BXFo6AtrKr8qo0M2mEObicYhz/5GnNvyLdUnBYE
Wn19ymgLALKJDrj4g7wkEnQi8zDaZ2fxhnj+dow/o7LEgmKZZHw+L+j+dNtlARe6
WUYNn7euEiUL6qvGemYLfZkcyr7nUHjhzUkMAZqaJ9B+6tj8sLikDsuJW+eX2QRz
wSdHbajYMDnsRXo10KCO1ShOIxbFRE8ReP7FKPkoi4R02PWOWfidsg61A8j1dPvD
xalSPKWmwd7vjMRd/PnDAXqiBQEpvdnLkvMRb721RR8QRJ7O0FJAMvpeJRxD2hrC
jTqsKFQ/TlXnBRrQl61t3cmU/yPUnSj4oqdWySBGcmf8kuZ6ONc2PaNiyq9RYeal
JiQtkqfLsR3QHIssvMcdUjDb4YMl9D+HqmNO17YxIXMYcFVxaYNg4osWHl/2Zwvy
1H/+hUctD12aKd+LdLfFKYLuw3BYRb7n4sdaZ6OlhInqKv1ODjf91CeqZTk1ZdTY
SoQaU6Qmpq4RzQ2R4auLZtEFmmaYXKub3Zj2AseilXkootVxXzRcyQVnu3f2qGeb
wFLJPHjYooEe1AgbW7yrUUxKbREWGxNk27qL0YZ2CGntMrXTx62sDFosnQhFOxoV
mWkN8ovcuQcclfuLtftnmdG9ZvRfZKPHXuNrSo+ZRMcJ/Pte1Z8UU/JeUDpZBGlK
DHNQWsWS88wETsLJVq61YRNb7fYI5G9/QxjClVDjDfbdYvDGam0F9MtrCi71QpHv
CpAWRFoLuW2RKxDnCxisq950325tlN7yu82oVw5EtQ0kfKtoPUepfQV4NGPs/oQ9
DMwIgCrvAaqlqzQMiqthgtk6GKEzqugK8AVkVyXeiN6cM23i7Ty6GFrlGUpsMWrQ
Y095Xa+ZaO1F/2vouJ7fuD+Fdfy8dJ6b9HvFWEI5jxenJvwFoj8KF2cfh+q1QnyA
SXBbJU+T7zZJfxgiM5MFhbmXYwCqBqU/hwzQAhV1NLGFXEQ0+E1Nnbp8xkqbnXFq
T+u5ZIyQzl8FS3AS64s5gBlMxvextnO2x2tDaSJCudTerIHLA2zhvi2NltAEvaMh
+HvFVNB9oYxArERgGchRCZbZ2ua4Ilbyz5s8HZ9QsUXuCE+5ZpTfGq+ToYCSNaLr
432a14euQoGQuSYw+7gbT6aJ/JhJ81wJkFwAPiJrg28G4AgbSpSRFT5t4WMMecOW
EcokygLrEpzRMYz1K1oKmCUtZShJtKCsvOakYm9xE4OE5gvWGqX3axvDym0P1PcH
okNtd89o1lzURgFSC6qNMhMNDeo5h4Ii+GKRZQSgov8IvaNr2NY0zyiAlz2OKgf5
DyOCj8J1VtOrgjcRNsWF3j1nJEjHh0ukFEBDRpeffufIMi5wYGESNQoD4V6u3luO
1cFCYzKWBgaDFLW7DU2m38F/UxsTlmoV179K4SDsdGZF3xyVOdBm10DoVJjkRnU+
AjkTrqlturgS8tSPZ6ddKd2Q2zcRpWqyNA7VYhLRnw6B33onyjh884AwAIhtud2N
xW79ETXORHHjiP5B0wsUfwsBJPxaU/V0i/0xPu1LONdyqo2rNF9YHTLfJylX0JuW
6QpL9HBvDpSbxRcD2EpUu1nQk9HFROocD8frcd3/J/7UjUncQIKzZs7/YonSABUP
5H3Wc8S+in3Cs/6LeZIKtAv4c0gd4kAJbr8JzyNuvADV2gVFSCiS/+KXZUQvHRb0
3Sux4GBt17w9qWqFCIMMDaL+aNw2lckWjfAoFQkaj/aqFzsZ93rSxdi+kpIWv8fJ
RbBa69W6BwP3CPNkeN6aGfwrXmensU+6nioy4xvOjQ5PN8kig4m5unpGl/3ybTeF
FjIc68deBkRibdieZyjhhne4uC73Y8qb8kS+p9rspsybjzOG4ZuBkNEj3hAMINhf
CSxcbX/u9WYkw3yhpFa+AqbVYJm3RFPaDgbMqnXH1QsMrXjoM5ci48VrtRpCMq6U
Q0fklUVvw12NESYHnCyvRwsTAdgt3SgR9SBdZl068yKd6fFhWmaSYjJHe7H/scrw
0AQBnZWOO1FH+Z8I00Ut2aM4+5OrsM5Dezy+28L6cjIJYPPSYRTM+EdcjW757WaC
zfEb9yOeiwdQcexJyLC3o3dgdOtKdLB3nuLdZxqEdLFoQwUvdIv0aAfRCXHuOKZc
ecouihyE8SOMVra92H9fVOPlIhhV8tINZHUBjZ7oTH4cKjrTurj6Dfb+cBczMVEQ
OGo7VFRIiHTJmirpfm1+IaH47QPT7HRIV2XgzRACJYy/Y3NPhZRyEf3p1UHxQp4+
LaYOGYmbrTlZNF1Wlw04Nsttzx8ABPyzvQJXsh7G8UcELSseSMCIsrtEs1tQqgrw
HaObYHvw/p6t6T8sFbljaYCBhGMkn54uetDWGszkSfBzCLTF/MEmPhHaMpTrmUH8
c2COJF6B8fZyEyEJbnW4BSSloWB4UC5CXGn2/Ro0xZQruljn03Q/73EqZCIeQPM6
pemzp3cc71qwX9o9UuYWhfqOAc6q55LIMOTc8X4+2J7T/8w6Z19GALbDEzfqTcD6
hzlWdo5vxtzR0yLwkiimTRIZC7boJ73LBijVHUZCS6cf6Z9OthKyC3VbeKvQeGqt
HxHMAYqrHxJdYR1bG2mdn+BJ+E8aWS0QOK5VXtBAOT55LymhlvuvcVtTWYnDo51C
eQdqxmuupZggd84G59RocjGQbHzGncDAVsEe/wUIur29KQZGU/01jPc+e8Jk3E3U
voB/Yd/rAj+f2cDyc9KlFvneNIXDpIcklehjhnXpr0lSc3s7c8Dx4rp1hM4Njthl
vr7JSr8nzK5UpFbhOpA7Y6hbN0zYfB9c23HiIR2lpudms2SPONE101NwmFyLUscE
3OiQUEweP3hHWpsuhmoJRS4wsGhuq1QTjPnuGz9cn5jIQFZFvzNHymEwo4B3b6d4
RD96bGpLRhs7k1Hvir5nEHNOu7jhVhXD8+7m976gH34sOgekx8noUYiI8PkeWrZJ
`pragma protect end_protected

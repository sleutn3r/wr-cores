// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nFVSKebILK20n0fiDhtLQTt8NNzrWUsWzky+fh7S10/a6ZQOllKBrznFf+Wkv9d+
EVe5XqS+HUjxM8hpu5rXZD8VVZCjbAhCkSNqx1Dnc1RyrSSTTvJcPw3xQAME91eO
KmoPkEd82Y+3+lNtHbyGkgVyaxxNX1Dj6zI1FmzLlgY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 34480)
pLIGMWcmBYbQsZ2K3I+LxMMyR1jb9YckTkntkwpcca4bEBsOq7+bTqgzvTeohep1
tbN7nl6gSQsAhaVXBT/WDPRbtTw8KiKhaabMbHfcbpVIedzEk6/OaQ2hzy7TpCq2
DUQp0++qC/s8XemtAC2g3kA7Uwz80qpbYpQYBN3mlPY4tBTPZfacqYhjj4MkmUsY
D6RBHWcFAVfKOi4UYni9e8jvXr13sLfnXm9V9naqfHbEDFswl3z0LIhcKTvk2ueV
aNMSoOSmeIuvNIma/fSIY2Prkjc8E80ZkWnhsZapnkZar3J3jwlJBy45ez7jdtHM
ceABGGxI54bwqNAziG7ehmX8AYZ0wz203QQe2QCwr8tU/A90eA8bNaOpTDbyUeov
FMVczMrPs+7BcSURgwB+uw+1rwMTRBOtb9+DQeLyzJpFrPScysJ9LzpNW0WJHrWX
cMYP1JAK4dddO8TjkTzPuuqRIU0xmnHoCkXNCB8IUmKti59eypk4ErMAQsE9K555
oPNbN222M2jGiR/jS+YEhYK9QBsW4VejOMAazPy0VqHLy3kebUi1oL6P7i5sVhra
t5wl8sZDri9gai9fs1nyBHEBNJTBnz7XKqIipxFZIh81nttqmp5p1xHFW2psErOs
XvnJ/mcjj2cn5x6+e3yQhVQGyWJWTpTGCL3/uJDjOdSKcachqdIs5e47PVPnfpxU
Q1k0xgarDEfauuwUuYIRjEnw3dekBLbElBJOQErwOvF4dMTQEzH2moyhgrB3G8oH
v8buUIDr1l6y1wLNTPHEIedTCB5dbaosJp2o+qz8jYb6k5tEJgPRkOBAC9EPlIyg
MPyvmjtdml9DcBa23JT9kfA/6uyzLAClvrNPN8KCFgmsG8CqElaU05ftbI14QXNx
/3d/CyPazDERTa7dees/1hkRcehkQoN+UKRUzxFdqMAodrvvWPpKh2EczOpPeBcX
Tx3Q62eIOABnoJDxqs1VRQQZ8n3qbNJb8vGiYXOmCZ23hS5JPcYJiXAyqcmbXn2+
HWLYQluE3fiZH5RBdURsDzJLfC5CvVtyqnno2xUNZKM4aUpUJFuGG3Jaa8f7jU7h
giANOpV+ZGxRZDts5F3VbmuSiXJOuyWHnIXrrYIrNnsd/OtazPD661cdS+r7ZYzj
zj34d0HTd/AbcrVkQPpbMUT5B6ayoKBfXpTokcG0Ms7cQNObcRYl0ncJODfYYwNm
CwJVikn+hL0n8wW+2/793fD2uv1DWtS7q3XGJaA38zEF42ZwqEeKwXev6y+5cPeN
maseNyykYYxziWjAQPVEUlVqXH7eyi6znT6mRCJR7NV6a9YhUvDsMcGRfzBoyXvy
01cA3DCbVEmnZS1mNaRXfHLeRn0PiM/i7VWYCzUYpJyaukGDd02T24SldhumlGdK
D+eh3WRS/Qhtv7egBQ8KFsya7gj6O5JDWfa7jpRm92L7d/5la3rJQtl7b9G0JbYi
6th6CD7XZ61iSjrO75RJwPANDZRhvHPAQlXA6EL7dOfZhYoK0rF4TGEr24txc5kd
7KufkHHt25+umTtquCKZ1SxrbzktHKqTTzaFL41kgX1CfjdMwru3s+wFbwZ+Lrr3
ST1/L0u3t6SCPgW0wpK54fx6BVqQUwhxjo7SJ8i/gI7fRRZw2Cy69iFWzCpTwVK4
DU5Y+RKk1IXNhUwgQ3u225Rxyse0tJmDQFEqM6t/c7KqCk6wu28l1t5TR7RQisRF
GE6xpo0VMiu5lMVLoHwU7b+spZW9QfYr6ukxmPqDqCRX0U6DX+HiWSLEXknrsvrS
xBmWdMKEY26938NHnZgJ4MitBNhdl2R+UhGdKawyJVmJVRI1z5RqL0rT8fH9MCFC
ePf47/T7Hfg0XiqPj1jC659VeYwMt0aTtN6HJiN1M7eJTRNHpetNsh0+tU661+BZ
Y16isBJGEV0s87T1H2Ri7XTnPNIJicUJNOCDjfjhKaEJltAhlUhPJ2SV47w4Jt7B
F7xB9Yw9pY9nwEtGfek1O1KbAZyxJOn3sfa11kS6ejf6JkzT13sNV00dyaZC+OiM
OHy5VoL8Ahsee4/9itTPCd5Y3HkMrQBz1c1SL3Ik+O1+TJX8hGf8vMOnySXI9syT
x+d3ip63kujN5YzNre8Np/JlgKCMCjJpEfudbFSj9ik+hpLhXhSmdeu5CRqUlmPd
KCb6Os7nSjcW33NAFvXOCkB849VftkDzgeN5VF3VujPk9wligcn2LBhOTKEpZ+MO
Uj2b9rRsIR3DErN1+A6732Ba0xfVgq+HIKHqswULstG4BnwsmTsJr+/nm4Go7975
RE1AQdIv2tdiIydieXFYf8Yxq3sfXNZfnCdBgB26O2Cv+9siqd/N6cuXN4PrzQFS
d8+0zCshWGr3xrNL5EpcKIBJgdSRp6BkxuytJC57h7MiQuhY2H3+JRTsu3J3+VkT
LrF2drLAnezvGG7kO9TIUQkDfq8+wDTfKCAMSdfn73PRB/HJOFXQOBU1o3FAWXHR
SE93ML1BbEBQ4DwLViolAv9JCbLplzw07/0tVjf8Gbp6sRxTYrCbGcWfQxVY3TO4
NBaKXVJj7/nOYG150jZ9TgOdRqPrxmrDn5QblJpLfsq5ClTz9ubmFDJTCt+9CpxB
Dk26ahPXC9Ubw+VwJUDXKGiTE11lF+sFncqnNoM7ZVXrTbYLmDfqAGaCxAOslT3n
xBZous4GEGLB86DZSXeqmC/VCXu3f2ymr8B+A+LXou6OwlIRkweMZbXxXozWBbg6
lJOgo+TylPlfztd3Kngo5aGLO81NsSVFulkg1IQU7njTHsfFwYCrjamutsf9CX2/
ZFz8/KUlnIZ4M2SjflcPMJQ6e/vqT9hjzKzt54dqhyVmNs202/fiVvCMsiWwsnlC
WTS2bQjPCIVe8nE4fLE63gOQ3uE7GS+139wBQKP3Xu0E8jMR4EPR3QfzdC++PPXy
Vuqu9SFi5dASY9yFoPjBETK/sjedw36hhSFRDEMha3WX8SO5oJuXUYxuOt9vyBbG
NBYfSVkWZOUUj3wFRy1/UjmPjgUmE5TSoDLu8qpijQqnRNSsgkNUedD89epgAXvD
2BQ9A1UUCuNLmzgJV8NKH0vVQNa++HNM+jNqNraMCKC3uV11S4UAdcGOh/6i5MKJ
Qp77+sBDQv6Z2Y2T454BvmDYRA5KV6oOBlgF2zcnN1UFWDkywb2TPcZ3lpnex+Lc
aMxYefBSNAs6PR8w9f5iIpCtlRuU4MPrKcbvvRtsRpWf5Gg6x+z2/WUMUmA5gEDP
tPGUkzrv4wwCfd0bzZ3dpi7bM4R7Kg5rvFxPBIMIpAFcQlbjq0c2XgXKQg5y4rly
BjKDBd/O3PzkHhcxt+CZYNSOpU7UF8ie1edA89R8kVZkHEbxp0iNG1rZNxucCPu/
Joy/nw9jFZtPfMiQlDtymbT72i7abAHzfLd1h8rIoyuiRbW5o/8AR0J6y2c6C/uY
30ThHFa/GG6Sv8xWfuI5d6dWGZm5cuARjZuBn8P9tNp7MV//wyMwOamZDH+bwQ4x
FKg+/akc9SasJLffBTzHF/tGw2dESO4J4Q0j8qc7Ujq5K51rERRKZeAf+CDsm0CV
8nX5gW9jchilbLUaJy9n5HF9Zh5on75pbMGe029IRc3VvFw0RDhcP2h0YpPhXkHx
KhLn9ASYd9nOJuX5ArtMJnGgr0E5jdt618GUDiHyLoGKA7640J5CmM2L1w1pMNJr
oq0w8KdFoq/zQ9k+ZHxehdW9i+ps/wUfyDEnXWw42DzWC5vjyPEyfPBqQzjHdCJ3
90SwIhwDsq36wf2OduJ0IXTcQt4GteyoOO1iWPe0kuDa9fg2M/TAZReQS1neQAN0
cHQ52Lp+OlH2qN309rdOCgFbBZHm5kI5cavoiDyer/DDhhm3lXKekfowIQMt4Fp3
AlO7s9lnDHcLTgURk+GxMms3JJ6Swv16gUT90jYZwMzGGUEOyCHm2S6hK/DOuKK9
2G1NY5nNQNlGk4kURQClHQEPICc6o/Wbt0M/wGnBQ3lHU5xdhh3wIZqbWRNLmvbg
M8+c+u2ILLVSN4LtTiJLAvJ210p61+GbBvtZYEWIVXCANFMnaJC4ksC5ZMHmJZda
l7CoqXEQp57lteOMEkbM+T0/00Sfk0nPF0UfwfIZUukVdfD2Dlfxegr1ZPxeCjY5
zSW9XT/yUZFBzY6pP9aLfOYUzuOGQ4kpeF7hg/dsjQdUYV/EYOgn1DLMii3XG5mp
zh9AoqGmXYQAYGxtmEL/zgrbOOsj/dh53nMxz8FjluGz7AUB/qYPOsLo0t9Z/e+P
vvkl2HfHzvRSehypvjGF3kkWE5KizHlNJg454y4KKH8Z3IypV8umwrHEF6bOpyTQ
5rd8YOK5Wjqg7qiNfmVaxT1/dRSrjiB6uFzPHKbq5Epjo4OJf8iXc3jhvCKYaP1i
mpdQOTk4j6V+iJtKkC+oL7Uk21N5mH6hZtXFXofMPF8x51JlOvpgDYd+34qJfyvH
dx3dm4PlUzgvxX2eLyVn4jXCo9Mdo/q4R9ni+TUcATf9mIrU66uz5s+WRZPvNmom
THIJYR/LBz0npI4fzH0hkJqdzCgeTIQYwLw+Bxbh/xUlR/fUg1O2dKSo8wtbLGOd
sx7A7Q3KIx8MRWpdiDYGG3hyDZ1ob8WK9UBhGpwrADrbP34ZUSsEDZ58V6rVX+f0
oY3uz8INn/a38iDvpUhAA0S7xrWsAbKzA6ghxWivdOomPJ6BmcR9iN9HVikurU3B
AbHC1o5DuBK9X1//Zl0fcjZEKZSMNGbSOvyCzkTNurtW+1zqEKHn5X1KEUT5IIY6
vCYEoTpYfLL0U/3DfF2zr5EXQFkV29NKiSS9DbGaG3dlrQ1IPIItlSMabTzgwM2U
/hzdCu17USyF+s+pxieLZ8TIJa9B/wH4l1xL0NIr8HY5NF+sdut4+vq25xcRendx
oEopykUrqfeVoEXicecUgsXre4h4TjpNpdZI0R7QCC04pe6bKad1EvLpQlLxoBRj
cMtUZBmobvVgPUpNES3SpuoiKZ9AVePbDvRKM/vhCGpi0Gtvn2ydHvL4c1ZHLXTV
jnR2B4iSdN+t9RWcY1bnIzq+obvIsHQ805jMrreaAAdpVm2jy5ZSKIiry2WmYZ3w
qBCbjmKeqmCzOgVoEXkCHvxW0e0cAbmMGpW4XJuWlVJLAlewEEQYVG5GV3IyHwYy
OiHk3Q1nZ01ULg0yUFkbtP+9JuC/4r6Ps+yZhZxy/VHlgO1fBHVuBR8JnC/rm0e4
93UQDGaFKg5PHC4uQ6RolIBOzmPisDVi/oL8jUB6gMsh/tgWXGn1O8pcyJXK3itr
LgiqbNik1j1blbgKw2hRFfydebdYaxf0B/pKPerGTjNoQNCSqXIMYusXwolFpJ8k
t1Pg4OuyR88bP/PmRFfLapg090iPuoSzlB1GcSz/DSRIqqOKNKBU/NSRNPrGQqUl
iB4EaquW3hT06Gspo/CNisSfc4yBkvUmcy/gnKH4zTkzgzhtp4md0JKAYmPhxplo
TZJmUcovzqonSuxYGzTLg4wLgp2DKmZFJoiaCmhMC/SitUmpat11sTVoyLJjOJvq
9TlJdiIaMpIayUdRFjjtIHSrGe64CKunPNsfiO1ggWDb3BQHXEbmnC1VcR6LY2N8
c5UsofVuO8dnQEMd9nLjvmg7gTvFDCvhPCiZ+PPEsfw+mutAQ/F3KlrNys5WyBME
XZeitC0U4Sq1INzsq2AFch+en62g+f3DcM/aA0tuTQrat6p89QYkYopA8scL+HIm
A1PG4RhD0PGbDQmgNGpkeuJZaGVSnTtGOKhOZO1uWRYd+UnL0MbDaU0kZ4M25Lzu
z39E67DK8uBgrn/WxWXHD4nME9CVsGZIKgJuIPZVWEwlATAEQhv7wwMabiukk61U
A3FOaav5T+HFxMe4mf18n+R++7IDAsTEBhye2DHKUdhTu0LP+eB1HMMHj1jeU4sO
1Nnyc/w9ZlQ+oBQ5uhRrdjIKuUhRQBdBMSOyURSnpCO0TK2JgAH0IRi8iubXgauB
L91Frch3y+XsemhyWC0WoiFHXAlHUzoy2TOkd8pZ9RVEtDWJ+j5lPh8BKLX4ZlEt
GOlq7e/M0g1zFgoPNP+D5wAQ+y0Jb+xA/p6E7/K2A2iFT3v1XXNkyQqsQQUUr90r
V4FAji+n+5r2Pq8pgc3OoGvsVlqzAfKA/9A5wBlzMj9lRj6ne8a6ESXTpxakoqar
kU7ajT77NtV+1phUgcfw7ch7jsIBoV4cNtTdIijqjPul+ocUP+kHlTK5ophsPUmy
oOqg4pi5psNNF26KjBlcL4fzfD/ZkOgR28KYcTtJSlymms+tC/aTapY6FtkMVWs4
h1yXB4kmf5bD5EXF7NJyNy7gRfyDUOua5TL5BDZpZP2TA72TjxbQqUccJNgtuTBV
xDLyIeryVjal2xYJXWty8Esi4CTplt/b15KraPzfES7TcHGT7f5TyQ7aPOhE2pZm
HlRE8kOQ67a4odS+o3v6wshvWpBM5lce5jt82rslL3nnJyXEXM+iFW3MpYTp+o14
Yjuw2yi2sPoRt2af5Qh2y88kpcrDkHR9/Zxb1TpUNO8+ArO+XBbQKAnNtZOBlgZN
W5K8T4upEygtQq7LfC5FfGyWhSLJxkV1NL0voexSjYMbrtOvUTDPrMcuDbQm3Ogs
JkNcTWlelpPCTIGFkkR+zjlwHkUebpbWpYPlRMngnujW+T/2Cts85hpWomhFVN67
joAX4m1Vcdgt0oEEgJiyTBrw7ePU9ye0eok4DDjASABIPO62dvStRA43KqpViwn8
1zEQRx9doQufZVnSB7Fh+RdR+SKZyGjOTlemaogSzzxlTs52l9A0TEo2TMpSahHb
4iO320pujkwPrjBgQ0Fl/3nbg5mepurBenkLVjFMmwdTZrI/xXgW0TVaz6d4TMB5
Bkt1R9OwL/5Ljg/5ru0XD02U4jFMB9B46d+cKG2sCjQXK8sYptzmMza8ui5G++e0
QiICmuODcn8n12at3698XKnHE/nNshpPgcfM7N+vFJy9Xdet9gYrJ8C1/aVB0LUS
lNVieFkIbzNwvw5whZGcao1P+eky0O4hhuphzw9dkFwlFbxt032aDUSz+gRBnxEj
E+UcwTdfChjmXucZw//bR7AacgNk8R5kq1wkoYZugTA6w2lejFw4VBpZeI6jHVir
pfQo7QCc4fdGJonEaxNCirVsEAc4+2pFy0R1np+v5SwyZRs1+IpvLQ+TrldN2VMY
p5PnJmZDD2E0Z3FXsdIUXxQ4MadXjEdeBC2Yg8Uea9KFXyFEQWkMPPSHY1oI9cw8
r6R7gnSri1eUHs+pgzaf6uQ+IjbQ/nIKLvvmV7BWloCDx3Wg9CQJ1cDquZyL/N3D
0WAs/w26xHxehkKvCRuomlHZMgoChnHnvlE8x9RZw+e9Nq5w7tBLwApxgsi0n1Tw
kpOhXV8Xy+aUHZbBfssrSHaahBIBENflODqTiAzfeIijuGsFu349hN98emmqF9T3
/hIt1Y5wPsIueMP8K1/+ntsRIJYoQrtf3XMR3vIGyNoFa6js6P3RFweuGALV8/F0
5MakNoUw9rbbmONJh1F4OGy4pWLmkO/xHLiOPA2FgsPz9AMIlcDN8ecK5to5p7+E
AuJYBR+spLDln6GJXc52Ny3O6Fuq5zW8WLfaSOB/GuhMyHbmtw/LDY2ep8FXWac6
F5vMlwfp9cp7d2KHgqUvMK4oBU07Lzq7uVl0eKqGZauPeJWsLzzwt3L/le4ume1B
vqX2vFksMH+7PUs/ghOv1rwUe1LoaudMC1gruo+XFhxcw8kObV10OGuDg7gD8ZXU
NkUe8aXdJjZSfgaiAh5+OemzwXZDWMOFPF0RCuVG2id2vglhX+fA6RFeePjSQlHA
tdkkSpFO5Nnlz033YFQDC1qPVlg/hKjWEl7Z+zYCkuxOCUeTGXiH6umLbaaD19s2
Ejrn/+qPMNb86PfIRhiBreg8pM7IKaNqqsW6eyQ3aozU1jXipSNOBtiPuHaeB8+n
6WA4zmCFDqHIxhqiE1ZSOKrQ+hN4xJZIbiUk+xn4eZWtCKXEebEmEx3I3T9DaEre
NDtV1aRVPNds9dufA2h0wVVOXBtmY1O8oOgzcvcjJFE5N1YsppA28Fmjqbzl1bhf
MAS6bJmMonXBe+PvIKw5fjhonloRGM+MVEqRC7Qp9mgnZzlEiZSKPl9O/qhlsAXg
v5BxiRzS6Od8Df+ixN7DRHRoJsMmSupR0gSGd0qtrqM4ydJNc9KflnleuBwbS/n/
tTzphvRTtOiXiKSaVvYIqaH/UCWtvUfmQjSFlXfyN7T/xaG40yJwR5DVGmcqmc+0
VRHKkVmzl3rJ+jgh3TSMAASkwzF3XJZgWJjxxpsfEAPHOWn9/gWxBESR4DNCsH4K
xrNfb6qW9U9PJVdGZeTsNu4FHZhPTMtJOflumkr+RNCik+TggeWjHND6xYaHFwjT
9OUPnwgxdtuWExBqhU1TeiExTQLXdz3P18wKChkVff71qHXZLeTs3T3Eaxzw9vNq
LWnwPayhYQ/KsJKGfgkHGZEzwSTGvY4vnD8crYZK8+CwIQBDQ4FD9g2KpBVE505N
mZQfe6J1153dM2WlQ9K3V/+5BgJgecSgYIE07Ga5IyyFgx4+vcwWfqVgfKobvJAm
FExFXrpE3p2ZPLr04f8FW9njdueaqemA9GFAg9EityXCwEvlZqwG+KABPCVk6lJa
AQpos0aIiNBTVBe4do/n/nU8mkebVR7a2Y5AGksxZL34eEaf/iHrabGlxxKyOZb8
MkqFGp1+XznwDS4YFq06w9do0GmqQq0pc/4OKx0VuvfP3neL4X1YlDTdCdF5HKx1
mjomtqHygxy6dKcRT6aVb1qk53vfLwxh4yZRWaV2wl2Cd1gHmAGUZdH5LgWLHvy8
xaYXwYPjLkKy0wvqJQdjDUTVtjsYp2UeC+/FR1ljhQ/RrH2Qrux4TewDNHfSCF09
xQ8bJE/3K11QSD/ge15is2tuIO2NloaceUrDXIhhvVLr8tHa82YXNlVd8TWl2zAc
Bc9cs3FoN4MuJTjgFWJ7mFpGUuhhgtGIeAfFDIfCcCFK1X1giTnb1BTji6udphpn
H3p6qYobPbY/04Fjco37jIIDrK04EtjK2u/vYEABMZbQ710gxM1phoLV+d+Tm0Lh
xmzJ0ueQNyCQjYEmMub9mZiwHypWRTchkkun+RA3j40avoByJza0IpaskwFymYJH
wqV5uuz20c7sYMo6kSFJupjEroQ7zQwXuKcdYZPZJe0b9C0SustmHwpWXPBXt+Sq
V7TAYZE4WFU/CugczlE27bn9SGJ/aSEd8EA2zyTZROsEpfa+mYb9fZtPduJqb5rq
jhjtPE3DrNTN32/61wsBKCpJtLnI6KxcH8Vx5to9AQxpwjaHqrJiPMtL8jGYSxBb
DB0ItcMBgtREMnOXKvaYlLnOXEp9p3rye8JdH+N3x6D4J0zh37NSEn9giEO3IJoL
okJ0+jchx0sMhfUJ92dKzuniQhh9zrhjPIb4ECiRpel/Xt+vOP1N4uI5nn7gO+hQ
8sf4ltwYcm69+eK8jI9SPyk5rJz4EqH1I69UdL4jNsOaecpRrvMukdoUkWFRKNWw
pb7f4YOUTTydC+VCAJzVdzG7nNpniQdHj1wJ/pA9kBgOGQ/QPrqhpjkDap6neZFN
9nCDndTzIWGe+TjBgUJ46/YDPYhhGRVYgts1sHbyH86YvDofwrpv5oipDN3GWLou
Tel7GULt9UiaUpOkIYI48AgWlWk+UzS5quGUz6KVFWshpid9zbYRxfbeSa0qrCzZ
oGmaQLN644GGalcsUCP/qZ0uZ1+MNJAIHYLuimqgdaJEUBSoJ8FC4Sl8KXo8O3Tu
CY+03+PXrT/wYJsxngHqiGmQ1IwiWFwP70xt5KxbqCHsx+0iLMH2Vk+oQvD3CIun
Bjfap9Ia3yWbH5JpYLl9qbRVHTcVpf2dONCDwStDoAkBMzEdlTETgDbbJlSiTbZS
CLPPLD81mPKYmI1jq0gGtN1zaxD0E4bo9fexlt2G6h/HKjIA+cB/mzcwRpw59MN4
+A0DgcAvpCAT1PW53wS0L+9PtwEAQdk5FeRjcHi9jm79baMxZ9jvJQyy/4oTMERd
3PUWBq3tTo2717+prgVJMR/l3hFlq5LM2t5N8CSKIjXk40iH2M2lAx3I3q8NCEjs
PbNm9njIhQkP0oJYQGuO+hU4H9qW7yy3fDflj+eUz46jZlABgmtPpheA2WDAKj/Q
7C1HbHiJLjywQ/m29CyyUj7nslYGgXYdKKfb489NAGZq4XXKTpC34ha0Fja7h02F
NWmGvutuyd9h2yEr3sOrmM/U7lwyxyizo9ESbtWHsc+DMt0uOevgGs0vtme1m/3y
YBaNnAvPaFQ2Y2okhECkr+ucgA3bVNC03Jr/aB5amu13ch4nw+KBL+N5HBfUmd/Y
Cgn1FIBwbJkEzQETdvpNxPOszTd2iWkAbOKDVMTn3KgtAMAFiF9sgEV/5DSDaLHq
GhdNJGVIT+qpoQF6COM/m2OeKM4yIwcC48Se/uliAaA4noa5uQXre4rMAiV8HcKI
48OEkBbY8AAdNJeBPNlk1m5BJnONL8Yr9fFl8QbfJLRhQ6+AII6S01u7k2e8ZHyd
af1G/vcX+okveww9el91fnYZpF2kqI1+E4NLvW5ZcxRLpcWAgfVLNOAxCaWnW7YV
gfylF1l80KF+3QEdn3tvIK+MnPYoj6SnRUx/H49p0UmF0mexMx3gU1IzgBEmoY8O
aN8s0ZPyhgT0h/rBnVmXYmsZ/p/ACPC/7DX7Z7OTaDj7JSk1sIhGiMZlVscgcYev
IAKbAhTbUE0LZ/stm/DogdJHe8exrL+EzB+yt22/36bJ3kI7M9ZMKqnXjNx7eZ+p
tT5EnjmMfpzVBIg0qm9nEE6kNKhrB/Hb0CdbQCV8ReLba/Vq12CH8A4m/XDPUOyv
sTlh+BHHnbMLlSoGnOYHND5yFgDBsdgikoDoeSD8qMTq7DZvT39aeVLJg8aHKUig
ct5IMtsAn+B5wXVVHB7aYQ3PLIWV1p/ZD9Wy4Ksp320qByw1is7SfXP1Gx2pI7OR
uq/Qi+q+NdP4YUXR07a/NaX0CN7MvhjwrbCxHI29G80/sL9/Rxb+Dm2NDIVfHm1o
nTqpKHpg/7bD/InvxoBIOiuhrsIfwPpRygQe8Kf79RlDIg+aH3WLQ1ceKofjKIUz
J/3ZeMIdBTz2g6JCCCwTEYlYiqLQgWtHJODrvVZPvD+cD2LFh8p3x5knu7qdYYCG
4hHfdTHEkENuPo4Vp3boCoPYZ/5yms16cH8b/lXzOEbFt+oacZcIXnhBIk9d13lF
9Trv9IExyzUu2ACRXvKmGpR2ls+G3y1Vkmf3s8wDgi9pLTF0/AOTQY/cY0H9Gdsy
AptlqGChuq4c5jb5WBPJvP7cxsxbke6hgl6XyooLkiImiA6nRKNVsa9RaxrmZD9z
39rVKeGA3WWcUJQiPV9ccwcJxqh9WM7ujBrwhgp6CucgEZ63JXZWOn/nROC/QZBh
2CALpVnD1NFD4RxavYjq78OwNfKoOJaXMC3CAeHFvFOp/y2pklHMXmA/vryst/Kd
FHJlxuzkAtrLJ7IG645S35CEiyYsafjES9/iGnHcp4u+OJHzHCH+voadUY5lLvRk
PdXVHECwj3CI/Jn9wSd095CU/3Bn1ZgjCkzDH/GNOgP2k7HztOKQ0bbKTw8+v7/R
s4mKAosh4yVVMQetd8Foc00gzbZewQ643JLrmBOnN0MACYn6TtuJrQYojxfr7yPv
kBiC502Xn+7Tc2ixLz0WwMo6QTYnbqBYGNhM5fXgg12Ze09Eurirc9efPbJqlUAc
pLLJxQj+IhR5OyEDFeVGQHIERrB9cDv8n5ek3vk96/66+Z1puj0nwd3ptaRLRYXn
mwhRjpphO8qFO4m7zfDtJVo6NFMxmCBi/WoM+x5lBs0qnHXwkp/nnpgXJkh2bgJX
kgi0Sdn/PKCAohBXidlQh4EIxAkGHDwVzxffqk0HsbM4zc6ehiUWMKvepZzGOY0z
kfa7zmL3yYmZNdjvS28hQ2ifYh5pu3xGdDW2Pr+46Kf1TXw4EVFcAj0JvX6sRu+l
7Lv7gaSlBKZgOWWogU1HuEoXjJxeuJIrE7scvqH0jb+8lhyW0XFLa4pgs2PhBCPy
11jXF8SJQd+j+A3+2tP20+KKL22ftV1Ji+wYK+09Di+7Qu/6u26jDRZizPzHCWG5
HGDEGoq20FUME2p1Sd1203gRTTTepj8wAYmHhJ9q+QcWMEw2rQNLt9xvAiby5iAk
bXct9UB3vC3Pzz0qlG0RjNpOngrPc6gru32QlpPE0M+oecAyb+8AFWSDm1Hw3qzW
tiuIz56t1gSr2Y2tQZef9zOoPD9y2Z2AK5o1Xm5Oc4uFSD9TgfC6DXQoo8R6rhSu
Cmz4BxqvrnGZotGebpMwgCsog3D6Q+0p/EfSEzRCYiKrhS6Ty/9KS/ZXJhy5JpEI
N7u+9kbDnOpYbPw9pTNMyi58+3grh3qERAfjp/R6zrtNDLF4QQ29343uxEoAPATp
KZJ6v7JovzTv83cmbkAhVNT39R9x4g09s41lYhSPyV++LE6y45TsrLcMUXrW5vrx
h+hOYBrk/sLg/QMr1p7HSW6VYAQ3VbRivJlC1Ujuk1jaBSu5M0KsTU6RWs+vMsS9
lZVrTZm2F9Pt8L4km2BCLx4f4PZyNF+t56264dz9Sx4baei3ZCqFLlkEusDQ4+dr
9vamq8YJ9rs61Z/tgU4nl/r6jqwKNo5hOCDLdeE4/WAGcgjBXeSWB7N+W5h0OmFQ
ZbDnGCmCxOyUbnnsrpqonYKS/71f4FOVKswlLPk/dIzPQCCTm0t79CDXsAGjfgsm
Xovu8ElrbDJhxyawgUvC9ge2Th/ZoexQMbASCm/MXpI+hktntt/Zg8yIX002JQvX
OITFh9ALLzEEUa0WLAFJQfG/YgvdvD7UxptJx9jCALsCWhUZhAHBmCNoNA6P82di
TcQ9mBQ7ZFuO44yMPkTy/9rFR9dQz/Ly0rB+txwuuZAVH2iQNEaU6nTFHcKr8bBn
eu3HIVN6rBAwdFLtH+IaJ97t6LiRhkPx1XUWSj8J1bJxD63W/e7WgXd4sWH/Le04
ePml/bcjNj6zLKzmwWmxmW5LYVM5dBUcypVaTiaGbutKaWZqGGfKNwz7yxzzMhaG
Hp787PiXM0OJ/oW3DkSJduRvTmJI8+I0BafZTlxn3nJtMVJp6WdoBzZMf1OQqBPp
g+kOyx7lM/hTPeKIBcWu2u7cdkc4MPhqyDFK3smc8mw6atKTjYC3S2oZGDlGh8Z5
7u+cpZAXhye1tJSVOxpS4NvWnIr+twjFLIHy3im/tg20u/WGduR+wQbtGdpLSYbY
1G56ORuILguaXTudEOC1vcA7xtIvbi3BGv6FX2A9wJbfW6SHdcqs+ieZRyV9+khV
GpGgemAae6r+MOZoWVIhn40K9ZpqZWYElmzK6Etid0XM0hGfzDQEV7NH8Ztf4gCV
7+Mm5xyK5DWJwZv1dy+MHP3x67GyySM6wwNQZvHHQKUSzduSH5dV8kB8UpAWjm/x
4Ql8/yc3z1A4iOn8nTPW8Zi+KO51Bns6OSvfD2EcOVZBJgfNnYO1Mt2glYV6/o1n
b1zmTj0kCFJSeFSfdoRpCmFjs/YsFETw1G3PxElaLoL5uBP68SteXYnYMdrnsoJv
xpPSYOhzAc+BMeOi53/r40iBu/OyyZVgVSaliU0Ky3qSSrmUIeaUSojRBnZBJK+F
HxSl+lwSqODTfCpI5RPDFIvRtBHStzyKiWwMWH8eVu5Agia2OPV17DM/9+C8NtGC
56+w4ZQU9MJFmaKFyTqzVmGU4qMxJVemVLkw2Ph6VnRqtDskxL5d57VNAgBSgCts
j0hPmuXGJWrVD/qbxua+f++bq8Q9kXJ6pROFkybqGFMdfjrUYesYoRIFNiKUhb/G
1Ru1AjAs8TWUspF5S2s+Cr2pbLz5fCmVTjzMwTIRyhSInZoJ1+TYLfe5G7jOnDDH
+U0nOeZk6SdF3V2EdNHRZbzqmv/TP3zsbht7JsfadKErkYqbmmi1d/uucWpK+hqP
Y8yZEWKfiHqJvHjH7SN99xozvMOo7nZYmmt+fXtVTq+mRrBDwKnkPnFlFfP57j13
WpgHRiza7D+4o0gD1uLmerWrxNo2T1l3/HOCVs+evy+3w/A9NKhcRWzPLJKybLUz
k/1emdYvQlhQKTWR3Lgo8qdFmiXqn7u+3sCXex6Q1knWET/HfCAu2hXBWGZZAmAJ
PGHUqznAx+PtQGhdeb3VNs9ApTe7ANRd5DI+3V3rnPhOm29a5SmDUjkrTcjiSKSf
5eRBuaYvmvIdNbO7BI/+sg8/z73vqT4j4zqIpl+sfCEjL9pPQIF38uy4JjdSPuXS
Fr/mSk1K8bbovo2iw5Uquiq7UNHVh3bf1OFBurgaP/QVaJdC7/fsYpkcpimGYz5N
rh9/tYWKkk7TadOKgiJzQd3M5+++6IL9eMSmuYTJW9EK8+Wa2lGp+Xx8qawuI3n6
G35BN4rvK7zqwWqr63m2JhLjYUJV8jGKOdWmq36Rc5XEjwMWo7S35rf/by+wv4SW
iFTBkaGb4I2ZoS9dxvtAj6FZUGgUXaKhhLSHD6rtNLejT1n8GWLwSmI/Jqvbrs5t
fZ1mp1SzfGRCnQdvatiarwmmUMMLEKBowigts6ulLiwoWoXQwUMKyiQ3XkLDHfS6
eTtJMUhE5rKHVej5HXNPMXHUOlLdAU9FWpEA+FaGtr8Xc4idDUePx3puT/96cMBi
Dzth4jb9gIMbVlyfzCMk+D9XKLTsGso0dW70dikSu6FWYVM85sm3TAHl0YP5lSwK
JolLCbafr0TBXmwr4JIXU0RG4LzTbVnxqQBM4H9Qjnyr41iFCxxUPVtFWGGEq9TZ
omtsu3LQnGhU8Vnzp5iOs97Vwykq/cMBaUOdPyeHqHk8bd92RysxOQwVuxd75VEz
Ze4W4sV3ZQWIQesRuENgfslVKrKqTF8MY523ch/nvczswJDw3sR5mIh88iaA8QKR
+h5NI2M4DQG2rT58WZh8tQVacgVelaknaYGYxu5y9iILSKUaEbKXT5+QDabzoZtv
MafkdtTs0uqiSMeYeveWscsbbZfzJ/cH9Ype/lAxwL2KjMtlFVuafTaUT5gi0m2E
/FoLN+gidQir6T+BtR4PJvW0FuhJ3R9c9AwJZBRkJP2LiYQVgTs6kMTP7RyUCMK6
aIS5EDo+hICmpA6lCd1FqT02841mmf5aeS1vtmF1rzgg4CZYRocE1RDFDsbSowkx
8my9LUM1Ugnw2wIzXspRSrT1pABUnxvNnJV9Mgrc65CSle3CU6AA0J2+xQhtiJti
mjiNNhCJNQp+y0mhDnNxRMaTj7Zdc84qWEiaTaLJPx7uiJj7j6IX10E3Hpkw3Bt6
0/jeC0h8OZwSqW2oFnLxvD+N3bJBPyvXzBTOTRx1nPeopZBtceeWmO1mavog8hwU
V8Cv9pACQOoaWP0payYrRDZutjoax0aWNcURGO3ySpCFSFDJDQ2WzPmmp5Lhp7Gt
BvPyWwWShe8s6XnI1Xz58Au4CfizTDoe1rVVip9oJW12EYSbPUaYcd6POwutCikP
9+J7cT/nTpkvnLgyJ3vV4uL/Q5kaH8Ozd2MwJvx0yuSRhCopdxnGvoMbOk7rLJ2S
IFuC7nnstjz6ZWNbwQiWTaBOTwbqWhzA5E9tOcGWOzChOwfuuiTIoUoo+AVzZA9A
RgzjxGdHP5Cochn90L7FC0gt2XiXVxfHmkPZFFtumoUxc5khlwr5SepC9q8UZq49
W4tIZAN7Xya3e7PYXB9BPWUpjMTYMhcxvoSaM7FVh9HH36jgF0lCbbm52r/7zPw+
/Uw7hoVoN+SyRxh9ofrR3TXGfRsQQftOMFXMU7Grm8uHfu+RtDsB6Tew+rZ3vOEA
3bkkdtNBjEjXKnDslk/Pl8+UWbFn6LDQuZJaQO+MG24LWdhJ7Zz8PLgP6/JMSClh
nNnYUtWkTov0XYHx3zTfT26vnTvHXxAnyKlQrHfRBgrx85jKiP7KNKwo4NbqhJLI
5LImno7BP7oQVPDpcg9O4EIlazpy3/WkOKMQqxpmTXBlngxwg5KyckkoqOSMwtvJ
7pR+JXWoghyy8jWdx2B//B2530AO6lpE0ErwOox1EFE9KL5ZAKRONiazndhxtr/d
GeAo2OwPnTCFdzBm9BHlI9mO5ds5Cptp/9p32pqVh3m3kI6jMAq2w2GbxivYFXZ/
8VwbTKjFyiux3MeQrnzv9e5fBjQgP9fQB+lr+O+rtsVL0oEAysGlAn5YM9MIm/eh
vlOJOR6egHD5xEqk250qXqAImzfamrn24FLDOoNMsajOcAzT6GEtM0I7inx0VKbs
H4xLduGBX+m3cQ4Se05hMWZKOqx50MZ9oEU4kWDAZhLIt7pchKkF4xvnw2VFUxhm
DTwzk7tiskFFUNHfyuV4jTYdswzZT/MKmadl0tLb6mjyE6B986iR5Z8iOb/zEZk4
UfamMdjNH4TSjVv8MQfJctLBgWktn0WF8gzyfDlXZxaZE0WkOuW0IZoZe3jrRg9O
fhyGG2CRXx9T7mEswZnEnO9fTj+iCoJ0Xr2rXDhmO1aVUYY6MX3ETCc2379lqras
1aql6k9SV/PMudCtCrUhSAViubDdjru2KpATp0A6zPSoNHJiSEU4/10tXrHHztDq
X32blKS6LfEB9Z1fEvzBAkz1VbkYcIvk3ySwkFiJvcTSFj7FePhPQYDg4n3v5plu
L/apQYMVIYRT3r0vdx2jNac69HCvS/zC3SOd6GrnF19M2maWLvn03U/lVr/eTWUe
iDTNFme8zMbkuw8BUB0vego96yOIJhcXLaxZweW5f7ogX7j+LOzmCV132OvZu9Z+
Wz5S1+6lvqrPID6pOT9US3TP/Ui1+5OY7Rek2rKCFpfTiQBChWjSK19lur5DkSpg
z93Wcz6crU/WlhnwQ8GPebJ/DZWKjmhoetCWmeUA5BteQmvEXb9WdYXFWl9QhseN
fCce1BAvVjGkaEIECaXF/gHY2aoh0OuRiWyvPmWBdDzAISJFrq3MhK/HhxR7c61j
HeZy5g5nxQ2xcLN5LKjBAyGm98EP96wO8CgA6pI6trs12wLlfbR8hdr6LRPZfgDo
819QDm6wO9khrSpvKojp/5T1i84/i3ZA3XFyAvBEMndOQqTwfCsp/vcO2ZMypnPC
HqXY3WAbS8iBzuIS6TMY09VvR6cXQxXkA4NYQsw17ti94ldIXo1bl6T9uD+af1IC
DE6DP5cMqzFvFLEuz7OG2pjMr1MU+InX0+kol0AP22JEc5gvHdneVqg+IGR7JQ2G
TQh+eN3i5y9oZBzS77z5zyCS92W6EBrqTkduB8bMrtWzL8uSXfT6Nwry0A0uJ1St
4Sub11UdgEcAfXt5JtrbW69oj8GOWGmXW1hU5kzJvSnvadAiUD+8NPsjw157qurG
eac1cMpwWmIC3O6lfOoeJeUv4D9XxepUVWPnd3oa0b4f/RTG39tYLK6ueBX4jODa
9+psHM0w2pXxnKrW6Bfsp4CZnNPtUZpAtk8bKqvCQmbklohCGiBPURTSv+m4Ky5P
Ag6Z8qj4HisGY6YgeL5cRWvqlSz/YHQ/JkZer+0syGhibCUo/vsNBK/dhgvpWkE3
Ho1kTa2/saRtuVljNdq/yOqhRMpE5HhERzRKvz00efwzjWpqCZ9mWEAdGLCJFBtF
4nTYdWqjcNPGuL+64c7LD4v3CbZDQ2DaM6UimTvqQqhgFM054k1FO2r0ykFSvr3b
IGGCBrp1/CarjUWq7tq0noeSwbUqWCgwuj4VsIq36SQH7wmvlF+ADXImUubjdPBy
UrCDg5yACdKTM16N6qy85w6cdapO2pqcOA2GJwppRxQJC5mqs+4sQkBcYhkXA/Oi
UVRj238h4k6Fqg67NQ/UuR0vgKfaE3KO2AQPezU+XmXrgePfFgXUyySCtOSmIUJB
x9gROi7ABt5SWCIYi2gRkFfXtUMCQL/QaSQPwqwDkOHpldpgljZHHrLqsDVDaPRr
4vTtZcKOonOXkN6vqidzhQWgYH21IUxgBaJ1/L9UH78o0OSs00Hs0epNf3Blo8eL
rdaiKUrwD9aoJUEfb4mv4KkjPV4ObH7Rq9c+PqCU1MBV2nCrmQW+C39b/UoJ4bmD
RsuNsi6OiplGkIFdLycMM2zPlXsxtGPZUtYS19tJbmPx9RM8G8wswKicG3bVs0t/
u4/QwVVVPgDPZZy2TW2KRPK81ssbGGKlnpm2uvXxWSAqMeUK0afDcpwcoT4kFiSD
ehPI/vqDfdCugY6cStoXgk4hdkfiNI1I38K6eaM7pBcaz7d6nPqlp5IGNhw3mgqX
QfQUk4tVSu05bb7h1NuuCMt+7/VnihsIvfDdwWDXelZhYGOlbhjjull5QHu4jcEQ
3jCL3fAMq/f+sllayPhbCSgBzTAeBErftbYTxIlwElHRD02xW1d4lTBMVUwGdl5i
vf1ZfVHRSL1PNQc2MC9M1D/xGHb2ton9RHllcM1RJhc4rjEqa71sA/7ZysBM5jyp
GOEO29DvEe3efTJzHjied+P3u3R3Vz7cmXrZV6xNMPc1d9bdD7+fNv2lmsCR9XS+
WklU+KfkVZzmaBa+0kvQ2+nJU3mcxBEwKoNH2HjC+W1AYOpERSt5ItisVjW0Dfom
t54/AgMeZ+hWDGUA425bzwytKyqUJ7OsbyT4dYHdIYXUvAxWYeIWI+Xb+wd1p2Q1
yGBwXkLkBdf8mUMDCYupPspnkO7Q0x9qDLvYh9JDD44P4dLr58DQlCLyfgDiTfr2
49pPbZw3AeC8cJbg07mqufLED0vESmeIZK76RcsO9XdgnuVHdSktUODg141gzF8H
N9reDAVfLNKYVfrwljRcVklQ71JeJX6RyWmKmpfWQ+gluWIIm84xqpFqjRW9BJww
bsmaExc6XDfNlg7QUa8xUfKKDOgVRNnnGJgbzuW8qDrHuLUdHkuoQA6rqnD8v3xv
nW8gDW8ULoDTkmoVYQ6z3cbBBMqh+nG2d4LabrnN37hQQrilthx0fDBR0HoV09qY
tCc5S+hC5i/BZgogr4bs6n3ghX8pamYARYhCMCYjqxTfGq57RMDJRI4TgH8+ocZ5
J/S+uQWDiRtgni/HDzAHvin6/H4t/KOCrASBn3PtwTJZgfAexeebfC0ddGtsGAB8
wdDWGtBLmFOZCLSZrouR21JoeQ+aXwzvMZacT/Q45dVVKTfaqXD+qTddHUu7yEcD
0QpbUB1VeG/D2NvxjkW3/28hWeM3BqYl5crptEOLEYyOxSz2+SDcPItonXdyuKhs
64dQXXN0l7Apu/5+Od66LiaRqK1kcaIEB2kMgf0hQD058YcEEo+sSi7Q1hE3VHBC
9UuhL5NwkqqsE7xPpn4VTmcVey8i4baPb7T7U1JAY3jCPiCVjtIUwQuEMMNvGrga
zQhRukG7AT8FZaxkPFScOHm03/WxMYPlPnUEcLGJGfLEtgfr5Cqhn2V8ngh1J1Fi
vnH85AGHFlMkgz8QY5Kmbr0ZBx8y+dTImoMJz5+15iRvCDUiiJP9R45+iUkjTOxj
CuyHCLHNkUXCih3Nvpm2+E2EtGAiNNtJpdV9Mp1K/1rKMWcaHgkTYny/8iopOpme
U1KWungPvr3xcy3bQexU1zX0h5hEhYz91mkTH3TCCvII8NHc83TeW+Pqm1nW4s6P
L/fHoLglJCrRStknk/UbMSdh2z63E1qEj3Nc/NPiX3o6qGTcqBjwRTqF+rgRbppW
vHVUGhrIr0PRqnlmUPl/DYPHEoHIC8gUj8MjF9DCwqt8ko6XP0q7jR3+o4eljux0
gyzAnf/TSTTjvrVjJTDN20hj9rWFxuKOhmPYRK2vZXTGDoTwFgV8l2m3Ctq5nwxu
rR9ulT1jGx92ewp75pqux55+tCmMN3ohcyLPOzJN7IaJjAt4CN+rbnqbzOsXO5cG
YzVHRN/4sZxnZqeEsbJxd9U9taS3tREv/D+XI0a3VGhu+piMM9Lf3bwEt/OQctFj
oUqzJgM9UHENEze4EEb33I0LmYD3xTjnQs51scRqIN23hJlUCq6xlgUh9iqCD1Uq
hOzqqhOp4nPVVmHW4R47iTs3fLmVrBZ1JDNH3w/7F7P/AOyV0g9s6lGoe9T6iOJT
ZHFNwbmkOYsScG92OV+gF2kpAhkWl+koxFJZQCb9OgN49eOkFSd+zWNF9DUKY5Cs
GASnbdwUW2XjK8ESt8P4VDBZfyvqagJu5HXRhw4JHz+uzjNHRwNKLX0z93hu2/DT
9PwzVcIusLxrOkTfSM9uirLsHO1GZpByhgWIjXh9aeGsYC9b6GDnGM7Dwve4x/AW
7n7f4xKihjC+sFV40XxkjNSrK71O3apqhjnHxmw7KjYkyqyXTyt+1HIE9U2mjjZC
A91qNa38O6sJpF6qekVh9V01nlOZHLCizlip9rK51shLd5/+59vQf54OQX6qKejd
DGvipnyXqLCclHxnatNqLL/Tx/pyNxWUBrjuscRki2nUdmfInALQfqhVUdUJXIYu
3+RE5pUDvWNeTsX9kjAD+JDfy/y9AWoPozbtOFHOsxrY7dLPlo1vloHiDZm9w9VC
eN5b6pr2aqH/35FCYBtk/jE2kqce8CM8VUqlaQTDjGM4lAtAbEef9pdZodW6EAKt
LzNY62PKYyl2LGLWFZop6jPVo32z/qC+DjefdyJkVVy/pL/OcHMsf7pzZMhyQbQc
BJ12MzPPN2xk478YRButObW+qYIPJ8o5CdnJEzP0n8TTJr0FvgIk1FsEDA50c24D
jvyNnCwRZ1WIVXJy2WitH3ZkPoDniS2vsuFibIyQV9phSAPl+3iuwysIW/blWGNa
CImtqqvFQgIlU7jcnODMz7sBu141KfkWUZK7Nr32UnGlukT+L+rJ1r5DTi7MyCuE
nazxqJFfPgLPehovQQIJ4Pz25xwA/pznCy3B2+D38McHaBTv+PgcVkzweRBbUZWK
43qTlUCAlHizflv6zMf7eMO5Ik7qVzKl+Zm8XPLVT841eoxIF9EausjrPZpSHeAt
/YZDyrygMU7/CXIiZmalgOBmbk+IbHSLDDBaL5Xew98cdMckL6UQ/LUY9SOPweCK
sQskMIFESS4bXNTBg/khsZEm6cI3NdTeVV/fZjcrjJwpmLt44ky0GQ0P7WqjP+AE
DXbjl/JDL5RgaA12kVwvyddEtxkbf0BDuJDeU8b26GlPKGh4rzUkafTPIjBJllza
aoCUso0BXkyVagwmr829ZE62iaq0XkvIyH9IUm3PFu/Xw9nksT8o/wQmb862qjHy
mDunwvwNDXn28gFbGoVBfoAv6FS3aipGLg8WnFwIfrzhgxO1JXIW81ZFqD+NzPEm
cSu+65WibK41DyWFT+ltPvZAwpL/6J9t49Ir5+uCJzlQXTcX+cF1zgpgcqLC2hNK
tC7YIKdNDSwCv3zgNnXD9FK+RIBsZmJs9W19BpwS8J55HsnAgNrbi7upLS0+JE1o
1wDICESa2aX1dSXOBZg6kKn+nsgoUhrjNRnfq17g61GJC1EwexDhcn2znCxDIMj+
VOsC332+l58uA62oMjw0znuobK3wwsmbYoWePw49Yv1QgVlw60Q8uHQOW8o+Aqi1
TuaLWCaN8r9XWHlngrYej6EyDL3xV235QF+cQDMN1GW8ECRtqgQc40F5PFqcmyqo
ilWv5XLrdly2zA79VnRW1PjFisWlo7Kgsmzqm2QxVRff520BWZwgzQG/9+2Dcvjj
JL5qWOUuwkjokgKVjvubyhFRYvLCMNmKMuAEL3KmwcIycKwoinRRfXq+Lvkny+rY
Rjh/7zRzqZrLSBCKUfYOqd+XoAsrpsrPBuYezLfEDZ5WTMe0iejcEoEOw8QxVppJ
B8f+lXthl1StZEMtjzlsVB2nvBV/30NCjfBQwv4KYVELiO8ilpklzYo1HyGLQ6O7
wJnn80eiqxjXpGD9sx2NCpW7KmKreymS6V8dSmQeaX6WiWlZ2PhT30RngaBFSOe+
m3Kl6gR3kqJuMM/cbn1K9hRN6wwtVjUBZJuni64eio2bEI3yw8ZV051zUGrcpdP1
Vwu2yW/tsu6BZj0dafSqVYNfTgZfYX8chcMwhLeiXoqjwKkbk4j8zWoigp8TmcR0
goZHAuvQHrcNa+mrw5u+wq6CGwmTJTGc9VD3MBMQwMgvFIxk+VVfX89c+CeUFDQV
kM7BWPh8Wt4RS8NsI4D7FFtzOdgyaafiEcaniuqd4enZWLNkHHV6tMpvG37tx1XC
zh+iR8KAB17GPJ7aei/gPZCO4+i9kZvVWg1Fv7x/CsENXXDqKDzDmZrswud9gfRJ
1WJzPHkZxBYtFJy/5JeISF5CsnIoT3Ea/7niwDnUE0fCrHekKqeE3XejkJILXm0w
ZmBojvxH9essEsN7/FNriR6ZsdZxQe+NfFimU+uVXbt7B9KfddmzrCtzaO6+JG4k
7LwBNlb8kkX0eVltwoXy4PQAoRFdZ5LUCUQM6ZoyM0X6fYODsbeUz3z8wy9gZr6f
Dq7x5/Hnxxk2a/HyV4V2cqaXg/pk1crtXiYLhLSO0wEZuQawXoIT2FF9Mma2XizA
dh6TTjScS6S4whh38iU90A9zO46VBFu6v53fok3HJf0IaUpnuNG57TQzizBci+M4
4HyImGodoeZwr1HwE/rnq9EyZYJPVNqC0fS9g2ROpEv5Oo+pthvZq5AeEKPb+Nie
M5jeTIW8E1Y8zn/1OhQDkbYM6ea4rsrPkzBlo+y5c7sypQCuvmktlHEUNPNxLzfO
1OjTPkPIbbfri4AUk3U8swXClBB0wOoXjR+kIddMf0tdSwFTNUGuI44JYA+l2R8y
TpkerYQ1NVbWXf15ZwJZmYVkeKfWw3YRyDINlx9DYts5PzQg0VnybS0RTlc8/ai2
94JUc/Rl/rHjFPwtacBIJxNYxLq42n13h/arPM5VNhKHzZ9yqKu7o47H61fMyep0
DE3gVDZaB88pzS2TQTEKtkW3QvQtecTH4/3Zy5ceClGMGLQMYpQhnfLFEyvcIJVg
43JjYafmBYmKUicYxsamnOfaUblnHoee+jv9d/nSPpfum0mekrnUVGn83F1QCTLl
ysTXjZYCFxq/KgmpZnGMCLI3suDBMeimwq3tuBml6tRWuExvDuLv9tZICV78+Z4Q
azbEYERxwWVlEsAOiiLljTr2/fNyRMBn9gQ2WoKlJKP6GgJTMU152BtGfQE7TM83
7J/SmUgNXQg+ynJZLAlWYmneBV2Gy/8mRZ4ExeDqzo3qtfJ4qXDoxXvA04yBDSuz
Pbc8mwYSTTrXkffs5T4uCGF11nEVNeTSO7pNM5CfbGEq89si1wBsYwTP9TO+ZnRC
ioXohnCpaFncWq60A25Gb0ErkXTMGxd3f8axMdJXTJUZ7ZnSfQKP9TNvYvCeH1cW
lO+PsN4X1KuWgxRemHZZM7xPmHPCemMDVj+9RVVgBUvS5pUHvudtnMiPp7hw+njB
bOCjXrZX8pgwAM0Nu+91asmenyV+x0kBRuUpsmZK3bCMMInodsZavZ9j7eyGD4oF
Qiz2ewq5Uk3whzfP7feGe3ed4nOVPOw5pg9g976+vHwLFA9tRn7xBNX3eWuYcnU/
CXjFOh4RAYOlcNiKMDTS4lCQBcgiW+QQBK9OPPVH3jyV5G435pl+kmcvOT8BN9/a
AtnAxOInJVsuprNIOyWFAweSnHK6FBcBdCJ4bUIv6ZfdyWJDVDf9cB2R+1Kox5E+
zu1w27gFOlwTxeveWLdQTFjKsHsBDi65zc3TNOB23t1gYUtSeTuYj/OTp0WzDeK4
jCdpR9k+PMVggjZGU7ORpW9J2NtChByi64IP6deRQxN4IK5pLNfgFtWK8l7A+88K
pyUMGt4dy0PxWN0g9yUaILmqJLD4qUYFwOKbWtm126Ws1awU7D9TqmPsiS9tj32o
Tc2+KtYyt4o02p7nRqPOyJE0HDBcGC/kdFqktpWgWxSH7qlYbRTARGnKTUMhwOxq
wmjIaSCmB9p4gATiKW7huHRPT7t6SREFEbIHe/5P0qhydf+C5Zx9ndl8J7ZglspR
G0ykZi+jcFj1eXVClDwE8/RHOwmhgUlOkGp5GJdQ1juQkF7Sh4N2m5+4pCvXVx7k
pALFqr+pYRnTLLjxSnwUNGk3riaR3GXgptO+7y23QTicmNBg6UX9WRFEVVFjdABY
/MUJCK4TubVfTUqV0VA7a77nwDARq1d6ces7jgRvTl9WOsCWiALKGdCECe1KeQSm
mc4hmEsnzMngWYaITgcdK+Cu+vsxpJugk3slk3B1aXDs4VSqHTI9RlAvk9hnLv4g
uWj+XGNhpKmVewRMbIpz5vHfqoRtKXEyhxeJVclyGc7devUhOJzXzIRJDOsRJ9hg
yusW/iKtwozIXvYyTuzMBNnr0O5tacYqXhuuhL6CbvccNCgDjWK57vlwyFm4cRFz
kDXrh75JOf4PYLo73iaYFRKNhhuWQif7vU64nLp0OvO9emG0+mTG/w4QI1QOpEBn
1p+gSnPuwBex7DgYlTwciyYXneWfmoCyMQaaATVwLXEpsA8hIlkR/47E9mPB9/+b
hKz5FvbBYCHCL7o53jnKhTXlcDYyenJn1qZefwAfqOD6Ao57Sa5PlsBzTcbeqGff
+qVCenpTzXMQDr72Ody5Ue/FaR4ycPiEMPdboWF+7mjS4GRIVvQ+Ila4l0buvRha
DBJIUtUM4z07f5bnrkmAzvFJjLkvpT5XCefCpb450sAUsxCKlPe4926rs3AJs/Go
mFTHOJjqPw6gheGZUkG4TNhFZ9B++bPyaKT5yH7iQsxTWco4i/eX1qKW/STMVVg5
sG1T+Kpo2OEZNL8qLHEHtTprkAH90zCftK8moKGKWg2creR6emi/cG2V2VzF/Uo1
phJCfKmWRgb6J1gaU7hCCyHXjveW1gcfb8j3d0TngyC6qrP3cNbK+D9xfOglCpnw
xRcATuP3RKo7b8wugRqNQG37CTVem4bvnRF6mpcDl+8AzZS9MImOi4O+nKtR29dw
0Xx+wNdM9ca4J8xlox9zoyjnPdk/bBJKZ+vKST+7nFskxfyIIqVY3Kiww86SRSUD
tndrmLkOXkYFUO3jKVY/Wko4UXm6+cGz4qJSUW5qKwTSLGxCbR8ZobM0T46aVcrm
J4t8x5QK9sCY8iOX6j1ie/D3XwNkUxgCQS7U6Wajlhd2Zd50p+nU/tMcwzVWV6fc
6jLywTBbk7DBvwyIv2gm7Ld5Jt0Kyeex4EnTMwV5AWE1ZUFi/bFKDkzUDvIt7Sh/
+g+Wm5or9gqeCHMxwL/wWwJnSqt96mV7eEwEEc/Y7sjy9QzEP6n0zxQemxOvOpXK
Jbf4iTlIPNFtQNacs9wYWD7/lbkYjt5kFfAA2A9/6OUHf0js9Pes/2I22X2K1ZdZ
uqWGll+bXibE3UEawprbSADE7mTQBKuBHqD03NH1bZOKL/JgsdJH4c/7BjlX+EWO
E0NeQMQeDJSQhzel3X3jkbEdnVwJOejUEc74ZvmzknMbpBvqqWYxhKPCGvBNwK7d
zebrsbF/7YDbsx/1f8wI+45kdUubcw13J+esWv9egmBp1bDCFoRTgpwn0xE/1sjH
dhuT7IB9hnq6USGlgxmqMvMLXSOqvjS/PHaFEKxF/VyWGfUOIp2g75ydEhoG0Q7e
Pc1cmorzwypgtK2Cs3as0c0Dj3bk/+uxQlIJuY//7uBtxN8dyEaaMZdlhAC9tGcQ
QCHAjGSq1UEpgri+DeH1LWyBYy0cEWEv+AtJU8+P4qSowLegCSARQuP9Bw+SoLDG
/yHN5Ia3UH342PbuBB4ksIQpW9hdFXnAxDVsmKadZn8AOrPfZ43OnUj1i0sBSFNH
y4pSSIKg0EIo2Vlnf3PLDD656+3cgxJ4wosUAecu4L/K2KIt4dUkhBeT7JFQhVVA
Eh1LjFY6mv0OKqj9NNe/js1vWege/TAlckHFPImIxW8/OroMiIy/dxABvjWQRnO1
oVPkWJ9CaPGk0KuqHknOrAy9AN45m4Vi/z3WjGI09bBHaYe8Jdmi6LhU6xOH5rW5
usDI+wWOGp/I+i8nnUBIedV5Rj7rdTsaaQ2kkiMLkJTkI/eEHzUbMzAozD50l3Ib
2NZ+L46TiJkFMpTRjhCAxKhCz2+HY1K/btoKHb7KRrtmp2ExLI12a826KL7nX0A0
hHrxKyPx7yS2TnzufKJ2pehQcJtdCWwE0sxfnLHlzankTqukk5EsKvQIpXE+moy+
fVzNzKL5nSWJeEaWkYq/Uds8MuQ7xVQwyBxWzOLxYiWsNl3TlY1TAbe4Lkb+fst7
fW54VYIf/EVnvxo+r/rZQzcnL7LukMKMNOV95+1SS9WqlcdCPlP8LydJZR40NsZt
fIh3uuVzcz0WgDmCkYOjv9Ja7J6kuRWB5SSBWEmUqfrnzI8jk53e0Rt5uLYNDgcz
EBDdBa/LlG8/L++BU/oGaG13C2DpCvAGUAtFjWmXR9GTLwbpUb4XY5Z6qSdrLHwa
hH3FS2VYIWTDMbd3rIgWXexQZNlRQbTwlPNVT9HcP5GPUjeUpjym4cdvIh0KevJ5
rg4pOmuUlpObYZ5HEtyqR4PG/A9+sHigxjO3xZNYeN84EvnmG1vZ1jA4gJIWY4Iq
Iz9zCynHBDaWCD0K8DXPUNfcJs7/UhE4IDzT/fwFHjaeN5T+L+zAJ+Kvzq+FNGdX
uAkeAIlwK4KPdA6J/lPCD9iAhRZp8XU/g4Z/8m7j4nb8wYKkdrHQWGtTfcAWVKqg
UJak09QabHsy0jYBw5OSE/W8XavPf4UvHoh/bHGhtCq9Dc5dJwY+JX+b2KZWPtjx
cxP9cIcdu2sHOFtkD5DL3Nfbpv5IwmBpmLmwftf4ZSxYIRgfzky9R0Zh0f/gv2PJ
CGKmd0RQ/Ux02am2ATUgXDOL49U0b8y4PeGHuEh+nGvQh7aUpV78LJeuzJo3N4F2
eYRVS7rrIY0gpwb80wBH1xCy6IVr0wSZsqHxmWNfRCWmy+VdgYLeSPSz63D1Twre
N7Ou2zy1clEQjJ15eB9zx63PANfDx+GKXdtvOCt5JIOrn7KaeITdbhqlnJQ1sSaP
d3PBtlA8QW6ZYVj1Rg+4Fv+K65QR1A60mdkbUOgCAxhT/oRPoEdb/nM7WCs+Wd6c
qFRHUbUyrnZg8LVG+RqGEyXcK/LQuPc+eHzNIerNa6ZvBbzh+M35g24XwfmgqUEg
4xerE0238wZOXVjbF6wlAhMVAxjBF7v3SMgZGhiNITJjzPj6XdABB3d/6hy5YyZi
IyP1Tb8WXDowaET9pUE7OypDzfR86AjM8teHP0lbcMw+YYEKF9VprUzAcostnKaJ
l9psZUDM+Xlo9EZQH6itsPoLpX2VWpwTuW2jT6IKTof/J/GT6f6ceRXY0cTFYYrA
nDOKBJsNp+Klh3tyVIL23ih5UQF2xjhF2XFCa0mWa5jx9aWfvaAulUVEmVFdwKHi
YViCJlotH+3yLxHHGYlKGKaxasQ9Y0MxrT8q/ibCQZsHZirSguoHb9///5Skncd2
VcVDjNSwUP85nWF8LwErmWx8LkkK1emD8Q5n6KTpt7WRa0G5n2qesN5UgyYbD6Ou
NiOe0subxmhvDxBE9yJvYkvcwXexSt4QvGQ5NU7Mx3PG2xvcu7o7Q/kZi19LbLCo
scYau4ic7kNpXuMTeNk8GQYXQbj3Mr0BcyODKSJCj2koW22kCwhMlaLt0Gfu/DvC
2RObnNEDexbjCf1kdIiTxWA9cZZNq6wFTD/21aYAaQo4/+TAdBLKVlsJo44gCHYH
UvZXdOJw0S3W3GTNKXR4ot6E4gF4nq0wtqO1+r7fFP1IDwbpFd+JjNhDzbZYlf+s
INMpDy7+/n/m/Hz0xrmAlSJkaaHXXy/4oUyGm+rRrgyz69Dz17Xt/GHT6Qij8l2O
NuAdM0Nz9f7DNhEu3KMqgohQxmtqQoO9JnC6Z6+Jy5OtkmpOolITiT3AvcOXfbA/
U9sXuWpcH215gnrEXjy6lKO3uHOAE/pLFIbvzTwpSOVFO62XwdegJ2VfyC8htZ2I
VMuPz5Q+1O1YBUuEc+rNs0Cpaqc5zSQcNv70d9T/hoRa7AFPzz8wKOx8Uu5L6mkS
6fGt0u6PE79dC7oJpxRYM0N4njJ1H8vRmNkE1lZYCKGheIWKVt7feV2eHZ5aYui8
Uj7OsBX3UP5cHOFhmOgGYE+NdOCt76jvQJ4LRarsYLof4LhHTGtAOQsiaRi4FwhM
rT8K6s8EZHcaR7bWPxslbNhDu+6l0kccCSNgLM0FAOXj3Db2kMOE7DofU1dMdbLZ
/WJLjpk3rERdolXo6yAsiDpRICMjytUOqcQB1WSbAQJHgpaWgbqopnARU3OVBOdY
w+YXRlvptT1mVBN7E8vk5YOSO9yloKp+WAldQgOCgrqoTM3An9FFTO/E54pkmUYV
cqh4rY+Gtza3VbALqw4cZp7qRshSwc4jb+OHcgKpg8uU46EwmScBS9vwVOVfLkG/
tb6yyDeujVJX7apCByOQltTxwN586+DIqUjiRRpdYBxppAqIV9GCn1wfJ/CBwuix
ot0Os9xVnSGJZF6iY+1qvzNlNtO9i2Hn2i6WD2TfDkQwj1swJPODOGxohs6n20pz
watwf78f+hV1r4+EWEqfn/mMI7WM42nMs+A3PxLzB53dLGoUc8kht9t0BgF8uB05
sT83SHNnfjA79kqWdKhRvrgZlD84l8YeqGJPYWymT7zmUiO282GfavyiLq09NsCu
1/S13zrYfo5ADm2VapvFYtKr2WiURtqiTHpbUdH9B6Xy83JrnezUscj0yicRCNzq
X1D6OSWsJEgCmYEQAyGuQoYDWJhPDvITB5ZIbr8R0Z/PRH9qfJm+x4k9omx6s8gX
oBZNms1PwvoONLZXz4cVL71YGEGtskRohtMhFyUidE+yukgUDUS7IdnQ6U5La8NT
Il5b8mPh2V1TLsJve0+/vUq+T6C0XkSWjiDLnOSrfDZI1b++l3POyZB9Trv4ApYk
IFSfL4lnnnOsGQGaOgMSC8WexLn5RYoMpVIgrROfrD6fn4JGc2ewHFrdua5qClzJ
s4jWT3FB6OJKzKSxQhRPmWefcd4CexXEtrS9SEDDvdv8cRKqeGOyb9SANqNtbVad
OmRGoGSVJN5LK2tpMscsd5XnrC2EZpsqWd9CluH33OXUnkOJ9P+fdTVX0wGyNEuS
g0r1iz+hjhMkVGnjPXEfQqsQ7YS4CY10VXM8aBC7BiLCNvm+913m6oHH26zAAJDH
xb7VN6CBh9XSQw9u+3/AqVkZBFeGRXDyxriamJfLHXhDFwXiunE5uazV7EWZqNLN
Jy6xiw8puMz0Iq/xmFQsPMmlQLyCkqwdtAY3C8yij0ziXEDfFLR0Bei/aJICd/WP
4U16QHgOoKMpQseGlfH+h3sGuHQulsifofh3r+HcbmlaDTC8gUxAYQMKlJCrPWsK
2Y12vZZx5iLmCPSN3jRgC1uE+3kcI+o2XUx/S+YkGKOq1Kz8skUBiT8FUE4M5QVW
1+cKa9zwGAE8qeQKizCMoUQZSS9rIue4HLG0PgPSUT4SOZ4wtbpGVTUb86z+DCaz
TnOGpOFha7Evs0ogTg+NYBwNXOFN5guOunWFuffCPN7r0IV2KFnSACeAFmGv8FL1
kK9r2M7dYj0ItSDSgQoE82o/HpjF4auEuhIAae9pJUS/7k31dYiZiX7xN6DWnNZP
A4E3QiQwhA6BZwQJH1jomCzmYoEs/yIBClHE7TqwVUhdQ0adzh9uKiOLwtuGErEd
pnjkDcg5+1Hp2UvzV5gqYSdHIG6pk2/MMru9RM02muUng3aQavcuCtocxtjevdhF
0/eHCww5imQXzqlDwPFDU3KG1evd3ZKD89yVGnyRWyekta6jGqIxuHd1Y/7B6Vk6
jbs+lZrf3ASonaf35Mqg38CkVG4nVGfevhe0n29rViLilWE3tB8QQ699tmtCRO8R
2cVqYGNM0SMqkMqE5IoQMLzz6nP8XE5gocMZ+ejU8w7VhohGmhelqe2KdRMxVtbP
bpjIlSMSPqUQNID3h1FyrJx48uiND7HAv7z1timxvlJG7C59rkkncMiy2ypfwrWs
D84C0vs1yQppLpAkBwZcimu3304FHEqhRLeC8qD/zF7MxmftIzIhsHThLaP2iN6Q
Jfs+g0Tv4nmN4mx2jSZVnmWzv6PTpo02uG7a6J747uWTi9f8VlagAwnqo/2JDqKP
DulP42A+VF0YvqbZfFMF4f7e82SRWgzl47eK9LXsDwIs+5v4wGY52sRgA2m82v7h
ZMk+sNc0zL0waber3BpIWxxVWz4hWD8vnW/W1ihzCo3nYF5hGvTStShhCWLSpYOr
Wd15H5tCQl4ro9aMkq5upldkneJENwvMY1kEfFszsVFjDY8xSRg2yU+/mph7a8+j
W8wlLYy4HRJqaMz7KG331x7rN7MfM3xYO5EYXfABgt9WaCUexl+AE179WXVWea0K
gYG9Eo7z/xaczZOL/hLo51V742ZVAHzWOQl/KZeoEn4QtkUSBE4tLDjFMPQ9ZkYq
KKW/iean9OtOG7qsDYYrpRXXlrdIVlC/h3tjuhTnc56qqmvG5/IvCss4zfVNXbni
39Xpr+nX9Av1kFibZF/msj6ai0qtPcFwJFZK+qg6O8GZp9vIepW089uyJ2ZBRG8p
RV9+l7OFfqgfa3nRMe1/tXlZbV8bpzo6wIFEfvLycM+98fyqQJxv6ncNPuHU++DQ
NTZLmVseaiIq8z4jCR+Hh1Z3JvIGk31tfKki/MgOf+IeFXiE6BA/iI8U+lKivyyT
2ticTlB9BeAw0ogplJ08cikknvDhzkNOPVQG/FfuDBNp9bF5ZnMItyX9lQqv94Lx
rT+6GZj0vnPP1t6atqb4XRsdmLqWH8gn8y/oemKENcVhhK6GX2ZTBF/6jdk/mNHp
Lh+RihZxcRw3F/BfLO+d//Pyc6XuqeKZnpP3WFo/J8E98Wi5JjY2QU5PtGEf4w1j
Adj5rabKsxEVSl1Wet65ZhsqbVDHLb+o/6BhcuuyOgDoSWxJAAVZNojlMbqmg7iq
odxGpZ7Ak2TaDtjhPCNV3HwSyFIeLs2RUqPAu5OMWz7HoE9317+nKptdZeclh7yT
4MWktNd3z8mQ4bWy5JWN3XubK0ZbZrnUY61sXMBy6mnokwk7ITRHMG6XnRTwt+Br
aJeLe8460x0DMAUSPtMvP1exyCvWaeZj+3TbBoU1gvKqixm24u6ESJkv2FyOqcQD
xA7EwnJuNAqaLQ6xEgIawxdH3nSXOQV4Nm0AtJw1NX5xI1i15PtnE/ciYy0e+ybb
4lOzt0kzw7nJNRe8JLlvxaQjo5+AMTclpRouOZzN02LfLfX4KH5eO2z0K9Y75P8d
3iWCqeAjrj+ceXX7QtZaxjtcN7WC5J6JcSnOLw81YnCbAuJ/szGpDGnPvM4cQocz
0V2ZPm0+5oDUXFOOhMg8W4DfoKBH7Vo4QqY7UjOEFNM0UQwbc0K0FwnI0qWnMJfC
34OSCT4em9zorDIUqNkEuR0EzMtnFONTXICftLGTH5SGs85zaoCm26S+u0pHQ3t9
egdABYH1yRTWQEnPxSCNXiIBX5NbJ6ViqrPMjJi+ZubVEKm2tANB6TP6+0uMOmtE
MJqJ0DudpzjIoeLBF+k34WAyQaiY1DqTIfP0oVSX6d6vv6vyj7iQa4P+9Sjs8vQQ
pFk/twe8/NsxJSka2Eo6PWrhOnznnBOLW4jdd/5FqfgHhJGUxLCQNs9UhvZ5rKG2
anKOOho9AqiS2pA1yoAvgVXuHmJMoW1Y3s1R0CHDf3rcb/gfNvUYd3y8xHCVm0Tk
B2itCtss0d7+iGsOdhJxaLytz/Q8N7GQf1tUTyymDdmLPz9R9uU8+LPOJDL6MwMJ
rH3PuRwixDKw8SYf3L4c4roiHuMzKer/kevRKjXHAsvEKQLn0n7ZCOQ5pnGvwbge
6zOq6evmysRlEiy4cS4ZA9qhm7sM/CEXECBOL5a93BazShQP2wP72axtftyLFh3V
AvKBH0zmzHAHHbZW92eyBTcmBZKydftQe3/t7181fmTWtUEcUqIAhtQwLl4Oz6k2
GCfaNHrUNCBIt7qMTsZ7u0SNs6C2lYmJP+GqG4mYnrqzgp0PvLIXeWXbwppARKc+
2PCkoZM1BopcfWHGtUUlbieezIrjz5nZNEylXolgz2YPGaxF+xHoQ2ymZZKDRyYN
VCSgpKbESzopD/IQ8C/LW5zhf9b5pMjfCVhVawtIzTuXRu82jF0gSWdIuj3KYI7A
VZqb6d0Iv9LCF7mqnDbuqoKiCN2g1vhSfUEOOYZf+ntFj+7JmzwydhltAg93tcqE
TcJLynPA1OFuAISaiO71Dndr8eTNJ6U/M/OXNZSwEXVdKcFNSWSw7HdFiFKeRnCY
dED5XfsjXJmQIw8NO3ssRstAj3U3pcANTydRcgWski/pFs8VglTqI2I/co6o6RA/
KQQn5AJtisJMy6oBghmW1+OZfozTmaOaLl9hatpsYoswxdXytep3w3d0CPAyd08D
gzQ75FAQAYT/Mu0mV8nBH+tC8SM6tagByzG0UcOp0HCXSgv5qD3IAxhZSjmKFinW
kTQZDdDiI6sYArRYavLws+fPiOJqI6a7kefZDwt6tV1Znkb52Y6tI74dey05SWTB
R5gEPltK8ow+2g3i7nnovWmOZqkQMrEPyZ6sXLkKNbzqH8810inAwPZDmwesILCS
5zvOj3OGNwU0evPz4mactoxLJKZvxO9vcl1HZpeDwQ52UKAbp3HiuX/83XQtgEfH
cDFaUWJE4mxM8ZPjqQNYPoaG4NR9AJoCBJfLqjSwwchLFv7nfEKicDQhoWjTn7K7
FACO1vV10tbDOLxXYmctuMwQBFglZbC0BYzKPYn+7r0Vh3yREl4vlsxJIJZFyMuL
smIEi8ZiQs2Lqr7mCoggyBElImuxNUKEOGP3r3xsR1b9q0Cy69fE7GyRvr9Pj9wi
8YaagUB7mK6Xb7j+aaoKr5Q3svJrAxbSE4rXUvbdm9wBK0pjYhUUHnBgE4VvHFCY
GnvpHAtvbE8dSx2walM9/g1szdGsre1J/vlajwERCDA4o8F9+zoUIhMbPERCRMhj
j4jA7k0vNQiLyesaAJGyUUdb/eIp3w6m0CC5VlXkzLNxmPTmXO+pNDpoTvbOItPl
FjPe9KsV8OyZHEAkTfjRXMJLAGFf42jskvgg4zNthSZ4ZizqkW2cDK9J+Vw7tc+2
sygXdDYpteZc549phtEOXzwyYPF13cZkiYH+NryDNm0szVNmEniMLSxO9BtRZZp8
K7Ny1MOZ/COW1sTWEqHfqXXX5RfpG/wF9yT9Gk7j2J54sHks+rRt5itcbnCCa5e2
conKz+2/W2dQsHb0XgwDCj48ShWFzQ5oX+gXlKjV5SmTDnmp4Zt9q5GHprr2RZ/j
v6GcSlpoLozSD3RAIr/Qgp1zVkX6ykg0UBl7RLZFz/Q1aD+X6qTa3Sz4JEVnOiNE
8lqPnainasvLLUIU6h0Iszz3ei4lKqR7zi8ZlcvDWWXA0FVP7qu7a80mumrDadJr
cRVnY+MVSOzZb9WeYHgzQxj9gn0WKkuyz+ECFIbKAjWJULo9JwXEy+v7o+85dVKc
Vl2Yy7T/1QJ/3oMiA+yELIArraC/y2jexjv4nooiI3eQvm+rr8Pz6uomRuFcpZoQ
i/kcfW8aWtJoT86h2Xd+GY1FmrpuSu/1ovbPvteNtR8NSA5iIf/+ZNGTNnRBjDee
zatY9tZJm40/q7ULMa24h19tYVrXEb+JV4SGLT8q3kGHSypkuVlvIyAK8JsHmLZv
FKfvR++0DrfLI8aK9ZaP14rKUKPWTTSeAGqIxj8ZTlb3X9coLDTIJXnc0R1q6Cx4
FqS8lSgMhsRQDK7JawCUcW6Viqq7BZwRzD2m4TvOl7c09Jc2uxVKQVP4FHLRQBK5
Xc/WhusFiVV7kLdjv9PoJtSCfM8pFNpRb/mMpfL+KyrFzSu8VKYGSh33KGoxG9C7
uNQZkrRtLK+VkFzhPIGUH4XHlX1ihfD2CPO0+RgxVIY+xWGqsJqBIiXBZfTxoftX
bwxr2s8mb3spiBzgAarAFXhH+ARSKAPeegL1mz/KoMJWy2aFS3BMsQH7sSY0dgvC
EK7mBPtYcj6dsFpMXAvxX0V5NCA5lnl9ku2VWuSeVkKtFrCcVS29HN/41bEjvSnb
1waPCyZIisUFzQhGDPJQUdeXxkujW3j9f4blLVzgiKk5qS24RBE3P41GYnbJeD0F
GYJwqyK1pM+AGPSub/3HqR+Y71khLNCUKbcHy7p+YeKYLlcNfcCK1SFsmcLiteB8
Sq3Q0zluLGyNSOlbObbXCNUtxvy/QpQM4UG+ofLpGBstSW6iOyR13uKtc/JxZDgi
Vc52ovL7O5m4QjGZiPAlGDhHxSBvFmP3SGD5mX5h7wy3lEVaMVgbOBHboxdjEe6N
Ycu6ayKTz1DSCWxmkpsgi+Q9R9FPFVDD+hYTBisdowfctmfEQ7Aj0YvLfQTwMNWN
s0RZH8XyxfS7fCu/xXIQojKRQRdKGK8eZhoAMC+X7Hbvpe2g0o9a8kigcrHOXRZT
tIVgahZavCx99pwGnszFNGJf0TXL8NlndSShARoqFhM9z1+bx/djWY1Yx/b62paZ
UbH59gNuYdrAPPcdWv04yg3jEZpiRM8s0vyqNyo8XevjRtjUNz8KSRxDaTSdFR/n
brsQoakDWjsf8NQ927yrFb7oFwNQzZCYMpOwiMFhDRmkAObMjziwyrrB2lTgjE0Z
CtjJOPdM+Zu1S7QBp7XchejXRgQ6EkN6CQuciPVnBrvfT1BXe43rOH+quwCp4N+E
/6QiVABjEaYC+MZiB08M9VwDikSWQL3y9o9eQfpFZsh/S7pXIn6VKbTDhb0lr4tf
3jFHGtVpi7AmMWlOKFiOGdQ46DWT6qV9kwwtevgOnA0jwWiCNOtjHA9Fg6I15Q1M
OJwBdEWe8PC4ZKa3UQWLd6yeHIkdAzNvHtwC6m3/ktjd5TpoeL4WLS40KGGaA7VJ
mJNNb0CbusXotbYrhKu/mnYjckq1iSy57MJD+UHdR3/nYOCHen5UOlQWAD5MHuwo
i5x8TkngX5+egP5NUjon+1Fp+qftN8PVe4rsxr+IR1q1doKTR7PDVxU0zTVqI/F5
yT11nMiYLoYt6cMuy10dorsnCu3cnISU27ZG0pJB0heoaM0Of+7XrBStafSpwRug
qux/Tn96obfBA8bc9qadtFOnkrSr+DMQkMN5FPtpKM+gm8vvVgLVkE46ihqcWBUm
Vca/mw92mdBSuxrs3JxmESOumjBXePGRvtE4PH9A+2G8yjJGqTTIBj1+nKGkGovg
1Dc98chEsZt9X7lNyqYPsds6StjI81q6KT0oUJY7hMquUAGaKDWO43yHSD/Xg95O
Bki2uT8D1HNBhmDHAZY7GxONR0b6+yvjxZSmlZ7Xc+yCR20Gp2dGzRA7Di7kGqDe
UihfpKVgap7XdQVHTwz4QJGOfe7YHlHbKNCW9rivv9KNPC5YM6Oa7daLEHsVGrBX
vzF67ouFG9kCQ3uZizrrnKbla5hYz3BCrth5Me5vlUUkUj/wTHJBWGBIbMrFk3yA
JmIGzZwSTq9zqUuFUtpwyq+s71CE9D4XSqrySbkjskEzMcw+h7Hc7kx7cpHcIl/o
Wpo4rjteZaZrTeUmolNsFFfU5/14fd13R6vEqNpO/0AAFAd47F3RTc+HmtaSYYbG
vQmnz/N6TKmx8ElYC1zYjnxTtHvrqCWMcxWrfhXeBk5XKlMXnTe/nvGcmj4LXCkn
36juc/jvcB9BjzIMsPkGJlWRjKen8ITc9rpYDEhBGk6ogMnMROv8TvxN1pUwRQLH
/E9IdZ2MIL7v3JZ2NGF8hy8JvYifCyesRjvzQw5d2PuEV4lLnm+yqd1P+zeTzJuo
f8EksCLiS+t5U7CV6SgwFKM3ERznvo4qtbRQIRECJW9jtjF5jhEcDPmBnlqTptZE
fNySjt8UvcUjY2W6OZcY3fmlz3dbxhEW7BLfyeo+g1wa7LMaEz051CYQ8zaiYWJY
UCiF2V6qNLC16gvYDtIqapv3T32VaZcmGCj+FBQbDN90cW+Qn4/zmZQheQzL6/Vm
v9KxiBPd3mIs3DpTzE6IA7Bo61vbNVXRyuVHElGtwVf4XJ4kJI1bgc0jIm1FyuVJ
3t1f7gDBdIPhkYu05On3tZ/qvl0CGD4PJnqZXAJIiwanODD5W0RB9TdQ7+Ysy5kp
QNKEy+NS+SrI6dlJvpsFEu8YrjNSAhRsfIUWAi9WoRcAcf01oRoq8U/zKnfPpk0D
4mEKd7Ul1g2Drdbn0z1UG/MMfufR0jKpBWwelcjGlxA5P33hhmtvcTzky8MVSdTs
BKfUey0XCjgTh7hZH9JATgK3PukaV1z34GrpdXmnagoTQ3qAbQYxeILGS+mrYsdl
7LNcvI4tGelmTJ2mKGk9xRxGYiVVl4CE/Y9q5U1tQXL3reU6wcurQZiD/fG1Pag9
fvYc8n0zmmdkH3CS43g0ooLktnjyz1kG2sc/AJARCKX8Z2xic6BY9C2jN7vagIug
nEqYNyxn7W+RdRsteSCP8oc3rzV5NjtrEFLcXATYP7+6UDWrgIxejVadiGJr5x5s
ppUIWMMMGPwhd4IBxxisoATkoWUmMCtBVANsyKewsAMDK9x5x2to7j051ZayVcw7
W+IRgAMJEfvh1m7mtS/ZyO0B1f2WVj8hWu1b9fWcMOWXcnKfzSqBnqSza8m9aLTU
2YfKZR02yxYZAXxCWkgHtCzOJC1rsPJgTlXYQxLbv2dAXdEsOeDhitoCE5ht2/0o
mhaCXTDfOh3mn4icBxv6cKrYRW+gmS2YTC+M34LnWcseGwO6LhTv2tcycRLhnVip
gVvYnZUMITey/Bwf/ZL/1c3eiDzWknUiX6OxBNaKfi0QgJDPw60Fl2KRG3vciEIl
/IvJImxkVQqaNHNz7GdnLTaeS6V5ukJl8yTwPYWgsFuNXXNNhw8VC+F2RC7BkMze
Xts09QPGzAb9i5ckICHDl2nhG8a1pydG4B1Qa0SP2wBKqdh+eisiH5fNk/jgOkF+
/bJ0ciq6aHv98oH+CZac5tM1VGBHzW9xcEX9u+7OIf8BuJUbl+gMhPUK+48Nh7SC
hf2IslbUWWYQAvuUGGcF5IhfIdEmpWtbwH8AMWlhLSlrftcZ8T9AphdGBnRr0ySn
8+1jVbGIcEWKvYPMH6+w72+JF99XQvuOylIkfbQEhaS6y3r60AV6Uvr4MwoGsRJV
PvZLEdYqD44ES0MyoEOZJzW/hqLzmojUPWpRgeBsCIOmXl3llb2NAkZzd06I5WxX
L6QSpEgD2kpK8WQc6s+sonIRJnYEczREWHzdBznjBBMFnZydMkdsrvtAG+1XuszT
jGqCw/OYKUmuv4FXGKqHIalzAGmTQKtDYCwII516hOHaobDVM+8d2p2ecSd5mJIG
MxZKdZ/le5paHszw49Nq/PwMqCeBMNrQ08lsMbbpZpT9LSXTrpZHvfU5j1j2BI2n
CmqkFche6aLu7oWN7p0ztWXqCgoKrWr/PoEcsDwzuABpA6uBhwXHSqPYFUkt6uKr
DDl0CyHT5K9WhOAmhQJ2oSdPnhExLG5r422zbLaB0ZguOWjoSE4Gesd1MIEC7AqQ
mF9MfLieU5phrie7oTi3tsA6O1KS5OZMENVkQtfn6F0Nhm1mT+v4kTtCJxL21ti+
rpHMr/UVwvkIZpnt+aSsZBpIc/cE/Nj05Jv5cgQKgBhbGM4aPUcnzPUGa3TTUcwD
7wCmIiNU95Q20ILOX5K10ly2RIBE46ZTei243Ux//TAKm9SBxHty7MXhLv8XAFDa
Yp8P4VMD+tL7EJkA3SMhJiZvI+STDgaQGbBKLKKmlP0rnCGfV2jmAWToTtrKQ1Oi
d5HYnHCE5R9aV7RueJslTNkLzliHZ1nMhSUDBEX74F1Ra9TsBVBIt/Ko14UTsNSV
BmHd7ftxPG1wyx0xB7cKZamv1h29H40+5sPPbj1s0f3ex+5c7GDo8+wXwQdLtNh7
lhGuPpMzk99tiRWGl6Gk+qkD1vbXv0tHE5nd9bxh6xfqru44KGZQ6nlEk4Rd/scF
mXjQMc9L9KFvsx4bJG6L6l5MgHitwhthwmzJJ7rzMMz6NEPNZbZRNWdViKQzPb/y
cL1AN7Qp/JtK0oSAMqwJsf+xA8Jhv15oBqGHwGUgPy/yI+BW9AR2T5gemMObI5xw
T75D4Gpv+qxNSv20anyexRb6+lwM5oKxA2p+k5O0drOwNGJaBWRSur+MU1fvzj/L
gcGwiG5cEgkjW1vMQMNwPlMiw4XMPht+NwFMLbNC7GOESWR/YDFV4Z9siBQDBkbc
pk6m6FdL8f8hCoS5XpJnw4E3C1pBVQ5HhTOBg9d3bxMH+Q3qmv+QvkSHUGgkVhVp
n5wXlr6dh/txLyiiepVaDrxnl1+M/gpzchdSkx+D9eZmYjRi6xU3vrmkrWkprgbK
iYb16CW1dciW48j8tuG9mhbO3Oyo/MnslrOcwDvHAGJzFJxVWR3CwB3UbQ+7RCm+
OQkYJic44fK5urkgeDkCsYIeA6SQfXP0tDV0IuWdRgVddMPPN0TaTsABZkjfoY5C
HQ+JJU2zexRI8gg30aS1xPa/t3wjU2oLV/ZCeXW8eQ5cX1R9BmKEOu0bQuYUPVW3
YQXiu/NBk93QglVyaw8PDKXTBVr0YwsxbGcOf95KQMaAjhlzZBZpwNB5jr8ZlDfz
0fDWlZB8ceDI2pPmsc9u8Qe9zqLjIiegY7igYfF4s+QPw8/3HpHTjaj4tNme0Naf
cTU11oIB5dcsI/TlqJApHKOzvFvN/PLisjo14X2Th3K4C/2IYgxpuZqh26KdVPIn
bPMp6jOwXu/D3iq39qmF1rDn3Mja6R/myEJNleXBOonJGaGDNtYRCfMfV/dr9hzZ
lNJisaEl96tFIlNz88hpfzyZDe4dHPekYTq+oZlFeh8dSLlg/YrYCIC0qy5SuaZM
7XqGUqir4fB/wUezDiEC6D2u/1d+3ZIybGiM7VKP+aJUkx8c9/hmdCPjcbkpgzFp
04UlLXMK+innueGh9bUChY4iH26YikLy8JThfUWTBD898FtK+wQ8nSeZLnXJQNfo
WFdB1ZCBkO8CO7dDDhIxqxqrTD5AsehpmFDmW2tupg62c//COGA2cGgAd/I0UkY0
3JEfWgBU39a62udUatJ9WWP5+kbWmKQ8YX+KSfWUIMcjM+jvdX0uQnTqP6dkBFrw
WmF3/qkO/JX3KloaF24vzrgCYHgGzzhBS8O3AdL0Z0jOAs5Ws39sIBZFYwC3F6XW
4AxYWBI+8WBcU7twmPmQYQZ7pmXqkGp1sxveqda2UGimIzqhyZSYv/uQTYEj4LcK
WlFHb1rLTE0LXYTPlOP6DxzytdBGJ0iX2bE0fwJ0ALR5cMTHW3HmQJ66FTBm4MZm
/9JiD9rQa4tj0+bYp2Gsqdl5t1fqkY2VjJRH9qxnDxkpl6nKdw3r2pCK8OTeRvR+
LyRe5RC3+xkEU+2ltVQdIqf52wxuka6zGkgLjM5neUTR8zZ5aDc+93daDnXj/siv
LRvFFecnyH6TAe/B7xQ/hrtNlb/mleIJRwveu1I23XR+S5JWvu1y6CmO2a0WBATQ
wZ+u02vFJJ792sEeS2VLjt/NnKZR/FyeTy92YFDcGSoyOE3dQ+7WN1OJZZGm9c9S
2jkrR+czIPy8v3D0xXewxNMEoOX+Z+nN/g20ZS33Fid87Mkk4opbY4jtQCRkPi0p
dnbEjijKoh65F4FPssFD+7UABwxwRYWY9f2I7fumS88lHRnSWXxYFnf6OY37NF0t
v5vrF66rEWa1gy49WnBE14seYK4eVJcXZoid7MtPPU6M8svSEpmayyg+x71J+N4b
oDvvD4XzIe6N/yZiF2S6K5YbibqVx70xbM8+AaKDQskNF1kkUqQ0Nn160s1i+GKt
nbCpq1A9GDi3A2paE947/a1gZxtSxPysfoAwi9vFVrMsgpnlmvKfImxwIL8Sv4uv
SECaJrJBIS0GkxHKBIABxWS6VhbjUP34fwQGYDUMdiaL7NAqKS0dbMDrXIxQAAMe
o4UPDcUywGrTU1D0K2t5oxongD83jMDlof7C+31DnwWmiMgMTf2X8TLXL4VH+SmS
J1+ok4zp9idiCKlQKQaIQ/MxH09MKBaerQuiNZyVAcnjZAYzKprMBVHTYaAacPHx
2pcSY8U0G1WSihmuW+BaU035JztOS61p99/PK5MLFyAPUjEF/qerAbP13W4dLyLS
IFkFSQv+2bV7VgVj4HzTj9i5Ukg/uU9mb8fxYJvHu3DBLAE2Myriqd97PpC9XxDg
ZpyCtITdaggXPw5cbX2Kjb0cK1g2vx3ME+eHybLaJmp2+dxaT6mrwPsZUYqfiwq6
QttU5HqrmXfibX4pCnBNdy5yZRcYS2Ap3nCXdJez6ypvGngQTApgT7VGGobYKDVT
wmJ9wP2HOdFe6SI75rrUWiZ3HsWXECz43vVWRhmiL1PDC8uF8JlIdCBKFYBhOv73
rMoykSgmaPjjSnmyOFlDFuWHcwbZOmpj3ztAojV5ssf/2uCQ+h7nahoX9weeVhZr
9hKuI++2pDXT6dDFx7Xcova73affG4MVikG6PNkfHJlG/tEV2vFLkd/xLhIWt4cU
xzK/XxbP50GhoqC9oggCJgKAvVQtnAXqodElcR5qbRpf7aYC9tOlNfqtIg0UcPg6
x153k54uL7TszGI9ppr8CTM0KdZJc211SPUDwtx1vxIa8fTfxsErZ9z7iz3kJIjh
uBN1XT1x/hRKyeQ3aInf50b/I0lsDalH1omgvNRKHJ78Z8E4+1PVk4tQrelDKTKy
39dN/hUZoBrNwcMT4Q3+9lnz9pw+f/N1q3O+CbL5ojoMYmHsABrTQtiLfU//NE09
wFcMfPGVpRlqlamIS+F/h3UlXQBChAW9hDRbyPIODSrSaG/Xduxw90P5lSjkcZBH
WTF4ovXJE8oPrjHO1FoYdnHcW6a/9YsM0VJVIlkfqW+NPzZSqRsZkR7ThvP7l8XO
X6ezG+6BHF4kSwgTr7bkmf5O5j8Rri+MaVMGr4g0AT4kyVqimiieKMMtJ/KZ8uuq
B4Guu7Hf3bHE3B/h/JMkXnySUKZ5OaPOX8r16CaSwrHCb+KEXM/0cMftF9Y0fkbX
mLZpHDaH6XWiw0+1WrMcSrT5iN8iHkUgPEdeMSKZ29wNl7V976c7m8ZsNrADpFCo
FFm36BYt5mwFQ0lY+OLaj0kt+Ei4mdMghb1F8eFjx0PkPtmkdH+TFXK3VwiovAmH
Q0x3Ez8AM3QS4Ok2lCo2/6ltWjeCI0SLTmJZud2RMsWT/WszIIw9YWY+rVhC8AuS
FXC2ao2+Vqv105Kls9YZrW6aX4MG+5x+ee1hijYiqWjEyKqgogYzHAOQqfF5tdaP
Qkp/dp5/7U7NrltIEk+DTOfMVgn1iKUa+YsWfdu+4goPSstiS5/rSHPC53GyjlSk
Ew03z3ls1eoWFRyws5soGF8Tcc+27k3A0PsCLFV//FMQiCzTlg8B74rx2KVWGIlc
yqFVxRCsOd1JS/96xKjtR2myqJC9+stV2xrGBGgpLKpA1VQ+ubCWG9b7Q8VgjMZF
Sv3WRVuct18yhCiAcQwn/vlrEldmdbnNJB1seB+fSFSR8kyCkrj5ZfTcuscXA2c0
ccZZAro+gTLNBvTlfk4umwHX5G9A5pudlLMio5CxgUWkhVNqiLoJLBRMPe8YwZH6
0y4Nbw+b97RMdCW67mNQWnCR/HhnCB98EzplInyWmYvqRPECUu105HFm8pReuvlk
gnvBwGHaZXZv1hUm9vzv+5IwN8QXDiV6OxuDze10Ojb1TsfzLFykfESUXEjknwEm
9LOKGcma4uY0m49tYBkil1+FbvvjGSiSQvulCX+HbzYeWyLcJBpMeJ2lKeaoYuTm
qn93jSzGnF7FjNTXYbTaU133FOGr6mcfLp/9eQefK4HsGxcuKM4Ln17bP80J1oVP
FTb6qKDvnEHg19jQH+YV7J3FBJ3rY+StHq4gp3yrogk8fKDFLQfD5x6p6V5KSpBt
aCorkS2OQ8bH1JeYTKpk0ThBmwwZWOcWnRC8fnLvZCGkxe8UjOIUhox2jhyVRiKF
PRgpm/M8gXDdTjMMZgG6NtMxCMpOYNSPXJ0/bXP93MakBbhkrqSTly2s0g3bAbyv
60xbzn8eOEEeSnHlVAwuRkPdZHF/yP2ymDVsZC+yXlsRY9q7P00oknPChzMEqalG
KlQ+NY/q7hDl5nF17TcQgAC2+hRyPjVER87WJoc4DxIjNGg6+gmr/yCYqmle2a19
/wmx5Y6j8iRsjQJkk+ojJ2YcdknFMv4OvC71HuN+Sjkku72MVfViExmKWcgbBWda
r9+wIjS4jhVHSuYuADe0SctD4H3EK6uxVUVHu4QEP22SPH16iFtN4jHt2D2NCy84
RHi86O3BFfD/2+UmmpuJIXbx7p4DAtHRHU528AXzrrMjyFlc3rrFTmTI/iumhBdR
+EMwF7isE+WXSChqnonkkVGez9vX0XPARm2j4IC1fud6OacTXkbmtJ1P2JSRC9fA
BssYnrqg5mUDk8GtbM3m0DV40hZ6DLi/PmuwbWNnvZI9NiQyGTQq4FZLIdIUzAKQ
pp5TxxiIhES8AOJZKMtKl/RWufjQNitzRVdV11yqIduE52TDNGP+HY+PjpRdfL8M
JXvWDbEVznxf0g5nXtNSnhucV7cHYhjo918lhQz/YN9ekhTKyeEZI0hfBGdDvsBR
BWj5L2yLpfLEmKbu3rsdpFw2Y0K1A80hRuhAuxfCie1xqnpkVjgCvSKXIn0UMT9C
zaRhSLFAb+xjt6fVa8lfDECeA5e3CKApJTAOH8QuUVgG33NfcSj+n0g4E6BQ0+f4
SNyCyRzV4j8Dqy3oT9dH/+juvV9kdVo3SaAH0vkbgeTNCEIisKtFShZeCCzeozAK
ZDNpEQB9es5dwVRCFipMrXMs5S7UHEQ9CACbM28ls/Wp2e8010jYOjqBL3H/aBWe
x8v+KosOZ/Pd/illeRJIQF8WQqlmLcYXGhjVrA5KtBmnPG1+sjloyGR587EWBwR1
7M9GJWI7VGm+tgz5pRwCkvEpeBUqfxGE/omCXtp8yP/9fhG2gMlUXHEgwOn/F24H
UNXQ9s8x6DRI/qPS8x6PCaLS1l0lVeq6EmOeEKA0wJY+n9jD/9f+UnkQ0FcfZHmZ
fHnAcBnTUtOlFzO+OnEnGklU3mNsRSjdjm3yMWAtHtpyM4Xjsbm+EJ8KqG9EqpQP
JrIbDgNATHO6mLef7P5BY6LDHF225ICPlL4fEF4QnQWlk3mWXSjbgtchMRvJHhRy
IGPY5Qs1/cBo5d0Ql+zqA0wFOemyFe3063P8CEcs63AxgwUW2wtL3LFSSm5gABWV
2l4aQ20OZKT4mmrGTVDgdGW+gE80cf7ZKlX1fom4kVIZSFVPZZu59IWK5ywrmhXI
OG1uePLkY7QP7W+pf1UGUi4VuJKNldY9FMOz2qd38RN/hFRbcPb4Io/qNks7JCSq
1odrIt1sqXDtTZRLV3fqY3bWnh27l2lMwtBrAFHkzgQ6SLHIri5zofodtvcBJTux
Gegdf2hbONHiQ5LS+gFyBywIRoGGUvIeOy5P5j47DaJjXt1FgAh4BAuCwMk1ePHc
ZVn/WsrViTiH77he6IXVS75aS4q8jrWlOi8scV+EBcSDvlELuKmWR5qGRbf9xGmr
n2kj4uTSJHx2Hl8IuM+xaxZtcW/kDjUBIk301pcdO4yWSXIvAkfKrjEF5U9jBhzz
vjJPmtyMM1RBpcyyuENcCoy4wuNz3h2zBbTFUk9lhgEWhmss/5YVk1rmon4+Eywg
XrzgqJSK1KUqPFYfjaCyOfV/YZNXKHkk5yM/T4Lgv7vAlAzsicA2faxVxUXL38pl
iFeMP4LSzXekB0qea5khgBtMAl5p0FZb0cuI5lVlY985BG6y7+4QckRFHFpE+ncC
SltxvdWTjMe9NflFGltUg8Fp6HVTdta61+z18liaCeqStGk4mbMIZKfY2SF1rpMC
3BuFzGl8MbSyZJ9bEcrmW54yOHt0TSEtz1PobL08PJUdrL8Of7afRLzI+BwQbo2P
ShjJTIm2uaTgoY9JA2EKlzKKSCvAidnXsOdZtpSyDaSATgF8Bm+YS+EW8HIx6aZK
V+nJ4AazzQhusIuQQpbarJMF2OJYz5o38i0t0rk1NGXUS8gaIWZ4ySfK46U4fwii
lMrD0hJDkexfeT8Ce+ytv9LknvFOkSjf6PCjonF9nzq+JkIZh1KeIUkAz7ntam0C
jkF2EoSYy6MdNiIrhIkiQsmQgmYvAAMCN9P2aaR8o4t0FxuBXNAVUxineOOCNWWC
8VEDXSnONhpGkxn5HyDUo4UW+0i3XDSmVdoaoSQjJfc7F9UM/ncyRDRTMm49XOUQ
wl84Pq0+gwqg6br8rGsm/8JHL4V8RjZBtAAUbCVaaq8e2FopOHbCxKYfAbq4rZsW
jxAqWm1sfrW6SW+y9fGRGRkPC6Y/Lbmj3Mgk9FGw6u5TK0uInKeCaOqhBcjxix6q
I620afVBV9GeXOrJEaifGTbppKi4bSAU5/nzrfUn53HrRN8IovPZp5C9LH48adeJ
Z2BbmqjlrhfCnnO/9yFUh5ygon9eZaBB+4yfePkKcXSWY2c3BAXzOzi6wJbJaxSK
H247b7gSnCf580C2VmDeK7D7eh2/6vFkLjw786LlGiIiogUzNxiUEk/5QxbT6ef4
PSKQBu8Z5w/+qDhBvodlvDNZ8DQqB6K9SKbA2DeI31FkpJ4ofnBO0a7iguVxemle
yyq7Fmud9rwIZq+VDcLxnMOuOp2CgnRqodiHRM2WfvIV2agO0Ibm5isZjybHhTQI
5V2yLdDDnUwrES/Jf2vhIKEWTRqTxWJdzH7cF5U00kpzbkg/31BT3K3wzpTOEnTl
3dy0pVeC/d2k7X8Ba3u5O0KsIieiK35JhdiX4A1E7gdZAClrbaaWWqHcbeyhILH0
J/5kPOsw6qmtUQZVV8GSmIS4AuV4Xx1pRMmmvXVV5vOSSVSg8ZI2adct1qwdeBL3
Ux3UKm2JoqwoPKmLia7fJT7Ho+UokEwY+QDaGowGPz1hdZcqh/EXxoHR6Y2D4ytw
z6kPYfzj9pQqutUrl/AMsyA1bUsm77F0oqB4zNSkqyfvf/D8iZ1bAD6Z7N6B0OJC
gmLWfAUPLihGpsOuwPO0xeRkFBDogf5iLxw88m2qf9M9mkcWM6KNXZ+GmBVqIUae
AYlmamopbDJ0s9bpr0EYiuu4yrHMlpyloYw5zT4IcyX4q1jYiDj68jd39g4etUbN
b3zzjC9cIpRzETf+7ad8ZO5JKes/xPkMKFfRvAViN1Q6T53IeZ7y4yOb011TeMXO
thqGo0Zwa2GwaWBXMoeWsdE0XhIguVUkxzRi0ujd53b9TmoFxt3ei6iA0VMx559K
wKXX82XgreJhbEAEz1nY7q2voiNOcw3myNH6QQ4RliiMe959LuPl9rD1raq4+Vr4
0L4YgRJFUh8Yv29fuxnxkKLPn7VLzxnmlrxVNsdouS2lJCsVmR94cBBI4C9b+n2a
vysjWSiICNIdgAtCdMpGAudsbH4yYcqYtn45JvRhSakoP7Brj7ofoTy5N7xXAUTJ
d2ydynXVDJfcAWmq3OCVPolK2TSvEz1hCTAylCwRwfx2gqnNR5eGgNbyDLmZBwP9
JyigZAxCUwUMwlSgyZqcasrhrvzA646vT1PknmbpCEfvYREjikPHe3lLBztmzmPG
V4RCat7EydkA4RcJ0IEZ/0mjOVL6yFpR/+HfVwycbKMunmlZ2mOO2cDVtbRDjS7G
CwXsYmOCaGftr+rWnu2Wz+x0h7Wy9kK14rFRzcFG1MZXBXlP56hMFAn6GcWBLjo/
Ww4VJ+kCje3PZpXx4CKuxGu4oyfCQsLciYyEf4OwAkwh4goQAMI9kRm6NYaEi8GF
1wHpC4CELQJmDMvdxpuF2Q==
`pragma protect end_protected

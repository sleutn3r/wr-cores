// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P33x+fvGw5KIDG2Qiu16EMA86tVCTBhCTRYn4He8tc9t3jPh6zbAr+mN739uILwi
mkAUcg6u/i4u/gl7ZiaqUO2CqLe+ss59oDWFZuw9CV6WykI4snbBNjhue5Jsvf8u
qLPqFbXC+0E4j5Iws1rMCq0gpdiyJyIm1Vua0gly+zs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13312)
z9cZjlAclVmI5cON46fs62mX1Whl26TtJb898unhkP2Fn907o72IAP5Wx9KrpsHw
FC0C3ZQfoR4psDFLrH5hGLTC9/hZ+SkpGVCQ28hEwEpBfJ9yaRjvtpG0touL/d0S
4RJT0sOMVvovgekKpzdXl5PN96elEKhHWI9QuP/pbEUxil30AymFjghXf2EzVQh4
+He9S0Hq9CER3Mz32YT373/ayXThvRj5GCR07Kgxqh1DqT5OZJ6ottSDuvztq7IO
o/0cEnFxxyPYdBF9h9qQ7KD1SRuQedkz5Ao1osUqR959bMNSeg4JBZKUx21W8Nbg
T1mT+/GbAG58TBY+y+FDKtSxxh+IjlbxpfzRsTDRhR75+HBfIQLRt6QEWcAssM3v
zte4/i97Qf2mfS00OFMTiYbPoA+wS0u1rYjRNMhz1GnzmDotDOstRwUlXhm32amq
JB1Gfw44HweAAWNRRSCcIyOkC0i1/8Z5eIZ2ZF/gxXYmf7ahMVSM/mfb76pBY6MC
9vz4/2CmDWI9qG7K8gzipRMvtILFxOQkzIpbfUOp5IM71Rni7A4G/WmjlfVHEt7/
2iQrMNWnEdAg8P+OxV6UqesPJX4JNwStrUublPI/wMDMeytg2WpDUj+OQgm59H7n
n2wugiR8h4TSbV1DSJjC9+WPzCXpDcHT7b48Rie6Q6Duxe3JuoEz5muQUeQYae8c
npNkxfvbcaPmZODe+K/cjUr4bkNJFGlmp3714Weq8SCEg3xp7W6UucRHvZM2hnlo
wETDe4ibzanC0CP+LkJjJ9lK9ZfMMshqODyUafUWCCgfvbSWMAZi4seU79nJTeG8
tkIBT7aU2WQkFHm9tGXq6cW/fbj2SXlsMClzc9J3J3ZTKM6p2Ib9fkO1u3Sx2cZZ
mE5H0IBLWgUA3Vc4JdDyXpT24jWD41CluGy3hW6s8Yf2dgviUB/K3cOa9BR/wa0v
EYGvhC56DJgZBJe+Y8ifaNWDq0Oyud2t+aFoSvNUivmqOCe/XVWuCSrjHSBMcEj1
kVtKSA7yjQGtzSmCtZ7Fz99OGjX7OH5CF2Yz1BWyMyLboD1oWFrp/D6GibpjI+Pe
I97O0Td03kgBeWYQjiChd7GqNPhqVM207spUe+QfjT/8zSJX1gSLcJ3gdhEu+s2J
WvSIe4rYuvVNN5LRHGKECM+psCknFQje+ebcDwocAy/2zl9j+TIv6G0y3aG9usnl
j/K4m6mm4gtx8rahpQqqqcCA/zwATM9KQOPCPEDqDHfMYeAfk3hIeweFNFP0yAqU
al6YmAc5KqgSw1DYpBKFWEIASshILBPt8D/k/qQoUOrfUxfNvAAmk17nwVxu2gXX
Qjj78dJm3AIhLkTZQqnkLre88DB61kMgU3VDkaEOInGrbsFcrJw1Xy58FexZ1dmj
5OfL1T1Smjb90GLl05UpfVTvYOD0mJKfHjqR9GzmtmyCnZuV9O8Be+6Xh720T4Y/
IGxXjNECyvFQ8ijaOgf9QsVUEZ/Ja06khl6/lTNlZiFB6V5+flFsXx/jaj8Y/Hep
tkX1bRSn8y1eeG8W0w6dXEpNqtOqcz6Coj6d/ETdu+i/LgfZnSbgYtOlEnppTKvx
rK31er7slauke/XnRDvR7EedlV1yHlfTOidrM6r9rybA/t5jUivpebAEKLPnlPfp
76hR1FFCioFb0kdx3NtKagZwXjtI6V625MGNpzXLlm6u24GcaI0COfE3w6Y8ECLU
qFnbNbeHzvTgRovxfOjch3woIEZpCySbN/gi5HelCD9Ns0aEHLl1Q7L+L2zxQat0
BLHK4JIKSlsfddDCpBr9h3R8OTnj0Cb1T3bkl2tLUqEeePOBdBCG1v1ZlXfHkxv3
HL/tmbXbiZt5if1tySj/3dTLdBoZt57k9392malGN0wdjyYaxCTuz1NbF1K8VLHc
nN6nZnq4iXUSMBcL1/vxfRP2bpCmJmkYAmvlAmCFzSlmXGurouQb0/pmyW1Onzt4
OaeFSnD8OReEVDbLD02kpamCJyzKIK6O3MY/UK0MTlOJMv4nre8/DDufXf6JTA40
VcszCUuzY3jAgVxVCmKqPrcHrShLWgHm1DBMuCT69XNTmwPa3ugT+fIafuDOj6+m
rpc1PsWnnPMzOZNgzvjYRjVaL5OH22ld15gokoDFU6n4OV0ulb5lJcWj5ItLZt65
q5lh1Rlz5lvE2CO3GpGzLM2MplK0uKs1V0uHGPNGF9JUp7TgM+5xLm1OHGAYgW9G
I8TecnuC4IXjqggpgfZdgDeeJ3zoR79GTJDB69oceHlynP7Wg0goLIsKTe5WFg4G
KheNY1vDJRVzlGdREaQHSgsSNdn4AUl+HMirlHSjU4iTDKtR48AqgDuZ+Ph3ZzAw
9JR1b7BWeoZoEw2kiGBXVt0zKd8e9Oz4bHDBJYHyGlQmUS3RgdwGqKdtP9OjEdxv
jiYramBvgQyzWperS8RXQc5/MD+DsjZX+lXba8aMLmamjWIi20KlKgMP/jyNkRdw
/3W0GMI+lX3UhTXdeWmhvrN6QtGkUp4wufb155rAnu3KT2/K/u4KDGWkEwVIVGie
vwNYPbepXHhnlqQYIygcbHGx6Jo+anR0Bo6HBkXzP5iWty2MMBTqrwfqk5DLMIXg
608iY6HdhEvVos2FCqAfat0UaK4GC06FdcHigSbzIz7n7XBmyPwrj+4KFf0vyTpX
dnIHk3w3FxeTqlUpNPD0B3mgwUQS/YXF0PRh8u5IjsMUvWK0ggP6ctO1JTpC8fmo
XupTNzTOSCsfvTOeqYVhgH3tEnP5tScK0KoeKY1p9TJ2MOQAB744ecKGkbyT/5I7
2Npiei2new1tZFpOtg073DYC5RFcUgK5b7QeLJuqOj6BdfHc14c3tEYM8arvNKQZ
w/I26QPesicDW3gDHn2s7Pc1grBYbNPJMsPZbMlgijtU3HJ/USxqevspKds7pm06
aml8aLpvEborKSPacW5LMFxIZnYqbjPy1YExTtCtVYw9qnRfd7s23L3Qyrghn0Ll
gY9f8kanBBOa7eZKQX0PAAZ69BnGrAMYhX4ktInHqor6Qxv6rQcgS78YeUyF8ssz
uN2Zyx+HkDRlxEtnLAcHBHyoYZz0GJ4f+nITLD56P53sJcb7lR13wJMhU6293HGN
xFmcTkD5xGgvd5AY3vBcaak7eXA5sd19uSwLKS9KaWQhhDTtaCb6NA51tj02yz9A
6XjwbOcA7KHjvGPPi+D2BHGDWqMN3F3Lf87BLRmrhGl94vGUdfIPYeZ8yuN4nOEC
3iPkn8L2Er/LMu8W7rGy1b8CvYCfvdUGItYmXDVed8cMcoZOqKeVzZbEL2JD/m5O
l+3yJwH8dk8Ipn/1sNNF7dliAn+Ywc62jpoCi7qR6OzXPkeEQ4PgFu357w7+ZyhX
n2SyzUciEqBTmhmx1H9vIgIKfF8Ie5xvO3U/1G4HYNr02kRKNuYMHZqIhXHzXhTj
suETEb1Wjok7szaa0636XBOuwDEfR8ukIrpX+yTonHzeaWV7UAVvY4WNBPAVMIHJ
/SITQ9Fu2i3U69a9KgczwfF3i47u5ASN48qh1tz9H7bt8qZ5MKILrHyPf/a/MfKr
xm3j5lY2B8R9FePISBzFdUIoAxWpoZkJc0V3ADN2MKJ9+ZElw2bvgw7EBOHz1xI7
AGi0fw2sd/cEIymYwsI1TfZ4NYVEi4bt2hvSOuUVCHT1broFZb4tqSvmKtpI6yTE
tAsR9f9pACpZKWP6iLJtZPpuNW/TVcKzHAs3Jwt+J8EToCB/gtGWKO3bom48W8Rc
P4uWTietrVREolKEF7u7FKgWH5RvDPl1/2ln8LQ6GNgF+7kLCIBN4Ca0H4gjIkOu
LrGwArxm6RRwVoEvgrbuYEISvMK4jAm7OgstxeaNcwAceZlPXRMdLd+8nn1hTX5H
/9cKxEdPswSCHKncCFe8gEFAXJbjTiaiTy459TW/eB5fkjseUrpYFqy6ujhq0p1/
x5ZYD1Fbz2Bj2QinbMge/4Ss3biI7icDClVrFsp8QpKKE7HBSEmHw67+sVFXq18C
OZHWvBSjxVezpaHtng3H1fZTVpNDylRh0Piaeo1qfAUXvoC22LtBK+TOlzmS8kfN
wBBsSVl885gVkXQzANcC1tRm4f5LsQnW+RG8iMI/wM8fiqPKdue8m7zX8Kyj1IDG
caVIkdclP+WNgjF2cS5GvvBsvFIdkBBwBf4LcsaRRKndyabUwCEfdk+xny0Fbcmz
UGeBOsVBPac6BQ6dHpux2KioGzqsFHxxnXteGkQNeXMTNKojIuei2cnodjm/Rs+v
xvYxmicNpCwaiqwvMLNQfxETHWc23ewAsMJPu+xrsAbqA0pbxuehGFXaG74vlJNH
M2nLlZtvmBImdPKBXAk5tEBQpfbzjycD6OcHPYhYKLsUAGFUAG3lmzFa392KBoLW
DwbwM8/n1PqdgZPZuXVnQJ6wAxKX5vcIpug7RblTsuZh1SzuD2ut4nQvpdE8c/+g
GUh26mJk/fwV0DqrAe3wL9XdnC4cHX72hP2V1ybaRU8qV5RdO9ut2PcZcxoBT5gQ
49XsPh3eCIof8wMr+bWle7vIBPtYlSC233RToB3DT1laupnI30WECdWQv+exMm3C
9tydOAdL/stijVw5ZEeHpK+payQuzI72BK66xAbIZO9HCHcB1ZN9k9bJ/H1XWp2F
mk1o74I58oqrCqn7r03lNZIVnjf8oxQ5jaF07wXl3/YSXrVhsoy02xi0XbVDp0GP
Gtz8vckepH/aE+tFBmXL812SFU3fKbHcN4ui0v+3XFuaj7uc43Wi9ov+k9GitVs7
qWzgzKgpuO3+Hy375622DSqBV2bmALHwR9lrn7WXn7MsVPRJCxkjvgNsAZKGWhFU
fn/LOl1KHN96APtZ56F9MjTvPut0ZlvVlKPidjp0ERvB5VVk8L6Gp5kgpe5vP9S6
bcYJRExywv22W78xM68FynWcTHySvN6M/jYN44Iu9vZpdsfzRJv46LsvFBIgW9fw
uihRs9XxciAFQudIwyJ5SWYVUQB5xPMTbEx7FePBIbYafki3h+2mUTehY7cE0cg6
NDVYiLmMqY6TdKY3Rlf+NuY83fSZk5lJCZ5yJq3scSZ7T6QSPGeEglgQVXOBaOwX
HWm1K2GhLuCuovHh1HW9lHkdqQt+j9iw5n3YBatxbFZYuE3c2q8lTaCjTdXf7WFo
8joDr/j6YCwkanPF5qfvAIDAhKhUrYnrkTY1x595qRe7iVEboS+61tiP7CPXTuLn
KAE0FQ/vTjLRQQQXIpM53YooTN60C+TePcchnzdWrS03OSlvl77WM+1XzOAIHvdM
Pq9WIgV074jgyaWKYfWz+BMFlMJmI3d+eR7QPMaOLEbnhqczhM0WfjPOhnRL8nc9
O+19mxSCOiOqZeyRmoKXQQSTxS1ETOzrIAt6dA4dj6nIOTRmq2iUUDzBCeMZDwpA
hmvw3fgl6fxSZWsKGq/KVHBLScpzHYZxtVRGWVA7jBuQOfMm9ueXDELeWZArfOhi
DxdorFatDspBcxqcDVfTSa4Ma97Wc8M0WSNJmWkDxwdVViUGkgzTOYFkfioBaTN+
PypbOd0cbF2dbKxwGVPPW40GMBEjTVdD7q76SumOByjrMqd8WnHujV36J8QudqxO
TmdD8ragAp6ncG1xSSqUgVVkqsRB+8y7lnN+l1s4zp6zyyogv0GBp+QIUDZdxWPv
G0WlQk/MndM5GxWoLShRR9JwxpE8BTn7OgwFOteEhAc6BhLToQ0oKbFyvi6pcdI1
qadXK//i/+d0XJK/0eg1ToHiljLAy7cD6oGxOZFlO7za1jGa6Fp+fs9ZENxJ9NJF
Ev3BbLBhmNtg7RQ+GT62JHvPFdcWBLsDAA+ihoYhoDEVVqv3pT0aW4lkJ+pO7bZb
H1Xmm5es5DrlRg3z56fwE8cAiOIGyXRFJH7mm2BnR3h2ZnayejEvgmVB/EXdobt3
hd2xpvKL1HWUZnMLPRJkGGgOXY8nLRTz6MSd343uFu8Pia8sXvHq5+TbU56fNCxX
snlyJJvSsZ+gSZgVMekCdtv9LsdFHV+9M6SJ8Kws8nEV6i1lMsh8spfuJMbU3im6
l5jVTAnGx6Zwi1khBJHCNOSZOh/ozUqyQcfsiOslnbKazM3EHihmQp3/os+KEcvi
KL9IfBBipL+PJBtYDK9h1A/abRFowU8w+bXGBJxEttcUuEnHQwAECfkVEYTU6JOk
Ht4wqNWuUTnGlPAo4Ori0Z69LNSwGxLn62tQmAKJMjiCx1OgDLBRkNWsN13jBnpP
2FueM0FwmZHiCMkXR5p55vhg6lcyCvxvcnlP1bI2nqLt850TbWkSWhitCrsiutQR
IC1hNPmhwyQC35MESdrcnG1Zm+JLODRgV9u+GpQdnArjPr3cq3N18Wmiz1vvoyed
/mITwnoDvRav3XLSI2sL5o5DoBI3kuMAp7XWlj5zdWl4M13mIifRuBXO8XzW7HBg
fdwIsNsNMgHJGqBnLP/l4CDpKxbuIkxBMwsyuQ+cNCIQPI98LR1pgFos8bxuH2xv
QwIlAuLPF3+5GzertyTpLuNO6k4UI4oCzwLT4OTNxWsIDd70Ka2jj1tJ8fQbLbb0
0AA8uc/qHe0945gr8QcBxSY9AOTmxcOB7g95fqvMnTn4N7GFZoHr+Wfti6w9OXuk
WArYsds50tmnfTnE4OAJuega/JArwRIbxX9OMOCtBzp2DbbGwsFBPDh36mrDb4bv
nkfAHKRbo10VahX/H7HJcpUKZSPARwpjBflGvfshCnw0UuA/luSjH3hnKem5bwMo
PpqQqUJXMyRkR18DBwoGJJUi3JFEX7OaiyFdZB+kDeTazeyZQFcZJx6iIy/Sc8eN
+wnpESHiU7/nR6Wx74jg/eBqjfXFutsQAcju5r19hFwuW0wgKe/185Xj4OBvr69D
7NbHmhqYI7Qfi/4UG1LN/xivHSEmzMpXFNIt1EG21iP17BGcS3NcEwKWD+digwIc
0aI68YK62bQNxqFM8N2oYhn/xmXyuLwXHq1S9YlPzvj1XUwXNGyrNuU+IQIuzCv7
FOHL5jHXV4YAzY1su4EPi2Db6whYXcfD9aW4u7S0R+2fLx+k8DPXrx78zDfrOQoX
lTStedsn1UmZMA+W5LAY1+UmPUJbartFMN4IdPAFTAoTqLRZ4wKDZAisrU0GpUYC
8KP/3b9HJ88UcoXC2qtvmr6rUxd5tu+M/1m+mKNFq2bMqJAgb4bcTwJe4Nwnsdnt
bjQuOcFhq27bahTfrubplM370wYBwx5mBDwIhSApwsRux+4iE/XHwq2FIKD2TtWP
dFsoF7McglLPsRnOQRP0oZ5EK/XdnMUFDzR267ZNs0VgPgnMz+lRTvprBVZifa+N
XUktTBbr0FGlbo9bDGfSLxwCfAFwXC19MorFxNopyhC1xevhk3+xM7DnaMQEwcZn
k1xUA/ufSMSesKqUvcDLWmu6wVK+ih41qW0WmPKsRoDAjorJMP/9WUvxpV3WKgio
kOBbNqCs5lZ5HNIHa5Spoze++WY7MMHiplniOG1gqO0mfLMJNVREAZQTGIcGPYSh
6jE/ePo/mnEWc6q0zir1rKApwx3EXLQl3alKcPeZQxXwSAtd1yB1lDINtfgkcCnk
zVhglpQ6AI7Y72NGAsg4M65thIWKJFAO3Pnpuqc9nav916UgitdyeUmQmafcRBr4
ReUA+KkqFziUDnR7j+V8ilUC/6Rf3/ryg1NXB5O3a0HVHyxjlaHZDUrzxzq7ujXQ
/ex9QBv6lQOQkGxQQsfuWoSjlR8nbIjuZah4rYmoURltTeeWcw2u7to5VstGajvo
KkwChFw9Ar9iMjzqnQuMgsHPXOt5n2WCi5G3kjDEQO02RestbjgFDTM8V13jvHxZ
H2D6xvZJQ5MFrEg2NzFE5ep7M2Tn9atv6IZErrmx0maFKpFoAHGwdEauBayVV5hU
2UDfY33JrlgopGy8ghg6G5M8VWeVRA2g+ywG1m71upR81KZt+i/IZjh2/EprKexj
r5GLf0kXx/PwhvtagiMCVFS7IndZWkI6pY3oRBehXAB22mnxafCJ2LLk4vjLau9L
H2C8EjpfvHkH2Ywxl7cKxT4C8QmUCb7m8DtIE/wnNXaVSc9BKoZ/iyjHvRyDiUN0
aihHQUqDFeN2lSXO6cxVFZE16njwXvORnTcJu5nf6jWoXmL1nKOP4Q6FrIX2hKX0
99HA1+PTRiyeLNSM2Z0o7NV5u/IRILHz2HMGOIPamK18MI1+K6U8K5E1PQ0QukPH
Uo2jdbzwxtCST2BoC62saGemm0/9hmEASJoZLf4A3lWTU5nY73YT9ZXAE61hlxQL
jzElwlN19VGaQR8CEXRy7VgLh8mI5nn/1s9M9vLO4fEkssWqtkJOB2BmmiXhGw/P
oRFoHaoKj7QoZt0dRZaNbCvB/XoIWEHknwh1ukxnTtkABPmcCFkh0kn5wRCGr8zc
xq8kKLUMSjFEpTafUQ8r417Of1wmVWjqZ0FyH040xC1YKncAHiymUkyIrwC+/Ltf
zwjSxvPESUCwWQzFtjaC3OLmHS6mmYCEKwO5TVjMdyTzBdwHlZkQJTv7aPKQ6Q9f
2KeVCvxbDlBh8WqfNlyo+x40CbNkciOqsSTHUVGgL++QBzHtx9xM1ZSIpaZpJ6Ii
10WsS69SgQJfIZm7fMZwbM4qxKR3ec6oWyWx3ivRhUsoVg5wj2X1L4y4OQ/R3d4b
aXV2z8YHVg+FJoStbZkpo25wQWiSVl54ekxgskkA60NTJ70sxBluJMdUKP7lw1WW
AIoSsy3t6jE08+lOfOJm4vB9+KooDZujnhl3o73bq4+8glEJeJX6RyZqeIX3EQMP
G3wBhLnsHj2rlpSd30HQiaf8+1vzrzBpwhkdF/LSKuSUZBdVwF0o19rg6IEqII7y
uecrdZL5TyObvsjyCHjJxyFFjOC2azVcIwce403fa1Zo7oE6QxqDKkaKi2q2zeAV
b8nyBxoetSxvqPWlgy+Q4BiUYoTItaQEBrCZtVFcJW7djtPoIiRyfshb4AJbwjMT
nRr/1RZAkLWi3YarsnD6wNcF/ePfh7KIfW4/HQwQwhK065y8DZopedO9fMj9Es7G
7prYD8JC/ZpS1i6E8E4GW9itwOOIagogwRBsDG4UYVci1kmmlUavnl/DL+13EFdF
9egybZ2ZztCeeT9ume+3z3UdBJNFC+nJcpmoOtwUdJPC+lYbfO2/Nh/HOQec5SOO
HP+91Sg6aZmK4f6zcKo3/mTxsXtjIpx5bZ0T7pxkbIsI7hRjI4/zMghYNmqEIxEi
d+ThdUYy54lSNJXX3w2oX46e1fkwDyvPfYuC39FDuZ9jTOyNJPTJH6r+xb2CRplW
I0nOPUTNVTmmKIUiOE/Y6LK366DaVwQa1OhHnre9aLm6CCLQjwygU/HcbE0SozW9
vTUrCbZBG6HVDyK6wKK5Or2+5WMnrugyIPtQURNB2oAP5tJMxE1G5T4ENR22gEzG
h/m+HaOgVn+l98pPw2qwHRqHBc3/n7PZZdSQel55ZOXDvXkse8XrW12nWYz96rFn
NwvMfvuTPPQYAy12qAHXB2qYE8GdfvwM/LyfcJYYYSkYUI/yZdDvKmCr0m9/sMwv
chf7y213b+McNTU+TAoEYeD9klGn9kQNZTtI2GINd2I6we2r++5C+KUneJ0oZ354
cjkjHSvOfpy+xu0vOV17GcY+zc0HPQMO4m4bYWfTgks1NpX8Xv78g+KJ2gqlKW+A
u57/gYEYJWIx5GYnt45HopwmvbVYmSLztIe2XZbo1O644YYuJs57cLiA0bs/ceT2
4kVgdsZ62qYvBbOx+ETRzglHh12vR7WupSqaDXM22IL3HcmEipCT24KlsKJ1cZt+
08G0PYAHRZAf3yloE17XEk0Ea29hFwlrmTyBChbsWCDFWv5lEaSPxKLb3kaW+nDd
cWntnw7catBRMSYz0SYR16n1YxrmBGMxUZH0irufVO1X7aGYKB6F5/ug0M5k6B7u
QNWc2KIdC/NIEhZBCCN33nIZtZ4iF99vp1vah0HC31L4EQ/Z98Vzl4/iqoqViPV1
1UAaCSBW2oH0gyM+hJ2OFbKb7qY3Hs9GwwfQnIxFhYtnx2BVWxN230kQqandrlIi
f1feS+CDluXCmfqvPmw0i2+WWZICYxjbjYuwelqhuXNYvKjev8FE37Y2CmPV4p78
7jZUIJg2Af+L4tuyLWYvHD1agocmC3pr8rz1H2S+sX/cf2GHLjXXygp4//PCl2DY
7xWPG6ipXl7BXIa14ABPHBpP0ioKoRFZY+OCNW0O3TJegp+ykfN7ChqFdYEgmpsN
wHACN7ln1pysX/KlanoOpS4WekLpiYYqZQ1uqIDNM5K8guiypRT7YVnGgvIo8Bqr
f34QFHn+04klWWzNczhdArzszSqY3ffOnTbf26W5lYvvCXDfXNb8nc422wLQhOEd
j/hy40MWK74P6gp2U1YfEZpLMysEjuuz7IGQmCKJEm0Ep5oQwPEsGlpfsSByuTf/
++QlFkzXcFG/dc8SEcgt7CtLRxG2IBCtvPa3n/QH3DYnD2U1fHrJv/4H/nRiDYYh
dBxUzBnr2qIpKAm4mIiOkK5IA1hbUtxZ61SQmXKSsPCsLsn9bSlyeF62NxMGBhM6
XiHDOd3nKT1G6jd9LNym8rFuy600KCK6mxqRK9c+ppjVjq3swG5khWtnn4lhmEXR
/kajjfwUg/FdQ0Yq1H2BGY3WrQI59PKDyYp6jQ/De3TzMx4UEK++vdZu1W4uAbL+
u4yh0EoFq75R9aPCgwmvuHsHOoN8Zfv3OxJlVtG6u95vccmNlGDWmdLOwqY4XlRV
66QydTy8hT44oDudnMGBLnLZ6p7/PVKxgqKUxwv5MY51yS44PTRE5+/F0McygVMF
Cds6j5ZNMbjmkPqM7Yw9z657Tn5eOyRtObSOMTUkI1D0cClOd/mm0sxXo/1NMbQ7
+NRf08uCjUDbhoc2KkVXal85UUQHx/QPRFgJP8mSRpuvdhpKtCAkjOpaJTVQ+7TT
kO+bTJ41u/LrJ0zZOqOEX+n/EcDXQU03DzA1yi0zzrMUAt3RvkhwpjSiOFDpX1gz
FisOWxaAsq620jyEZCOyd08ADjN6cjsGOEvksrJubtHkEkqHGgBR9APHG+4rKpfV
wukdmPsLCkJaWpilEITuKEB93dQHV/+x9ahIH51n93wrCQkuXJXqfP95/65Pou9l
bvSG/PKza5te6qr02wwtds8DVAUB+QSdydx39/yVGn1EgYfSIlLX5n1G7/h2aNRC
JS4PSZm3+QCdv8kf5JMJAo6fe0HzcVIZJO2KOSSAwDFyXZTt/1G0QvhT2Pgef8/e
0q+OhuFjTf7YeiqGzivAeHNt4tjAec3el2SAyku3vj534u1DYxWU/fcpQ4mW7LZB
FQYhIQ/31ByXTQuyqyCbHJa3wjqf/pzeMXau9tAF4MKDG+Oky3Fe0dvkbuKTlbs0
yhDYzJpoVei9u4S/Nfzla4WFCyYNHAPfYfyn1HoY6E3J+KQcMlNjFRzpBHzDK+/N
Y4kgREbZdlsW6K4eNhBJJ9Lkuk060MzcELgvrZr8ioljvAJAIP+QyCb9i1rEVmIJ
St2eGWubZd9YDHhN1pt63ZILfb+G4of+hJ22JVtEAWIM6DuT1QZJtxCRP2bewckT
bVfSv7AlLcb1wQsB11AeWL/4c29C4BaFh4fPzA1mPs/V3dv1zNl1ruBP+4ljsOoT
afLsvObDS/DRe0fx4MM/zZH4AM8xzOtwV7f6LzsYSgfXaR3t9h3YBjj6Ec1OOvBU
VynAvc4NyPfD7fqrzcV4Hbs+uMPzDNvtK4qiIUNajIlRUHjxipN0Or/r+qhbtreK
4xpyX4I0xfnBQjeU9tN3Xq+ykLarNjAVlQTprzPqtXrYUzssU+LnhEpw7oXod1Dy
GUXXj1IqEcBwy6Oh51mbdBtQBI0svcOzpCnjpmzTyBjqsDh15zYR9+Q6cIveU/fL
BUSNV+z2HJRAyDYXaM6Xowss2/2VYhPEyhIu7BkIPXmuiaFUiqSySCaEYX61CrYc
7okQ3FsuMNJkaql8N6pCw9Fnl5sysO1qp4g1/flfkSdZtbcRrgBFY/tEt5vf8jMZ
G9QNpmFkkwWF/9T8Wd+Dkv+ObUImIxeFrwntGHGF/OtToW5yBtsZF+xGYA4O56Sw
BpB9+922xRaDNOeMKCsDCLzAQ+M4FI75zBuKwk3Y9ZggcAXgPO0Rt1asI72x2nQS
xZi+/+Qfv0ujgoBsnbuFcpdP4oXl7YTOLbLcZJnuPlt/zO+4d5PZj4nkie7aZI1y
odKVzZqPAWtp7oHKB5wrh4Z/klQCiLDamzyzqElAmxdtgbTCb30j0vCAuAapxJe7
cCTP60BWU5JMQP253HP0VflfBE7fN/VnDdKWQTweC9uyOxIwp1nmlxdjf6MutV9O
M7b7bcxPbAzdb76pmkM9pIvO28WRZPb4ZepF2roTxtHX8FvuGv+D0vD96nqIvpzs
NmmJA7malCy2XHTki5OslzFELNBLd0fbegntnyHtHMeAAUmE/ADkK6+x/i+87hpc
Tuc21eX5MRIFQ8gFJaFtvuzRLqFqA2i8dMR8DQwhZ4+1fBKITXtv6/iL+zW046Y1
VgOIPGd5pDTARPMX+szYm9PtbadOh7LqGRMhwkW2sDDUIdaot3NtEf5G0qpPZ8fn
BLEGTvd0gcfjDbxb8sOdXptITJiYykbHX3/Zos0SMV5JmI2VBjXDIBNwbU6eOg1O
0jI3NRdI1EXICiPAtffWwuIM/8oUSOGhAhtf4pRmaz62fvbQJgu3ij6V4QodQygB
j9/vnQxQ2dXDNHBDoX0DqlPidufl8KXL093KuOel3HjMX3LFYL7ADVfL4RS+Kcey
TqZecL+zmqlb3smYN/nTTgrw0w2IiN4/FN+ibzpak+vRDCYGlvX85VeoeIzBD26M
e3xud/4AH3kEATybBbKmvT7qpaagj9E9lCdX3FN2dWOUOjexmwTn7McjBQs0DEBA
mptMNrhpIXRmZvMtwCYXaLTsAyh53v2LU8PdnwaPaMlzpxx+/pTqxifnec+7fv0F
mAL/5Pg94e1NnbNBoFIciakwqU7hoxJP8PFz9I25TrnOirALh1RABtmz44npDz51
vBswrEi3XXatlM/+m4rYfijh/RaUn/FsjsLV+BMxglwpxZWvJQMgTfnpWrTkiMBB
PYi0sJlgLqpOedlWmWw7IFlSlL1CTw1fP6Vw3SzO580Cdq64fGh2CjcmVtJkwQhh
/wGfJYqUmr2dW0PVYzeJ4NSqq4BKUWvboN7Fu2e/WsNq4ddx25zgnugOCbPpxrNW
4irb7hdXuBX9JAtbt2TXUYrMCOAmrkUEQcZ5dggdn8jUhtp5XSYYtGKQMNpnjWE3
YW9kyqheQg0IZekmGC0JXPCtMXz9uUHJKeFxd2rtW1DjGpQ+M+pbtoqigYAZCb+o
jQeCwxwPd03lwFjXQaCNbo8gmaWBl02IrVGrJtnCTzPW9SfKzPxVKIcdKfVCGT+p
Jyi5BUet7FN9rWd3YMsbSsgFIkPuiqq+F/0JNC09U9RxM35S9q2wakOpqkfgbgyd
Lv8Wx0LgiGWjxaXVEuIw6Y/WqxWFgcqDSmGk5iTotwIvtcE4lVGCMNiVIpY9+yLc
n0tDP+3eZPGXd0ILo7yAusYXcWxSaHkJmtDHmGcf4DTlwDprgT+Zn0yknHN8ef9i
0toVTElwLJ2Xr2edNDunnohYiXt5Ko1WvfzHNHgu7R8xnAeAGPTNtUq/rgr0XNGb
/IfHlWArBPlPJKYslcwJrE6i95B/EVF9qdxEgnv8iPxr0VlmaYZLCRH6ZfLeXysc
5uevNDJxS9NUXuRgwtYctug+hoQASm2cdxhuwDMQOm/KCWKrjRVzCopvxVpkbQTs
XqPY5y8l3rUMxi5dFCIbs/mtRoV/CSJRTDJ5Mvxvtwg8EzXlaw+TEZLHeUKWpfId
8geiRI/TAOJRf8i/MAAwKsVbIxXp+kbRB2jfbkK8NN41AJTzVyL/pVqztNoFWEwG
7ny6IMyylA42Ac9mB+OTj+WG0ShnxGg8MP1oR16FUSqoo5obs5CY8WeZbFnGd7JU
Qw2153bkP+WJSa/kropgd1RaiIchE4BlFcR84LzS/7qu6Q3Sd4OQK5o2tvwC4o/x
k0hST5Ne1aB4SunRbsSgS2cMw1PR5UP9bdYzKlIHA1oF1c6kHJiIg1qvCd2TSG/s
Hg5TJRzPp0xc9DHcD7EJC0e3PZMCqWnnXwQVH/JdF5bXbvc+HpRf1y0rnhoKuZs/
E9nd8bvaNrRK8QoDIPJzpPTH/YWpw0tWuF/12zgnaaoRDdBod+qTTnSbSYagHlIR
RvE5EUOCnGMh7/Bjziu4XEDOBnZhKWieJS9m5DhPyvCLGQkz5RYbt5Qp5RgF5A9Y
KRoVSVMVMQUpOaznu8RKpVqXFfvsgr0iMwV6sJdgjH8Efb8rME681gklWF9/kD1W
ZeuaJF2Vjk1nwzYO2IEv5WOGb6akxhCRg+VjFXAHnV3vkvtoo9U5TtxoXYuosmtY
pDRfY5qiI8qY9hoCgqm6xXimW2lAXyn2Z4KCc5lDcQGit9I+BKPXK7j4NXG9Tiaw
Y4/T2Fr469dj0yFDt6YFBYo6833TK299UHdygDfcVJ3/qwMRSDFxLP3kSa9N6tH6
YORSCWiKPCs7JH7eutQYxvn/Tx19jiA7xf79A3GGhcngasD0q6Mpaq0r3BM4zToz
4yGcSUllUr3/ZJQ7QmvOjOPnqKoG3Aw+lPsHpj/o2EfHP+vliK8JbWVfDwWJIUsr
qd9W/DZ3Z4f7p3KtOdxIFoXL4barQA0sq9/m8OMZeLfKIIKML2r01xbMVviAUXwO
Tpvyk7DA6rqy2n5erRZYGrtLu1NockQdBNupJ6ybomvbSDuKL04bEn/l/n2PEQcH
V8Ln/VBnMeIMVlIXVDV9aHyV2mnnxXbDSWzglZWUtHknPcngyjIk8/EvTLJcLnoK
VjZVGb82UAehUqYNixyPbIMBeqka5tNixuITv+QWwLgCc23aUkRdbp2mZOOQTPCE
X/ieODQ/nyZH0Nz8viLOgtKTdo/YGAM4yIWWLM7/YEsS6VdIYTDnI/po0588QsI6
88YEnuZ3TwSvz49WW5SrzOXdoHCgwNylrfDmi72bRdomWfhk1nAq7FxKVQJfubMt
1tCzBt43nGd5ATYD0uPEuiutCzwdk8ib6IFwqe7kMfMfXonsFL/wKIZsetZ2+b+E
Fu6IIeyur4MxHAE9EZUqkbxe48WhKfILVkxjlWfSi/4zyiRZCypVepdBDickakS/
+5NseDfHwR5Enb1gqGwu/tnCKlWo+UUmGISmao3l3crSB2MqeGjuk5O7VIlO/o8o
ULfMPTKzkenzXN25TtO6+/N703+cqinP/p+xqbwDM6y1KqAI/Eo3OdBU0aRl5a86
OKQd1hgBCzSjwUFvj8PG8hZRaGhqdGIUV2Nfux4tXTluRvtH4CAJ6dOiwa+/peWR
tpyqJbkc+7jR+V72jRzFd5msZDaWQYQXHG0yFyYJpRuxMhuHGNvXz1hMSm5AREPG
Jo3m0DajSUP6tFWnTRkoWdJcC5yXB4gWVf2E6B+4tYtQ4deuzxinSpYM9M33/9NR
r5B13FJuaPZxUTScMV3NO9gX8lVQtq7IX8MLyt+7gWN9b6+IMhhmBdqTJMYS1VZ3
Z/nIGIbTsYG0vX3Q7JhTpc+Zu5k1uWWrIGk8UsVvh18QMj4tSUkoYum8adGk60mT
7FgLqfJ3abK0Xg8keCVhpZVkUCA3qzsXo733TeeEQYDVN7mt9D3nGwETl2yaZmWG
Wj4veklv+lL3hR3KTH3jSUaqq2sLMNRHA5Qhhx230Is2rPElHorwS4trwZ+1PryM
H2T/6wM/ULbgnv9iV0+eioaQRoFmDwB86eTkN6aD0j2On7O70Jcbnml6Mtf5uKA4
Xo5T3WpJG+vrGbuXFteS/sSG0trmRoCj6FHLKV5puatJtTEZYxu/l2WipaBlUYlk
+HjaeKmKA8lONIBY4kJfAQnzZiNpdsEGez/msYHIkaiQeyjP2XSOooLDzteV7A+W
4iyyDmUs4ifohkev6wpl3c9U1bcomFUnzOCWOgtLECmLebtg5g5/2OzYwJ4kp2Te
TSBEylRT8pBf56qRqjINLp5BQGgh0g+MAgvIAPzFkKdS0LzGTvRdE5Qyfw3HfpIN
Xcj6+4GBVyzdI6gyLPPnpmblY2BVsduLEzmrXqsXMk3+hXCw166ROefN3pSoiYdS
+z0eASwh7wVXClEztWvh3qW9UJ0AEzOXZzzLFkrokNO9N6kzw1uB7zc16tjgGBrr
oWvL101Yrs55ea8vRra0zSZU3QW2pKDuzAvbDW8SZWSla7dO9I3K4ffpbA+8oIgg
dBGP6vS00WCPNKL7ClVvv/4/KEVTxelgCI7GhM0USS9sIP48CK5sfcBuqXZsLqNK
/gKFbp1T+Pfr/Ti8Y5pYpTrG1H9b42ImadnVttYNwjSUx+yHAMTk4ZTUkdPO2qEd
H4SPaD0Ds0KZKsydNAY5sAJYT8cSaoBOUKlWNBb7fJrhoftKSFpUOx/kvkYPMLV1
+/D1eW4oYUEZOLb14wW5sBodpTdLR1emDy25fWN+lfDuVygUEwJNoTmjyLofYMBm
9NSv7IELOVeESKQxxRlAD+DC8brQNjsEPJFdMrFNmliy63DnC7wwTY44TpeQunSK
Z2VRh/BHuXiSwmyPAyUmDxPzoL+WX4/c296D3SisNG+d9pTJ8R/tPQlE0SkEHy/B
1Gm6hgMQ3+IrgYoXtg2pSf/kDiRuIRWQJ/jL1jHqc/mgditmRwQSK20noSr3ZE5/
PdasfQZhQDQi7+UqAwK452u0pGhOwMxK5uqLidzPss/k8fSIjHpRcYhdTiZ3CtSB
9Pk2LwkhSuS3CSVsv9twZfMHJEl1HAGVahB6I5/5MNYbnaLcVKmYGFh6EZFvavm1
aWAKty2MLT/Q335oAJUW1XhTMr0yz27C/0AWj+aHqfTXiSGk35iaAwxzXobh+AFF
+09p/kiPSfeV2gHziWCNazCTfWU8f2gElrJsPy0TF242xDDtrVJnNNlGbO2DDEB9
EnhEVrGwAZIiUdxFGWWCSgOOkgAYFnn1fnD61pwlSqN8+hIzcBCyU6HGq0rg8lEA
dy3dEAB7wJt9O4/lOkSYXOeryroNKNMyL3Z/V3+M9knwhHdXrJaPGYHqNX/67fvq
2il57iwsbvYmChT3cRsCWZp2OmA8I5rvlMpuU4SUACWuGRBOQgdqlAoYLKK55uBo
wytzUvKH1kMvZRPg6RiCPturbbqkHhbmbalhaUN1LxJLYXCjlfSQLgeWvVuDr+Ho
h+QrpUe8c1CkToa0cGBM0/IKsd7vP/kNZFGoskOj5WMFwx5uuaNWsS48MBIUy+QU
hTpZGh7Rd852onsSrfrw73cPwI147e2aAhd7ZOU/M3EqDV0QpbB22Reu0hdK9Pz0
B9XgDmx4NNuUDqRmF/Pr/2KDTBGmFIxzs3amCv0tWuuBQab4/32MYosnY+DJB0K3
hoL+DyOMzokhFVRJToQob8iT6LiZ9N7dOzb4K9//NFyMO0HWmukTZKOn0SHthiHR
/AsZksUU0Bebz+W+I1Qkkct6JGOdfEB5yqSHaG0eUGE9fMXFbN+lEQj4iQzqb3hu
OEtslfDZZ9ULldcE1W4w7m1AIhLx5Vy7OqpTNSIgSHU7msa8gUQYZ+3nBJUO220g
TU3Vp75QZLHeQQiLx7xLYg==
`pragma protect end_protected

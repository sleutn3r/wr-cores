// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sIgdV3Eos/cqKd9+8GdIYwqb0rwVIHsh5daC2h7XIYXy9zxmcraXlcBZehVzetpT
/+E6LOSTKpIUZVP6OyVDFL3UJbrDyAWdwr/OlwqlSVB93ci0XaSI4BM5Bh7gSqQM
k0+a5B+5ZuqgMFvJiT5F5U/yO9KM7lfu2DC2ouQSA6I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32064)
5fLm/tIwzDJwv3RCiE8Lv2gdxY7NidZJfxCky5jv4QOMTAaSUVAiJECCEMs+hHAI
k+ff20NO6jyT4WXSuC1G/NhSSVGO6RSp0g/h1YLXclFtEah64TGrOA5MacGAo0L1
7ehWWfiQGRcavMbAJze6vthSBaUlEKKn3+tGPQBi+kQq6uZy7v6JVAjz3RYpj8JV
4e6v/LQljs3zKFfXcf1sb7aXfSaUR2YL9qpWaD326K+ZFnZd7nZ9uWJZR3KF6pjh
abXsURFCNCgbj+A5BlA46pTHmW6veiU9jlBh9kDuxIr52AW6c8JhLnnQt400OL5n
SpHj+MB5tAnq3gGeQgUdMDujojm4JqUIqrpF7A7Z6Tz/LMaPOGgrliU81CeRfwVP
HkPzrsG6zZPo4qG9DrN0xlifxQ9j1+GnNZLVNYe0PcCR1Qd9z8KSMW2DPt51+DOZ
xaLJC3T6HLR67Dh99aIIJEUwVCUrUA3S3l4gSKz1zBeruLET2afRFDnoreQbxL56
obsGz0WtGAn+vlCFxGT4S/6XRyj1xlXN/Z3S3YQ+HBB13vf7YykAk5E6rmiyAOPG
a7wDvfeAHOIkQXWhOz9cdtcr0wtlkFYyyKmRZEOlpDUdyZ2b2/mybQCEghtNCuP5
gGJ4r++AbYLaRYlk43WNX3t0tdN1ACpgti0CTF4UgV5G8bBbNNVZQPQUhXngRnwQ
yGfLqYkTSM0+8WqXBw4i1yO3kFxC6iRMv9/2ydcnm3KMA8MFmplYwCTyNDeBFwGh
XlWHZUL2jMaE0T+3Huf88emHi8Wpm7e0TAHXQcHyVohI3UaFCD0ogHeisIK5BVQ/
UoIJoX6/lPVnJuOTVRRUJKu7MtRdkTS3+HzKPIxrttBeZCzhJcirPc6nkapKcgrv
TM8A2xH1znn9UQ5wh9TUPewHc4Iax0S3GGqmnzBtzQM3RXY66Q9IbMMpHRgWlvYF
Ce6VsoA3za1NMMWGzoY9xFFekNNqQ888s/Et4nRLHaJAPTEWG2eosVt7Fe/cX/wK
kI6trRR9WXg3k2dQFsFhajRRCtj+nhZ8IIrQwz8srrWz2saFfeF50TTNZNkeSXy1
CqBeGMIFsLrLi7uttoI4CO9/iNdmGaqnE934Ih1zypXfgsS8q3fNp3gQW5DvRm9s
H2ZLPZn3HIY42twu/vaMTacxPu8cKs7yygP9hrTJRvHqtQU8ODCl2aTQUvW/yGJt
49fY3gLRRG4G/SFh46skzkBhG6ORLHgcYqOm9ngKiOISp6pnzgxABnQNHUTqqMoZ
QFGB4C3rD1XDOGtAn7I5jquHpWMFslZPK35HVAFvLCkSg+0UfvZSPMr8oSA6Quxr
tJvrB6PH3iHB44VfdUyQcebBboXbI1KRbrNjO8g2qiR7hG03MIlNIsgM37cW6Hue
HKM7S1LTnefZfNvmy4xRHFxZw9oQlJf3EPOw/Eg+l9GGccX/6nXJp4pHVOAZ8g+2
IhpAkqUoPMkQ1NkxtiwIIKwraNp6XwbgUDMXGHnOHZ9IzXH49+cc8/QYnZgIFfW3
uGdkojqRmlJUiYFCI43TLKGVoqeVm8CRASP+EFePg56jW/RJxc2R4B8Tccxv8c+g
9wt/ElDYS54plzM2dLIVV2hxAwnLazjps0fp1yUm5WI9M6y4XTG2e33b5A6t6Bsm
8X1GY4X0qCUre+2S3cdhvz9cJoGy6HTLCtL+m8hqfSbPbTbqc+XqAmH2reb+sGzk
rd8gYx5Z3wyM0cerCYWsQiOh+cdXnAMTbDiKuWYsO/c8if3zAEqH7WIdz+vR4/5N
n1XmXOHF36DNZph/iapzL4bN3qkGrOZGkskxCGcC7t2aDktSdqKBFbcCdPWc4ryz
/pL3AidcaphZUFoRgDcIh+ASU8nt/v7Bt+f0AZ0HeIxssNTQkUz7IkBKAcJQzHsw
WV9apEQAQEgo9junypY4DkPVb/N6tFqoqkH1W6FmKmAMYZxENp/OiDlXQTCunJZB
ycP1l643/WGfmk1DrIZV4SKjtw2KSjCz434PqAq2a56aL5HE9d5+Qum2z/HiUWWU
KgNo0HR0Q45gno3uoHkHy7cDBW8mdKcZ9g91KS3x4z5zZ/edziEFTRCOj9i3/8cv
6qy9SjpgnNh/IJGrF92RI5gl58/LnPFcw0PqKuJu6aJVflONcOVYnO79zGvQ/IKX
tWUSmp5mKrv4NDm/9sMkwV4qxGT0RHyB/2wJmmiyJI+Yeraye2fbSaKOocrg8GN1
A16aVctx+mAxL3Xrac/4K5iT+2WWN8a8hFNPw6vJBM9ximcdi84NdphDpODVd5fP
IpAIOaV2k69/DwPvXmW8aOlFMmVRM+SaD2FgHxlRO+YSGqUk5sSYNyE0WVPiO7Kf
KJT+oL2Bw3Oj1LKkrORrM5wqzxPXp0ylAl/0lgAg1rnatn3/Anf0je0kGCPa8iHl
IEpzSNRhf+yt7hd0EUh4Xkn9AMtzgVmOjhm5zGh4u1J2wlgXlknAJPeAOIM9cmwe
VfWbujjlVVqi+UUhAOnXiGQlgOq3bP9Rsocz/bMP3cihyJSeCvcByej0/YzXS1Jq
nhWe431LGBzoWje91+brrKVyYiDVjDKk4nG8Mz0fbS+SID79x0Bm0xdnvrfClITC
/1WJuD3sfb2r8eHVKgupow47qVPtrUHBkaEAemuN4SIhMa0Xs939Cj3AW/K0Vqe9
xPkU0GVuOklh6OWRwCR/fKoLnXyiZAOxs9exwHqOdEkVaKlDdjmHZ6z6/sku0sbX
KYevnqZx6ftt21tcZ9BXVCaqJRevnoeSt7BoqXYAvoHXP7bDmGoAkjG0/mvrdXoR
/jaCFcjS9214a/2orWqi67nyihX9exH5reQAinVAraZrbH2jGS45txLYQBsaKL2/
pz7zPW54FLmB/82fAi3PZxni1wY1tmzuUcxU6L8fC3zGKEMTfRz3leMMfFDrt5qZ
a+4Cb3H9EqaBKzxJQIn0oQdGDIkoNGyKPVzH/zSmpAVaCimGSAd9lBVRi+pAZYew
5E5aKDUs1FONzDOzVQa04aWau703IcSTB6SyomyozF2io+cHux18/T2DJskSkOFL
drPlaW744R3ufC0rbBgFaxw51i8ROTOphqz70pSWQ8f86VmA3h5e3uqUVc38QrlV
8wU3ky+9fx+m+TQtwKDTKSXUhH+d/Wy93BUGJZ5g3dXeuobptIToH9PH/ocFq4Q6
Ox7sxCnaor5u/TafHRcVvDaeY1nrJViKgeMY2GDP8wtdGwu05h771nEQurhR6jxz
IckhWYd1gQPl/bj1nDwAVfPZ7ONI0Es6SiI+TrhUo/Rt0AOlvl3UbyOG/gzVQrdq
ebKdhM3zwZOz5AiVdpXI+a+12x6EZlJD4p8uKMK/unuREX76p5kGjqUrG46zrP0n
nq2bmzxxmz2TQ8T3XgkHBxad9zMUYPBYe0a2rYi4r0IbQni3/kAksZjhhDo8lfZW
wovjE8F8HySF0nQnP/g+JEwMTcO33O4DmVF4ncYjMs2QGWmAtd09k1JKpnG36zvz
6wrRcqRMcRgURz6koK/ZgnBgPo+fYzRnbKR/ZOLrnsgD451a7JAGiYzcnqwdlfHD
tYeHLtPJEKJj8+uhGTUPutTyQiQkFDGPCYCzBeeP7e+5/aOnfM+7oxaKWsDEegN8
PsBcRGISFXPvDW2W94pzMAEs785mfoLwynarqTqtw9OVXykPVK6+FJMZ10VH5l11
B4elI5nm6KlhqsGfQqhYs4MY9VRBHm8vD56qyVh6b6k9gjhtPQ2xPF0n822eiIlN
+LS7GjWXn+pQkmwypKhnFWZnDJdTAH3Ye/0gaRWvq9Y+2AiedS6k4z9w2TV2en1v
2iled+APUmHOqgkq4zMx0jXTC5/p/q9ueMzBiRCxg6To9T5OlmjtuycbQ4rsVkNN
Swy8XQNsS13/Tbxsj69zBIaeOJopuamaDcpss54cH+m6qnhatPco8AN4Nk10dFPW
4Hph0JgUUwOxngiTvikD+qhjvdOaGRXiloBtPDTG9Ag378pwgCh5GQHOAl4IUry7
3/wV7uZ/dix3s8o8ku6bwAdOFbfE51CVH1fFZ70V66kpueHAA3Jc2YsNGcbmIgCK
efiLXTnl2XJtWNScVWJARzDVNorj+eoRmdeYz7EDOpXTvenat3umEwieiRu9T4t4
ZtrnD87HQf5XhLV+Z5OZuCe/F6ZRT7HK5ocIn3n4zs6+3r6nHxpvdyaWX29yK2na
QaElpcZwHdHPZiLdhfxfSDAhAN92OgPdk7UsgILs7Z5neniloJlA8OinwjjV/73Y
eoa6wo3CMR/dv/hMLeqKRs3HNpvtipHEeN3PtKkw2TQh55lk0PfFO5UakfPKjxxQ
LpNr2dT7qGVfaF6DyG4ZeUYpT+lYs6XihRnk3pn2QC5UFY2uVHHn15jYJdaGvzVf
EYbhNM82Cx9eWIt6Rfivl1g8OzILGrcEaZOb9Q1qRUcdohROD02g6o3CN3vZT6+H
uirGotixshSqD8HyT6tsF+qdaBPKU6YfyRSCTkhZOYRTi6woawPGhBdWRsXr4NHu
1kp0cvZrSpBF4HIvoXWasaaeVttFFq6dz7kcAUEDkrW+NwpqULVdfiBBE9WAgkJA
VM9keeu90x1Jjw5V8QecaVn5YAeMEiUGc9oUpOeSu9/AcuEO1rMpCKg+VwoNo1sW
YA7k2hBpf7GWYz8oGcDDjZVLCF4G5Bcdz7DiNgP06M5gxAOdku6urThQxCAzObAw
rHThfxvlPvIBr50CgoanajW8dKIqKN9zKMHo8dkLwd4ROehlh0/3JdW7Wibj4TrZ
7Wm9Y9xWbwx05EX75wBNXHj7Lbf+OosNAZsDCWigmlh3XAev53u2b9khGtWLzVo7
fNRIuOWxlzLAjdUl76V14/JZ6oB/2ZYKK8yMjbyP9D4Y5E0O0WNXdXKzjhFCLJSH
Nd3nrVqIBFPg1L8v/3xOxEBV+2kyzHGbOk9bsYAeH2ZD0PBfHgcWcINoKgM0PUXQ
fM1nHJbHTz5tFmEY6BSz5YWZxWc35U49gIGmItkimCC/ay/UmbseuseDlcfuh5Ea
/sx2EePbRK1LNpJiaKkgfuUX93zLKxzEYao8TTXFkndBqKBWt86/QLwwdmJaXTn9
3qB9FQOf7iCrU0qfaBTYBphTA5Tvj7uZFcnKCKBWVNUH7EOSX7jRnqDOKkIaRigp
djfvjDV75wHQJU94kLl5lLWhfj4aTqjAS5V+LCCwcCDlvf4QMoCJ+HNTqDJp3NKH
qPBnZS47pdmxNElPb5n+D8fI2a4iI5asiv2VPRvo8RWogywuI5NeJb0FHfLX1DA5
wgzW1Eomh8EqFRABWxexXtjd+8dXmS9F1ZIM4zKz2Fbjw04PuiToB6ayqFqXbisG
CbkT62vICS9iNvWxBs9h3TTvx+I6KXIr7zkL5+K86g1O1wO99kEaw560xI5cCpim
aQ6YLtBSFOMwiAcOMMN9WxVHp7ut8lJbxZEeZwnGo3V+1astSi2UYiTnJ9ydZ4nu
ecIsYnl0+vObbVUCTEy13HdyW4eHAlR8LtYB7yHgOeH4JRPZqJu/szwJdkkafa+8
M3A3W5rB77T8z38/vu93MKCkNdDvAxdEPZl+8qeaAnS/ptdIBeEpjB7XZ7nTf4IO
auusSigwsX/Und62DINAGQPU30qC2td8UP0mOMbw2HLQ2djnUfSGB4iAcfqd5HDs
alY/kiub1h/ryoncRQT+2NCozsLZ+GEGSiTJHI9Oa1UZ3ShF3oO65MV1oFpQ9s4p
ybv14l6eoPTBJb43v1SjyKsCL76FJzGaRWDvnTUK5C4xqneI8uwFq+lygHyxy/aW
iNh/JiKuyJjq0598pjMaoAm4smUEhXhrfcVVUmO2Uc1M9UJbwzTjtenmNx2UfoGF
O3OYfcTPBUlpr37O9or7Amj2gws++9C97ZcpFFNQJ7Y5VbeRmU8Tvt9Gq7ZMFWIN
YPXMR0vDzd3zWjZ9qMVbrgH/Dx76JJXYYYJicKjICiaamFdJWkTDTWfquMHbZ6iP
H20u1/CR0gguFSmBZsduayHJiy19vHg08p/ax6T6fL4BY7ZBHdKOQHI4pJKBYhLL
Fy1x8KFVdMqILfJgfA1BvqEBowf2Jh2Qy7Ko+ezeaPlv2F7qs5tcIfL1+lu18N9x
TL1uZDtAtC2nXQMclu7YBY7TfJ0L2di5mE0J88kddQ83Y2yNHQbryZCoBR9rV/BC
u56rURRAMJzD3aMlBB26MyeSYCleHrk5BDQnJLJlfJ+WjiZoTPKTrWSf8OIYf6AB
u/y2RzKNiWJW9fNFhzNZMUMgPeteDS0NjJMQ/ZelFKxIzt8pT1ulwRFJmOhJ3Ytr
+urC4wUWSBrW+jSJkyV4IQJhnR7C7YrW+7WNpR8uFe77g8g0MHrmuJU4PCyj6l8b
XGnDqC2oHC/DUAkgF5EG0rd30Y/ec8kvs8ecw/m5xXrT/1S5vPvUs9BM7ADCActi
pjSAZDBX6PuG4zq5BttX7WFApZLB2aKL+TvjFONgalb4enFDz11U+/21iFbIkfMN
wC0ma0v/1/oKhJDnk4+dz84IStsKuFWDqHRyW5aa+q5+G8vVzG1RH0NcnVajW1b0
/1joUuhuquhUHk7uib7h2M3l+rVMqB+egwfabFfKfz3ezGqFq7J4ZuYeIGVWeOO1
e6mG2QQAx+t8LohB0ekHBAYamfvHNIsWh9bYK+J1Q93uSgpL18I6+Fyh87+Iiuk4
xxWr1co6YZVitypABHqXDzIo/eJz37ODAqx0LsRDJ4pypBXAQo6kO7pNO0Wz7JqX
nvhUrcIdIgO8bZSy0UhVqspZ02SgJjm5TWid4vIedCGd7LN/kYxi4hFiqf2lqskp
qJ9ukCJEf2dDF6xdzlaI89rgkEqYWki7a6bdesDxTzKQRuJ3HgF+QzypLQ9zGs62
CmaV/iuKf3h+lmJ7Svx96UwmBeo7NuSsmAdzZeRW/fTje/TKVZRLfM2ofR1JfUx4
wWTdgssqwAjSzlMbUS1AsD0jjWsh6d+Rtm23Lq3YnxZCvMStVsSHl7MevKfQjUwn
Mno4nGZF8lsB0mRpfcg4xWN63dW3q8QiG1IVnquM4kOIsNy67b8oSQYLP6dy3iTb
cHMXZEm9N1QkE/TcAkrjqYngnFUR9UMcXgM0rOOrceywZAyMS8ywFw5XZeux3oDs
y0Kjm90rrmFBKHltZMrXICWdhAHk5pk+htO0OboiIrIpAhEiXpDdNxssIjACvXID
i3bDaOZCwaUScexSTZ2EilHECM4anektMtbiCDGJhfBsOP9Nmn3eCZ1306iWUj0l
FY23lytcG39d5I1Fd1A2S2/XnShCQ9N2hIDhaEgeYQR53GKmojiNWucf7GJvwP3b
wfIKN45wCSRzC+CrI6NPGmT13pl1hVA8aA8Rp6BtVk9QzVu8S5/DtXJfEnXP03UU
gzOkEh3hPGRj6HF9fXEEAfC1SehQzLrqRoE8LD3LFNlieT6WvmMGSfLJk7cLZVH0
XdYHmRfIWmyDnsTdMwWOHQqPVeNTgVQXTzTm+F4m7eEARtR65gPrH4IgvCcETYN5
KEbtVlJHlprn2vpNSY4RsNmnpsClCOT2dABy9E1uSjRle0lWkKbaqX2ZJE035dtZ
YgePBISXGdHKwqwdpBn4gYcOuAXEs3uzYk8EP4fTnDfliEwkxRxHpLGA+guzpXaL
OxEgQlmt4cXECb3U4SV1YJY1kDXKJYs65vLVuYvJ3Wys1mDiVeeeJ6jPD3Wm7F6l
XuU6/UY1dIh9wYQ4C1q7LHE0Jx9s1N/1pD/u8D9sLcO/1FWEAmHkNcQS0Ixlt2oK
RaCyZJN4hQB5KTw/FAnYmWJqg+fP86H0zCOFLwkRtWscXhyf7JNom8bGOKqMNzn0
6NjoFL9dz0Jc8QNYWsEMnhm1Lp5MaVAg6IRNx6Lu7qd4nblx+uAgCZgmd5dltCP8
3pFANjZxY3Nrzs0ie5PHrZkLE1Kieih70Hd4sYNuLUE5GNM6qlgUJnTmR2nEVWFY
h302a/sGbB8xeQL79BfSV0EGaD3LhgQ9b+kUT+mhoNgi+KXRE0mWq7iho/oBpuYy
52KIC7/Pv8kUHuiy+jgzesE2cVfJ037ZuDynLUdztsoKajfPxy/cpvKnXJcvrKD4
ibNx83bQ87F79gvqT4b6oNGfsMzyM67Zyb6neGH2AdO1dutZGvQudwmBsCg6g/79
EzEJY2QIcnlDVv5DlbyBJVYCbO2YeOz57Hu3t5fpNYMY97PneMB/4LXAXyGKroR6
9LNiq+FrD9/npKPPTWCX0iKxQ9LX7I12YeA5fAjgGfSRzK1tnN5nhy7gdvCl0F/T
yA0ZePEIplFpyufuXb/QzFEPYY4DB07I2OxReAmaihWBolX7ds2gMFyulxK/DQLo
+pmjnkuGy1FNtdmJes05z4s+AmLTIYDXDZZu1rksMAINOhKrQERqDptxjpf3at7t
/ItubUuX7NT9L1p4WZjAMtvauiduEmebuXJIdJvViN8uvO3z56C2TqXDM27ioHoK
TcVfATvF6vqMRntVSXAQ1C1GRVlJ3HkHTAWJwbfR9xFlg4uVAU1mAcpAzZDsylHP
TDyc73RqfEPLh/ZQrrYNpFkXbOHfQu6FB3LOZhLSEQw8bk+C8Jq69p7kI0S6r5cC
FYjOWdBLSwc69jT2AvJdTm4kGwnlo/8LzPkbdBx9wQNQrQ1VYdKnztp1JdHylPW9
uI4b60qpPaITslBjTxSStuRF+XWPXTeQBE+TmbFtrd5OolsUq9cERgXPgBSQaETz
wqmTFsBNIWQlAs1QoL0fyk/QeZvhypL9Zpmfkk1KCkR+Wmsj3LLgwyeCkyIi8kol
Uv5NklkEUnc3uwZS6X6lJHVCZE+oE3fOIlgcsHGhMldoF73o/PyL//u8TJ9BTwGG
LV4s8llspQJkyXqa5YlpGYKGqfUEWVWvrFOUnhpkbkO1iaGophqoNwomqKxkTiPE
VW66Zxva+S+poEOeJLVkTQEGSrL9Gpf+AHNeclerioZFMsm0gHTeYNwpE1ISNLrN
la5tQx1l6X2WiPJ7YnCyDvhMZGNRzkFhLTdnwLYT5+IFh1+RtKoSBirZR10NOspn
i37U1yvogn/+o/OSWhRyO/lOkhqbdA75vWM5EiUUbbBAjZoIzp9tRazLhW8PeOAP
wVne47S4LfKE5C+2Oy1ohWS4CK1QiS3oxA+f9uPo7gqtF4KBgOQkXTp8Gq0nR8kH
LitN9dS8sOOC04bTSkjlhO3Fr3AhmXCK2zpZdwSlCvpMrKY4DxE5Jr1NWAFSlFiv
0k+m+sLp081znO4lF8RPmsp6/BKwdv6cC3mzGRl4qNI77UbOReR5uhvSjdDhZgT9
shWPLS7hLzgjUEoRAgQ+aejMbjhmi/VyOqJKubrWa0+oPOsN2KLU89v1NY1bPnOi
gLRsLRBUfsWBDt10c3eKrPoxJLJFDvuF+hQNcQrUpV3+vL2+36AalMm4e+ii/tx6
Fz+jxPOuzbsQIlR0ROnkYf9EgL5ri4BvMqUCGUOiaWZ7q2+mZk8GeVBIBklEG5zo
s90auOIYxRe8o5TwpCM2P5T7PDLe1e7N16GGA+SXVLZ0DOnR2RlYT4wN5WaR38/A
Y3Q0DxqK9gVE9E/bc1GG6IK+SXcM8RkzZZWSIgN/Pwdzdok5Q47Hlt802bBh6K1B
bM5SEFWFgx/5FP43XHiw85KnatGF0x29T29K0CXmiVgIwnd4xFK891au6hfP/a1G
8kUDxNMieDtVPa+Uz6DQBLaoo4m4Jvu/dtE6PbfnfDQHb42JRTQte/3CJ+IR4Agp
E5VXmYT3v3Ejx9HHeRnqiAGUW4CUfhosjF27YshcPu5ErTfthk6rA707K2iGjdhw
r04pS69yiTydKZ453/oqMFBaPIPNs672+Zu7XEtgC+UoFM05e3TuceZ1e0d56EgN
5Ic1N4ipbeaEjd+hnzXPVSisfnbxkfDuFk0uGxHIGPFxGzyNE8go20rAChG3rGlJ
fpyYK4geTi0Tubdm41kEqHDtEGgQjvrDRQw4EItFYN8u8ZU23ohPDNJxXBvkGRvN
LcHylLFh8Fjhq3iwj/SN6Q69NvXboYfC4oLFnya4xHWPJLYLH3FTlocRTbbfSqBV
EbEDFWh3y3P8L7SpTh597Cm/I3hk2fazwNgDRLn49edqoRXoh672zp18NjmwtF+K
Znrpv9EIRn/1csUKM7BnwaTldA393pXyXZLq377XzTQ+8KBKAZ0Wj9vBRMsDfgEp
8o7AE0vHOih4Xnhws8MTon+w5PhFrOwMoc7T7byBwjkCTLmfg1YPzIrJyGWM6J+I
H9xSV3eA1ETx6CsHyx4kf73+CgcednS80DI/C8cnnapIBBz8RwCqeO+PGiRoU6tA
rqT/FWyeoPmTEo8KSAVDhB9kaQ+dAoJRQ30LAZ7hHNpeB8vE+DEOGR0KN50VprAl
0aHDhJKPoPiG3TSACYuVEwuOXOTCnNGsiJ79nheOACGxPZfriFyDAGQfMK9gX0Rt
QPOVDdnsTGOouUaXe6O+uiq48HJv12S/fHWOkOb+s4s++QW2eACSaRVHPeyjKwgt
QGQCAukbEaGPqIVRXA0n47iRLO2vcxrfFcRZvxtogNwcr1t7mAQK9/o00huYWdAH
eqLDUpkpjxBDMJExA2w4Z9e9sihx5WtQasjm5B+3+r9b31iKYlCIZ5dtyhFo8SWT
hU3vA360iyH+p5v3ygbZPes36HUiR7bfSupx2iqycx3CqJCsz8CTRBjA7lzIrd9J
DL1m1nK58yqZluWN1/W00LsqAajE6dyHTk0Zya4oMMqmOoY+aEC+ksHHlwnsrzW4
/sLiDf/kU2pDo9SEX3RDOlgDNPklno4lgy7SamNq/5nthCBLgOSjGJ/+J/m3g81F
zG1lCB86S1lMm7Uu4OkMUCZeUzxsLVizhxLE+eq/+Gt8F1ltaVno3TutRM7rhM/c
afHn/gzQ+5jNhTcT1jzH6MEfQKYn0mw/C9hQXsY2+AzFfKsDlPDNm6PdCojVs1IP
GR+dTZN4q8gs1ehrSW9+DllxfwQp+9O3VEBH81QOVpqTBXHOEiPClWFpUU2WDCZE
75v8X+1H5ERoDvC3Gtrf2XFs+yYklFf8yazORn5nUAQ9qhZCuqgk8v4WxdMVk4Cp
O54Mjdrc99NJcUv6wqZls4uHJkAwLpBKjCzbXmoaQ6Bx6NVAhUxo7Kb2Q2XFyivd
bpWCKD2Y1JS3yrpOJhE16QN7ZJl2LgGxT0EXqBmdexOW6U7SpVAr/NXLy7oVER+t
SgzebzpYh1YF9KbF5dKayeAJO69LEAMnOQv7mwwgUZeqVToZpJ6teLkoud4w8sRt
AZUWpGVgejn4GnaeEgo1zQycfxEftOs1r9Cc47HDTZjvC84oAQwPLoXX40btOqB9
5Cxy8NTlatILu4+IK9w+rNRgqTEvUiNtgqIS7fittgeeKRH8FvxTJnAB4Qzd+c78
NGPI+HsFnhZftSxWDSQ/j6VKn89g/lnBQXDkJLBMTr8+3gZKSCS2XArzqvRAtCRR
mtTVM9ajnPFUz/MKzsDFvYSbrJfV9OA9CqAy5nTZ9WZlSn73ALCHvCQ+5br8fg4u
ZKBndyKn/yLF/6p5Co4tT2oOYdO/ZzGh7zK97KK8Y3urMZ2szdvwizbHNOAaKIAW
98kSv4UbyYwCbBF4ElhQNkz+6XmZRJFzItL0l1d80vQ2w3GiqpXlMGIwRxwxhyHo
y2NihXkynKhUWgt3sGnseQv7Kh06iQIKdCYiimXVEffOt8eC2v0UclUTHztZTTPT
u1Wwh0LSts6v2M8Gonv23YaP6/qb1S8RezuuN4fGNGk4nFDKfAuvaXS0wAmE5eCy
/g8Vo1kILHKzRvMfxg7YWcVE5vFAAjUvGkPume03scKA9od7G21cTQW5gOApyD/+
VEc5tXtVzctEzWcxw7p3mRO8v0COo1lHA3yRv0sf0HkInsjXkc+JX/FCfIwt/yUw
caeuRocP+3ZEYnzDrsjP9XUmAIp9ThIfNBYnfekaW/EcIZynzn/vW5sjlFYJ+i6M
TTcvv5fR8RyaIxayzlJ3JWHDGFKHaPlq405yJH1h8a8aAD/Ed8m1tXtXLndvv8Qx
jvfbTw2R/LOWxaE8Zeerq/j+lCh5+0jTHPj2wfOZtz65aIyLT3i/h1AD3NttQTYE
yH1G7f+X46cwrr4RB3L0FbO+PFzy/TjiY8113uBxihh0Y9bQsFEWc9g3RBPXNoaY
FJ0K1WjjIFlY5qmJBDqHpwAYwz8cozpSLVbkikeJ4xLTe8C05YX7ZMkBZqVxASya
nuNEV5P/UgFqEeYsseJjqYzTu0fR5pNmGpPbBHcYS5mqegsMCJLW9T8jmVjxGsZ+
MTUQJeZn5zTtEwOkULCEB6EOG5SCIs33h0bWW/pZrQr/0H9rEQw4NU0bwDBzCTmN
TCnVOPeNdUyPAa1gGxtDTzjw9dl/rhw1oTsLlrMzI0S5p4+EO9RjPSzD+H/06QMy
FvEUNU5uue8BVIcLmMCRfy1txNWTd7yo5UkbiKdpAqBa7vqnue+G0ABdLg+2gAre
yB1zcOEMoyMy9rZRafZw7Z28HMQtjsd180mCSyDhPOQhscB8oNfdOAO7fb757ENN
+y0F4G01lkjvUslE0Joc/4lQSo04Kqxb1dTFMdjdNN7kJA+i/pLhCcaq9ZrdMwtc
ooQUJ8jqP8jOzvykOdV4MC5MTc0xeLKVQN50kedtoHmxzXNmJ1jIJIDCFGvNsz74
wa1iktMnOcy20vvqVDqGX9Xx+MPhF+MDIUSbLOjyS4p22Ruzyd5E0V8sfbpkvGaU
TDDXCmnay5ASZA3F3iXhNnC6FroPiifNQTKnlEnwuODd2gtGsO0FJ/+2lncavCjf
0zBtqt/NdAT/LDrw+Zmw0Ik6Tw+rh4Kz8Nmmun9c/IZkxChyJifqw5bPdIcP1VEF
m7WAzGtRqc1BNK8qOljyIcjH3CN+OBI+rXmwqn1wkOF1TWmRYecdReugI1zVlUXr
gwcCC2jvjE+svMFafd/SqJNqwT+tQB8zID1sh9oM59HczXS/T0GNAMD0nbmrx/Yn
sG5C6tI/U4pcFAU9OySnmNdg1otF4hALBxEiXjAskve9Jjnu9i/zaUuF++/D7C5h
DzxRTyXYWMrd8bmJCAt33JikjgsZzwQT++1obAm0SZKNyPqoNX8afBkBTzHdGTiR
La5rtyO3n34gF0C/87iC9uooREG/vekQP1qub0NurmMFDZtMgoKzfNGTKphnuhS7
OuSrUuwkHYUsLpmyvLHkGM8tp/2TA2xeaLY2f383bKf+1NuReIbzJkwlPcNu07s6
WYBdyLpXXt3baF/bCrIdfaXvDb1EtGaoqJ+Qx+dfJKNKCIyUdIRs/QYo8yFtGwsd
AZr7PxK/XsUI402ech6NTQeesuuOLcbvC8ebQ4XPRm60unubBPJo3uzug4TET6DE
eSJSrtRO7V+Yhwk+uRoJvLuIjav4eqMSUmAcGnQxFdLRgT4g0+kXw0HLoovCLFkx
bSxW/IeLoAEGHu7HqZ/lckjJEdGdNhaMTs2gwVfFneQjfo7WkSJE8aX43bsqD+D6
T/UhQd6yEVGSU2g5c9egQuKSavUG31JrNAxo9/GYycxTLLUTWOHWUUC1y2mIkzJF
Nnl4n1j2L/HZ28y5YrxGYBhKqHjXVuFOkSRFhr8GD+vdfutBAprG8moaw0XI2Y08
vkeRN7ZXfj6DsG1T+1IZntLlIvbXgux2i+66oIpTNW6/R82H1c4atDuNyulw+LDn
Bgy7cDUVNRs8I+4kgWEKIsla/Ftvcn+1/bdnOBoYVbtg2JhJXf5sw+sWfA961GnP
4WqXCsfpgpaDnnZQ35FZSEM7Wg0UU4CrvHPnz/trijAmQHfhaS3taKIGXsxF1y+M
ywJpr012ygOrriISh0EwLobtosigtRlpqkD1lUjugW1YVNBMDWI2+GMMrSwWegWE
iL0nQ+892oLRUBT+9GYMZeXo0sJVRycCw9xMyk0v927jX2vGdDCg31NRcQUw5dRo
B85ikk19D9EMIiVD9Wl5wn+pYlQG5vRkI6iOoEt2RuJKsK42MXM4CZgEu0uR42pM
oILlWDWRyFvBldXboby9vFuW8bp4JNqj1u3WeQFLk5cZnNQyJoyQqqz/zWKYiDkY
rZENXrv7RR7aCQxDBIsaMweVZU2DxRLlqbv8GL/CW+XkW6Nr9kpAeFgLQyDqE62s
n3DQRqJR8yRC0N7pLVb0xOslekfwmgFIVdWRjYCMQED0fN2JnrZ6Ew62jgK7jCIO
OIt8Z9TEvcCoFhqLyd0NsBRtT4LnJLYKaQ3drfKNw2StvhrlBUtGtXab1zD2Stau
GgEE1ftmfmAeP0qi30JRcBIToshR0JpCqrQcdLQ1egQiS0op2Sye64UIIeNQV7W9
uxqBgeOK1hnOEA6X01iT4I30E5AKgpJ/ldqYiZqt5iEqdkbr4DFzBW/OoDVsH/bd
mD3XD6ARtU8od+e5ITjdQN2asbrXdmosslYtpLBZCp46nqM4U7dmDectr2SXFqBP
VMc780a/uVBedZCsvo6fZxn4PWB7miPPM3slSlhobFzjMFGtqweFeQs10OT2w64e
fp/j0Oppq4ybOaCFHfkT9L1Beff0l3bqb/zD45BVa7iD7LN/E6u+a6iRzbcbjKH2
FjAZWZqf/38ctcNG3y3WkGPO5xUVPGXyR02fKEjdUpu37Oa8sxN611T7loI4uUId
VIgL6wVbptQCE0dFfOFXu6DqVR5ZdNxe/N46bkOnOqdqjiA6VpUfUXe67Usxhb+E
ZaIrawUgtX9CO+SMI3DvI9vJcEvBZYQR6Y6ROIIfv0iNMKXVlIW+KUMHmahDa1Hm
XzUNM7hN2QrcEbX8ZdmzaYIlYQrD+TIcYqFwKXwbjVk8y9JNbmTzhcss+oQbGFyQ
VPdUZ96+OIJ+D/7HlMPQ8L+vaOebR21id7anlM5dYGfr09OrBz1ezejhiWFg4nhO
zWV199KuD04ktJJVXw4MfLv4I5MnuqCvrQqziryeTNtlDLPcNH2K6T++4n+EU9tr
DzS+ntDNqle3X3bkI0T6wsNnxEQvtUZdYbDmiYV+NPipHCA3i/yUc08JdGWltJcA
u7s2gcrijmt0PJi9vthlRSk/XToONTE7cq6wIkvHVmILpfBEopDYVDsXhlYWVIUV
h/TiuilyT4/WQTbP9eQwXpAOS4qkPKriTL++wD7bYDkRcNSDt6+9BWpUQEMn+rI/
bCwSPStvaT6cxzIdFRkET+ZH7ndP5HeTXLO2vm2HvvSbMIm729MIudJ+Abch5RqD
DKW0gnWe2eTnO+pge0C/TuDRHn9kPAjtIo15T/h8RNrYZVxdGEVemgm1sTUa2hVM
ISNRCaLftRtcXlHSU/1qCv4R1W02Vqfb9WbBiOVJexZdVIQRk0F6jHhdkhQ4Ulb3
4I6PGxt5CVaMoy5r4AnOuZ5W8VEUAOo/bQNONJSwQauh/y0RUuiYIeU/Y91ju3nV
2GVsZ40y9Wc77+WqYQl2uAq+QqTP+0OxgIZN4SsqbGpp2XHS/3er2wCpq4t1bsl2
ifrUWNS01T27iWGdCOtFrIGvm2yD7NW0/4+99ZQ5VXOCc3IIlzj926+EP6ZHmPQK
GBuWriuoZmW8e9IK34Y97F07Ha5yEB+fi+GqUSFdxDiyXPtffSNgKti864IWINx/
GOooxHftVURpjSx02GD7X8WnQE3LhsZGOvASBDohoeGC8pqQKHHEHQLDIdXdwqNS
OXHP/D6raXnkLJZXqmu8E31Y3ndTNVciNjbp7s11uF0BqYY4li7TYsSovav0OU7e
6pizLIgfT5TQU2zjfHJQeZ9/AqzNQ8FtI3yqNzNxaj83Ut5EbVwT56sW4OO4eGuP
guVqK2NkRrqxgXF9pgoT7mL7eEIkH97fqvtTdOXXD2jfND6kk9Ba786NZRAn1GWR
aPL9IG+2C5aHRFI8YUdU6c1cuQFWs68iTr81eU3lle9lS4+6bZXp9XodM+dBzkG9
FI+b6CgmVMxd0ghPK8Zdqlaz6WyqAEZ6nCuj0zNQIeKcP+kow48WkYb5t95qLduw
vnDW4srhbwfyGCwSfNCrAAsvfXPVvdw003S9QpNATwr9huwUYJRSENsGh1barmil
meqL2qvmQaDjjxLcqsjNqX2zxh3K9pzUjFTEmUMHkQdEfa+hhodl3nX5qK5UDcgg
h9Hhqb4jkCP+5J4SArouvAaNv6rScbJnwrr6L9Lwk7WkHhiE4AbUZ3/x19ULgwu6
+OXruL2e/iqvSLqA+5cqT7n8utFsgsnmfT9d2JdX9UJ9RJuS2B/JTGh5WZlmjzV3
zEv9T//LOdQaEM2q9sCg7IgefX3je/G/KlIqn/0ZLqRfsVB2KPRHSikCNgWBpchk
aoDOq58Ntu9yZNQlf3ki+uhYtmPeztu7j+sPJNZtZmuDKSiWpoODRBL3dtFH6ro2
7Lm/JZeqeOaO46MH2CCnAktAl1FPJ8DJaNK51A7DLwM7g94eVDPSjuAAQG3TYGne
FupdglaHEmvQfdnX8FE7uXxkoC4yAw92kl2gZs40lOo99Q/QGnd549YDZ7AlhSE0
SMgnK5cHI1VPPv+UFRvHWl+qrikYxmxAr0ATgcDPUCjKEJqCRfts1V7UV6+KezoT
16y0rTo/zyuaJumDjuYm14pVg50aL0vgn2LbjInCHjnavTz9qm4CHQSEl0P3ndnP
LvOm7jIzSQIa1t638I2ZQlqg6eyxf6MnJTHvD7L+rWMSRb0dhGDO57RpRtwqEkWW
ZM/12elS1XVUJmzHlRFJ2vchnA/YMPIfN2qddBoRK1xrtQqXQcFjigii3UViCpoM
xySGK1O72H40BmMMk2QetrdpxkR4HyKhzssRk82MxHS2t1qcoWhz4u9dUel0m00G
rZxh8L0d9VHTyMqGYw+azQZpkGQwYjHSnQ1YVT2YcbWCLZtEZbP6HaSeQ7m4mYrX
RkcVqX8Rx6KhMrZVPFkJfJgWwbFKDAqJlb81J8kuxcjH3W2DlauJWjG4SSFMydPJ
MLiVrDrPm8AvmeH4h8mPz9KkvmDKwe4UYKfSCygw6QhZlk0Ot5r1gB+Se3Hcc1g/
STOnYuRUhgCVr/7utjUd4dG5ShgPih5XKSSQK09xSM4lOoiqc8WAy9px+WCfp84i
fQUfZ6FZxWI+ejv/VZgjfK5jjDExmjnsGbLlnzeQGeYxTpuYH2OYMnc1WQ3Eb+eO
ftAKfORue/kAxC+gsN+irlzg3NzQzOYWu2JIeRmHV5QH70mfvQiQhZb3P2+isih+
3YHknPnF+jzTMIrN0lrI8ACcFpQEeuMRg06XQ3Rvy9xct4wVxoQKSBeOEaQYqfjp
7bpZK4x7khHh1AVRbqAqxSS0iycX5j9Nrn2x4INidpgP6KKVt6zbUkhEtP0roJw5
wxNcnj5Qy7zrNdnhBVTmA1R3yivgTJJh6CIsWkDqw4CeHeao3twZ7TIxlooTmrEV
GLik44ec0QOFd9Omg/rCvGJv9QjXI7SC+pqaqmMO/vWhPIghxRhFUpf7jplXiQbl
jvp6nQO74fv+kkXviHwj9J9jkd0Bh07rrLXUQCCRfAnXqzQ3/B7YDpEaqEqiabcO
rApnUhL6AjfkIUo6k+79DOtxikr36dRcSPqnRXOiA3mrMnp9yAah0t04KP8/5R2f
0vSx5IaymYNnhPIYjeR6Jcle/JnFxo5R7tz7J6eXtUcx+Rw7prBJrBk0UV3c8luT
JllWPwE3i2et2O8lTilWcf6CXIk7Fbq1n5htY3RF8XrC57fQGEHKUznXsYCIdjzQ
glnRHQDCRwqKlNQnmLDfDQo04WT4srq6JPhdfX5SFX02pwPEYLmxl3F/6yS5DNHG
TFiXtNPsThNpbNERM0hZuBN61MfYjij2/kb00iyc1F2oQ9cij5CQrhqt3+WoV6ao
qbC+RayjtRGBagGBS3c/o1p+VU1iPxY6YYkVn7ncbdFWRBLG7wlM02NkNxSfs1zL
NHlffKlXiXSOfK6gpdoxCHBG01k+N9Jy1jIoEXOmIv9RaolyP9dni12chfq4/kQo
I/iRiSyBcq4bJzADEbO+VcM8GtdEOMXdVZLpjluukwsoV9MLhpvSJp8FzKmcwPDM
2cT2k1Y13xlmHhg435hIicZtAhN6qeAmLXA0AMKPvD33+q5hNiViPJXPnGCvu8se
28pcwQpNxQTAZaJ0y0/ucuDaTOBBsnNPIciI6urlolthJfiwTuaDBk7ffDSLAbAH
MbBKo3cVp1FmrgC/Um1DBjygK5XFJQruu3Nf0rKf5cUkoyv49E89r8BymJC97oOv
r8jl2CW28hHp9YiG5YvQvpoU5iX5oClMgi8PSeHPsqaCMJFSGiX54lLOkF9d5f59
6s93ArfwmPelu1JUlkJSrBGtTKZmYo8Hp7rozgKOarKRhAzWi7QHo1ABP+GL3Yw5
lqA7MFwOOKPzIzvc7uiLT+Mgt9BYM6KrW/7En+x9ONuebcrq4uZptyWYP+O6ppxT
DfoqWIBN4MUw0seyj8uptfCnhAmOAt/dCn1kfxorEAc8i6HEdLw7Fe1t8aqON1up
csPMz0b75nIemUa3Jff9L1OIs7lDCRKYDLmEl66P6f44aLcykHRExeXhjP5xDhbA
+vWXzipX3TeydvUn7Au1xPMvwDfiopu3Sn/6uAoYrXkcJmkWxRo40DIEzCZpHqJ3
V9u54NydBPCd9fMIGa5F1rnPrEqtcfcwU31QJYtzXNBGsbYaqWpfKWsoacTxQyVq
dGszBoFpH6sZKajbMjt92KHeKMwLBsaIjkET1iWZMDj8p4GjQnTAUcLOiV3eD25p
czNTD5W2naURw3Fq0RGKpaS6wAkmyY+wdWRsb+n9ud5Ksr7jQplEQ7LiRX0fyqJ1
iWrU9wXO198WppoYyhwt9rOcXRCz8MoUy1Zfn4u9TEvbnLUAM0ZElJ+c5aTR6BFu
CCzH6uhkjHZArZ1H1ayiDMyK7lgx5rpYleLeT1F8GfdnNBsx/wI/982RoWdcYI2W
KAzBe7mb7VM+ulI7DysgjDrzbSqMSBGNAhAE7g2paMJnvFaGa07QsWQXdxI9knUd
EzawZszyevkuWrLzm/i0TX53MhO9JffIFVTL2Di/J1EQckSaGL5rQSNTG8+QG9rr
nDQn8cpbZ/D1bxh0mpotCc+1pdCrk6u/j9F3nuz90TaOZEmMH5yzSfGJVopF5uxs
n2k4JD2kdgTRYWtoRWe6ilKJfBs0/oR+rkEO10bMvoazrakGAfHP5pK1eVlN/nE3
yMLtKo0AN6I3yEJEB8W/G4Ss6kitnkC9yCkB4Es+kADHaLkvq5DcgajeiTqZgcPo
efwwMkEQqCTzrCkGPY9gDb9YijzkV1NhMF48dhqiX0UbkYeXkqYRCqtkt4iCmkad
mrXKMqeE61oT8k9p5Xseb0k4kcQHyZMGrcVu/fi61so+myxHEoAoQEp531Gy0Kd4
YNfb2YJbZg/O+2GII/2zkMySXvHvCOrhrN0r9M7QdWej6FzbXkUIVxuZ0ZI6RQQW
ZAunKeSyZUShBQ31hGDd06nxoMtHxYMWFygvWC96rQMIpgdqH3L410g4b4H+K9OS
hes0MGt+FosA7E1GC4ORGV7JilcjAO39ymKhg3mA2eYPpoUZPDyZqcCGJXSf6X1T
r01OeAxvZavDKr/0iNHXYWeEjmc2HwopLYnfQhkhhWElITECiA1XQdyaJZ59ZVck
3RWIZVK+Lrvt0WP83Mm4A46jqhP639zJ0Ab3oj91HY27/veon/LhIg1Jk7iz46sb
EHodZ3YhQDB5Xf8ymyMufhR5gDZXzhvuLVwm1ez0ZVIOU8OMz+krubs5VUACW72t
nDNzH4xfUpkogd330HejMxndBSZ8D6CX4PKhVXPYjQTu/I7aXfMa6SY0P7KezmjJ
z2gBVXiROaV6OJTjtMcQljcPxKdun8Luyc2+DBUmQwNRGKQbJBsXm7FSTX09uloP
+TzhlN/jyD7409MhZudRW1e7Ik5u98rg0Zy+PHfKRZKqmlhftTsGJLEGuB20Ocw3
JBzIJ8zSm3L9VWtTsig3seieUlvwmEjRaYhG4a1fV1kVuhCwCvDpeGn9d7MfgAQI
NE4gcM+GF7HM2Jl/ySdbihpVq+wW14wy+K5Po+OSsTU92DeOHy7BNkcgrtY9nU4N
UxXNHhVvan79X32VuSs/ECBqjiQxuTz5VXGTSCv3sSau2k1Ho9346YVdaCoeeZlS
g2IxD9SrXi7lxtqNxA8UFNDlAhq1nWAZDYQ8eioWBxZWuaCF7IiO+s38kNFL/J3z
oovP7mBxT6rQmHPQoMTN1pQv32f0vVzNKsE5Hy9xolmDhRGyuuwTbZrkQQlS6fNP
SXjGH9I+a3DW71URJxJQsc3dgogPzBRrLNu2XWhKyaZF6kUtPcXgXjbi6NWmRVgP
xhOjWuXdB7NfbBryPvCOkkdHlVnxarO3rXjn+yMeLRB3j+WQ9TUHRBnbNItyUfFS
1x2pI6iWeVJDnHaErWDkFPlzMs/opNUJiTrrgvTE5OeGRI2xFGKfIFPbZm0vYD9Z
W65AR1arYRxNy8WVAhOHdP6o7Ps1XrmaLR+8p+bKwBBpkdFC4TwMg7wLXuXxX3ct
a51y06v4/XWWyV+G3dERFdMOT3jor9scu1tYg3J2DaF8sSCnv/T+WdhfIQaC/ELE
LZ798xySJFyUZk4/D3swZnwrtiWPZ/Ey4YxTXcUC+Xpdi/6cQVnuxFiAKmVBR22K
zCHhRNBr9ijXu8yp64aTmXYs1EkIXPF7wRLCeAlwZHVCArJryACNVDXyTmdrG8J8
ZywVxNyOmb65IvxwuE4WcV28XTnX9rfjiMqyglCUewP7bEBMTcNSpwjDodWJTs94
tjM94rYFfc2D122gRzKVRZkDFpHyZiruaJ0+GOavC0SMCGEUA89i3qKxv4eECO01
gu3ItXjY46197DDgUrGDuqlWxvnOv8MPDCvWUWRy2KQ1FMbe5WKptzxKf3bicWca
SIz1UosIWICI6qKrcYEuAaFdJbF9yqellQJ2gO1SP8Ac1qxkQEPAhLN6/Kwaywft
bYXKldItAsJr/kJD/3/N4Sx+N1wzABp1NO0TUPIcnJTpc6EIWByX9mykzUVuhMvm
9yucWzOIEits3FDPG6d7J/tGCxzuR8RM/xe+Z8EGu1o7WG+PAxMPf9OgpuGkTbD7
BypiGHlBHu2AIUgyzSZ63ei/epI1E39lq39if1hqpIr0riKJ4mlIXB3GHpAHGE3i
m6wIMTgFdqFOmziYThvVWCbNFeFVTmN1NKsjEZO1t0E9pDO+qh/wP3teSvEUjzPs
CnlAUBOq60uXJTv8RQX9sQDjwuI6HkrRk2e5Cz4k1RH2Z/9bjne2UNJCtI80oCBU
2Rl9YfVyCPmhhHGuzFO23Ye0e2jqSCzReqSFtJN1zdRmyNd6eSOFSQRpO/I+4yGA
5mPRNM36HZVsmCPNHynuWn04XQpNv5b6SOentuPSQVg2DiBj7FSKdVWH/OG7QKLy
9yS8o6VFi4XBAdQEzQF0VJkClpe743HKIwOjv3aNMU81oe84tY+VD7PntgbQwhiJ
IQAXD0+EJzhff6AxGTuvQ1h+s01uL91OnFcnXHdRhn4yiGQV3P0zqvATNLBax1w5
+Z6OjNf0Y2meN1pK8wfdjpNPxWXHn3y6fd/2YxsusWc6kr5KP3ijbNzg1Z7dtvF2
gbbsGWbP4/TTZN63D7n0ctZs4FzquRy5NSrDF8xADJUoL5Pd0Ln6TK0vnl/DvQfM
yXxaGklINILiEhlVrhVRLQm8BrGXu0T+di/oZ1Gm3w0qAqXn0NcEXIVrXjegXhHn
XDWJag495gtmaLAfbQPTWsRtMPw+yVBoIVBRiZXM0YLQXtRTMbTCjaRKzVTQwkfD
BTmnF/329slGBgEvCzWr2LC+lsIyZcXAgSO52AdpTFGHISOng0dUWgaPK5+Pgwhg
gVAzhPOZczn4v25w0SZNHyX4qc5oy13iUCqfJahTDBE9FEgbpNs7lgBGSclzNl3f
J3HGI5nSOHvtRGqI4TbmL0CoFF6+azQto9/OxAjy9QH4UZt0ZyAifpaPppYXsyBv
3Dgww3988CF+s2dLGuKWONlrunIYmz38jvW6Vsj9DPHyerY70qKZGCwDLtnPMwGA
2G/tbupncaxlgZNs0D7oJ/7W45QFKOC+PQEdK1JLZGvV7a8dskQeE0aBgW8c1ER2
V1HkXUKNbpHqEfyeSUJV8Qrbt6ju9QLD8PxLmF7IK/wgUgzUsil/Kwy8aSuBTey+
td3F+rOAFfpPQghdSv6lLd0N7AqHKA37Qa+YRK34gq/c5A/Tmuo3swU/Xf7ydNUc
lTqq4IQ5seU0CHxeKX2G9jT7vtOKxxYE2KpusT/ayWhGf2dYNqLGg1O/7RzmPl9P
aVL+51N3b3deYcfZO7hcjx+k8wQ+MGPruH5O59HnedwbKLAUkzLCJsPCyFyU7qDZ
8nzS4osonkBn1/K3yF1rvgNyUNcuJ8fKqbjJ6nwXlO4GFUUTOWlGJI3w4ybk215I
m5w8v03Mvwmns9ggpKLmzQ36q8w+gg9KEG76/s0mU4VckB8diCcPwT2BIMfkqWzl
+wa4ttHn8o/EwVr5AwtpTHN3B4Ij4PVLkhq+lyG4kCAJMWLZ1qj6dt37K9pm+K9g
JwAZidQdvFW3+hYFrpolmYcLLbR2oAHXDxR+BxUv04thWWiDaZ0q8/vl+TeLepT4
zsxjsqqEhrbX0/gI7pOCvGV4Toms7ttWcNKIyO8XeH+yTD/Q2/rhoirgznQygyk0
gfPzxu2hTXN1+hwoGWheDIaxwTfTPILGBI/6XSVR+xhHFdHLawNBLNWcXTsdOJzz
YRiUW7N66OZlyIGKVXhl8k8Ct5aEqVJZquvnJVBQVIu0fuEa9RxfAmnAsR1f422P
FeFmyG21jNS/Jn8sQm/Y4xrXH9OYNEQiEQ3OjgG7ArTWpsHG8awZ5XSQ0YBro5/2
3h4g0LsJO5nJZBx3EaRy2zoOwvWhGLzGYplYFbQksmvHD/fEvqMYXrdWTA1X4jJ8
40eXzls1g2a6c1ykXdNKhtW5zSMc88slEhiDfGlDj3BANGHJl4MqLeFDVvsR8ekb
vVHWJl8ePDauPiOr6ZlAym44ZZfDCoaIIkpA7GhqtnId26oJ5AJ6dc5zlmsUopl3
4zLY1h/dHoynH/bBXSQCdawiw26n9PufBkS3QwwlcoIPy2BM4kZASETfqSzmixwE
VTrEyjCaZ81NCmbgGyXswOTNOhjPFXQq9eoj+NIjZD/4yhX8bzdY51CnQ2Fx9jpw
NA+FYT/cv5hCghMRUeciXAU6NreKOkpzhOJZqvW8Lid1LApZp9ikQnN4xtCJXiHW
8WidnC/2TzVxG02ZJhpn9yvbFwRpXS8hvAFfThSlB1b314xf0/1AaMza+2guzQDR
Q+exgfGS6AaI75aWVbL1rr9lkpL5iAVnJIB2xj11r5O7d6baqn+SP7ORl+xSZebW
KWeoOBgQbiCF6AUE8Q5eJJjjFO910pCwhbEGKfgumMDAZY0nFkd+PZBgr9XX8qrw
fInC94Qy/ive9Q7c5w+PyTSxQ7HL7Bnv0jdsag1sVQiwCc2orHVY9FEyeMYndELv
qYDYhRRGz/uuADOuGWIwjMrpqpUvpODQ7yNuHPcK85ag2mkTuoY7aVlI+aY4XfxY
LZNmaNziwgsBiDinY+jTpf0nEIDjXoFhPxgPVXFSHhG0ClOlF/Nq+oJZfLwBgezF
MI4RVEXL4SAHrVWEPqX2qE8CsHHxgWy95vPgbbwAxzEs0C05OMJuDPgByy/+CwoZ
9swsrSkBTrBM1uENSMhHFWUrl7lYa1a3UBxwCjKetoSUdsd3X5Aw/mvpdx0af8uN
VexNWt+I5A5xp1uMbi2dtTyNOQV/oPVu5BvLEE78a1qQlwwU9s1rqVdL2PRiIqNA
RkGNq8YJzRrkaCBTunwfYNRUjH3+74y+iIOb+kXwSwrqnVNvGGkP70ob9+yVisN1
RSQGa2ungyYFTGZjFPgrZz7eOa21VFbP/owa4Zl8FWJ49U3LwebBCI5JIl5xVl+O
OfuJHGrVCxiqj+zc19z7E9ryfcoH1ND90aC3Zv2j8kOyCTU2a+ecVFwiOS8ZYtCf
S9nXzLghlZ1MDrsWCztr2EpaCQUGnOV3d5iHRZrU6GvkpzuwQGPsIJfjAgq7tdlT
Fxga97jz+vPeTPdT/8Wv17N1znvgGNs9ZfUi0KK+l/pXAmFSQTVDF+AThTMO/Kd4
tMXtpCtCg0ekSttIV4+GDtGn2j+IwM7q/eF0HXwXDRAthGfYM+n5u1hMWEBZ97af
31Qw61FdafLT078inbwziSGcDU9niPLBS3cruzceIP9UGAS4Q+Ox2+QMk7N16MqD
S19zj4qaT26knaemG2ZiV2L32VJcUxV8+Bh7wM5x8P2q+OCIbQjEUugcgweAmyUk
evkd3/4JwuEuBe0yLgiQubtb+MTvgjE4LVoZxs1ktpd4fVBs5/f208FdQwvP4aT5
sNZ7cTlumS1FWYct1VT2PbaqezLPvtLTfP4sZnaSn4meadRkvMTrAzRzSH4bJckA
1cgj5/o6QBoVudoJNmYEVHVdVqFJVB9IPjGczsURJUronE7lUL5cA7GUvgl0qJ52
2hEZIls8zQ3Fw3FZ1wKAhLckMtIdT5XrFoDBMeJOTk+PTgUsTsAJgx5/E6aAR7O5
CrygPAnWO1qBEnYykUCoFSOkQb1SOdlpcoaJFE3vy40wCLiMRvAShSVAWdeboyar
nuUZPbvlUCfjc/sjHLdTppMB/sD79vAR1/1lajswO3ZXudWru/PE1QLoIAOQPrf3
RUtrBs77a56Y3vVAvrjxtWXhbSG1eQpMr6YqGUF2yUHBh1Bz23q4S0gpv4hjuIRK
eGVBMtG9ndBb3EfQvYNY4Buo4YXyC+G7UGObqOX4ilQlHyFO7uDVsEJdx43RFr45
1CiITF5QNOh4weYWq/3YusK0oewAfjCZiBye45O54ZTKXpMDAr0W1FlyI3aa1XSn
ZoQwIl5pi/JnsVhbeATpG6zPfk7fp+4PeqwJEdp0E9hcxeR+92jU7qMmCDBJxwwa
CxAOOjogdj+nChDLC0y4jSjUL6veikbtaOuc45PJjHJRH2KjEYIDsLP6jJqmDcsJ
UWoI1MXu//F3ElUmcfgFxpZYeLj/Ossg/NmYF0L/x/oqNZyeF80hx5OZlFosF3lQ
aOQezPbcQRwJs3+JQAAbHnC8yZq/BdaiiGbHoRTD2f/SX1G1sKN8cOYV3Ikgp/VB
svitumU81OdiSGBFYiknsjru3GJhDUHAnrb+Jo/aJBLEyKeETSqqdwkhHZBrZtQ2
lLBgs/if04xdsD9h0Sd9hQ4ec09imoeE1pzW2aNwfQFhpzSi5EwdQAWjwoVUj8RE
GQIUNk9ktFuYNX7O48eej/Vy5akqDUVQHEGYta0SX2keDapeMXH4If0Yj3KM+/ub
IdonctJ2ThDqkzpMyHO23fd9pJoGKxmDzcnwxPB/pbOXmtFsCZgc3SVDDJ+pdF6W
1crFxF12+ZmSyDTpfJXCTeTWQEkVecRz7WYlfAImDILySFYE8xyIyxlz+Duud9Je
WeJxn9SXgQDHpjZrjzKm3x2nWvrQ12oOOxohYCVOJSRJePaTX2FXuIz1kIspYEZ5
KQ5fHeLwGt6woOqHYsbsrgDQ1GlEGsQtNwZqNNmgInxcTA1XYccw9jEnEUtBupBL
b5OWfDcPUpX33OmMxNwmS5KtGrn1WBnjvGyuiu1pdKQWBkcBIvPX5pYtvE3yomTA
EJcxlJxRY6TyLDlQyG4g8VE8GOqhPNPsTSl7brpN7UWlETp9J0wU/7Ed8ZNF4eVI
DBMTHtN+HYV5/9zd6aB5YrWcWIAps1oCmFDkEnvbHneg5G+aanXBqiOOVhFuMD6R
88EaU4GAdI3du+JkH1Ja8tiE+1sUBrpOao4vAS5gPry0vkIHOQ9Tfe1PdrADNcYA
7XA8AA1kONgjxZbPgtxBZUGGDoYtYI1kjk3H8tFYmCZ/Qsx0Ijf4cMYZevxmN3Qm
zRo3PGQBNWmy78WHkJWHbYBFqLNwargr5PFg578XINvdDvU3YFUxZlzWwrjoSuKZ
zuuVo4sB4IqybggeMM3plZB4+ald9+h95G7Ble1hkNKE7hHc166BAhUAVtgwlu3k
DB+w6Yl5QKR4aN9yprLIMo28outQqlCzuee7CgLds9U3uKZ3EWZO7N9vW8ashOtc
dLGJuit/roMgzbmy8/gtLuwZHaxAkzOzrjNxSItyfR1iAqqca1sbbMADr5sP0Nsk
BhOxkt3iGpYlMNDybubhGr7olvodUMlG2I2YLpW5ZH/+uo+B8E710M8uUb4w7/3w
WC5Xwal1LXWXKs/x/yZkyRVB+48Sw1pOQtFfskZ/lzQvI3r0rxCavlFlveqhskVG
5wDgbkjhS1ZDwc72aX94GYYHkzkfcfjmVp9iWmDKTD86SqJYgG04dG0L6xpIpOlX
kdBfzwUV8VyN75fmpVZtoRI5ec62X55KXKA58zM2nMFu9oltQvVAyMG+kXnfKctI
jkTC8I0BdyKsYG8RH1fdIqDo4HQiErqqeoWMpqPhvpDS9xBxmsrrmYalTSv/FUCS
+a85HGRX0G4vyQPRyBO/MRdZAtLCoO/rGRxmNpVhTEpcOUyWELiy1Yx34dj5Abh5
dDNHtrELh3HtYphDslzeVS/cWiP9lN2Mgfb5NhDUP8YhL2En3VB6szx/XawkCzvQ
ggqkXgKlW5EzKlO1EUkIZzLmrwBcMkDA9pXmAV9ZJ4yLkWqZ5BW7jjRkVFJctO+y
+jhqbdFvAatSKV/jKO8yxFG3F8lg1kNGIyDnkZLoxWTs74iPoNCrexJLh7cvrg9w
GpmntspUeyP5qOubOjOi0T/0KB8cLTyFlRwoxzNxNKY1AIHYCgS335FsAg6CUCqU
BPbJw4umDdVLkXFgGJ2x4hPev+BN2EUxy9H3M1nCXebqOjNPpK65Jg7HFcNHE63y
RHZ1p+sIyX56acErG5nGd1M9rup7sh42wl46zqv/9GD6lGL5zq7naW7MzFZyK10+
+eB1pnGqvu2RTXj8qu9IDfZRUCBFMedcv09ach1wFs0gQxFMLpIADwei/Jch8y20
F2PCubUezuIwbR5Xcx8RTXqSnEDJobm985MO9U2/oTpriQn/jTi7w2j3LYBDjt9L
3c1Q06AH+M/YzifONUqP4G2fs0kKz+kDtNG3vjgWCo8HhVhus1SW5a59YpNuAqrM
OwUXf/E+2BYfeKZEXO+aeOyd3iKZg/KifjdLnCUoVk24KZumMaKPw6E0BldMGFzY
UWGxSnAuLjxRLC2rdwwZxKs71myaME2OMJ7od5msh/0iO8xO9tUFYBGoOfJb/r8w
hn6vsOj5i4eIhkHLcrnAnXgrbGsf8k/IvZI522Pbk7qSs3IIOmjxTwTJ4pAHvAP4
piiXgUcQv9pKMNp2WXeE9uIFhn/tLkVHFLEyGJNIoJMHmsKR8x+wm9NJqjT6TBZH
fgc15kkjsP4/KjjU5g3R5yRhB+q59kVdy6FBPQveAKpeLC9Cndy8RbckcsjchkZf
9yx83Yv7Gg/kIXjp0IjVTebUaGPebRt+PlHM7VVQd0Sc6TuIh7Q55OyGUmYodMMU
6LLRP91/vyyCvY/30N7EP0hOaf25JlhSzrnt/friVWGZHUbt04Dbq4/KAGPnjBsk
IhTdatBXK1FaoKApP76pCzAYiMsWBU5cdzlXMzdRSVUs1q3h1/9Z2fldqh6VVBba
lQvYlGob4wqm1TftN5WH0yhb9/MvTDxdp5oxZnEHP8Xm2xga9b33x1VwgmJfq2w6
4oTH4s5UDJmxOVvM+vTv5tZRBpWSE09VbExGF8NRhpBgahhCTdh7m9OgcfmsAmbO
DJe9RramKpOlze00OgRA8vSiwWVhISrIrg+04tuJgs46ve/un4DwkWQaX5V3vWrC
v5kElJn/yx/vIuVbrmC2AR1jDRrUNwOfijBCRahtUK7IRzrzEpUQDy4W3W0AsvA8
mrhwls6kIie5JKFHvdpcl1W8Ek4sf4qmxRDPliJob/gq8BZ/ZhJ8G+1mfOW64gVS
hlnIyahSIVO0bPFBCufwglXBSgEsIouHlom926Q+s6pItJWE9zQA+9OPCOzPkjCS
w2I8VLWmM0nnAGfQLb1X52G8xIZm3rjaZaYdapxKOm/kCu2mhIU1GL2NE0ujLVzh
Bd7O4Jm9L9qklIS4gYauUBEeR4RRUF8MoqQaWL90vflREgBbKzYQ9mY5oTG+RH6V
aDaKimj1u90PZ5xiYDW7dT683SnXfrOaaOO+w2juWn2LaPG91NEguT3YZHrGzZDa
Fd5tRyzTQMybhNFbaXNEx/6k4WFPmecZZT5w4lMxdCnQtKJavWMvJ9n7ThNGANKj
jiuGn81SYFAxkYaGm1h4Gdy8u1dhsykjTJJOmaYMIqH8p69i+EOnBc9EPe3rTlcO
g0M1cwnwWUkUncRRHsLTWKmv2K7R4sgXcG4ihZrAq0CIuPW7htCV7UF333Qv7c+1
InMbZ0TnrYF/g0HsnsU9sSnl6HFwx/Y2FXbMANAYNZ4uWTQzxbWCdhKPhWv3ricK
4ngJU9W3QTD3ZFWyTCFL2R99gnD8j5mxOz4AxE6+h2aZ1DE364xowMzBjBBcAgZH
nb7aMmu7zUMPDzq1vZoTdC10fKMUtQQjEThb5MTugJ3LM+OzSz0QhU9C1djuBRFF
JNOaZGoVh14WwIs0xm2EXQ58mdG+xMthXDbaZln4u/YLQjO0kxsmq9x7L/pKBDRK
u1CCRq39FayvpdakqOoy6wCa+FwkS7wh1enr0nhsWwilA17MvCMr6LC09aEN5PYh
l1xJmfhKllCeY0o4l4Rw7z/asxU7WQYZjJZDi8m0vR+kBC2hovA/zuMV1IP9OEi0
uEf+3Ba8kso1D8nakn8n0yJ1PVvfbnxpPNOcqJziu39Cnk1OwWj8Rrwn2R6tJH/2
cHZ7erEb2SWZm0O5FTub0jmnzgAhBFIUPKSjZGDRNK9L9rnRXfglO4I4SPNx1LUX
xOYFDkjtd3YaZoQNX4yfmF1gHgYkcweesUak9+CWoSrI4mH/hyX+zP3+KAaxX7uw
dTjrQkXoqgsAW/cE3d2KygoPoaJD7KlH0y7/u0JijPdCBQf7DooMFBQtBK0LTU57
K/J5FIpmYKYzzQik2kkpLR2Ja/oEn1vJPW16YVoBLkbZl0eAfziP9zqrpZ4+3ACL
NTzlCbqnldbw3Uy9ehCoRR3IX9FHhnrl6+Jl9A2ALkVDEMd7fS3Dn/r1O2icp47R
xw6Q1ewneQK9/XAp332s1OtRIbW4CKMA5xSlNMKOM8kZ2HuIqBpeiaEgF3ulkTYP
P3xbp4G9b2RGim4szj9pMQakKdJV+wWh0CRJWiHSeiLNvyzsS7zebjstRNoaMiHC
ExFlyUgrwYCG91rnB6pT2TKD/t5P/ohWY0kUB5MLyVTL6TQsGtNQ4QQb78wEvDnl
pvq8yxq6EeFuyXEGQ8sT7DCo09zkt/vKqcAx736kFbGW9tDrJ5CY79EpVwf31umB
6ey2WsWgMv08S3IcwMPPB3xi+/EWYhH7irWJd+h7QrgDBQI1HaBXaVidwpUcZzb2
bDOhknw1jZpkbHp6kUNfkh+8NJ+juJfRdkEMi+57sgv9A0KD8WW5/WzUkQm0MDQN
fbGoWx4yNbdOoY6zknMul1/glXpbu/65tplvJBHzECHNrHhuDzEPwDs6V0BC1A6x
cm0UxYe/5qZ8KtypibWt1gVjVzhbLmy1N+wWo0TbNVn20M/2x7/ojJvxwhfhJ+HA
GhESqWGtxYDJbPf35/m3mVOCPLMOuIiB8bqAQmq8oKa6rdtOYas1qWJL9yICCUD0
QJUAkEimfVHeysKg770f4XEYt2+aZ5L+YAy/YVNJ0tTTL9UBlrLSgrwdMe5zrM4T
NNq3c6iT2S9WdQwT5129BPnFWTyipe+bxJw/C7dTQGzONkeqkwRa8pPon0C+17Ck
HmRa2MUc4lmWTXVaCo2tqwg5TQbpzyvftHDyMudj3Elr55hPWNbDmizyZ1vIfFH7
AQZA1O4wqg2uEzljqH1xVzU73W01RsyMsXSBoC0nh+NcHfoA5LRRrS83b6/JnrGF
LSiPNOSn3oNCiUVhwy3ukU99lmFBYIoksfcx1QiyWWizupex/oOHrVbpKdPYOd6J
sE+/DqT2a/xbPPH69LYIutPjPADKt/Or8IM3MqC8q7VZ7cOhCxFr52px8aI/znPd
BwmLiDCCZcGgnDrzPr5BzH910M4CBvuriN+4FB3+AXl5Zrb7gRS67JdNr9xfXiRz
OKgnRGJ547pGSg/GbRmMRgYO4fnRpgHYz0V4ZzFh63HoWEgSl8ocBh9QADgWvaQp
RQdresjQZg6TrBriGfjhSzVklizdSx/5WfYW1sMaVDsAPSnHvURHoUmhSwKf3RGa
MVUmJk2hDc6R+k5+Zirf8rS65nQGoNxGCoaRab10dD7wp6RPnra6wrKFPAD3WFVM
OGPnZDogOTmWRyHtK1ajfoeo+dCcj4jdKp8a4RIYMyJUNhdkbIoiDkbcdUfbfdTx
IdZbJKiA6HUm973hdd9+Wm6UEa0OzXXHoZ9aVeTpyVXzPC8f4dZ/+Bg9Q4+4uAz9
eDWNc64KqFTTxn23R5fSbbLhCaUOHYJ2ytFE5yXMWKXtvdFUKL8rsORzZKk9+hfL
2EHYD/yKr2WBFPvamsFWIx12OG3pmuVG96MN0RHW1yNo0wxVWyugc6wtHUW6Xmb6
5SLFAxc1cJSAkKhzsb6zUrwA9qLWwmdQHRjVCJpQed50DZeik3QB/7n31xNPyRqE
YHQUcg87zORZUaz8wDzV2r8u20dUB3aRxoM/Kk5ahDCAJFy2mVvzKGffeD3qxx+t
6WN7GKGMMF5KxwVOzb//Q6gDEyZVnNMF1qGx6s40fWhOg/mcfFfBFzvmhdsvv/Uf
HJKx1UrgfFSB2vzYhD3B0Hn5irqQ8Ks1yc/tV/DtFarQrKSp1BzGjr5Q3zUlD94b
+wbqk/zpFpIYFTULPos8celBT0tNBmf/a06jX99vYrllBWqGJRix2AFufNaPlRUW
ZBZRjSwqekm82UYRreRBY09LjtuWyfbIClNSeyOG66xyx366yq4uZC1dqWEa+NNx
qhbz6hMkT2O9eiVVEa4yW8Z8sL8P/7VaPfje5AZJo9fsUVDba7oc8omranDu61Mc
ahZwyGotxC7K05O0JHRce6IaRfPe06Nrgr08DTLIZ43FAR9GinwOVjDTypg2viGE
GptII28cuo+56qKySwR5fOOrIUpXi7P86IdOqe2hF3UOr0groTZiNTx8bss1wpG9
y/dMZq/ehM4cNSGyDxYGHA1P88nYtoahm/WnDyv1RfvnrFreCBgb1yuXDP6qCpk+
CsuiIk1FI0Su2J96BM9hatfyjNDVu2po8DI3fnJvt71gFSybyDbAc8ZlbFMVSdy8
N4ZwdhXLzAnpdfN6IF44yS8o4qC72MwskVRSZYYNX2cnVkUoQFgUJHPwJdNGvUGC
91YTH6XJ/NG68EyH36qyGxAADpkj+5/M0TiS4yJ0R10ACZboBM27Ypk9muJSszcO
ctpRi73tXr01hSHTjiI9MIadyX7ALKgorBBZ7i36hPhBsbyyAGCHZOOhvZrdJGzf
jOqnAAUggtgM45GGLTADFf/rKwpgHdQGEsEbciOxy4i+yXNHuoS1K5uIul37b1r1
b4mkSJC/wZ6jlQUOqICFmEg4QaWRF+hBM8KKVgDJsbRv9/wGZeh66K28F2c2a6c7
P3qKkJgBU6He9ShGpFxx23bKke8+3db6+5wgMs/NNlyjQsFTQnid6re0IFD8vtxy
22Vx/OINpk7CjWMt8/hszuT/Bpj2oEEtAeBfaDwGzp1DNDoeZ8P7yoCOhiyFRNpJ
ELpXqmEWm/xrW7QHNMwUko1rSY2lg30j1iZX7tYHnMcgLmFNn9mcUf8wpTTXtkpe
G92OlwuWQNoRNROvOjFuGzXxOrLfGUFmD1KZRIlwtowPS11Ybm/ZOJ3tqbmRdE4Z
wOU9S60N6jM0chZ5Ju8tmrnZmhs/JQNpBi8jrDpwrnlz7Ev5Zla2kC1oSxB1yocg
4QfFVRrA9yBtbUYeVVfFABLLRonwjj6u4gMYAm8M1eDvliKmFzZbVUYVwLFEyCJq
cwHKs0LDOzHFLxfNsWACjBIH3pdwHnNM8UcY/qZIy+EUYOXmqgd+VT2BfHOAcdh0
BDIPCbgtF7rU9gYszRllB5KmY9HpWNVXdgvWkhF4CwGJgfYBZZnv/g9mRwMy/aU+
gTtQ+7ZxvlLUOXqLgfGziFT0rsdCLkb5SdYfrgMZXY+wShjBxPGCj/tWTifR6zxf
Wo+wZ43kY10tn+pI2RmLjHAysJxghFhwEygioTi4NrgUod1fqjw6GJ9jBt5hFmav
ehgEnP5a/sZFozdZfn1oSatH8RkmYqTi+AEQdOVMnn7s4NZuokdDxzePcBEobj/s
QLRqighXYytuTlv9/Ge2D7UCbqI0jAtpSYMO41mHNJ4eD1iYGFoVUS5hUpcfeshK
yTLEPxEFL1O7uqQYq30ZbsjHm82pJ5TwPtk5ThAaOX1lam4DHGxC34NQX1RV3Aph
CqssldwOWeI3qaaWEvIKy/lQoT0GEiWO3lTqn+a0IoxDHiRPapRwfOqLcIl/irgJ
1A+YizJYuTTjWwTnYJkRhnaMJTFv/LbQtJaGTcoKhJ4X0vZQTI54xIGbQy1q8sBP
lNW++RE1WAoNZqB1vA9i81DOjyqIi68g8kOtmhSQ8x9P2d9syGrhWQhpRVIICtmP
VGAi+aXs83EITqFqnwAJzaXiMVjCzeeqjRHt9+4aB9NTM4tfPrcCocv08hbQD/D0
hrc9uNiCTCUsyghdcExXbH8IW3sSjGBmmZmVIpmzaAVrmoUEQNJmrII67F3h5buL
H1XdkDpBkOHQXU+wUQ3Goo7XkAPSiNWFD7ptmCLNrIfDxqoBoAoZ7qsoH+JaVZI/
XwgIimZvkUDcH0rl7qJe1aAgsZaayu2CbbAnJNn6ZfvqfWecI5RSN2DSCJ95xiJr
9fS6zRBsBrHYSyQOORpQzEPySML50d20cz8YhnYBXAbhMO1nF6qmhbWfyXTcWYis
LLlBm93Tm0OGvw9VBspMlTHFSZO/NHay/mEsbCLGtsN9yGZefVnMDnzcjljcwPf2
JMP6l0jPTKUS0WRyiWWn4r+UGlI1m/leVBddbIWzUDIsUgGxyTos9++nF6b7D4cX
RkTplVkndHqgjjUjZfHcaZtas+VvisNCg1nhNafLq+EbNWYB2q4Yf+MqLvlxu5gs
kph6F77JpAnlGFsL2JeFi8sywUohFWzKnVf4pUrRjP4mlG2HcnU5ke4XvRx/ZSqR
pdR6hoLMXY8pAZy6+zrLiDAJsszear7EIWa+bDDER9KwPy1ZOQgRB75Vq8z/M5I3
gM7YAPUfNoOOROWqn5oyI836w/60WDKKIYC18+ISw1CsB+tGwfay+d7gVhtZTOLK
beqFnkb8Zzv43tEsvSwRrE3kyDzbq+0B9bVp29wWdNtMD1lUK3cleu/c6s8cfmem
r6G8jY5B0kv+O/cIlqIORo7Nipb0l2ZooMtL5X7u/ExS6mhnPHzQWVlC66gJVgag
mSxjxz/JjP9FI6xKazI/QuYwbCDircan+15xFVwuxj39sdITuaTroKE526KC0oSl
UEvHh0DjT6YPIDKtSQBZHQfARThYNhDRVG1YHg/h0oNsez9cPrkgEmj8xuNtZFV1
bzPJRTIUfnB+RN2K7+nDQXweN4u2HB8h8e+CFMwywBXQ8sqJGo4Nls14MTZwdHpU
0fn1BtPoK5txwGSdpNfK5iEU65A814xLXae72zBNMZ700WV5aFzXm3AwqpawdFa2
+Dcp5OSCpRkbNWdTnUn6dPMtXwfazMkm2lbislfFxsO3YTuJOAivt0DHjcIx9KPM
DnsLw3xzykMEUaMj3opTulsSuVaCnCJX9GiL1egrwJU5c2xpz57VJere9KiRrsxa
HXMrTs6F2dFDRbUuNlzJuFFFfBQ3NjnnssV+ZWofJfgVjGg4CMjTILBCCxWDt4lo
zBRbXOmwdN3jetSN7kvrB9KhwX3QPn1BNom1p5Ozp6mDTTbhHx/InwhNs6PwMbWT
VqqdUlaDj/LOGd86TCntxyKM2aAWnp3SEBTlA6AkU3ZoBrOK5IBP2aOyF3xhNdR1
QBZ/RF768jwrLXF6wdSSRuG++zzvT9xrvKbedNJG4e+ePWgG/IrgVAO46IGb2ARN
t7JQU1TIUb1uLDoaolFdszY/dPKSfspiOz0WZkGtLotgUWSFNNy4Ax0L6RKtmZTE
w0S0orF36P5CJnctI0BxOwgTeRPimCn9j+CGvDYe+fLPourlVtxXD80b4XNsxD3t
NJmNsay8GZqyGJFayVy3hvzOFF1+qwY1p6JsHN+uAYck1RmeD1QQXCeNtZKGHB5z
yKsNnnTVuRvkKSnYcS37QMlKUkKF2l8GvWuDcTGv042EWef5upXJQK0z+wvasI9t
kCbxUt7nC9bCX922zyQR+be9GqbnjDg+UBLi6MAjZwqrhgs3x1YwRgYM85EoeqZ4
8TBEgu50tMDX57Y/Tno1RJwIS4lb00RXEaIx3+1yXM2hRoFdyn/F8LeFLM5Tu477
x5UxR2/CECan0NpiArFwHGraz0GF4+vRBCzqxTs1XjsjqSoceIh3FIwDTJpDbiVH
LUThBn1zpO0oxX6BNhYk9YCtvg5F+y3sCIFdBGyIUZuCHOMOfE78vVXm1Po9+k4T
DUXrmaSZb5SIWSjmmt2UliX75OP0uwTScYIiRlUZT0JZyFiDQ9doV8Wc7dEQg6R7
7sVDNCGtsaveV7tZimy37s4NaHNzfjMrG2JYqMNHO1mbSHNp4p9+8Pi/y3y49SVU
rroqDoL7MT2pa/nNYtRJHBwfWFCx1Awxp25QohQaHdYZQEEhdpljeQSHAk0FJe40
BaFiYzegkLuILx3kBj0o+J4ccc1PijrTBiASmpVUnM633U40r/dObZKBbsxVqSA+
yq94csN9LvW0VJ4CJRzs/WxaDZ5iorqeX18VrREbcJ/80ZQvjrYEmkmIOI+B1eM3
l9GN9PA1/mZYxze+/EYRDXbmyUzlYqmztL4qoa7oftbpzT+gzcfSLrhA1YhqZpgh
KW2Nv2r4UvHuGWBq5FougBuMxmIwFuUpSGuQa7CL91U+ev5C+qJBqTzzH4hU86up
gqEpQHMVl7SW+1wq3AEK5VVpXSH8zfmeIVoZ67vNc7n5gXHNNh6uTij3qdECJWDE
N3TjimtU/ru56NrhvcltU5iv8RdydWig1XSuuzLaWFACc2x3MIN92lt8lXvwHJN+
x8wf1U180AhtmhR57ND9ySdV1G2rWAalZvNGT27+AiovmuuNDnlHyeamVeZSrfRf
XkmAaT/b14mokwDO+x4AOzRaYd+kGNMnRlTG4YJIalFQeE58s5wdUAlFi1Vx6bIs
QjQjVa6loNsEl0QNcdEKsfySQ+Q+HnaMC3ptJVM966KmOW3P3hDbpLICGjyzU2Si
60p6JrEGwgSWv4oGZJeFXfdzgnIx5ckZ6bQVww9ghjU29nLc0Lz+08KzAF8cyrBG
no7VvPIrHC3wG5Z/alWFFq3TTiOihope310zVKyF27fV6hS5eQ9w6VCL/rxvVCqh
UP+/9z8PyH/VftQCj2LFwWS4P70cTo+ISbZzyxrJVrl23iIaST2Yt2gFwYSL+vTU
b3ibtrTHxl9ImyKYx4O14fBojms7ecgtfebXHGA5TTv76VneiaBYnjpFAooHHgik
lxN98756adA+gKrrPypuUzPcIlNncUySGFK4tLFPtnPS6BB4avbHvf5IWfWT85l/
7xYXaw51icj5r3rswX6uHWzCxPS2kJ5VffBdilItMVt4VMWioIFvt0k/A8JwXXGJ
j2oM/dvdm7Pd4QNpiu88kOcVanGfzYcQvdJ6YtIXpfKTrhgaQO7LP6l9d7qUmay9
qI1CKZla6OHvSvSq6g1l31v6UQ6IImVBkRdfOQ4X33FOIGYkNCQh6uSlGnCKsPwu
Q6kqbri7+Xr64heoZ0eNpiqP/OQgbiV/7yjES++hEv8bPEo+ROO+Vzhumzveg4I+
Lg8FZdGF9FuMxbX/40SJwTRXsR+08F7Qs7DbI3rMRtN0bpdoONXdIGjQE79GgF+0
8N9fggXD0koHXGns7Rn1OGrlrjjZIiPGEBXn4zhqxhEjxCpt6MgcBiJUZ0KfRoNG
5ZSRdMpVYPrx+dB4jh2QHsSMuBq2APN1Bm1srAn3pC8YVWPOsaVxRnDHtqc61VuW
Do/40OTxkYP2Rxt5R2VICkg2aRW6wTlDIjkyzuho6bxZSYsZk2sy+Hp+4ZFKzKyi
UvB7bciYcpMotYig1Wc/0l6aq/8suG1cMSEtiGzpaJKfBC4aPSTvtql+yFBK6ujx
nk8mGeGoGzOxfQS+oIsmn1Ij3bmJdc34JAlZCKOsnOql5pwy0y3kHPXCepYh2vTY
8b7M+ETmvNbcSQWEpEvOjggwdd2Adh8awYSXEx5rYvDr6nMd3CKgmiIdeOjC2h3T
7pLD4FHeTZe1fhVW/YvQT/a5jnEqOrKSBg+EsPnCdsDCYgWqxPthS/F2gWOqNRTT
L+2lA1Fj3cOSLG2r07U98iv871rIfZKjEFBi7EOC4IjLOpa+uY/1sL8zZQs+rU3F
ckiiqNW/o3PjuYjehDyK3qPg8rIFATfNPR3Iqs1ONUSHR5/KJ8ilXWoTrwCLkI/E
63+X5a7WQPralpN+uq4HQgiUSZGTkI4lHiHTY0XlfnSLgSk68Nu4uAtefz1nNTk8
WVZk7EPSBfH+veOs51DX72K5pMUCu7f7M8ZSyXKKqTHSuZgTsEj80VXIFHxfhcNF
Pzj1rdZywn0gDDwyQiYuhcMS+4D2LVlCsFFZBXAHM23vZ80dSspnKW1ynyXS9an+
OcWKeCc1XRvizo11AaCb5ATl6Kel6ie68v8UkXF9hREu9sMZH2E1aV+EswzOfgSf
03UqaZcxCy18QfwoJK1BzU+geQPmtDyJ4Ti+/dVZ09ZLmloXJJUF+U8/widbf3XW
c13Ly7qv4PkabQDWeZiaq2hHTss/ZJPUkgILhb8PhdaQ9enMFCuV3AEXOuk1kiTS
S4IgYgufItgifzk/mzieAT5enxO/cbHvBbYN2J9Oye62ob/HTjD/doCTj8azTm7J
9NMeywO834IJF4IP+jNIM3cFO+8MmpA0aTihGgQZ/hFszQ/qg8HWWwdSF2xJgBNK
BiOD/z9sQIXmAsh9JiphwADzJFgvOmuHcT7Bd2TzKPwSySQ9Uke3ukD4aVX+wv0I
V4WH5FXVFzcM9q1u2ypYl4csXPc+ZBThGQri3b1e0zdbE3lVHBA2puc0KXa4Dea+
usRmFN4mjYBktHp1nb3vOe3SzBAE+W1E3pm8pARnGDHaz9EeFgXhB/UjADeeV69w
vjgscoPhWUQCwEY9xznlcClB6wxKZbmccLnvGPGO9A8Io+L5RBbGGqdzQXwEZfm7
QOdASbA4EkPXDsaRitc/nIkD3rR395qIl/OGsNRtaA4Dx+z4PrDPqO4vyFVkFYa6
cN0/ZaPDgLJqT11kCAhtshnNo/kGN0snK76Rp2/RHkropu2WOJb8vinxT1GiFUWJ
Y5KEGbQRA6OIqXKoRSO6oMs992zt4QJ858o19HCG5yKyrEW2//Ivu9xrEtUgEBMi
b6QEuFV3S4F1toDzx9Ie2sE1JEErfdPeqwdu6pe5BSIZ1aG6yHvwjdbrngsE5NC/
mBBzeUIqEu13Ze/64Z2WBD0kliNjnWOu3UOOVV+7iMAblUl6hd7Qev7mXn5kfOb4
sbusViqPym/rN6miRPJTXf7NnzE3QfP/e6F9S3kiXK8aveo+FnTu1shV0im+WMLp
wjIxxuoEs85BkVs08B6yUtxVptxZCJpdTIWc/GM34X9WQXOcSCL//NwzOGT9qevP
O1S1ijz43qwY5fUQdbSEwp5QYjE1YfR4hBuN1+TVgVqXOGvYPssLZv+jyLZT5YoY
52wYRCg65uXNFNgJf6tUVvjrVNEXG7t6su/H2nVdyUHHZtqNkkXAnGOhdi0/SM9H
0MC4btSzTlgWp+pVivxeZoNocqvO+Ce+vctV0qZa3INy3twROjLPmYucLLUE/0dJ
EXWAypH2vxtseCjYgqe0DD6STGouKtQUzG/uHT4PJoABHIY/Sb9X4Hpe7VbIU+SA
3oNnRJGs+8jEcC3j29AsfMhtUL5Sffc1lWUtzARBokoPFmg4TmLyNDZF6Ympse1M
9tvbgTTF+vNo7v1vwFiuPV/GpuoT0ToOXWuJ3IWsenQ72dnMl6/PvBpM3HTwkwoi
liL8HyrVhK47bAgz8U7cJ5WMGybhDE6MVqWpTnG6wdpD1c7oh8GBChQQF06MGISo
53jblatbiQGJrXpvoremqaJxJ/HN1B2VAZ602vWeS3a5MJN1Wr+pDUG+lM/+27J6
eQlIlJLjNfiSZoo9bTN/mPEisSgYDD9Scu/6psUeXg/GuWWD1M5jBxEC1Myu7vaG
wPMbejYy96bUxSGRDfQD8RRI/FaMurmrbtJ5ZV+fyVEcqP7CB5EZPhoZTOMv6w5V
JuEKYvVKqZNVY2uezc2aHdNuaZom0k6x+Wvi6ASzPOGCidzPR3vAL7Eaf+b9oKf/
XPj5jvhmiOtVja/LmHhOgECcSCng8U3sX8f1ci3aEyDM7BapTwYvXpzu60OjJzxG
dmcfpngG8laQNiwmOEIvnzc8jE5/pwoItcoAzAbp5UFB+Qk+fLSCcaw4cC9Tp62I
U/YCTONvPLddrtSUT2BLz6mJhbVgHmSyigD0+LTPhPSHaeQ2YlW4ZHlcyeAhTGhB
R6VMd9BE5u2TabsH/P4TrdvBZQO7Ajq/MLB3eVeXAIr77MfaJBNMf1jMGsSmSkjE
98/8NuqtuducmNJPUY/meThMqbkPrdWXWluKnIl7jlACgCy3uT15BWzgnWhuOTEh
u7O0S2Rw50x4VAJAm+4Uo7IFUBatxqVbGLJv9Ae5Qk/Jx+YfiRUblTrgER77+e90
bv8iPKSuM0BwbsCdMbMqoJ3XwX/0Vz8NEspBjBUtprQrtXrug/ABzsRv5TzihReX
P+kzet/WXF9sSzn//BAddb2Xsd/NebFu/sVK37ZZW9jlb1RcWzYpa264T+SxcF2P
V6Zgbh7UClXhe4jDfgrXAvRWjJv2SblHz6WUA+aJPPTJOTTbhuvCe7NjZS0BilcQ
vWOBLNaMf4e5A2mSgsYwcpywfaV9nFUQVG+U4XV6L81MQ8kcq8b+oIgR/hzhPH6O
kL/ENdIzw1HSUExFXmGcaTUmdc8VSJaG6bNRUcswOCshbGbasIrR8HmdXy4Qlnf3
PWSHGZw0taTfwEndIvu5v2cbhZbpSz7b8ZWfhF+08lBseKz/Zvm8UF5YZxK+p/bf
Ax2J21+V2xi/TcP2Got7kVjQHwXKao6Y4wTaZqYiEyj3a+9O8ruTtTZqLFezVPHl
Zy5WO+y4IjuB1gpCjW1kPwLhMW8CABEjRvvzu1LP8PIoC9k+00s1k/X1zwa52Vwa
wXS5l/e1haDObh0SUMxEYazLNiw+h4GYBpAqmBUOTOXip/VJhR3ouE9Yzq2t0PVe
HtH4pHN78eMHSU92i9jOrlyO7SXcJtxGqDKx5X4BReP3kuMj2AShxclxKvb7MSAV
qsR0SLFG/19JvAuVHQW3S/2UXoFwAO9pW5mhp/FjiWY5Zb0MZ9B1A3x41iV5kpaG
LK31rKtQrsHYfqjFJetOZX2h3nPe1MbDRp7vgVggo1M2LFLdKUs8Kw0QZ/mV+Kf+
Ql/dASIzhjBwI1EywH1yrcO7P5sIQoPZZZpNk96i0v6q/G2XRGMiF/19Pzw72EKB
LqvhJjf5/P14LhXHmhFg4uR9IJ6TnnXxdq9Bj7tEeeonMqrYmV0xFsxUQB6vYAty
neBPH7N5zKjdkwTUNi6mOdcUSlWVohA9sc7FxNIdtyWF1Yrl6GrsJ1xTGA4bj0LK
GBIY5VwcrTzpn3EyNu0g9Pa3f96srfyywwTPAnfkUJEtsU3xGSK5FjsWTYJuwraI
2HA0GrAx5cIS/2CB5Mjayh3pvtFJHap9QV+ceccU8cMoMwQjL36WdRQX0keilKbc
zrKdzHFCP47J13evw5Bi2Wp6yvtGd+57ZesehK8PBheZKny3UGrl3LdfTd7ox7a/
NgmZ/OFjAHE3jxb5vkh0Z29TcU7LAztJu5b8gUKjhJ7m5JTNOJ7SIqdHPJptFVct
pjNt9PgRMYoi5fJRubRrKe8DqWdns65C1MwvhpAyHfZs/o6JvGJXAjyF0MxF6d2Y
Z0kcTjgiBQp/9BCtOSPIe4uYX78RGZjBsS7I45jz/L3dDQg/SRSC8P9Q7PLF9zUx
QDnt25aB7t7ZiXabgLuFkdLUskBAF/AVvWeWSHfvy58phWgqxtJX4Q/F9XkoJFVT
EOlv+YwJe7uvl+qcPZQ0gfMWd1POEq2qXwyziC2mUDBTc//0HKM8xINeM8JSXYb7
86W7pR1oyk2BRI/kxsEtkzXmQcnry/dKI5oAhlsnBsRYlmAJgT0yHFRVgI4YwNV6
oXLLQENNpKZYrDHkht5c850rhCiqRdWrPwTMoTdRhJVR+iYUtcwOQY4ih4s5QuQ0
SlyI6DGDrorDyFsgaw3ED5rDLS8FIAtC3ct2u7cuG3xaaRYeqilTi4WYFIHIqnsF
gPel86Ss3HYY3Kc8f8XC4v8gHChZcr/EP0ESihDq5BjHAlBTogmmJUfz7z1Aof1N
F2xWNfbThJ9P/EAITWV7XO/4zhl/bzA5+8bGu7RiKTuAyGhX/v8/0nqwY7rqKxWl
UX7lwRsk/vRSnb8SE3L/Npf81dauvP6nRjGIXGJediawQpUwf2uMRZHCaPxaRoxm
ovl5swZeUBlQfUhIxjBCxvFuWCjpsl3eOXN+E36z0r4cnvZCfn9TqYmfUTKZhaTI
NKghg0XZU2CrU14h5w+8dT8Dv7t9QZZ/Gj9/j04xqtwTfSrnrAecRblXXkay1Rtn
t4C1fd18iNAKRMo4Y9IKG9lPooO+/yEaXIgSDycDZXouIyvIEWmXDgDgvTGljJcZ
bI9ROPje54FNTLNfC2HWfY+dDGMOsU/UmDpafjUToUtrdudySJWtrP9ca2mIXzWr
522Uk5Dd4CssWAAlWlzs+kRJQofcbqaZGaRgW2e1g68fpfq3G83pXbpA3Qi/maMJ
54eDTA8X7McsywuVHUS0DQdXAfrYKVd+s8u4Laqer1pkW+wvZQAM857VFeQn4zWj
cFkChqka2VuHJ992UFjx/TOggyaYISxdza5vyyayhcx5dQN6Gcxbhh1IcW9YAYMB
OEnf9ByRXTCD2/evTPWVKghwbAOUQ/cGcJYLHwQKPnouLHyI0QvPczKWB7kCp0VU
hprL64S/ozL6sjbrzDkU0UwBrVMXsw0m5I7dC5yLMq/R8LHh7bLDOlHCtsrFIiJL
Bhamzq9a4c79xBOQf1UzVxgVbH4jqqSQGiy3pWDzw0k5znKutsQW1Yfx8v5kzpQB
7UKl/1ejYzzBjPDlmOqQNHfmM7pN2Xga5AkkaIdfHi5vzs/ReeS0ddMECdjFyJWm
TsJW9QEiGHxxsgP2EDYLFjmOxxZ9mgFDSiiK9LjxtRHurNI1CLEqf2o1x/FqA7LK
Y3wXmgHyy6GFWy3gCZePD7Io6Y+wPKRcgRujGPIZJHC+XmvCWZeKutGugSTtSUrC
iKoe5RVx2JjI+Ts1ygLWtTPDYQ+hZPNL+gCmYDMw5hhsyTqtTA++OxAOhdQXoZSR
oAFNT3pkHTn0UUHEXLT8YiyilOnlOCnfvKRixbnEufFrb6o0x9d2WhbyKMLO1haK
p6EpABmqhrh/akOicF0JizmIiR99gRVzl9V7vMGuGvlZ/ZHkhY/Exfaij3qBwtxk
RFZ66iT4kaPXrZrpjYaWKOVlfkRZ/ZnU7zGe1tRt7Vb/TL93wEOzZtHQIt8YIZsO
67e5HQk6px3uYrYbUreSJ+aS18Dz44tv0T0rPkvy9QvIc1QwRGn5TJy76+9pLUvl
F4OCR7Y2jExjsyZgCO5cUSIQpJRBfCWUFXTOsze4aLKt2hN7Qe74bhY3SFXPDP3I
BnS8805/qfwDqCKcT1EVtm1mvd5RRB67hGzf4ZbOKWFQ8asI5In+P0OZ47HaKNxY
+dquntr538jaE5/zqR/fDOnyWBf2I8Nb3dlM+8z8ndO7uk/NVqPXotM+a9a35aJn
G4Luer5h9sVEiu4JYSl4iBtQBlwUW8TuMlBQsHnKYTo0hUdFbGmpuS6pakc0bLCl
y1L1yqtypXrLKVmqtTVqrt0IhyF3d99Gxy/KKS5bcDdhm2QOyeer4fmD4x/rGJA9
PV6cPCd69H8f+i3m1rMCfUuOdZHRAfCOJs59nFjGeDw+pfKq2kRkyBDVzzdc+93N
ChSeYyvpUvpJ76LY4ZFCXmsn8Y9El/rrg8B6PORoQr3cblrUNkFIuJ3wtjdOUFq2
JTePx+kmrOl9U6rNpbNgy5GfjnYwH/0C2sohvkrA0XPDUEO6soN5EvAtSmBDyxuI
dfzZMgdBczv8/Y6Q2YUrg0mXu5petK7u52JfFf2HKOwoR5XOwZ9u3NWZeMiD1QnM
SlXpuWGEf1pGYQ6QXESyGNJjig4sqduvfSI/6EMx04t3yFIAC2K2nehm+mYvfVqJ
`pragma protect end_protected

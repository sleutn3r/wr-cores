// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OLtcTZxBwFHWqRcO59eQDdn2bX6IHJSG2GL9Cwcve2UNHAdy/PtfNTh9UXY08mfp
N2ZowyZ0QgyC2inWPEGIzruby99S9H5iXOyWZSkJn+hMeYLoLej1mm4ETma/EZFH
yv6pNtnV33Pwuiw2KRnIhmiNXUj8a3RuZ63uDxLVLEQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13104)
McxRT25o3IkH01F4Z4gfMxD6H9t/t8O4GpdDM79TKXFeO6pdu+YZGPXcaxQdtiH7
4CF06IqkaY1fxjqtoZ4aGxg4r5glO/39eFPxHHWLe9uM3st9zFGLivde+OnnbbOt
80PCN7Lo4FrQg3apdE+gLq0J6UcDY3SD8/Qz4lgnqUguknOVoOVQ18KxHeOHQD4O
8hmsvduCTMKc25T/cxbZuNU9/1ddarGPoY447EdVhbkWLM/7d7qvrXDw5DVhI8CJ
i/vDCWTTZvYEV6/LbC+vPvFiWKckf4EbaJp8PxVNR+G9zYIn6Lk6BBd198v7GizO
4HtCtT9UP9dfBe7SN/0iDpDd5h/oLkYq47FZP2Lq4rSBN+UcDbXZSSdnoR94r+/b
arQB7/oGDdXRkH+Pi0hj5IoW6aI76dtE8JywVD2CClow8s4lFCnFK0Anh9Cpz4Br
XSgEOas5RMGjLUlKH8JqusRny6lVVsjDkegZ34vqRb/08ZtHZg1hHhvcqJdJ1mfT
zTa46r/Jw14cXQhh63x/41VnRhtGFaId4h/HsIaMNIxfcLFA99ZEXzPk/71GQf6M
xJaJGvS8A7W6l5YTvCqsq3Ibq5TGG46YC8hkUJeLTl0u2w15uz092NYCYPDb9i3p
/eI9HEQqJ0pmllNdqxuylZIhfc0l+7y5TNppp8wshv2o0q2BNFwkXH//ux54cZRA
NWPlDHFAoix7dmbibHkD16BCcsFezMDAfgoD9Wl/B15zDr5AsH4IxxRQEA0YocIo
ev2DA4S5oZSv8I1m/kOY0h4QqMl2t2k+lUVsN2vb3PuNRqBLlZwjn+rX0iDSam/E
KW27xyDQrFEMeV4zIyquRiiXSXm73D8HZJYW7XmjGf+mjj4nwc8X0kGS6H1sOGvy
nRSSC5sugSTNzUmcL8ZaQzFRg1HAT8/fw4HJg/aHgL3HvCOvXxhzlfDWDYND7qAi
336raVlpels4+wQeKZQjwQFWklYAwcPu61cSluLD/x4RkDQkmNxZ+2GX20VpRTrB
Caohr9CXtr5/wqJcMesiFjeaA7UCvYmcx3KLKRkQ1k2aGgYA7iDGeDZ5gTAChJEA
sk95X/HcwvhSkVg1vp+8lYf7iK5qCO5FbCw8EgvJZjfwajg5UOIooCtyFHhQe5c/
Oi3GPy5RuKgqn24Ienzj7kCml5lWG9EPfQkU7p2P2mbgcPWLuwyr4d81urMITJe+
dUqQN2DhMh1dZ4BbHPvC4Mp7mii25gaZRTYSKt5YPASBkxpBehFdggALJabl+9Ph
3QT1hfJ3ZxSWLbsJluGlF37hMBu16U3ZG/nSa/pNjK3dB17ntDcWpwy/y+cGhOHT
ed2dddmszOE8g9GnPWno0qLH8KwOoTZmbUwowUmghTNFOQYvPjH9rlA9B/ybhLMB
WCCKV9FH1XmqvD62NdaAb1++9YIlMWV1PVKnQsKWJrLkdXaKDFbhH7XRyF45qf9A
h5aRR4dCkCq4eOQBsGKQkyxo04tC+b2rdODAomChVTYgCIcmpgZN+tAC1DytHr5f
gDK3VdEEOD2VjF9jLzmQn+OTowoVpvYSLDm6D6hc7WWqIAW/PzZ+GA74yW49lyKQ
ZdURjqZ986CDBRZ8rLW5jnKlK1gUKRFt/Ts/OIQJ0px7dmEYHPmeT69Gc8oRY7AN
MO1Idh53Dm3WsIUWwaq3b0JURIb221dIiu/aZtGV4XeMjUAbmAiI8mItH2urWqdi
dm9mPKK65rcUTd8aalLvKYAAi0btzgn/DbhbJwQNnJbMPqu+lw2oNRKCGJp71zCr
XqH616iBH9wM5f/oawH6kvxhC13XPsV4EBTKAEGg2CJiMjyf3DSVWnZJaxz3yuW/
eD14grt2YHF932PB4qivzMMNeewz1CNGRSFs4qLaDr7/f94moGMfMU+GLLksT/fy
JlfWdL3TghPfzOFQFRFAN9yJZw4NlajJDBUudjWfDK3uZ76VVzo5if8hSja/IVJV
b2gZp61caYIFR1A7zwUKimrOp+LQBBT6/3oUnsbFdmyeDwjOLk5uNGp34uGuRARH
ASARmeGANuwd9ECqB//96+jROzRMoNKpLQaoHIpGJQ7tyGfRhxjZf1i4vL0MUdMl
NvKHT2tyJuaTsC15gN+nmLe1WSme5XKdnKyNQQPF54IwmPswKSPQkiUY/DJfp6pJ
1YEUe47ltnqPEsYwDKWstslwB22tZ8LXrZhFfA5/r7iICb+9FjQIREHkzcE/nAtS
F86uj0PUKkUa5uGvb0WQbPSW58snTVhOQm/0w9uq8cth4B3Sj8wZkKOtTesnZifR
kE2zb6x4BQpmJnCM8FmHQnASkr/tjRFg/lcE7Vs65t1LXUgTcuSfBNKnAGPSW/EG
qifBeh0XLhaDLZDcnxXHOdnFDjis4qk/WoXkbeA/54aW4t3qB1eA1CdIoqvfRWmo
Wot+51kdGmI7HyJTC8gf1RUQ9h+j/Qhb1LZ9hrXiniUHJFTxRkJvLw/dqqENeWf2
RgVbA3o0Rw9Iwker2yWbTBVAAc1Se4ds0rYDMmyCRJlqwFik8LkRss5pPCt/FO4Y
UzbGM4NCO7a6Rt7tpdpvAgXR7jmQBT51hfthENFt/eP0HemK8SnmJwy9WZS5zrhB
4eR5zjzdjXxADxWBlbKWT+VUKw1FVFBjQ0z/y/pcca/HQZ37dMr3nt5BR8czixW7
3cRi6j56luATQQHxaZwFDBz4swxQYw1QjlkM5MDugOWwYUlJ7hzPIe3WSqh9PqJ4
LbDWSFBBzEdU0+DllsiaLDjt1flthI+JfYtghmCMr3oAMycVG2UuoiRCFQPBwYar
kMdgz0MQE07aNkYDv2KF5HrNuYjZid4XukwBtjsK1amMHEo7oSIZgl99sOrbWjdr
DxqGeJa81imnhidpI4CiiWkH11hR7+97QwBNzm2UrwyPt4wPBO3lIPsLqrUahVdK
rm3xGKl1Z5l+DS0esi6dpxYCUWkJiE6ifn8Mk3nqf3FVdwG9n6CmO7dKrJoFyeh8
Kenoan5jxwfSb5L0NtuhFYLy/0S3KO8rJlQZFomzeKtSVyePNQDZWdePnMNw2Uy1
RBJre9JhDdX2xjkZD/ozobsxLrns0wOnL/I4L/D6vzZiQn8oXXuglC48GZjVUe6Q
Tw2Fb/BmCsXUVs/MGYM/QE1IDinNRJHByyWeTK5PCRZXf1+4RabaJoHWPaajPL5i
ThRe1ZXW1hrLgbCeyRohzHjwLdjt/tpAqdip+HuHEkEI5PPaXQPaOIHRQI4yYVwE
FaPFx68TPdK/XXHYjdm95ayM8lpXKEP9NKiU9l9IKg4aAWe/3o6FeqVG2v63PPWe
KOg2dbccTK3rskWSII70mIWf++OCH1Nl9L48icWxrS/lTmh2jO2cS3dIsH8EWvML
etvRmn98GjA09tLv7dqE2xvDiGqVeIe2kio67A8Q4v0rIUL9/6RwpobpPFN3554t
oYs6yGS2k2NpN7XyWRKOcCZCZb5sPlZgg1+JZk7zJ0rFWbcyLH1t5RsyTQPwPR0J
U8rMZrsT4BRrR5euLGmyeWf1sHk5KjDw2SecKJvsq8o209ykxUKTVjxEMHVONcvz
6Hyo+dIgGWuhcCAMx1igxx1LBcrrA0OphtFmOZo6rHQM4laX4nnktPnVPRJwoq86
U+NgiWiSJzVgs25dW/CPOdgSD5ev8E+d+fykjUhmnXDbG/Oo+aayC6sLi9ez9t5y
Mzydn87mCZVwG/OXKVnqHhbJoevpCDKuMt46uvK0wyoQUtcVqNFahJvrckxKtdyX
Jh9yKYODT3VuPR+LwFcu9U1ybqcR5N2w+WshniaWOd/SnH1HjXrcX3Hl7rfOqsKb
5jYItWuRUlbjSkc+9M1Keft41ag2bjRGm9FS/MtP8ZyU0PWxkb2EegeiTv4bGVyE
0M4Atx2XgknWOFmTd8JnUpFmIppYHrIuwB6tCQgJpluy09eYGB3bJsjIcwrbM/8e
lJgEaM/oytxTPbagYv7JaQ9dWUWMGNBcOLQJH435+O9iTD/JUv+oV72+6DodJLc6
pl/ySVp0XhYUFYcSdUjT4fbii8Mm11WGmJk47xjM3J8i7iGLGh9bO8WlC8yanvb9
NFJbRUr03n/06vFo6Nt9FtG8Fc30SCZR2HEv5oXXV/E6X2X6mHl9lUZGYmQP6hzl
pMZaGP/leEqRbEb+FDM2e8kd7VKAX+QtgfYnzLZLMAIylRKWSNBd5ZiCODzwRf4g
Dzw7Csy+KmyeHjvYNlSnE94TEbw0kkdep0XMiUEcD9ezVj6Ne0LeZXWGdelXDpDE
cnLSLncvYordanOHys1S8pc4Lg89VZbnaVdQrGNE/ImTyLM/mPrQzibg4ApupA2n
1RbfZPrez51s1s4WTNDlhEmXwfG0GOdoWm2zI+W2TgD7+wgblMyXFtwaGZMnk97L
UpPySlDwNiP33cFINjQJLtbcQhnmaNmOlq4vdEKtD7y4KKbFB1UCR/WhsswLmuUV
3lRoRe4UKWISWc7zCgGBK3QMISM3PA3EQfCcOyli6zD4Ekh0KbWidyuihGvoNQ89
olp2dz7eemr4bV6VBnjx6URpulO5WDJ5DGIq4+4TKzO4mxwcWRw8/N91roODutoz
X4u1oaZkZV8OCIrjKZG1ZDcEPk2sPYYzt1CHoohSnE1pGMzQsJSKhWVrPgH55HjD
NT+uhRirMS89EjCWe/VTpLo5/OMZTAyy6EKNxD4rU6nz/zTvi/tYVAo3iDaOUivY
RkCp99hoa0t3KZcjVEKRq9TIRsOwDNCKjAcm45EChOIbIiqmAb86WzQXED2suKMq
rRK33taM8/WPKVnRE7Qj7++AqhR+79OaYJRK585iEn3gh68avDw/Oi7dNphJXeLG
/4mdoFADNNUiPU70oWliwbTexttllUk5qmR39wyd0Hs5Ui01TQOT5oWdjTQ3X8f7
9K98cxXoshpdNr0XwkO6ZzVhYftAYRaewOldNFzbgYuzHsjznA4rbwX3qVqU7HHU
Dgb41bByAd/Djn0jkMonjPR3Z8xI96PwuWk2fdBjXH5Y+xdAfUtqaLfN8h1iduWU
5nKPZblgwUgwV8UmY8Z3M8pkiQAz3K807DcUmfUPb/936ZoSA3K/4Q391EOl56YL
iUHHNQe6ZkVaC8SiBJUTXJpshxgD3G9Kp/0V9WwbQAcjxPlEAHoEktVpW1TDmcM1
MMmuPB6ntq3V6nWKx2bd0BfhLq/0WJVa45ExQPXRmhBOBgkXYV0+p6GIe/bS3gIN
S4baPTYni+7RXwzPLSaRhMT+y+XpaTAVJV2i50K1vRfdtUaLEcbIyQ9zyVN6M/fD
RBbB9PK3FOEsmLkgZlgxa437ZnJrAhHSmkLw1gZL6xk7y+rhabEY4GL8H5jTQDjd
VXhQwESG0LkyRblpeaQDiBgXfDQ54yj95eZKKB4XMlVRBXVIUSO4kkUVs1BEQ91+
rm/FJEy78ySIbsyDG9sxsdLcAvTbcSezfKE1vlbNsRhPcJo2T7udxc1AS1Oq6dU9
2DhSaEcd+9j5GHhxwc81lkD0fmbgqXZ4xfVX0WMViD84no8/WYxU7d6wGq+/crJb
4TCORUD5V9yHvUuDHYEMsI8UYYq1/pE9vCta0652iRuWrsfKnIWai1BmQfGuit6Z
LG/JL1UCQt4lk1kM3hsmab3Bh/mGsM9ttlfBjgkQ8UhkMTnIERZKaUduQmUoWBfg
FATelMVl2XhUiXXbg8NfTBlnmM6xVS4X83wHmnhI2pyXiqrSzg+KFGqFVbP4wtOo
tJ+3iboOWvHV2zS3jykmp3nLTQmCmyKff+saZN/WdTWlVnAqcV6NjIPuKGBbfSwi
1BFT0/ZxOegYcZOwiXhIBjCqL8p9jghSDbWOmeUl44KYgzWuEV1w8yzwf56rNzNX
gMf5gt7g9aBvBG0vvjhH8H6gWp1WAykzC+Vvzk7GOlvd6Jkn2hpH065Lk8GFaTun
9gtxhjlOMxra92g/marforowfA2QQjj/S7qZbOSB99zeFWU23IBA7ZB4cmLZmspn
m1/O6XsuAhQ2RPQCU3GNRXKvuIPvtWE4sxKuhnBcM7hk53dBimVzaCWDCxrMmVeN
FgOCFP0nRP2GIo2VUhOxDm0rgqko0gCMAB47viMlFTmFpmEBE5xsLQfPBES8jAaW
ZutH1LJoVCZ6FqFZ2XIDHbHa/+YtsXJ3tONiPiGQ9ZIaxo/B4gm+jZLj/VmuEJG+
G4yEJlv4cr7d8D8TVcO+1hFRRN98I0lfbZqnfkONBVYmBd7p/Dk4hFN/bFKB4I7i
5Od0tvBO5r4SIsF1FIX5f3Xt3/4Kf1aQoxeTmC2pAUaTIY6DACCSf/BUx63KM7Lz
u/h2/2vfP9/XKWP/YkBdP6eFkSA6W+RKBzQF4bHxjN2nAEO0l+dUNV1r1vquzANx
y0F/PnPwXOPJsKnhO71EJKM0gAWqeNQy4M2QjNbmqZSRkUdg7ilfgktd/cO9ADn5
m56ssXpJBJPMOibziNGcfdIgccs6UQNsa+ndFiEhz+hCngUd+f68C6nYcCY0y+xx
caSinEqxtaajSGR3Y19W/x4ZXyHCfXkKDLYGvz5xh7SlCIB2Vkg7lA4BnoRqKPZl
a/4/X9pGReezaLmWjnoonKhVq5bm+bYK/UE7f1EbQ9ITxwcjW7f4Ff0ceiFBcwwq
IKfAIvN4k9FrztCWQGzsSPEBzG1UE4xb9Qpc17P1sgN7AHkfwSUS3udc3zx7VH1V
8vD0Yg1OoPXsNQpwk/xL1YACe02IErYe9pa30ym0yAdzpLB5n5Htl/xaRWLwTT3I
pgggv40nFGQn5UVPqrH+4zPwGMrqpn29Bdb4ADCrIWJS4V64+e8s8cdDDt5LeE44
fz4aSGZqUL7AM4VYDWRNNTiTH9t7TQmCZUpg+ony88Bwkx4ujkvhpfq1i+4D7Oat
wh7md6/Ir/LmOvp4y9t0UkMmYace9aM4Kk2wM4lcMMW8j74V74vIpCkLx/tJsWt7
5mdcQIxnC3Aq2NQlKbqVf3ndGxw6CMMtyTg2fZDtHEEkTdNo5fcYBxGynkQUAY6T
Z16120c/8KIgPCuCT68ZxoKniD8SQcAYHKO3ngzlS3Y17TT383huPdzesmp2X3Sx
EUTw1DpXNv8tWvJR9jh/ZdvnlxeugUtdLK5bsBRCVu0xmHeIISNFFehkhzG3IpWC
vt6GnXgcRvUSM9RsvJ/osRR9d+OWYtW3VNwsNZmFkOicHxWOkVOUYqwMXlJzAki1
mpdjKOqD7wiJGL/kS/D6vsvC0T7TchjxUVs0PlDDY6Ky66QJikQjDeJ9nqva2ScW
l0aktcd46MyTO8m76jiylSVYD4NH58YdoVfQQEws2EZdAVYrGSPxbxFVihRO1Kwb
wXrUe5OdfKDFzn5PdUyRmBPgaDEWUGc3Uze9I2+f+q2yk4BFXZ8nYYoyiKblnLCI
2hweyhTx6uFqiuCaXqa19/Gwpwva3Qh7uCF/Am7Xw9T2oCQLOrcjtuwKjSHtzmlr
nqT0svFr6vn71Ea9jMl8jdCfr2M0YnvhGCcCkBm/nEnC5z5f7J/ep1bq4wbkMIDS
R2c547MqAnr0Zu6Dmrl1zsI3+Q3DXur0Qq20PlBKx3OjzCCjviCJTXFjgCdP8xgQ
vhf7BSiKY04ukpyatLyMvpLU0Q8H8N8ftLuxoLtvmHu34SQqcXIly3DA5t2rUESB
4WIP494o/yLXRxZM9k1JWFu76LPmFewnhkuxuPDfGo3V/K7jyESYfLY4YEBugNfO
KdI0w++lP1C4aS8ovfi0nZ+vdZOHbgfg8LZjQ9g5iS5Pyll9AHT1nWvVk7TExouv
Fau5LGYTKazk5yZ7fKNrKDyXZomUs2YfHcvJogcawTNFFZn8aKFhA1P5OZEk8avl
AbeW0HVKGVuZFBiqBQ6/DmLKipJGlxAKev4XpA6TJ3b/UuezKkJXTkY5FwTGcEdB
AkVXoDzHkZTPPXcVYYRsewPcDUpm31m6AhvSDBRq9tDQh/gi7nPQKFTlAkNVvvhm
4V+hpvYyvN86L3WElKo+DoUPhcJqHhQ+NBs2LF/tjf4Fxt6/fGo8Lc+dM+k7VHor
tFFlo3Xe8rfxSoDCys1/FWNIrFcqwyo/GOqbMOprapnDI0UT0OubMhG/jAfbK6AH
3uerP3vSk8QWu+oOYkcTUIJcBOFagLlWR0Jug6cCl/p9LmTe0J/rss0CVzlotVn4
uNnUpw9SMhVHZVWqJhUCJsgsImxEPczNzSJoxc3NtRcO4+zkDfVR5Hhdwp+O3aHM
7Za78NdFE9TwOxPZYMmGl6fEe2aLVZJEj069xcJRXyjcIZyMHOm9mbP0Mm71P/xk
3MRJMtw+qlikfiea68fbC84tsgZ6bA7wA4SM3yhgiNsyBlDlKfATWlAN6gQvcRnQ
DRm+tVRWJymvy7akSjPJumTrMdt91xqQR/Xp92DqhkQ/1eSY2E3TcgsVJvsLliy2
XV/IOAkzQPSnn+GjHzGBIQ1YSITCReRF6ApPNorjPTfDCLc2rivXH42+OcNhiYlt
jqM0m5FDGX07bvvs3wX8KU+fsDnr20Uq1Vcxu+VGwthn6tC0t1VumrxYJp3qCbQQ
JZrod8ktafyYmdTFcx9+mYkQoKt79Fpa4eLF5NI+wwZ39k1mkDoAtFjRcLziTjYO
5QW1qFCaCDawfRkH0yk7kyfD32j/7YvF73OFC/GazT+9mfzcDybJqtitqcxnqUAr
MJqTuy9MHXkytmbGAE+gGnObgL4MmVG6MuBIPsREMz4vzMhVQ9Z/upsDyZnzpTPx
JIdOoENVCeNU4toM5torxTPdYW5mZ6Z1Etm1TwYiBzNffc5+JhyzoFKXCC5ob2Bw
ZIrmSJnxvvO+uVug7GbWH8kR1n9HTJkJN43naBatXJJeogle3nCLqVfs6FdLYUiw
u4lgs03+/UQ1UXsBEdumFLzJsJwyWliPTVA9KAZDEkctaH3I9q0J0K4AzXKR5g9Y
k1p4o2/gg3vusduOjbFxD6fR4pugPyCLC3I0qmkTPLNCXorsGXtH4A8A2XVtbtO0
PqfsT3mkHbI7scdEGTlPxlUdtaRj2OFIjVzTSqEJ0no02X144EothMDc26R9Xs3H
K30QmoqCNBThYI9QJVeuhDloALB3s7lF7DogbiUAI3hv69sHlCffjrjx6BmBwCUN
Set3GcQv2gqvbjT6C9ryFEb/q5I4eVCcFR9cP8nDj8m0zdk+hX6ohQCRWWIaETls
ojFprpzGQLztqINDtfXsaXvYb89OTewsAnnucYdWSCijYqy6QzRi5kiGiXmJrTb7
oeYpr1HoUOYheIM2tREEfxK0TZKKPhn/FJPR8m+W+zPeedc0+z1sfw8AFqKlMyXg
nFe8sEwDmZtnCZcvMnslOMZLfwbsy2JYtB2wrEm9mIcBBfeocI0Ns6Kyjhow7YR1
9WbwCG2sWKGb5XZHeghGJZ2lBMTuNc+WNqPTu66kbHFeySK1k6HeZ8fFJq5elejX
nMMkfbqY61eNKmaFxKS2J/KrgbCnlNmIdE3/gIiuNrxpIRi5vv+IhzIEbvwh5kYy
NJAuV93+XfTkAUtYnPJBXnNk7RufUD+0UxpnwMXJdPfi/R4AwQEl0Ka1ciPR+EgE
SmKm2mChj/0Z5Vixgpl7gKRaohk8T44ltK8xnQO6Lh4WKTz1EAn0nxk5OgReICf9
9EegAprmUMGQm4RLOhRYr2EMJ+dFU0sx3nKsHuxhcDglvz5MsocFigim/13Uupb2
uDK8mKkcV/gLkwWSVRHNWLJVlL06xLy9PGoxPo3GNAVhdEQhwSMGVoQFx7t5MdIC
4snSZE4Zo5SkLnUGR2ruV4MIZ0/bx6QCgkp5vYtDi7s+kRPh/WY4hAcm/YuamD/N
ZTP4jgFapEL7gAcdWniVoXLRnZUicH3NxwcTYjpI7ETN20aN0hn4P5QzdHm003qQ
UY/MbkoNFuhdoAV4G6wEcMVOohH5rQPK9CZNBJNwPVijXvnZz6V2mxtPKQtP75xQ
0GMwCsr9a5V4Df0uPUqmgWZxaRV4qn2xNLtSoBe94rPTGGWmPG9SWzflUT0xg0rd
JW+sZgymmYlrXN0aI9sN/foT2j2vj8vSCM7ozJdZ1yM+Ow0PVtfkjrUCPMJqI47j
ftULojyArwjsg2QxeeCH56xuazvKWziARff5HHp/YBKhC9YuPx2p8IBdvAKsAysd
wVj9sr+n+LBwLandGp4wjXRlBK75KcJtZyUKshzYGiN9IjlKvZZyKglc1Qi0jRP0
awRH+bR92YZNqiA1GutFNur+GkvMSXwwc7BM8YjbjoZ2Am6dRjOjZHPxUmKzp8ja
96kMblADCkwnVGzDWqqskpJkB40CXUZnyyLnmk9MP8idPuSrSaAe9nmQl8kQkC3U
srheZDjBRSiyf3gFd/bVkvp7zfTQAicqK5eZG4TNGOQeyhPRw50oWRyGBg0fsxiC
BY6LKsBhy1STA+KTUXf2Xdu43kMJYhh8FqcxYbi/rRDV+Z2vO5TBj1p4wF/WCxTv
yXucVjFa3TNgIkXo9M0mWafFu0WZ6uMhEOeq/dRlgZyJvoQvTX/PYbYXK5xJWZTi
kHAj6k3CRdUtZc0suVd/mS9NMQ++3/hAbDBkFYyE0DhNGOk9KOWT/KqBWu91bX9+
IB2muR7cdhAT4gcs6T2+EHPrpRmka/pFAVNt6MHFDyFpgJrMfLpWCjeaKe2vSxpE
WLURg07eYFZ0rB6iNgQ1l/hFVt+tH3DZ5vceBNKSJASe+jyNC8NZId9PIpYqMxRN
kDRZ2UXVgFc3cMenmyCWLYEUUC6mClQ6M922BoGq4EQYvVeWjXa76qe9T4t+G2xD
1KqZ5aKDvdkitMFmzuDVBT4NTeX1OJ5KuhDRtnFjhplZhWvS3HkXIO/c+gMCO8++
fWIMb3YBw3/CuTj7IWx7ktbX/UljmyBIuEo9OCmQCng8kemPTnfYQpdWwk2dM36s
6Dm9oqJTIiZpeHopHBnYHNPm920lVzLCNzbimTmSt0+04Gpm4Uqskmkh9v5EH6AO
GaYb6HR+YXQ+alc51icGBYaWbtsV74c1PKE0BLkRuxe3I1Mrib66SB9IKu/5HvAw
fUBCfpzV5ZV7xr8EE3hIB18Fudurkeao1n9gUr5M612ytBtAnNVEyzomULDZYkVw
YkXj/kCbTG3v4+fKIbo0ek4v5zjrwzzR6ZyweiRBYjafLRaYcY24IuA5lSmYn9nd
M93OutlMPm7DpaqlKKdtuRxnVGNLAbA8Gy5j3TS+13d7d0zC3gIMd2/dvpnYqpqE
Grg50kLKd020syR6fs0CfCAk0GsAkKlMTuD/+htrbJdO/q/u5HQ7k73MP5m37TMX
udJEcO+KDxuaJwCTEPACNiLfFDgJJgFVGWcUNBD51QREJyZu30WX8VMg4iG9tfMt
Ff7cdaMbJVDVgH6ns9CD35liaIFqWyzYhKW19kMWni8SOwavwoicelsxQvBW/MBI
3b8186GKnWWrFYChmsiEd6MHSiAb5mfyZnhgQqNv+d6jharjImxW0tQp2Csg+klD
TZ6t1ex226n/hvoWzv4F01C60P2lwxA6ufC8lhHE4hOuQeFRSXkY3JLmNtU3i/7o
a3oO9QLMVDL2H3LmPzB2IQ/KiA9MGCAq6QkkSP6YuvobP2KGLf0kBlLok51a1o98
DW4j1cOW75bA8FRCnNEiklpFEzv2sjugLnfC4zoG508813Sc1Cf3M9/sdWn9lHsU
Tpgnd6lVP6nwnMi3dezGAAq9dtW6pioQNLrMwTg0XNexDA3yrQVPb9FBybaIOS2e
Yq1kUZjW4pGOuuuPeaJCU9sqiKaKRivTyhyNvmsuBwnLvu9Pu2uk0OSrpQ2taO8O
CEe3GqrNz/RSNo3zRRLIJ/M94nvO8Q5Iabl0UMJhHHiQBvF4Tuu6V0EqC3oRQrsE
EwjGGlvlS9NwGB4hNzNOtmAyYu3R/53pZWaEG6A945HrW9zAMcwGxKalWwQuTtc8
82LttKZmY+iZ8Spu8kK6veqqcfMSQXPlEVrQQLRZS19xHLVFxJrRnuIHS+nXnfpy
B4wP0O3dxm888NRJC0jOTXfLiAZ2ElFzjvF+//FbM+fKOfmcgDgH57p6ds0WC9te
UyWsaJGYwfO52CLCszRPEnlSoFSn5Ihkd6G1T03u5bolOErA+NdFZ0jYuRwBKJ2W
frynRSwlCAsoFnqlczfh7NnTv02GItligg6EaOFwQxNu+EiWQ2J2KBRlu9g2ICbA
CLP3Z9lK6qHb4uv4N8bTCP3B8TNkOfG7yXiRjDmnHd9ZwTlpIPuVAN8r29nS2Wxw
XAQ6mzo+GxQhYVCM66ZZusPrtAMtUqm0pIcEV+u/zCorgyHlSdZEY20DWJut9fU4
XrgSyTHrYIJcajkBNN/pYoVrZXT7u0iVd+glCADhpqOkV5T68wgug1EY5uBFIXeS
nNhkMoFSFtuYb5YfAld8ldVOOB6vfGfj48OhTagReV4LdWGSv4lZs9JmJGkGvIWY
4y88gvU31XfrLCrCRyhafktBxz95Ygv59VEtq+2mD7qsHzHELKviDwsIRbQTqaFg
zMRp+kJ3QlZWxsTY7a9o4StERtAZLFN0/DncoUTxl8pFubUJGV6NGytbKRY5GW4T
Wecy8EVkKM7lnIGWNfZJ6ll2+14tUOLtykn/QcM6QH8gV0Pt6sx5QDmIdFRjVW7t
lQ6DrTWf0JpRncSr2woAl1k5aTkGvacKjd7TX5TAqyKPYTKBX6TJQMpu5pjbHp4m
V9nKQqASdHuZRGefm9hNdsMfAjGWvcLeFjN8Thwh+1AaM2tEkzJo2t1FqfS0PEX0
IYSppXfhFbIsDtqu4mpLSD4tKGCT3jFpZF1wpr2qCCPE29Q8TzmGLvjpZOrhBfm9
SfDRjXs5BFEnbGpytsJ5K4mk1o9hY+eL0L+8LvcZ6/WuFDdpIfHFL1ggpaqje/wW
Dj8rNRge3lDMX6jq8uCZ59NAiuz+0iyMtU3VVQZA2eJu/dVDqyWP7diBm9oPL2Zm
i6Dl8jhwf/v0JV/4MjY63MWtI4jcSmJoiCgODYXNxh3aXODH8tXDhF/uBZzjiADh
Y0rZhASe6AWJTabfqj3STHGj2DrABwazyhfS03SNfID8jBItcyT6gZ3XYz3ABXMG
36/J4w7m9KEpNrkEsU7V/+aIqv5qvWrinDqpKFqRLSrsk9z8HugXx1e69zKo2C2I
x/QuCG+f/lgy/muJEQ7veYJaQ2gPCFkWPG0MlNTmgo4sHSOBfrH7lIRUG1k8PNVI
/Jz9wZveXjrY0oZazGY7Q87cYWxpMNzFX4D3qeZunqzvr+icKjh7aKJv19IYzgaV
/EA/HLMN68eI0rYa1fli8JKIFIzvdoYUkt79za8q2oYnOzAYDGIVvjcilm65CFU/
NMWaQwEuN/TqI9R3PlMgk1Ik5JuDXRzCP9aoCxpaMzzBIyBFfsmrHMOR1mbsBMa5
VeqsYG/3YaBUVd5xd6vNXy0CtgD1WEjEtmfS+G3kET7y4QMk19Z3SjzPq5oBHYzm
zAn5lAANzciM0xpGEBz3K1ZBNw3FvJyJlyRZ4UfihGA4ah6fBOTUPkeTnCTV+wQq
wSytfYxp4DUV3GFrAjmq5slzpwVY8xqpgVq2EPErPu5LE3YZvuVBhSPKT5fQczBK
v6zj1IzijquF9+wqww2rcCGDvFuI+FPBwBeNJxNvA+iH4eWVMc0OPstRG7Y07mgc
xs6g6mAjlnnupQTOiByCCaW1ozTNgT0WatTTeYuhp8JF483363uAMwMxBPyBZh1M
yEobbCo46oSgnNDhMazdhUqpMj18K/0Tb+Yv5WdLbZWHZiEoLrGL715Q5i9kwN0A
44JnITa/fsaF1vV3iM3h9fAVjJnCIThQh8bW5zaXffr7kR5gR/NwCoTF3K1C6DxF
hR9AdHZcmCOU34lkbLOZ+jQS80BtJuA6zgGndW/vhHlKcm97E2MIJ6iqL7crD+fv
nm9rJKgDvVcQ0yewVKdObnvd3yMizzeRbjFjX2DoOS1EcvU3dD6EIztAs3644MpN
/VaLZ7yx+wUsPo0KsDV45T7eSpWeKAWArFxZTKr6yLHywQPFK/5u774N9mHvPo/p
hdTkRFTQG7Md57qHS6VGJACK9OTKDtM+eJYFVnd71osYGu9tDLET3j4+wVQFWOX5
MOm5neQ7zJAlZ/xIsfWsZ03Zv5/TzYtaS5waRH9IblZRaxtr7WsaYz7qPfl72GOx
+gI407TPITGOyPm2bCuTJaT7sJClzdtJ5aiLEzHiYqFv7A031yj7xBfw1AZFnx7Y
rUKUKyezAQeL+WOCAjz+GbGIlfDEcncw4O1xHM/YCkgB3/iApkzCAF/rtqjABvbg
po7oddQFWgalEb/0gHH1JcO20IVHH0erUxQ1fzdBdsMSr38FIhsvio32cEU/r8Le
H7eQBY79bit+CWwwaal4YhBQbhQASt+2STio34YffBFsmTVjIrXK5kz7ZwWMq1pN
jDz70vC1mms9k4aiM42DyI73c9sulTwYMjNz2TgnHyvjxIBwEqS3G0Eo4w/AaFBo
EkZAFRRAFPls63TCW9gEnWJX/ti1NjAqhSWmcoRbYXj4wTaGlRlzIdD7+LQAs2ul
deSAxwjrpGau0XMmOKQ/ogT28duF3B+kBRpbY6qY0ew6mpyY9ndfQn7IgMNGtesZ
UP6Y7EQdabjbyIJhINVIn5VujLgo6lCaQzzZhSjLUJkKh+sp9Xe6WquRn5KnxeEE
vqPBWgI6KdTd4VdSn10kdm3DhArOudjxvUCGKSWVXEmGy/g8gl2jHJlMz0kqC0jf
6m7a2vTKknj48Vb+FobLuXW8Oz2lAGyb6CtJF/lt6s+GGo0YHk7w2YF66TDa5CR1
AhQqqOqLXNn3FcW6dzOU1lpf6ALfTCEj+3PB+JhhGUvmeOup0nFpv3xep46HprTM
luossEnOqKE8JSbCU9QL0FYFWoiC+/5ZVkmNNYlir3n8p4IcFd9NEVMn14sgd3UX
llaHzbGG5Qp2Ab4ugCFggTTQu/GLRA/aTbKdLz2Id7Y98gwBtpAqii6lZMeEn3nS
cZ34/g99m1pgXeQllVOH5p/P0+DeAc0wpboKwFrVmx5QQIosHoA/75n29gLoZVZ2
8PqfoutY/r/l12NrOQqL+KfRtFS1NhOdzXdvyVDWyQ2y1+v5Yv2pln7XCUvNHD1F
SUUS2eNYa7UNubEzOzpd/WNQitP1e2xkCwj4ZYl/nRle9DJgPzY0WqcEBa0X9Ew+
ZEnMn4y6XPeoPqIXXu8TwQVNtQSUUB8d1WXnwvV1QU6e2hxpYjEN5460aWmPoBr6
y5cA8r3JfojC0GIGumxLqC+Ga/5d693/bohGfEN6gAPr93WvjFuxRCEu4g89xmXy
PazdynTuzDhqmL2rItEUFas4elT1+7tIxpMmhOlSTqyuL75NwBLa2bHAKwLg8IQI
TqBPJdaFOVBOymAAJK6VNYUtXXsciOxl44pjvO3Eh4njdeKyhRXsb6ZRKKst6lKg
S33kDRCXUfTgHy2K5A3VRCE7HWfZoQCr+mrJx3eAjzqZPBhtC9JXYNWMG02yRT/4
w8xMuy946NEGuBcMCJqEjxnHzgKwwagob6uq91GyncLy0QzcoDxK5icOIkxgh8qd
suQLa141+s3LryUskPSURpmsGOkoChElSgXDUHI5xjQ62AF/uNku4XgdejK9N6fA
o0wijKE2z7Nb5lChfl5Uu20kcK27pHTRz/Vmh6W4BleVjEVRzzlwOJBY3xA0gIHQ
OlrkM+SYsKXukKtsEY2iWsogd04Gcyqb4BaQYYYHyvbjZWavLVt+kxCIF1HQulHS
8L4uWL/EC4+fPvkbEAH78zCWdFVo4rfLl2J3LhnvKo8rCKg4sYnOPRm5B/GhqjGh
+CX5foVqifmT69Orl13zKhv0Yy9Hr+oj43FTeNu9t0QH3tDaqMUlKAkTuBGT/jfM
tCeAi4foHagZBg8jBfol0+BgbuGHDYGMlOzcK3rv72YCNwfn+dSBJsTmcYePwG9I
UfyqYywew3poK0wlynMugzE9AZOPIToGBNZvfPwjL2zORaADbXWEZyf0cwY2JPme
opFMgeUNk3DzTFAgzwg0t/X/TiOnUYm3KzLfNc5y9y/Z+4zvsJtCFZLHlF+YM+Ix
iWtFzoPxymB+8MQAQkUyDS1pPEMdrunPE8hIenzJcqsSj1Q+iywjkGzRo0jaWf9r
GwLvfZwReEdsACOnpyVvg+kxe3ZGMWu5PIxLNJn7BlijOwoWG5/y1ZOAvHtrdL6T
sxRgOeAUBPw71rrfS6QPHpxh6ExKqBNUne4ZmTJ72OSjT3Gm846U1Ivr1jx8FD96
1gxauOigjkgtztlHBCMYjW3REhPiPUr/PHDVjLCIRQMUEvBC4dgqHvGfGQwAibS/
O0H2/RRLc6UX0EFtnqnok0LX+qodU4ztC7t1G7Pcr6U2mK91sWSHPYiu04lmyU3x
HVrlAfHfpOiz7/8A5tRUR/mGM2t38Z0AZX/4SDUQow0v5CgvgyKb9pLA/vFdfUb+
jdgJqnuNLLkOgwUuz+tDGPoaPWWk8EFPuLpCUapb4QyQQC+k+PVogVgtt/JO0LT+
nrhy4CMREPhUgom5mTaU5LVwFd+4o2WIAX5rLklv3BBTyEyVdT1J3DVFHzj8gwVH
5Kjvq70/WVWL4Sp8SxgZETbYMyoDbrMDzj3V+a2obM4d+Y4Bbay6Rq/V+9wOl8Cz
VMH0+gj/bIneMkrGKXVMySkcuY/QQAE/Q3wV/sMIoqi597pjhoNnEdeYWrB6M4FJ
u5BRNQ2y5a1G8QJkXqcERfd+rlCaUpZpcbxdaR49k7x9Knw8qvLxn5Y6/zraWgI7
ReI4WG4/3WASHnCje4MJrnbrucO7sCSj/2KWMmJYIGaSJo+s8GB/TtJgaazXiwJo
wcgqAL0F3SRYE/MT3BT+4pdqnwyHBQLQzt9qImDOg3ro3/KVjc0JjEMtfGzcx7on
egPL1QnwH8n4KMMZTLMACMe1nu+87i4GQ3Rz5TF9TwDQc9U3YXLRqeVDJwqB9SK0
k8BAX5ayghC0Xq9gUlUsDPHKpIB1jVvQ1KtTtUYvXkYVzVVBkWkd8EKcWXMCnoMr
iN/7gXxLctcqeZgiLOZBHbmuTyXxwqwz/TxUn/4W8qSVDn+U4VGnsopmBq4nhI8i
dBA3CXzEjdM9E0qivcr0u9eCP3pJezgjtDO8KMUt6fkuAxtBax8X5NVBgryEX85L
V0AQYCf6HRQtEFEBbstCdztiqx9HLkRb/9vzGthLHhiUsTMNa87GDGhkPykecZXH
Abf2a2cpQXioM9UnmmBhux9/AqGTQj/KOz3Yhy4zd5LMQKOeanHy63I/jl/N3Tp3
69nrYmi/BEYHNkSJnBA1piD6QG9y6V9+AT0Tj3GsXbV1KVsaM4cv9P5QFcW8Bt7r
CVUZXRWBb9gT2rbd8nBeHHowkomprphBt4yI2Y1VLJBJmuQiSB4qfU+gzYFKSXLy
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R5oNVC86PFy6tWK9H69io9+10zhHq8z/2Hg8a+P4L7xIrPFq4nK9KlbD6U7ZrfmD
HjtCfzB7G3PA3ikyqPCfvobYnL0Zxe0fV+9bCs86I4D2J+8AeNDsWAE6X1LX5Sgn
9CS1J1lfdeX8HwCCjGMnyyrR1PTlICV/n+YgKFd1axQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5632)
wgwZlDmrejlq2NDOgHIIVbCKEnEXN5JjzUKvGvBZ9rhcSvhOvq4Hi95GeThopExR
VmyYJW8N22ClnUErqMioY1YS2nCeOb1EKlmgYUyym/l+6BMrr9chHhOu9+opjjEH
JQBHktId2RKYI0HFVWxk/F+IypfHx/7PagKMGgpxQN4UKdJLyN0caHdxak505nkH
J4l4WaBj5sb9sPHzryifpLDXuWO6tBRSbzcuymQfvYrMztg+jIlXxgKvVRqafYi6
Nzi0sy0jwUUSq2/RD41bnzKBmbl4+3H/KXcyXZ2TmtE+6fyhyy5Sb/9TDJBn9Aol
KZg+FKqB4WdJfl6YrYA8asEJ13AJIgHZIkj3QpKvoW2MyE31pUrR1O1wiEx8IAX8
n4L6iHMSBsdBB2eBIOWDnZwPNubRPG+jxXsFb+oDQKDmCIRL8Saz9QZBJYeqYM7M
TcW0nYIt4mNA67NVitgCCtlifH8cx+T78/G+egMcMshKc4XknseExjhIDGLvqPDj
6RsthORLjaOkSleynuhgDYt5pz0oYcwQJ/FxRyAcMxFPRfP+AK9rkj3s7j8+KdNM
K0tWMBynDXv007M6BSdLVPHocMjpvbc3Wi1NGgk8bvXxON8c2C9odjXfYY875QaU
V3xm55mOlDKU20QddPUO+6vVXiMl6rWOmeuxCv9leFpE6zAVwH3nz0ljvbGJvSsL
QsNpAiseQyyF79WSO2aByD4VPWewnUxDto68CEMMLtX6r0/pP9ggCmocl8hnBR8i
fHicZd5MmcSVXrhsVi9kWOTsOKmCYCpW11a9vq7iR8OPtbPPA7gVHTXqgVc1GH3I
MS0lbl9k8TZ/ZFouONExgOvQwnE7cRHtiqrljYLegXJyQg0CCMS3YKRf7nofkgxg
54g33AFfh9hNWP20hgvWS1GPWH6eB/+tXRrQoqwyvdZwAZPfaDANKfkXQb6SKpEA
BNIOqW9KBN8Nz0JQUDd1b5YXLg5Tb6hmQmI+v+k9c9PoMm0r5F9CdqBqVtmM68F4
m99JjZyDjGbW2VM8zNpz+891M/7SNgKZRNtDjNfULixv9wafMpYJGD1+1v8otx01
LB27pfLG7V3U7ziLQ/szlk47KsuWa9nnBXN8pG9bd+CTchGMGbIYuLewlsXhKkbG
ipk/dQuJGqPPx8fNJ5m91gu4MFAEKhr84bgQpjpBLnHPFgHo4dRKC8487wox3T/T
4ymXEwVZU9RgugAEs1aGVBZN404v2/oF0J6ncbc0IvQXVhWTmeea9j4jff87IiI0
3fmRzQFnhesgeXaT8B2cPRg51q7Ud8M8DSk0CiRH53adlBDcfKHTuCJJT2xaiVcU
LrTCLWVt3bcdwDwIUz7/lbuuK2iVql+EQ/uK4RITg358j5CcTUQHjO8AtlJVKsky
wtpac8x+7BQ1a80npS1WmHhyXJtwFtjLpS8KsKqmdmIorRwVghgTPAZjBCvlm3JT
h6ZFFX86hNlEvHY60illppv2AjL21+JH9WOENFnSmRhKYio35dGN3e336o5kDFGL
0rZICLBD8s4v1f5AfqmDndHJ8PEbzKHaditb/OXYho6DfSJOpJkZN41J/xQEmYxQ
ZEqVA398JXwJ5RmLIaXNL2bbviUXOELbnCTG6tjhJymI6tox5ii5ZmPLrbTn8qSO
NNfIyaxS726zSD9aTlVuQjRfi4zEVTcPE6p0Yd3eNA6CZF3tGps88O6UbrWbAW9o
BK3KkKXQzzENMOJJCNkoF/n14MtbUyZLhTs7lKLWkngFBd3kNCWdtY9NmV9NPobb
hIOZvuThG6hnc0QrEvTX0FnUiRJKpqWXEeddsM/0Lmr+C/g+r9ubHviM/iGmROwZ
UytjUIPzZevxxkLGJRN93U3bpHw4vDdFgYlumfN2DSs/1ck9LeWLom0zw1eo+m75
zLckcq8hHzLkLuBVNCFuaZ5OuZMwyIdzPeQH2hiikCWDDwQoixobkiEWJ5jeDn8K
/xDEYw72xgWJPHF85Sl1SqCi0OUm+AmsyDomviDfyCC9wQHMgNIJUKk7ED0RaKsy
rU2C7rAsrJLjiwjuBTwQqAuRpyJifxmI+N2sFgxBQYH++mQNegcQIiO4XeJH/f74
pGnz4OjfYkxpUqL/HEeuaRlEa/3csklNcFjIFi7u2eVsX8TurThgwO4JdmhxHGQ1
W4xqqkghoPz5hCwdgIUikyEChlXnmlDoFhWCZdLFnS651ODgJ8EGmpoTbE9ei01V
/tp0nclslhQqDwoDMyxhmMKoBnv1SrIJvyy4a/miiMZZSg2ve/u73CqLxqM6wK+J
Of6gzJ3kSujYaCiv4cLLmyHcFeAaM3OiL9tvt6KuxPitT/kZiu3217gZmge82S5C
8K1FfSEJRqriksh2NzN/x8ah7ICMXthH45qC3mspLTmNR/P+/nWAF65hgbihR+9t
Zm8C3h7cVcU+K4EOAyQHsfCUdVAaLAiWWISyBOxitVsYwsh9nn6uvyCWeKZFmazq
qX9svVItXPNmVgGvVyxSQSj1vdz8DAM5pUyctRCxqXE97Y/0bkM8ppGk6fUHJRZu
nfGsHhaPRDwTh0FvjQEAj8+oIQjxqPsOZOA0INHUwclPAADNe7ZD9JicQDCquAwD
TLLTay1HU+tTbzgXXHEE9FULQcC1kHy6MK1jtfMbmjAXAw4tu08tF8vOTaaO7NL+
jsiKS7WfQR8nti2qofnXnE0ToTuAshTIpRlJYCBuzIbFYP1kJSFIFBqVeZjBoV0Y
Dk+TvfetmBjU79Rq3Xi7tZLtsAnuFqtCcnPptkJF0LZakTrDApK3uxjxWXVuMWip
/M90lxOxMZmBy7iN+C2sNFI50nhIM7pYgp4iW9h+hEq5QS3IC4MuCXkHyHQdPF0s
cnEPHX5c5j+WqHzyBH31fpKNFM/vLfydKpOaBcP/LnFwEcmT29a0g9ThdIPFvnmf
n5ncF9lNAe4FoKNnxW1QSDdl/ZpfqDehiMIb8vB4PUwJQyfS3A9yGm9YRX+o+YDZ
+IEb3UHO53yf4LbJafNJBL/d5D4x5jh0+5qOonOcIJg27vBGg5CYcP6EazVMEQNi
IHzhLult4eXZ/nwjy7lwEi57hqfxnPf1Oi6iz/GJ4jMoQAWooIQ0zDuSAEO6KyeU
EPDeAa3kCg3OWODjsWiOxpdbrXuraV0/iQoRJpWPGmkBb0ZnSJ3qZweC9fAPrwgM
Uj5L0vwRN8mgvy9jqKVXPczo36IGTfuM370imRV3vBYS/VD99VGh3iAVuzYXRpXa
eU25byIsglyW4LFjxwYr+QHVryRkeOt6OyXEtDBs7WzbfwwnuVCE0j+d7YR/rTG3
Ud0asA74cpqIsWJ+t+44ERm8K3gQ+BUutuIwZbHB28gTff7Ki+9DU2BLaeaK/fV9
YOngFaZ3dcQWj7XvCCbSpJTJoyDIfG0usotpkpDAOeCM+j1fbBBwH+wKaFckVnmV
E+qVdoUydK1Ihnn9ejQUJlSHhTsWKn+Hygn/L1Iek0Yx8JlqpWWd04NBFcxdm2Wr
VvWKtQpmcY8lNJDwT/lUBHkxq/en0NwW6ZMmsJ6Kiku+RRd0Wy/yCsF4Q7n8St2a
hbTC8pkO65z14HkULH/mK0wyS344X52LAMJK6NlGNXsI3yu2eQ6iBs17zmdJBqwc
071Uhh3rUUejzHqHOq/+MsMfC+uv7iurnBCFcZTB6yparRnma6T/ZnMITubSaMC1
uSddGWD9DrGvyxRvp+KvgyaZ7P4XGedNrMSXz8YYa4qmW6UJTV3TV3AQGhe67OK8
FlE3oiwyseIjln19c6kyWMoRvTx3S39EKhFMibXQckTOgyCeTBcqTK4+bauC0Dtu
NpZ+KmJyc9we2Y8aBhcM+xAy1ucE4r412+/rCNKI5k9dr2nx/zYPf7agY/eb8tl8
pEj4BlnAZFrajsB7Sh6FEG5RLESDmLfdJa6brm2Ij7+P1weeIKjSxooxpHQFb62N
9cWJDqt4PWOrAPjtk0ifB+0rD0GxW+7pf1j7+owggw3mSBunLaohzRBXuPlAiN/o
jiddCEAuJ2NFLE59kx++S+Yn6I216vbG/7cDX0AgzW/vbKzDyrBwk+XTDcM0AOvG
ycOz3ObgXB2KTigXHxlVHzCkpviobDe3B8wtbMcPp+9rvC1RQfG7NcVrFuWeAOE4
b5rJ47+VvybXxChHN+9NEtz40vAU7N5aqcw+I0DitOXAwDbI0l8nsUlzJi4izhly
T+dD/boYM/fLxpF1ekBxQyq6c+b32rcgE4Inx/WZEzybThBKh1GVs9EOg3VhSHBG
rw50YyX2o4gXg/WxtR/3CenfVkM+Bu+0giYrry4MgnIbkPhoFXE5nKC7KCm2P+cg
ySLokd5V2WlONTBDsGoHQQoFXtZaoWnq/c0F2E+5rL8JEw8NFMQOm4/EH7bpo0Cb
hPk9B7AxofQOGkWL+RwCOj8V+b1rq2xkmLAzhnhgrKcZnNI6Gr4APzEVDOZPdWPh
l3vWkpZmzG1Jf4CuLj83yFLVu/kO4i3tSoznQp7tzpmiKZFvHOa4MLqfWZ81sg80
jxvHE8RdsQq68wtJBIIkTFHZXbbBzn/LXicErH5Zsc+wzCyYfLQFofO6OZWnf4Qq
E+meblALd6LcvrSNUkcRzLIWkwl4pUjt8wQiSpDGhI+hDHhExbkiLqGrkaTj5OB6
cL+SvS6eN3w1uHF3D//owCwVLK+aoeLtT0Icog9+NYQBmjhaGGTgBvQntMWI5Jrg
6UtO38xeX0FC6M3WlVWoVbsAIqqfCBxjeu/XXy0C9+jBRRz1qHJCga9YCJIuKnCE
UaeJbEkmixkBhHVOBe7mb7ndz9Wr8hsSK6pHikhxCrKXGcV2q7VkZYlcuFAGQOlc
nHy/bzQ7NPm6DiqTvCoGTjJmKyKKozIJ1exlgFVI9Ml+zSrQy5YBZJSkKNqWLsdB
3ag8WCPdr9fbu4+uO45m/fsXqzS+KiMVfcx08egwUFj4QAnxjtzc6TW6x1wILPMl
eJ3fwapRsuHZmerp01WXJgzIEslLxlDHkZa7gVCjKTqlnx7SXdzRHfit8FZiV1RN
ZnPpj8jEqGB9yvhFmvjwxVGrA/QjTXfHOUPqlCkaLrhW+0ZwOfbu2Jr7LEu34sbH
sKx+OaM9tRJTL69vpJ+6ax3XMojfu1zezxrwLTN4IKadk+MKdguEIY51+oB1yyV9
lzTRQseMlLF8a14QcnFJrd82bRPeq4iBdTaU+9SvKzXYLXxtnf+KoNNFM+uH6Woo
DGcbNqBOlOgEoQPGjVE3PKxa8SSi36ZfxLmgtaUz4XZK2z1KwhJvfMSgGJkJyxSB
VEFPZasyMF+dqBU/qOs5LBB2GioU/3dPgq9r5ljm3htuQr55GAWK2q3C2OIwSh4w
eW6NFfJF7Sa7iYrnq1WMXoKQlgoT4lT2Dqgx8pH5V3z2n4OpeByFh0QXXaPvAe6j
tjPZo9MixHhMTgvBUlF/DTOQe9EbhLl7xbGyFKSPRjj5KwL9/fO4tlNLX1vuK9je
sAKWXRcDPz3o+rnzwTg5zRTqiW3usQGoe9uaxao7IuquiLF321JOBRw7goTCLIps
QlEsWOBA3jINNsb8QCWaBfkXEz9corI7r1SmDdlFrmgVbJt2XrMRLahkBMmtv18J
vvYeeoSDTLqul90WAPTVSkPjdYiD87jcadVh8E0yx1kgVD3g3XWL6EoV9ovlgq7o
16GLPUSBLQpSuYD3alzGS7fGyc+F9TOkxdH7SI8n4nESyiTMXgQzO9gyHC/fUill
HwRwreFAmM5HwOXpHIqvEciNgMBINEeDeaOSdOAJrd6nsPcFrwL/eG9/FNJHOTD/
DhXoELHBXHRYIxTSFJLmkFpk+W6dEIZHiNJcVOkMTGceCzDOEO1D6aXwhv3SIYNB
4UKL4LU6eiMpMYkZPYDkuZyVmK4aRtJROP5xz6+4YnlsNxJWjzV/N/RUS82+0o4H
lHTwvGqXvNm5ghMCc6BO6n0AUK+pDkTnCwTWBmEKtt1N6b7OiwxapU2WRUjQsixz
lwbMdB+yu0uSy9T7GRJUpcT9crCtFyp7cm9MmlNilL9vR4u9NK8yOQLnc/pbIvEZ
kHl1g/hPkwo8ApkEQlIKni9prunWEqhf8M+2baWoslAAYk7I04dqh5E06QL+D9QV
29y+H2i9Bvdp+8f9t2n6B5EfqlsOl0H+yt1gkvB1/20jO/RLxjBlKRY0KjR6P0T+
xL6x9lz+nyK2eEx4JKOn+iN8qvrojXlpHnYct6sme5zUT7k0Ldq/bUyko9BVB8ix
qDAzSp2Vdto2LyqAXBDVfDpWV9p+E0QWstg2BMPjimtHEANiMMzAyfWrj3uVZs6G
N8YMJ5y9LnwYsbLAwE2S1XJ95UT/uUHc7aqIUO5grHdStvFTvHXWIQp6EFvdsAH8
aJK/80pwXKae3mwBGH4GBSjvxrtmmBTlCg31trYwRQh/SUMfjJPNQBq+bjV9bPZz
5m2fOtV8vnL/NpsuopTveipdIa5XvJxaMqOhzgQsDGwDSYlHbvk88/rAufZ1a93U
ggXdUuIVosBB3Y6JMnJneHiHkLHOhmJNwGSJAFG5hczksU6KGflaUImPJ/3aGPsq
GzAxncrNavTYBfBXOw3Q0NofpkOh8KBa0H7wyj6e9cp4g0kG8J/ltN08t52tnBUt
qFcVc8l6ng/o6CgjmvWX/19ImMDQl6wwxcg4PxsgttgCd3dMAw9Vr1oYQkXzRB8f
2w+sF+NIp8c+MYyJAmarYJ5F4KJZ+znoSpQwOyAcrorIL79DxFCpyFUY0Nhooh1m
FmhFz5r38s/8+5JhN1Zyd/rpYPzMoPllFa+cxtcxyDX7Djnlb76H2UhLpBs85oV8
70rMyeH5VP/0B+jqs/Kldhpxoe2PjvcTriXgh6frx5tvVkAGFUSYFM8d9vUoFXN8
/lAKh6gZmL1iXJ7rtv3vKvYqcMGzEad8j28YhHgBQmfAZUdEOG505DT13R1N+dRp
X2uKFvszqcLuXvedR2qN/fhUCAKSWyLuSYG+f+c5Mb4VGnPPXtLMgfJa8dxZ8atO
QzdU2MsHU6ZMv4nhzTCTGzKVh1IoMMLZWTNwBJ7cZljg3zUId0BBjYd64T/pDP5H
67Yvr1lUB/k0bNl1n/4gDg+J8P+nwYBf0RYsHKnFImVdg7Mdt/hdLWxm2XFmL3OB
exJ5wJ2OLRFnxjxXC+jFDmrPTXvqgfh+J+6BUU2gYDxr/p6yEihb/B+jI0GfUcDd
nQs7Hn+Xq+BoSHlqEbgZRPBZHLh85rwVKKTDCV2SmQ7xh1v9VucpMOYfRFxIy2XP
E4j0EGzbJ5SGstfNNBPtWxu3DVjRB3PUGcKDL88wFJN7gAeFPmabV5892M8YUITf
7eNkCjND3TtOJrbLNXHe2Ycmm3zk5iL3LuvChY9AXIGeGdnb5LU9Qlh9rHEDfz0o
PENSgp5jvd+GAriqQydhVLLta+rN7SKllphstCUDE2D6EY79hXGtviQM1fc8j/h7
bv0nmCBDXYQyy0bKjHhYSQ==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LpBWwA6U9bnPRYghBDq43cs1IecnRZCHzTdENrm9Ney7yqwJ1l8EYxZk5TgYx0XP
sdexB3BoLiyji3ifsjVpX4gPRtkHsOpouCQb+Wq9rLfpYcvSh0jTOHoSb33RfA0H
kodu121S1FkKdr8110XlHtiCTEDU1tfSrQ8FJouLGCE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5408)
odbV0bbmx46HmEHarot7BulKZLkYZkCD0A3EN+pmlLsTH6JQtnMf7Y3sWX0r4f6u
aREsgbL3l+DHLLtlu2ieH4RKmwKn9Rf7wS9gGsTGNYawnqi3UIvV1dQNQ3Gqch4+
d+OyPzIWvLwHP6TcMyoRX0ffhtwohPGTkUDNCWlOUmuJzxAvyCCzsX3keIl1wMrI
W9HtbKm7xL5hmSn3+zvVllK8kTy+A+An8e8brFrMnv236pNMT2eyVmQWQlpfgjDp
Lp/NDoVVKXIbAqlSgm1GTMDf+1xmcojOe+rGxb0iKRNo3LjNKOHg+8MbML/+KGB9
7JUc4WjyaZNG+vUAuPxk3ET4xLzRYtOt21O8WjlT9A9jfYlkUB1n+3YqogUpA13Y
Fem+uEcivWjHeka/Ie2cl3ZulpSJSxoFbqJjDtJypDFcdIr5QQ70MkElNJeOhDOQ
kE1bAPVnMQL8nlk59/FlwB3NwzwUp+cLNnw6OtSh/O/JGeb3xx++VE3kaxJyWlkv
DWiIudIT/f3pYnpMcE01/o1AXE9cULN6vgM6WVZDlAfBhyZQ8JJ9nms0165cUeZG
c03aPQCO7dKPjXzlCISS9R5qT75X1DD5j1RRkR+SXEQoAGaywYZdbrQGo/s/TQat
J6u2VJ0amyrOKxlfdGEpUhWX8FpAZM5R+1nGSJkioOvFYJSbFfU1qM6XF71z73qK
zXgUKPs9q+scFKQ1ap3BWvRQi/mBgNs4SnwwL955Uev4kXMIGPaGaObpOGdTcJZ9
qFzOuXUiTrd09+9DFKOSFc812q3SWWMhgOtHgQKTGgjx5PlIQ5vuXDIYyQWydkSN
mGq/LkQqBKP3Tq6UQU3pVFgnD7/OsooctESOSoPQDznQb61yGu0OZIzpikApGzW7
o5dJjI26oh1vK5OtgMseAQ1Sg1Sj/WuW6sAaMxNxMEWoN4cPr0JIZW85yH7gyNRw
C/bhU6ppv5zbX0pVnCHQXNT+4mhRuL0YJaQd85o2UY7MRsSqQalX8tlF2S5bOVmX
kM9P7i8X0PGqbP8+3EfYkzudDznt/NUF3DjUBm/gcbJYofb22rVkTUgzlvSXfrln
a87LD60BlEJVK/orZzbe91uzowWTjRjGHSUrJGUZdl4ajlpDWWFF59dBJ7Vnvl01
FZAK3vj0dQdiS39JvwX944HB5PUWApurdSejRuixOSEgUL93f0jPlx5K9UXUpatg
0XBUmGYc6lVwqAg3BvrUPOH8TdvbGNKUnsnHB3uGHENWFpt64QIx6v0FXDRQMbfD
B7/VlTaii+9urvZsbQgiHF74l41q+Dsc6gke19XmnNzN/hWzpZNmn+D+wgJQQrDu
V3aFF8UKhfTAZL+P3f7Nef/s4wD2q7FPD5aXPpMjpX6/BXVO04zHH2ZAjtOYUQzF
zKaGoL9RGqy9h06noPIz5E20l0RQMPkkxWMnijxYJ2ymp3yfhEzTZi6P5aE2VrVs
7rTOG8S+FZYfavkx+V2X8a4xO5cYtnrKjVAxVWhLChnj83uaNX+HvkIW22nQEZgX
irSxhzR20/MjW2+BMHL8kJJj7xf/jiL0WkBr21e09DIfL4Xfrr3mEIUZKzdTGcIR
jqnwSxYKTJffFMmUibQ69XKqfxlNXKrg4JlLb9p64/qiRxwqK33kgeSbnPFdvL9h
gr4J2KLbZE76N8vfrhMn2LQmC2lOp+fMv/4grSeFmP9MkTEZvVALay/vaqJsfbGO
ZAYMYCgTVi8vmU0ra1LLQtJsvgVgPdQpnZOsHD3sV3K0T98Mh95cN36xKXoTl9k2
2Xf0+oaRH6Uy8YLekQax3L901TOZEbAvvj8rD39PAxWQxA9wNvPmQWCoS61zwsqm
/EHma2YtjtgPWKrsCqOQPqBTfgWKJYPGZjw1WPMUsBQVj5tDgmj2L8xjIuQQi73x
Twuw23RteOEVodYJYdjTTL6EvUOgXk4UgNqRrj6kjWedJdMJmwrhCbafbbdqK3MP
ZejURYlGvbW6i5LwEZxWlOG46kYoEIlQuBoLCGSwXHqOKe9glb7oCj6g2o79BiHL
oI4s3PKCklyTkCGXfpL+U31htT0sdYjy7OddrXavsOEk2SqM+p//WypGMbM2EiiD
x2hoIq6uIpcmKEeTKLxTHbuw6qYy/LoG0cekjTRP+9WivJ/LLljpznsqbW6ZKAzG
fHsYoelu1X0ji8DGDCEz/nATuqlFq4TOagCi9qE0MfY9sGG0wYGs9MAApNhsZJ/R
mj7fnXNulhNQ87ztLwmEGjiCEs7ZYAKVwRYpch+FuPbSP6LICbuaGl8iqNjESZyc
lfRx6jUphs2LS+dJglLZuBofdv0Q4XcW2JzZiPyUi7NiaRMKMmkCftV19Mini6kl
4+x1P1Gegd8mhopAOpx+e+Zh1O5eB1+unRBXjjZiAXR3JL1sejrF8dhbfst2NfES
o21a9keo8lyK9KaKFFdDOrQPcs+Hr/VujnMyIiLi9SYprFvIhEDuiqBJ7BsZIgCw
aksrTQsxeTjtWcTIvqrW+Ftboss1DelwTFKC/m8U95a7AFHvkcj1fNbkU/kfz79x
udOyjM9+eTbV22TGOTV43vlVMW418tV9lYSfjAU3sRbq8vuetdl5xieZE6kFzgHn
6klu3otwGohEGX6nMuUeinE0Ola1vGLODk/IULFby2EJRsq+7WJNG7772uCmj3R9
0snCOiYc+uVw6FbcSPMIGfaacwnj2gs6LhpMy/PhcKZlTNEou9PnQPjG35YVoj6L
y68baRyVVTNMM7bPMNqgSHxIG/88sCI15ayomSUE+NtSE6QDG1gmDycVVGLy81VD
N7I4P2NF7jPh/xjL5Zxk0YuBoivhkSs88PPweIbDsDUf8StwONwBa7HtWp1GlerF
t2c1wbrQF/ZcoDZ5fmVYEM88agphbsMejxADEEXvs412dmq1HLmdZ62hnaWhQQnT
vMlkVayy1tR2D3XcazbB3j2FUvk8XAtJkqxfz/i8JfvrKbwZutgiyBWmY1nHNKFU
Gpdzh8rYQdjA8esxb+tR8VIES/eWr/ZWAmAK0F2iV04dZPtUDTD+mEfudLmT1aaT
nfH/RzJVgBUxbbP9v9PnA2CaeyMCaloI5W6iB0H10aDtMKBhChk7WYdrVsNrRKvQ
s4pmwQJFbIzpiUWInWQNcZKuJElREwSmMsnihuAV/DZ27UXaQ1PEVY6+8IPw6HZi
V3Tz/TZltfMbm82VsLW23bHIGg7TBsLVLa1EQ4UiLdOgF3zb6roin19poUTdKMDs
BZM+197s5yu4E/ImZ8I/uGRteZ8T1O3aMb2+brz2a0UMEOBEFnafagg+PpLjnwnM
7SBnnnhsk/J0SvciaBqP/suIWLrHiMsPHuW9dHfd8cMkyHwMo8mb4BlwALkJR5wq
ot8MXSHGvC92aKmcIbnBnm5VLRq6RBL3RtdgRYAEMNZtBMJC6L5tXwqmP12kudO6
nrOohS3rNuzpB8Py70HDovBORh1WE9Cv7m26Lmv995etq/kn4pzhaD16AFqvSJLV
IFRY84EkmFVXB3WN2bI+huQGZP8znnketM2pX3AKKra8Yxa57ONEE4LIippVhblB
JDmpFKwYbTs5SGIx/KZmwOOqgHmG4klfazUaaVBLL6QCqIN8T+cSLxBWt+Oe+W+6
u+Vb/Ib3z5QZR2HS/GFLewO157WLLpA5Qm4BPM2sNnNQKKGqmxBdu7YFO6ALqPza
z3yt6wlsvtqGcgKuoYMXIUj+sGDreGgkuf3UXmJ4hqc8NaVpQMtcUQmq9v+GeAwC
rwnUXYWHloGcr9GnekwwwCwffGNxu+hsMV+4hbqk8aGhX9QTDT2VuGrizgAMehJ5
djV0j6G9UmESQn7OX0qA5JjH85ENKYFVW4V3fPKTRUrMhhQiBI0dItvo35+RcARy
n0BF77tdWACKgvgCQHhwntoGu/RfhIpkfOYPDsp2AHpGFPTsMqnPrWjCAmUMAXzw
tlO1p9kgqRoyAjYIAS34njcqvJR3LYnDotVKONvwY8sj9llo/E2jD4l0MPIeSGMo
vJnn59yAfggRwgYXK9Pgzd2oMwhMTFHm4GmzEcSAgsqAe/jHAbXszLpte4txVL8P
7d5u4zMNMhCYekMxuogJGDM+u/hiNKLhndzES+391J6hpPkzNJW0WFFouS7TjN3N
m6s4qiI8dljaUkBrm0+NsUSl9WUfSUR3EXKKeYR8waQH8COBbTPVf0ajEacA3cyY
BGHAJiGTm4icNQ6R012O2tB5g91TpZc/v/jRFKDPXFU6dFhe3B7VIlYVnOCWAsTv
Uz1wmpVowoZIkMxKhBQe+V3bT1oAtib5fYIDf8UZTmLhvIyd8GSquGwLIifQC3F1
m4wB4xJCmbYvVl3oVaMZrBB0kqyEwjGs5XlpX5AOX8Xf5yR1i4cA7SNaYnP/WumW
EUjkci7pISkvsfGBX2MgYTV5nfd0ipGytPgQSrXZoRAnUghmpWN3X0y0S3O7jjKy
mQEUuK8vi/6ajS25Zt2Rv/3stSX6o+kZyadbkDI1d8eXV1xv0q3mbl8iyW6K1uc3
tOyzk0+jeIpQAHLQmgFe6OxZ9iDdBsNbQrDO28Fh3uHmpau9v+Fx+vK6JZU38GIm
CH+9Wib1o/RIvlDzFnIl9+UsfLbR9tVmpNckN06UQmrlnG04D6pAcBEtBxivccrK
a9en5KSzISEvM/iRDBc3PR3lWCxMpzdJdNsXyFUPZvUxk9+E7OD6vwnqK2SH8JZl
MRHGDLr6jtieAJPstOAcJeEAjk0Oyn5TW4PT87Q5jj1D5PeUDPhcaxMJA4cr0huT
znFrT5KsTOPQGdkS0YjBbeGXYXscsVCljCx3N04KgqQ95DkIDf4wW9Z5oH/tOSPq
w2CALgnbOWsoeEfCrOPORe8z7EKh1NQC53QBuXDap4Wzigo0xixlTebwxi9JikOo
Ff5SBnN6+sWa37xPsFK3NNNXrqRo2RaaMF2t1OsOH+Zk7FSF4yOBcd852KuxqBY5
35XftnzbqB/7GtXxsc6q9T5K/N1otBsD1tuaTVZFMT6trlWkrypoWnizZe/ztf8M
uWIrqbI5dxjU9NnduEXZ+hHiI0Ltgp/eZ0pn8totMsFVZggCaQe3wbHB8lfP30ja
eDx80LkJMF3GhmVb2E8Ot0A09aecKYO0bfNOa2JjxcUEaxxMNj/cTaFHCHXXUr7I
aFNWNFlcmz0TDWqYIDwuMqZ7mcFP5hHk1GRZl2H789B33is9ejikSfn04BMj+EjH
fcWkYr2voYP8ms4cNQltXyNjQkhxNeuDypyfsZlVoO+Iogi+wdSyBre+GVL4nII+
mN7XlHxxZrJ3igQJk2XPt8h68Lvgr8Ac1l2m5LrE7WJ+19G8rDOEWiAUZxTyXKjq
CQ2Cjn0ZNIs5dIrPlaPULbA21Fz+OnRHGjMTo2214BPL9drp9Q+pd8CaSIgu2GfJ
8h93xPKrCOeiTrtuvY5CRtmyqG3LaQbXEnK/3iCy/ZvkJniw2mb1N6uk+Q18Am/R
quiL0RkkW5eveerOhWHjCDnfwrt32pBuneSjD+1v1Dd7PcE9P4/SqIJjjhoP2tZ9
CNxKrrpaXoO9esd/ZyQzv7HE+yGgW64iWLgGdq6Ja+2ti9/deE5Utx0tuSdp3AfZ
zkzCheb24zwkAw+An4cuXVZuo+589dweRWCFgESPEj26HxW3BPilHvP6RiLdgXe7
jX3K22LlumHkRU6F9Z+2vBkhLaOG7u2UtfHEMDzcjTVig1EBzmB/izUyp/rfViqG
2IAtRMwS1d4vap6Bw8SMCSbLZiwSZ7ajACzz3+AsNpxiqj9LyoQacC7kwcXth52c
YwUDlrBXnIL3rSabThBtoPTIRoBy2vyHoJ2C+3wMfyVL3aDmvoLGP8V+efwg/Wuf
t9EKItKh6B1I1oEdQjgpENvABhh3ftxtopqyMQFXvqPg+yrIsTnHCGxGyOryiaYM
28JuuQXDrVLrhEOF1W4UVrojCOKS1VjGwFR+TIj4GPxyoT0tcGGQ4gfA3MYurwr6
2J555Py63wyLaOg4Qq2BqFhogMQoxwNxXwJqcK+GHHy7Qd643KMj6NbTbfzO6UV9
MQaL2OVcLgQxg73RJmwJGOwy04pdRfW2PFA5qCXd3AdNlTCOR+Fwa08Yas313XEf
SNWnPLv/oV5SJaYf8wxNTLeS79prnUrH76VczE+6LgYr/Ed1+nXsZl2cErSCBzfP
VSefn68j2vz0XpEDAeLCkQ+EIbf2MnvvA6v4up8C+xTyD/8d2XEbWgtQxhRZRVct
bZHvWO4IQJibG93rozS2mxwweHQmNICkLUsI71el1lpit7wZB33XZ2cOS74cC9Hr
z5JBmaiiqBC66c4z9sgCpPhAEyu1t8MUDOmuGZExwQ+DgCVO7pRCyTnjm9IQD6oA
EU6i3xhYXlu/pxerkw0VgP35cykLTwlt53bbgjkGPJth7km/35p0vpH9YrqtRwpl
svnixCfaHYYwjkZ07Ac41VXT5JElJ3lKnFGhJWJjbs8kJb+/lkWyxp1W11AoJTt5
A6KfHmQctFYQUbq+MU1Stme0PkbFZ7qbHxgziEyOoQD+QYdT0Uy/bk7Vcr3nROmR
kRnMU6nWs1omm8rfeC9oV0A3WYOZ1P/T6yXG46cpIEaOF56o7SHfgq0dIVkLr1r4
5n+THESD96+PJTmFBHjUzUSi9vKGdeqR3IckYqvdfO5ROToDrFI7eDRE1mhV02oR
XHqynQwICxMXnGq3HpXClDN6rMGgCBWOq9zMByZb4QVshwkN/ET/l4JNOIUw7yxJ
llk+tnd2dNxqbZblaN2ar4+oPDqeRLT40o1Z85mNzaqgctyGMfdtkTkBgY02ffHZ
VrbQnk0AsDROHRKnBq7rgaHux0diLILxofDQhGloUIJnhjQ5MYz3tuJk8d/y96I9
RdE6TYPiWUdKoQ8dwkG5ewUh+VVgyIQy/n7CTJQH2pFWVCj4L/7BGlEUbIE5/v1I
nO81+dMPYMBq3FfeNO7X0j0Z3wqnkTHSEUYrGhiAaTtU7dB7WQzBySB5WpYFExq9
jDExMYj0Tf9NJW2xPekWp/Hs9sSYei2OldI42rPinGFp86Ho79OTDKQLXUEEd0+X
teIvfMAigumfHF4YioikJSC2oK5yBKXWPPAVuTJ+FGOz9UO5QiaKZD/dGuf9xQbT
iLKeWlSzS2gkPQluKM6egfOK6IJYHXpefNXQKwQZJ7Q=
`pragma protect end_protected

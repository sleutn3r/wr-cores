// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
U8Vzj3F/Qo3QJUD2pms+ebzCFB6nHdZuTbDqzikh04EJtE1afxF/n6PqJQWcNneV
O/z2PxqITLntqUhmdPvmHs1rrXwFo08WUi0GU9tx0OVZyZjvoKtXkskdyogB29+7
pbYTpD5qof072EqwSiOIK/b7Opknk8bu065xI5ZTfuQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11072)
VV1+oTJ9zKctNqx8iX9K5ZwX7CYR1ie8NEGohM75GoUIW2PJHf3v+eCwvl9wu+Rl
fZal1cKj7+I243Jk40DFtUVQJc3gmw0zNPhX1TdVCy17WenQUr4hJgDBMJQ3S1J7
IMhDBzq5Ugc2fKW6EAlJ91bx+njNQsjzjsVFE3YOtdyYoSplegFysG8f5ymfFRDf
oz+KRbDri86gLWPzUe2j87WjQFdkjKLpnkuocd40h7gQ+FygYlHlltEseE494pMy
xIv2q1+xLnhrZFi2Am12jjsFbZZnvto1up2pxDCfBtWhlvuxlqQsWK5Bve2NxRZ/
/Rm9is/j92NS4JRnbYaXGIQ8rrWWnlxBsf17tnWfj6iob2lr/0glsvSxPj7aDouL
xZ2QNL6qJ8Z+BfT1DNCdF1GGExthOZTv1HrbH3kDYjccI3Qee5pJqMPOAPkYswKQ
hc4K767IMdRzD4n/cjjcEJM+0LvMz8BcCbxoVjY7cKGlOUH8HNvwFrVcH29126ty
mCYiUkkfQIiTapcZQl4vXhamHdOU9izLu8pK8HVngOuUFP3NJ4rm5R5HYfZkSDYl
+hjWlFaPWMFnE66c79IEwsyofbm0oNXNkhVF7+0PjvQXEoV1hae3Gj27u0h5viwT
noQgpqvkVGj7TLV1NQtvg4jUaNcQKCIbf1svUXYzr/1T0mFihp+fahWeRwX93tWa
xvg+MNG6W0ZHjRE38EHRUpWOCkBtGzonCLkCZBKb6WjynU2eTBqVqIZArx7wOCVP
7Ws+dVuazLQkurGhS8l9RvsoRbcEmK/fMoC5TPB1BcieJISC9psfy8HBPi4jGfWn
VnoqnhH/1J9JXUTrOtxFDMYmsA6efywN3mdmEah+dQ1KrJIKaA0gm8rMVfJhJvS4
qNmRjreBDMIufKDL9G/Fs4obgYwr7eG/hBHB6RrS9VGz9h82yjVHM0MhpbP6WO2R
YqtHLQa2oER06sg99y5qUCyv6W3y+n7l6ZiKCNsakBL9i1dPe9w/koEgboLPv9w+
EvWHS0G95fDfaUlY9GVAuBJZ0EFWFALS53oGag0mWABXPGgVGoaTkSKS2asdBvcw
IqH49poYpAnNpqkFntxwtC8Uu9WMNd3mpH+qjzS/dPBOLBWf5CIFEOpXZl8oNgIT
3Qp98AJSrSin0U6aW8z6nY+VZ5wfYRCLDo7dm4B4Xe8V6h32m4FnbbinFQPU4Xz2
CXnJTrxLln3Eumf6S+IlXYhWRLb0JvLpdsEvw6M3/36hu2+06kIn7duTGX1jNwXt
jGzsvW4c6WyTedi8nTEK/7E2QZXVNKC2yjb0JHZY7vdjXT2ePCCE9601354v2s8e
6Glo7Z0ltRNjo1S6FJQE0RR3TdIS7OIzYs3OczFjWJVFylIVm/Rge/9YCmejVwyo
HHHFw8uwdOB1euwla025Y++rGKCNA3KbRzdkux5vJy0eS2RnlKUfHcJMGJm4mHHu
DYoB6wifJvc5WJfK8W6RFEnCCcd1SCuNC2yuY2QgO573gRx60do1nBcg1d+QseSG
N4eXeizub5ftGSst0xEkVQO/+mDu/4z5+M4/35/HLg+pBco8746okXYcTecBNvmH
dgSdqC5/cJhj6INNHb+0ZmfpNnR5WtS3jZTSovMTy0+VF5Lx95eKnKZhPekMOzpd
DFOlKa46nWrhDnW1gmP98jW6yzsXigoWeoJiOGVGXHyMy8E47OehCL767d6alYL/
5Jf8mrO8Sdt9rwo75JxpmPcF7Qzk/0d9a8Pfr5AThzkwKcX1PMuP5K22Dj5RVoFu
wwp+87+u0pFJg2oYfF0vkCmEwta4uw5fV0y977vKhzN/iL2FjrAjsA2jWT84u4cK
0aL0bhbvTq1KPPFl1p4zAqtisKzWnbu72UxxMcdU9u6Y75I4Z90l5j4TIJ455hWB
BKln+7AN7MuzFHTIQxOWKryP3iqqxwYP4u5t8RsZtqS01ze8bjfARhxUaZqciBeO
IgfjHZwYRbBrQSJj5m7WiaVwjh6tKPDc7IJSpBSAiwUJ6ARHIf6RGKxs6ms9v65S
oIouiEgPvyyJY6zv983Sv3pJGj6k1iFlZkm3NlRmBd0tSLpp0hoq8IprrMFQz66k
5ZojdExu43riAWEqNJ12ofd+vRft6ZQjvtvuG+zjwjaAJ4xhbPy18jiXHO8/MwWR
3R9/hxycY7vSb3dkYcT7iZ8W5Dzu/5DwwdrI3UZoFeo/5k5cIecvwVaF+Gosll3V
j4nHKyCMJ/gBiRQXDOwlGIXhlOnqH/Hs5urTk1thbTIDKOAh1w+MvmB53ofusLm4
2LsemOWroZb5LYCgKCWKZs9YZbyUTz7zAMjnpDcbfQMgqI9Uu9ZsEKwR0ByA9r5G
/wcpmvR4kLpJ/iyHt3b26xHLet+1oeqgzqT4lUpobABb9ZxZl/qLMhP2m1sTXPK7
1VbO76KxBgT5SiP4wYJqCLFiMqqWM+Ev1QH9Ebocq6m1RQl6qzx40CxhPmYSZvrr
ChIKcQmYOLOrjlOOedJIpZhlyuwBhvw6DfXeQGZ7m/6Cx0Ktma9zIBsTrP0l33rR
YLNjV8TM2u/XZpV9Q0UDpEmaoeyfbJ2Vu1WqXuviJdivlqPmVkJenMAnLsCYfxKL
ztCnINheZEAIhOubUem3b+xbtI6g7NG1gv4LouvhX9qnM0a4oRYgEAidU1KjvOUc
i0fffKVKq3OSAjubUqoetHIpT190z9l3vRVQwVEXdDcs0k1NIrxIUaDt24b7wD4R
Y8PQi9XZS/vuK+bSlnf7CVfV6D5kktWGL9BRgLST5ih0T1UhbR3e4APVAaRWSgUN
yp1QqyxNTVjqmAm43cPxGeJzBp14ts4n1Loq+VFjTVuKxbiALG+iQOgIZNJpt9jo
SMvbsVxJ7vp7fCKBU8dK6I4F5HDfEMoCZkdmRRpZBaZ1lFJ/KM7FL19fL31PNTtS
dSZ8vVUU8rPMXtkxY+xkL6RwnUrm0br+wMYLCPuZruInMZJFtjYlx9sesQ7LP8Es
X1iAi7S9oKz5KNb5JCTS/1N6aeiHx9gIPdd7wMsznTgsoHuZTkjbwmWc1jffzVcy
exMCYH/81ALNUdawd29lIzqALnXTrAEI8zYLFZI14VdH4IAXNevxD8+kHv9dp85G
xZM7GvlB05V4bHBtjU22FLZsj1XMQmqiaRE2R/sH7l1Nn7LQU8tc1sd1MKAkXluM
Fa5peiok5+0wguUtsEgQCUzJ6YK+Y9qpc/UVKDX1rDfM734MWh8RtXSrn+e99OsR
1x2qEL2yeUUV47Mo9hUlvKlQWuDe1RWGyzfX06dljf7CqogXBd6AW7k2U5zAZKhW
eqPu2Tymv5lzadEgE+ACRByx+ebvJqcwb3xlCmVitTB9whKLhYFCPlgX4HlyIX5N
3cxFyoG+YYHd+iI1MgNfeB5+FwK2zfOdeRf7t6B/9v4T4Xx+mREBxzj6TPXTILLB
2SVyFW5Uyqrigk2DJR/LXyHc35v/vnIeMRwRV3apuDb1lG/0WbRniThZJzQfv6/b
bTCrbASw8oCaFAGTBON0DwOZroVoqzrRmLk1s3U1BBFGi41n2dSDOyMAkKOpFED4
C1MNGek3gggOm+BVr/Xm27GKhbTW8/N0uctn3LsjgIyj3yyejegClV0K3cV2RoCS
o3+EGCAT2ziicYB9Yxkt8P1uc3Vv287jI+d+acQZ5bNRseAVjvsGHYZ0kbtxDaL0
LzgHef4HO1Z6cbf82jl1Z2t/qndxHB4jd5O/Iycm0+OH5arUjzm820fdXSpI5B4Y
DWjNEWMxfRWLwRihYO1YKxTd1BKAV1duK1eLah5u9j3Z+6VGI+VUJHMfiGUF+JYa
DQm/yyY2rxvAs7aV7xHmQK+pp3WrpNmAMGnxLbZpihX8T6APaiPB6zQg2rymNaEs
5/tD37tVNIPELcUXdGkTd6DKRfRWpAzwZ6R2dlXJLAH5G73iZ9N45XpTxF6Mri0I
QF9Cf48wgRQCiEAFVwfttbEFfHBXJRvs4lYDqAQ1Y6Txfdtwi9auV9K+/d8dsVIT
h50FLYX7hHIwQqlZcMIcif4f0IMw62N+swella/eFyCu3JdtvKuJ2Qw+dHJB8c5+
A+Tdy9fqxfZVwsKRl+Cug5xg8dEyXCl+9AitaRGm1mnt35ryPWR5V5tcu4x1q8H9
qeQzQRj0nR4FquyzSho2B3p1vIZySUTfxL5tQbt9/90+Lk1E2igQDkVtS/UkqSlv
sEJgFTcNHrsRvIPrPbPF172kVv4YjRltZbZfEdyBN6Fc5e0mu/Eh9SHoe+XUxIXH
fBNvhgAJ73BjHIFJAhK87g9SVDSHuRGVX7ffoe5ig9nR4VtKZjtYRpHI+N/KlJWS
JJJfHd4h3BMoyx4JMSzmtpZ3hJr6QC9hv3LhZhGuiD2YMLVM9n9yGe+EWnPMRd0U
VjR7UCjcDnO/C7hoG4gPpbzsXBxu1LLwJQiA04h4Kjdlciq073maUuTHVJpAzvLW
comdLSC3aJsLmbWCBOubh7mofQUJq3454cyynNyBpV9WzQLbHDn6ka6iCRRdtjVg
st9iouYIlIBDsoYS9B4ekYQdnMxPvdwSs56VkxBdg7rUFyGhu6bRhI8tmaOqP8Qb
VJOrDpiCFmFGHHnG6obVUfVPX2UujRlzBD6SL4hGVt4VKU7k+v3J0P/EQgqneTJp
2el40xbEk73jjuuM8PrZ3b/EqIgaJYlqsAdcVehFQBPx926V/Vytam8oSyHo25SC
BaizZYMEa2Id97CC9hgbD9laCcZPF7KSeJShMPwZwZsIsTXzSTz+XhNhM9rwM6Uf
JPXLJZ4TBmwCg5dg8kIuvyY/6joEW0O03uCNTRzN3tarFCnWqHVsOj4eVPKERCrO
ZR4etwaHQ3DQah2DP5oVL1TjZhmcu/qSN/ruSo2g4EgAzdHtE8hExIuwuQNQotqm
iyXwjxPjTT3CmPcgTHo3p5uTVEFtQ8ElSYf+BR86c4VArP+P6YFCoyHScFEq7Nyi
c3kYLsLIF+gCNBve8mdsjL3zbtoMKjXao7KLATR9vLmX1KTwfuXLl2AUfEleU6aE
VFCfKH2dZCyokvjgDgLpiCNgWTvQ4ttkXOjGFkNNpI1mNebJ8Gn0cU96ndnOJZRa
dh1dOexG30zkSDtEJyqisIFqQ6LCAmchcusKw9v/T3b5Xryql/alRi+iAfwQDWMf
YKRCzuLZ7zEDoyFWuHW3JPWKkBkkF/+5jL0VUGI4EOhozpkbigYTAQV8d3rgewyI
nx7TwgyHqdj86aJs1GxDvLE+BaE2ESbDCg5n3AroInS3qKORKXOhnDfDpUo1wHVt
sx7r+jB+RJeQ/bTN9GtuE7uWa4zzOA3NHdtdMUf0Yx+EgOJ3BtXnuCHCMpU+Zkwt
E736bjoe/QdjVgUar5nO0KPU0XDo0KbUJ1UPF/BezbUkwEsbKbNwhwji5SvMk906
BH+s0lPsCTg82gWSI35ooy2AlZ+Lx8W+AJ9p/zT8TAul01Wga4S0/bbYhgC8yAj/
ooJAWyf/9TNrA4dVxSoIbGvpHUMIy/+4am3mhl4R2175kZwb6Dzy5NDIbAD2Ppe/
OP7YZaAUj93qG5hD1DbGRFnVEO6cpeJ3oLKRjueL0zb8PCLcXTv5rqSJ8BwFWVn7
gJpmXu2GHEdQ7ZOrvNtM9kbwy2PJKjhuePCZV+53s4qGsTL/Xs/S6IIao6tgLNpe
Sdmrneyoc3kEnBfpAED8cpB3lmqjBQvnXB5bY7cvl+NPEdi2L7u9yiwulJjs/3ax
XNTC13PqURwkapsvgui+d0XlTPvENY4mWS9FcflIJUWA3g8cRmPqxunQD0ZP07ba
2P+Pq7ef2idYZv2kme5n6TV37fnfWFkvaRE2dC3uwE9IXhaZ1is+Xtoupm2XE0X+
i5w8FFsMRejEwwOTRNxGMrp/NKNRptGzL47pBezExTP+jS+7yo4e2VzDnTKTV25/
52JDAQm5cKLHnO+JRiYAJmuNu7YWRyP7Of/8ku2fzMfnR0s3a+2hrSUhqnOJ+Rpw
zxIurdZevwRMCGFbtv2rmjL+XbTw/aczhlQQz/+PJQ2M5VLMbCJ2eyYFk43RE5Wm
VWwarr9hMoRUydpLfF3rQzVdIB9rqBikXugbd/ZkSzPnVdfe8t73JXWBVawyL3uC
LXEYaQx0mTm6Lhws/nufZsn2y4lP438SdpEBzEYG29U97QrLjNh7wUS61O0UEL32
mS4YCTpyzgCer7m55b/6I6HJR4rzcuiuM1tCNQgyuR/TFKEbK73L0bgP/kFiIYoD
kMrGi0AKJ6EkikEJDk3pr2rEeK01a42kcVVVDSHqCnhMGtGcqzN06L75Debp3R2H
qQJdP0kBo/aCWMBFcyGpiZ4Xnk0cZ5SevybKMYp15E3Iyk1mj6TIpWxapQG8E7B4
OXv6qidq6BZU9nggyj4+jFmv7F/WkezTsT5dygVkvH9zqGd8EbiIpwwtl80j8Jgo
NCNslSqlXBXU/wppMnsupvQz/QAjmbO7iMd0ROmacAo5RHfXWZmWySvyD3EY+Btn
UFocDEaFTo0HpTeRLD2spxE1r0pcabM9F81N+zSGePMgeWqXIfxVUtofXvVs7R40
BWbYMkpm0s6FeygwvmNQgWWYA+gWV/RyV3S0S+mxK10Dtiicfegnjb6sQHYomGdc
U/f/AEmqtQBKHGoxnsS/MeNf/kjywaa1XLxhFt99l4mmD7q9IacdHD+39BDJibAu
AnZ78tu/DrVMzmxhVfnpgM9Qt1+/uKfUZYLLRiMB9m19NlGgaThghgNAmEQJKLh8
b9O1xL4vN1X1dFbVwfpl3y5wEZF9ca6N271mxDLKHjrndLQPNTrE91kl/ZXLsuuJ
W1KVdJgnpB+AwFsZblakjku5qmLCw5ZzvlNKXc/K3Yd8D6frRXKX/en2+h4f4Rh3
Rqq7ylmDGZ2czpu3lyFqTBJ8zCzMPUUD5QDe+7oeGWERp7jWgkHi7WkeVWagqmDP
9OCbMaBGgbriAqn2W/TOoohbWrWBw/Hj6F9wiQZpDkAJjkVeQyJ8JsCVKcSCkAp1
VoSyrbhNBmIKFPd61NUYF172VjjSZmF16/wRvlheHxMFUcFS3nmJ56k/iuo4QRMS
T2E55Oq8B+Ken4zogQYofN++GcTxK3jgjJsRjXugf7YMzS+v4ptpXq2j2ywbSokk
sZFRQFtwoD+5NpmtcX8WnO5arIAjSW4NijTrL5FtI24WGJJl9P3mchUgkSRickZG
Mq3cZKYa02aPSfjwr1cFQlpEo/jnO7wkbHcmzBm4/Dng5fmWto/n/+53wwMUptsU
6yYi8XIIQPJUtnHhTq9UuL5XOFQT9hpzMe7vdXbXTfas/nFrTr4PXAgV2GyBgcMb
k0SEVZZu6ZeDxTeQSjD7J/pStFgEu9MMhq5icpMczkToPgRH5xustSwkliHSses8
y+pUO6wYjDtLj8Mcf2Jv3W8m1r/nwi2Bt5KAmHRBh5huQTx80yg76HIk0JRm9x8X
Sm0+SrHW1jsK/ssv3hSUd6FBa3lNvLwSVoBR3jml9h/KaqO37lm7y79UhAT1dV0y
/vRnPdFHgFaGFhGIhM4mMzLWHs/qIsxN/aIacsGvfeC+Ndwc+4TpNwQe1SDlRX8e
pzCQ76xoMTvRqFTslSpToOGtwIW8KtMwj0ldUER5Ivuke+TWHhBWA/S/nELu39Qo
YsZUyn9+N2IjXyCwFfno4OmZrdjBVexYIomIg+13Ghkjx2DcV4gXhDPFVPayvJai
g4QbVoRHFIka6ozlvs68UJOvFCUR8P3cFNwbMVABpggOXqPJwpvn27G/mt3YQA70
hKNXn501clm5zfNdYPtK8a06cV7Cwz0QRG0clq9JFsCqULawUzisi7eeeRI4lrMi
/q0wPoFaeDxKOqDp/hAh4c5OThv7+LfCSkaa7dl5RC6/IBrudv/GspmoxqEX0c88
IVegiJyGMY2R3aZMphKnIO7/OT+GypEEnxpw5ioL/6ouiL4eIILv9DjhwhzUbl8t
QNmYuvPwM8a7ApfT4mUU1CEmuo61mRvaVfUYR5UH5oS+buUpmDwvsagAE/4xxt9R
Qwwe9CpHNqlFFv+WPNDTUZIUUBdWROWKsRNjYO1E/Z4tp8oQrsMaN2npvqKEoV4V
wBvfvlCSWOD0M+Hu0I+161637D5njWw2qwP6+TQ8DZJsQPq2LZhCcFlx4yrfY8/d
1CAx/RKfr0zc/09ym5cPvJdzStiMsXMjqQxGIUm6FxfmDlr3YzwnM9heOr6modtd
2HHXTrHS8MOAy3u1FCQKhiYuj2JOAL/liEh6Iobp1U1/ev1tPHYG7HIZWyIOCGAJ
Kt3KuWBKeo/Aj56eSmGMj9X5OfCvyAF1bJbCzMqFypqE4ODvJ3kQqdfyCk/0vAMr
trQ0QJltAWpfWZ6XfvFIXUBKLDzg2JfTslqA/VHleWqO5H1vvgHy6vkFDkTrW6R0
OCVxCseswcNpGju6+P2NGavN1PA1B2PRLDKga+M5MCzUIZdUchJwaXmHpR+GtWJ4
c8SrJOZS8ByG9hfSE7oWsxtgfr0reCcL/LzQBhLS+FCfI6f6zJvI5EVZoIqvdOXU
cIkaablW+l+aUOK7rhQcEgvTL7OvAVsZdQiZjj9uukkbwjygdB0vlRdL5WlmM+KC
trDOdO3/quRJDqYujrzGirz6T1OOV/IQKcsqXjm5AuqlYImUvDh25bLLtnbD1+2P
Ky5/nu39HJ7VD50NuuZWBZmLz3/db4NGzw4SudHqFx19S30agvDBtcJ9zApiJhfc
Rf87IgDLJuuu8tXAZ4fqwC5FPyAFWLqnM1m9GEb8YwzubzIyI4stnnGjlegx+C7N
8as5QBbAypzUqgg7UE9aL2ckoUU16mLlSt1GLngLUAN7WuhVkE3u3wQN/LvnuF/y
ZVx3X61bdfZX07rtJM6Os+Sn7ktdtgZNJiNpKeOVYBuSD/OkZCJPOYcsU0lY00I0
UU5KIYvt5gfFbiN4e7Qw9uHa82trK+2QTraNBxo9yUGyn76y5mNj6ndFDgDalw5B
rNN5kEfJMn2sPmiFkEqIn/Mk8IgJJeyo6l8i/AgkiXaoPj9iESDr88r77eQUmPS5
NEjx96nr5jcqqD68hnTkQl0S4D2cA+ygsEZVSlJ+H37v/bfJ1rwdUjUWoZ3SdTmd
FjTBHy/RrdsB7FDylk6vMlZX67RqBeS9muba6oy3Ek1lpN2Ju+0pMvsKVFRnWM63
oQVwbGWWWrn0aBwxI8LceHRHG4MH0OMM3yANzeQPGrHewoyCozAXYQ4J9TfSBz8Y
Mm8C5x3RI0BlxuvL7BM0VFmkkWa/fW4F4vWLgeGJmQpGGgt79w4v7GT9/9MdYXqT
ZUtXjMic3yr0xyZz361RVaqXG5Age+efmUz4zc/jgdebXi5zVmgxbM+avVPpHJuK
Oota8OzUsQoEvJIpBGwtQAiTmq10K2VK1GZRzIOUA4IJXv57CEp6Ud6wLrm/dOdS
cgzBftreE4wMzSSeXvsdPJVuf0z/VRe3VNZ6JttyiDb32VOpQxOwW1q2n9ObYLab
JM2ykXkkcDSIuO+1+wglwHCpJDhnncuvKLiiWmqF+kp5/xtMw+sLTMYfIPT8wH2r
lbsK8ub+LlATkoaJnizda0Am34ngsIyxsSCt1YI176zy6tiLSXUn06q10p76y64V
KPUSJirbiAOLL/4qhdqp0X8IojoCJk9iM8Mq6gRH5QSTyOLnCLorTcudrERudch2
3JHugbw+unM02TB+5cgRT9oMl6Co7sEm7cYuQsXVs+wuT6IMD8vhOkhixFxrCTgw
fV2hPj12BBzmJny1tR6G3tFSbosk3C9RDJ1YrbT2cMF7eVjf4ekyuOyfF8g1uTnF
xim42zOrd9fQqglzAsNEgj7+baTSKDYZUDRZDqvB2MtaQgnQu1y1TkLQ9IdrYxmJ
hI/3VJbc/xlL6cJpOxZwKl2Y0JQQ7djJCZ1rjp8qY1Bm9Jg4xoeMs8CB4CKXE+WE
I2RtystUumdt2MNepAZ83nf6C2OjpxmbL2WeqkHGYN3xv1LR/pD8KUQDNJe9kFRw
KekMjs/81gweKw3CG6t4IN6qQEZ7WDYE8lTHyzCByqxPZzuJijaAkBuNJAawg7gI
vEFnbRnXTr2OAGtdZfJGsaaOj+WHFJn5AMtuGBeyhntrETlNnI9mS5ylSbAWHbtf
DFSJyI0KiNx7e8GJDrB7W+twLSasETTnay4AS8DyK88X9ZKceDCen5O374lHP/eP
vn6l07TPf88b5IUDljB58U8R5LocdIcyLZRcIhyHBe5KeHk1SFvAtx9hdGJITCAx
ULPH6iNJ18xgfT/eJr7qzwlQ3OpNWgFI5/p3AAp+M5cmP89OzL4PylZI5Qw/b3wM
36Is1GLg3ivVqaW0L8Qqkzvp6ZRsDTLX2xGPcef8KVnIHBhsLKlpQQy217sB9QTh
1z5wB78SsEx606KLM9aJmJ75PkytnFQbtDZQCYJywUCHugla2/eKGw6RYsyRXW7v
cNNAgDeVsIMx/MtX0d+X+dEGeYOcJw/agnQzXLYGKbgnHd9dQJOCumt8ffoAVSFL
r571oxuMB/m72wFILbPWBYI+DoXOgTNgKeg9WvrabmxfbEc+yaywYlOlYHhIMcgn
mhHaorVmqGb82Y8dlKNLjs9mFGQiDAQ7a8lCRyi3bS7tXNPpl4Wyk255EdR52BXS
cMSd8xdnS4YvNEiPOtX72eC8hIRaZV/j45Kt7TUt/YTSSwtcHHU9dJHqFKLggUJv
NxlPuHDf0swuGkisqoF5oGCDkxrXIbkOdzRyFVtCe+KRLMDttJ1YnzZ/6rHX5twv
BjXdEutenRqX9sXq29iWogizWkJEFBPsWGmQ65B7zyuuRr5e7W2hB215BAZit3rs
cjadn+sMq+BjGowqQtgwmKZZQbVkNPvIDgEuIagdS6MwGxWRRNHyh0UjlQ2n5xGN
+NKfAaVXho8uhEjLbEVbsxlgl6EqhcsRbYkvD0ktnoe2FrdqUzYuJsh+xoA79Zdm
qUJBRw8SxNNucXrXWi+TFqpS4uwFvDJkgEDHHLzCsla/bDUH3nRf+E2kCUiIr4QY
MiKX0uw4jHWNHt1i4jiU96NBDSuav+q6zugntXEeQuuqkzr0XT7c6VfGdMkROaJ5
eHUaoFxovCppqv0MyAV6a9iTNKWx4J0suutWVxDRhdoQ/UapbL9mZA68bEKWpTR+
F12OwEFkuBfeM8PmZVgF/o/+id0/InElHGTYESVr/fVdl1fEwpL6HEqWTx7NkOW6
Vou7UFbg6I1am7sDnLscdtSBicCPcgtWTC5hWJc0WAqN/vFo/TC1bnoGtnjp8JCi
RnQoHtyCDGOH/5Oj8SW2QS/B2uwBRoZWz5HRxIfQ+DXQtjRzlQ49t8u8pcnSbpUH
eh4W4lurXyQUf5g+HfouqLwx6FgDS3Z89IhAARGs50VoWcbdsFyrStpROeafsT1I
AJOrN1RWaO0SuBqabfg4DcBiPz+7IK85zxznOzxso5n54l471IxkjPG/VkFojc0t
kDzTlglOMDRz7eLHmi6+Ss8FKDGGYad7OEK4dskRpX8EhXrtD0DktDAsYp0yZfoD
j9eytDEF8rZ6RXvI4FcRr6g9SATiRVjp/6TdeodHv4pjzYANnvAYg6ayIhRbT3XB
OPhaWT9awRcU45QNVFREvWow2ryeyxlduXDrIabWDM7bwuR+ubSBBQAPZEJpYQW2
meborSXCeDT6483I/I6/TI3+aXVzQjjE/uRxupdRCuH6dbYJOrhuobDtMVEdNTvl
8soCVX6kO0VwQEAIKCDTEWEEWmAo3V5FIEYRuwPw2zp0AoJAAbEUArERkdHtLwL2
naGJsRXGIiHQLHycWCGnb2hVbobW9I77lijum0DAmkkgs3x7rXF3qZcHccEZj+h2
J1ZD9O4WQg0/MkArS2Hcm6EVnkNNvEMGYuB+WI1j6d4m/QeRmAP/DwmOaLBXOtJS
OBxK6KHMayAnBoJpdSynGihfFc33xOF8d8HvN2pwhoOAEGxvH+oKEsAvGmxGMNCz
WIl3nLfhmHOMPhW16/c0ZXT37uOIO251tiTLbpx7B57nCSoyxS7oNDWrlk+ExsAv
yOBSLfFCCiQea/4VpB+E8o+5BobjdciMeZ2Zirg/edtRpieVyx82g8m3F2RYz3QQ
VJ6mu11Bhx+CjimtIpDYRjtXZRE3o4GoxLNr8VZgRW8bmA0dj7fnuGTmf/T8x2wo
m/GmqroYJlgW4koXUHcttQPYS2I6pr6aaHb7BiH60hLbJBGINuu83d8zR854xRaG
HDsNgObk5kmCQqOhVxQj2UtEWI4a5WI5bcrvoMKmwevN5gZKtDYUTAnDMeNbtiUD
slz3MMUxFLO3/owFjjCiNlh46SF+pKYzCAAkjDkCZqqqGrLM36j2rP20RuDLb9yU
qDe98XBIm7KhRtJbPc4740sbGFFJlZmGQToM9w5HUQ59SehFPzDIdzJFyM+7cFuv
kach21++ZD9H5ascNW3GQe0eIsUaKRvp8TqlVX9sFm0vc2o9UalqjAG2vDHyjNpj
ZOhRYDY22ADjvNTW6oauHRwdyXLAaHz+Q8cQyYj1tLYpW8+itMZ13s0V0GAMNNDo
dflRK9WUtQQBu3RqnDvi2dkUD+LpTvTCEW6icjlpwVsGzj3nBvTrX3VmgEOqm+51
hWbOkYxgFyWTU2ztRRVVMjn8Tk72sY52HmuPD5xjORohSaR+A97ksxPvmvGkhnAn
FSU8IeegK39BBxbVeK9Dzc1MKRqPhQNQoi30Ux9wra4j6qj/7rrcPMJ6v/XJvDln
o6AEHKxF19ixiWXQpKzG7iPNRz37LuY4J6bnO9qrRRAUl/u1KgW7mzhiikxC9+7Z
6EkufiSCrkGcIKkRiRQcIgsdkMArca4Dd/QtynInizGhT7qXhhIAFZYJN69Q0JvK
dKYdUjctiO3UL3isD4l9RHzZrChYaJJ6c9UmvGPcIZAkc2jjj/eHJ4dkjOcb26Qr
qWrXTK/GE3kyKBDCjfisTrBS91oy6uJkrERzknWJOyUReX8wf97vcP/qyZoVAitk
xu/lZNkAGBsXb3CgMfnc+kKQTmxJ/RWvNM3zuLfbpSWD9NeuDAj5V0dH/tPxzS4x
W0SYaXTi+u3QI+diBxKZ3NsjLSn8A8LNL+P9uGn5Dmq91PWQqPrVhGh8BDat8xwX
jAStldXi48bN1FCiOy3n/C3Ktlnbyk92o9KSn1m16aMGTLkLM9no/9P1fKrxca8p
X9ojOQ2eyVPG30XTLQmGoCRicjQyZC5+BTqShczE0HbJSDmDC+LirPTvXLwxLY6z
jqsWLAP4o0VLiPmtV5KtEJls9/pw0cb11FnQtGTBFuH/5+PSTIQhUTdCxNusyYxy
RDS2Mb/dr1vyKAR2lBfBLamgtIZFUi2wqnbQC6yuX6YJVk101PLmv3WMF1riIsk+
Q0usjOf9U4RCqI4FaXDm3RrgRsr2oigwOG6ivctb5TAwrB60K6+w4ohbagsgEglf
zJ6kHccrwA4UibotPDGZd3VUKHgczcC8ziTz8UIFfvC46wcIX8IQd1wnsiUEFSSj
uuIm4n+p7kM02BalgoKWyqccm0RtPFROR/zsF/dUf4MfAvXxP+dPNBnhmVr9TwF7
t6SM04/NHn36c587q2Ld9CgMIInGVKzfjHI+8aOHmRGCz7KNgkHbsq99o8qPzvPi
Y3FmI1Q/i9E7PpZ3ZxJ3ARsbpMwyyi4XnCyS5avWnMj0cAzNER35xZIQtOuCHfO+
ukmakWpx4tITttdQzy0Bb2qgMZbg0/fnA6StAXS74KmxJS+0W5DUHXg+4zHlOx9a
SW8NYDZiXCHnmcWuwY17TFwwRVCvQ4v1JsgDC3b9ndHQzzp7cEAiEffAxtzY32hh
bTCXZyCfkqDmL6SqHJvPf9KAT+c+YmE1sn6Yqm2UkaYrmwxzwe6u4wilr4CP80Vp
gu4UAwadxm4UFErWUAK8IiBAAoqdxRBi1QfCP//uKxjXtn6d0GknWW3gYCPe5XMv
cjEoHb2WtzsE9+Dk41o6VyCCnOUO11rFJbUlrOaEfG4QVBjnsX+GAhT6+ps1U47s
j2alrJ+wNMILXFutnql/fMDNqWHWzGHvQwT3Hu4EH5YZvIUahp10Qs7VCwvcrQgr
/muwJG+803bXaRAXbtvm/3MxWY13ohnTQyipsTN/aUJOzjXx8I2e9DW73hAoGgaZ
JSEVjkfZuZwuhUNtMqGapjXR1P2os7ugvmKOUfyg2OSXPprWmlxltrG4kKPfw4f9
wwsDCUZA8EL+W5a1X4EklL/R9NhSGxZJGDmEUO7Nqf7VFpTD5HySGiWBAB/vxGh/
6sCZXXmccApvEWi2AeeAsE5GVVx51R4QHOARjMs0KaI7qxn1Qtd7ohinoDrbcoQ+
eBLeBMgkj7GJj64/l+e+0GjXJIAWjbPz+S4M39w4NHlE377idDkCUMvVQmexyrhk
+ABL02Bv+FPeRR/3CNS5vhk5lI63ozuQ89AlNVKC4nNgHGfTqCcwfSuMSGx5WJXV
9zwHsgUwsH5mGM86qhx5kDGSahK52TADBNt0QgsnD30e5zsKRi9Bmxt1NmTWeqZ3
r1AzNXGOB7o13lezEqDb52EQzRNoHoNDdE/JHw9vCgHEXDVY4WOW75DyXweBv/CS
ibBW0BIjg+ILJZWqGAWMaMqlD6NBZRVPRVW6m4vGVqy3qFqUjpg9i6RQYK2WuqaX
OcDYcTeeAZF0KaPVmcdpktqNanzgpqBr/ObtViJmXbQ=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
B4a6SZ3sDwwPCLxJ6mdpxFwBwcSpzU60Cnw/LtZQw6Oeq/GfnlOjE3k6tfL2c2DK
9dobu3w0XGAcH3Ai2d23NDYje/I7AGxCmzVQGlV0bE3BCuY6aoBNnHLE65Ya8Q5e
QKfrzzvYY3YxZZO66w0UWxEzkT0hDBOHBCLV3Q7yQEw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5472)
IiGXKJ3y3G+BHqd5C6xJV/mRqDO2YF8+sdzx02QyFy14CT8WpFpT5DcoQ6ZFgCLe
n45Zqc/KliQYvlQe8M2seQkJ2TxCUUiw1pP1ti7h/vaBNwfI2PO7ngvlydaa5d1/
1Q6yRjk82sob0czhVTxuGQSET3rCCd7T8TFgSGNwshofaHDkcQrBSlqW6JHyv69u
l058RljZPwlB4xngq8YCuOcNmaz4Yh0YzxVh9w8o4ryL2rICowH08vp/aMEUUiPy
Qy754/D3MQJ1RzVKACh+gyvz+OEO11AP67yV3mszzdvA5vgKEhjihXFtMFATDtD1
3bDJkEyW1ethIXS2JjA11qXkHuRR2jd+Q37EIgFYvQJH6XI77Kj55CkleUxVbb7f
/zMn7oYof1bsIF38U/GkuiHVqRGFt+RmJAhISgcgwF7PEyQcH5b77ANc1cEHUnx1
oOXCIQMR0ORwVl3VawV45TEKoddPeGvhJqFv++EUF7iKOvuwYAOPE29dYo6o1vZk
+IId9HH74wge5qg+tJTvvpsLfDXrGqk+a6jHkxX1Z1n1HvSKmBeoUvA7p9Lprj+R
AT+8Eqbk7867O4LToMJMG+zQt91ITnrjPUEis1xOt/oJiRETWAURyMjMorPMxs/H
NQ3e/C3XAjVed43mcbLpfWCwmN4AIVbHlqTSb2g8IXxKLd1y9b5+4lIeOcnS8o32
Pmt9Kp4ZdA1+5PnVRGY1GIKRggdg3hRkuBKXmKLEquwb0GbdgBQU4SEV2cxciHu4
YHR+hlg2CRWkvXufTrOhErRnhk/2K488FMrzvQhIQgJyzF6/XPsciFRii8oWYw1f
fZK6YN7+gAgUsxdCLJSDj/XRxwhGfa+K1Kj72DqkMHFdimy6uBAOmJykHrFHCJ7E
DZRUigjtz5043qdYgc8UwxxdFk1huEUkEBglwG3YeNQ83PEssoKSjVwTfOvvrjoF
+oc1cWWjCL77ILFMHjz10G3pa9bAK4EerGnci+1ugVMrc3W7dddz3/mCGrMiJPuy
HgUVhBCg4dQZTgmAyH4i1HLfhHgKs8UNnSe3K3Lb5z0A4W/FW1e9fw1LP09qEmUD
C73S6M84GQJDFFmKBOyX2eqJ2ExJSK3j6MUaWn/LNsJ1S8d7Fzv9IilJpwZWyifI
OsNtOKirUfq5PebVaq+c1CtrY/vuDaHWyW1+KNAop3i8lslBk8tnRc7/YyaLXS8g
/Y8H6uLf64rH8pE5JZMlRm/2kyAX3VRxsKbctslGjuepNfG7BKjfJzHa5KMXLAlq
coyV54Zflge899gJ6ff6XInHCSv05RrJS/gnN0zOJI6+VAL4hs1xgrel411gy/KU
j5CUf2bFU/atg4FmPWNIFNqQfItV55oc55wztpJ+m9KMQRAWR1Y0W7qH4RTj1Quy
F5ApH0baLmXSWpbf37CNyGfeZ9Ors5K8TdyuIWBW1geEuq4ESL78TzvKfcx5x1su
tpsrq+gzqJpp873YtFSkMdETt54sqyLBrzd0VpFTEsEFzA7JbQWVpyKk96zJBqUg
W/tl5Bij8iff2+prH3vTX/cAgHOkP/D1FAZGgoAN6U0y5wvuulfjqughib6UdCPd
m5ZuQefvw1zDkOARe7CokPViWlbTpXqqeqh1FTJh+dbq1aBxOT792A5Qj58N+m3v
PQy9vS/JPgLnPz/FOtbj0stxhBWaLoCDFYUt5I68oGGqjRW8gewaZv3Hx/YL3eFv
ter9IXkqjl1DIdSLhHtbGkChofFOg/hf2XPjs1XFdX95wu6owuaSW+48+N7tag4z
LdhCaQiXVQ6FvjK1ENMYnOG8xHyV8oVgRGowGsg5d6S4WdZ4Q68N/KWYLlz8sSlY
bU4jMwtP0Cnlzvx/Kk7h3CUWSjERXc+30CCZXtsdjJZDRgnE6QbZv5hIPV2maiAd
na6n/q3sMqjaoHBjVf+rIiWKxIBw6J0eibsIqxnr3Bsr04//9hJpNAEOvQX0mXUu
0m5KqRMTa5lgvQX6WG/oU8jlAArcdQr1aEz1YGpLIWRqVStKS7Mn4/D/hpTnEJFW
9WIezxi3r7iYk5BeViMzNr1yCxMA+H5PXZFnszW3tDeuJxaa8iMUKBDnUxYtr+fl
dDyw6/bYOkUvfAGDttm8wCx7IbrxfVSvYQaOOQgXKDjruH6H2guJUtmwFHS3awmV
JvGDMdyIKcq6MuyEopv4Q57suv0TB0A/dZg2Qv5RnNpXdRsF2Gyp8vaIG3v+xokK
j4AqO6ZtcU7ZRdZYTDnhy+bj4Qt5ZM00H1uG9dN3TWYtne8g7y6ec8lM02mIPZ1d
Aqg8yXYT2y1v04gPgeISb72yFgqIQsjKFCyV3A2CZuXb0W27sDU1u/80JJQEsT3C
iEx/l6yEnI+1ZoVKk1OHtzBvlwvcr0G5snjA8HCRUNGws5U5yW578zW5MADzekIH
IQ9PntbDTuE1neHrpwhbE/rXluOupcdJLZmd9VBVtzinpWS8uf8cdAULGvd8bOZH
bRLbuS91Aa1p2l+kpVIMTeMZ24GbybD5jFV6rYOv+itYBGfNVqbBLXhG0iWGYfpn
688b3XNbkNaPIIAG0lVOiuh3enZOdbwOv3vshAj5UOtMi9F3iKCjLR4SfoiZbYfM
0d78vT1Tck/WEg7NKSaupNBP2j7KLTIkp4qPHjplSTHVH1TLHisfWz2dW4N5dAiG
2YLTkkuSSATP7DlPrsDtnXcUV6MbRe8jgGPLkcoX5cdSWHBalVhW6eCQ2IJMPm/T
X8PN9XsErd4e7J1Sbx7sVpU9+vYTtaq4NF2dtkv9EsNKvAK/FvrWpMKBYGaQAnWM
bDMqC681StUYZ4zRXyYVXqwKqMxv369P82Qdcov6YxY13fxhXcHItDsk58R5lg/0
panD0tqZpIMJEED3X97sF90hTIgw4UKuIegnldjwSJfIAyzmO8X4GalhP+bxCCf5
Qaz6I2Wlj1S/GOaaCa7SW/GE9gdFvWSs9SvGZH+O9oepV2+9HwAcDbQ5fXp6ICuA
cHjse0kSS9MCEA833V84CbXTHVLLPTOJ8aIq04KyspqTvq7OwMuf6H5Nx3vAYUlF
GA7HPzCnvtee+OLTeY7K7DjSmQ69HTJy7F/KzxHp5v8a7U0/jpQh8rGkalVZeGGC
atcsDduKp+81QNFKLcRTcm85zjzGWXd4ANtSnkY4gXtF34bDmwVr7UCmCB5Dt6R1
V2elp97I+ua3fdi4S/ZyAghmMabCWhsZz5PZF9uX7qKFrlY632Qi4fkIrfvV9Jg5
AuahT9iRLDhVw+5BY6437OHuc/IXeII8E738hDfxuAfSLGhLr/wLb4U7J2wEo4S5
puvlnr5Q/ltuNaCrHmTSe7DS4vCYDXKo3yfhPS+IBrY/Mu9y3Pz9hUVtkAKFLsNM
zIi2GM2MCNDeP5vGMsIX0W9KbpBgHaIAbmpXlwEWg0so1BB/jAs1Yllvd3sL2QQ5
9tD4GTwLHlEaiB+I9UO9uEQZXM5gm2Czflvz50yk7TQsderv87hh/AFva8npGEY1
98ZUFDCvp8C5t46s1kapgnGJiGXeHlqpq84RJIO1UmcZylJUfYiAzrLhsv2ncVEp
DVD9itGjjkj7b4KauJwingCjEllykaOPFio+qbdVASnWgPBXjWPiPFCGIUYbjFAR
t1P6CmxopvVfnaKPamvdNcCOmE07+MNxo+FGDDolHcI+wx5KQVno7lkeTzsEOJ33
ndEA+dhugxJmSrkaoGVReu5X8unpJbRPaa/qL1fiMJ376BBRvK0K6yenmMVo3+78
tQ7hovxEP9DgInnG3aeBvyBfID+kW/h2QQsZS/Aqi4Dk1lTavvkqQcY3N7SMUO31
exlm4nSBpVBq7IZ6bI7lEBBCI1QxSwNjJqSa2/waHrbn95TAFWcRFQuKq/SS6riF
s16exF71uhwMlZoIQr+NdjzoZY5e9DHfir41aes4JMajBLlGZOteXN8rWJAKpvFF
gbevLnGdbmof2PhJyB98gfJdj5qei4CsI23prWDLozS2iC3QAzUMltXwQNWnbEdd
5To38rBy4z45N62BVk0Lv4C5IDbLiUwIRhDRG8CvE1s9pfPgW0d5s1hPuLWPejtT
+O2sNNZKhqvxhYShqchEGyekFDppnjY/1OjXbe4WHz7Ni2nVye4LPQAa8cSuJakr
5zgEm5MqdRsuv8ATke0bCrJ9toW9P56zyAFN7ybmyynPsjloyjLLwuWyXOzBzIdP
hvjlSv1L+7/mwn0mivwLClXj7uGq6GjGjmMkxYJgJnpFzndj+AKZi7/To3BrsvGw
MfnCYroe9GuWbyQTC9bsDVhJrS0k6X5/hZ6YeIBtrjmcbTtHb/0mI0OxZ4+X5eWv
OJ0zr/RDhIy6gfD0pODThN55AMJNCeQuXKCSPzQsAy2bwrxX8GsPzSwlv/0lLJX8
EQaYDdo8Xfa7yZR0JDRzdTRHHgPn6n9La1NmHKI/oJVfXbeCE8WwQ6OsM/QCkXmA
NaziX0OBYshvmaa7QEuuQSjWVkVxSrLejJ79Xu9JXtw27HupvHBEdUm3e91T3Nvy
wYbZwOyH1GENl/j1Ty5fu1B8fA8LjP426I4M9ML986r1o3EXGZ69Xa5QPxjqonGD
iJOasZpYbddQtPmqO8M42I70NiI7WSm5ZsSXqLQoOpfUbBCVjD9fcRAuLV2R/Bu+
5wKIw7T6B5xrHrZVCPtz3L9R0Fa64moyWt74M4KWmj21nfzbEeo5lemJ7hfMv87k
rBGJJ7NSFZx36sZqw8mEbIwffr4syzLkZe9ZJRhrvQU7XvXCk8NWxsQODOmNy8R2
Xj8cDayllhd4v2W2UJHtIDPqffb1deG6UpQ5S4iZK9bhoA31ng354QKdYLp+VkYn
W/7wP2/uB1xlGjwheFn2gQVIu69ZhNnNaqsj8X4eAckm2YZw8GeMntagrocJ9Y3q
GwQk+qdrxdDW6SYzwVE6QKf+8qaahNx5VbbTQfcJ79wYzG9UK7EbX6E9aMpTpYsn
4H1Ky11rUI8fsU0B8hbNWAH7DrjLMo520CeZEPfTGhpxFI7Gi85bTvoLOKCnENS7
0MqWmnpE6EgApgQht+c6FED7C0PkmgpX4JVT6SEhulqBUMjEuCJk4eWu9e7akuXd
CC8nvz6ujn0jVux/68zNmf+j0PnDcEGNkhCSWuz7wTUuzsP4NT5SWCFViG1HEtQw
QLwpWgOqyL+SZ+1uxGa/TR9tpfl4chb87Q37pU6nul8gIhtdHqWmR4cxzM0LoE+o
qu8Fq2r3eexN55AzeYpsWVN8wO343VaaLaodLzfuP51YQHYcGna2jfojzLigisYD
te1hvB3Fh+r/IArye2NsgLeeYw5zcyF9/690TyNqK1KdWkwc39UcIFJfW3qBJNex
JH3ANTFDO7FK/LAVt10McIIMOELa/fiIXtSE7aVTMWATQnJ5rDGmhKwScAnhC5w7
yRZ2I2PXfC55L08TRJNn9aCV12wUHdwFlgtKkpS3MWtkuitNecdrUkS3jkXesK9r
lJuiDoytNJo2apOP6htFj9quYKvzYJT/qVzeWoUhyBwUk7hV5+Q3I30RKu7uw81S
LGquFQ9wAXY08pib0dGcsspcMNg2RYUASxjPmGAEsK+/P/ljnEmVhBsbgh1d8LZJ
8yPLiU/UPyCbVxlRXch14TCHYQXJmHvSlYP/I9o9/pqcRq8vtngfZbuMrgn+UvxK
wr5Q/qkhuotktOUskyvRo0xQM3Zzgdq0Mv+UpMproEokmiJAMFMhEbExymCLokGo
+v7abfA4izBqbwbWAPVHt+pVBjo7TxpIb9vTq5jiKCDCw0+bjMjVVSliG1HSA3wF
bqztuPUMhDU+uxXd09Px3CEaWbFLaCv69ddtb5Otd26eOkK4/d9x40OMFUbqHSao
g0gPi3+PiT9j6I3OijwFWmjaGAAd/tHFTE6OCp8q8OnJRVVyZqroAq1YADLALOag
bJUgfAeziga5SkcBt6XKS7f6sKc75W3x/cIOUrTGu9SKyrIGuQjza2OtDhLQzFQX
TC5TE6rToEEUMY5DSddfdD6u9PX8slOhjC1crSRauEsp+gw+iKg3S5NsFJ80FmuS
PMqRdM7mNeqIIR8zIw7W07o2C/sha4lq0TGXNnDSZCcYR96E2o4Q1+92lkRYHxaQ
wkzJhKoPKH8vpK8C/o9vBU8S9h8GbufAQFs/hvlFpXljV6/9IY8nLjRR+G1K0Cf+
K5JAhIdBjN+4Ig7VJadzWXq7kiMQJYUqjAJdUGQANH8QTMmGDl81jllni326qebC
1mG4bLFyaV3UQMnlhlBpeAyIcA6iUiS6mR/ocS8R5034FckpAY82OJhkyR4D4HJE
rmHa9w6hByKDJPTttE8UwwEafp/0GRhsk+uX4fZCsAokghDSPHua59LMhkYg1fM4
EQeut6VsQNV4p+G4rtu2bgE1elOkxvmq++R+kRXXyccSiGbbVFErshcyjFtpavHW
5qiPH34B3oKQ0KswHQH0EtT+rP7SdpZu7EXvB/uv5hyEDjjsAVCGT/GD57hJZJVB
rPD4Qmv2VLSBdCp5yvT14yFi0ID3omAV8PU4mvJgf7Es6paB5VyPnYSP08w0afcY
sbksETb1jO3Y43tQsO2ZiNJ+jvVs4/OMgXGTBuGHGJd8/ubaGx5RC8Lm9imPKFdv
ozBpEiwbUKLwc2VcSoI/mfZ0WgCBo6NoV/N8UEQVnAn4lNex34VPiNDF1PZ9lsgE
TcwymtSf3/Xq0hUIHPDRN8Zfz8PG0jcKVSYiPNm/IzdOss5unkrSidilIAoy7J4c
WAJ4KGqrN5IzAysS72Tsig53B+9e4/OLRBR+3VAy2Ve5VYnfpHeudenPfbIe0c3k
1j816XTZ5aTJoZV4O9F2VP7Ln5xKb7DLAhythmjOZ4ghVSivl/a8s5F0TlMknxw/
FPfONVt8NvVJAq8xcKlCciBAXDFgHuBp8lKfLkSdGilg6kosNyjpGrw2NAnv7F7B
MnoUC6rncY8HAbP7gLIUi7oVao40v0+K503H2hkqquseRxeWnqvofdbqCHMaQgKt
WAGfVjRzWr0xmjvJyNMB7MRWROtTT3b5Wcw0M0pVgthke8Yv8ATL+iPj5YjL240c
n1NGvBp7sUcgPFzIhazIzHYNDnVlmFXQlw8bvVApjTrcavDUslCz3HW10TamNaJR
r5RZ4nJC9k04vNAsZjpgL1hZrXy+M0zj6OkJFEVi3MRlpzZRVRgMF+wHQoYyKW0z
nKtUGZO4JobYmYFYCiCir+wTrY9rsR81V0xfuHudS+SeEdpT4fkFoLa8gtjoBc6A
`pragma protect end_protected

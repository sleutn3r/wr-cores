-- WRPC LM32 RAM initialization: --
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.memory_loader_pkg.all;
use work.genram_pkg.all;

package wrc_bin_pkg is
  constant c_wrc_bin_init : t_ram_fast_load ( 0 to 32767 ) := (
        0 => x"98000000",     1 => x"d0000000",     2 => x"d0200000",
        3 => x"78010000",     4 => x"38210000",     5 => x"d0e10000",
        6 => x"f800003a",     7 => x"34000000",     8 => x"00000000",
        9 => x"00000000",    10 => x"00000000",    11 => x"00000000",
       12 => x"00000000",    13 => x"00000000",    14 => x"00000000",
       15 => x"00000000",    16 => x"00000000",    17 => x"00000000",
       18 => x"00000000",    19 => x"00000000",    20 => x"00000000",
       21 => x"00000000",    22 => x"00000000",    23 => x"00000000",
       24 => x"00000000",    25 => x"00000000",    26 => x"00000000",
       27 => x"00000000",    28 => x"00000000",    29 => x"00000000",
       30 => x"00000000",    31 => x"00000000",    32 => x"00000000",
       33 => x"00000000",    34 => x"00000000",    35 => x"00000000",
       36 => x"00000000",    37 => x"00000000",    38 => x"00000000",
       39 => x"00000000",    40 => x"00000000",    41 => x"00000000",
       42 => x"00000000",    43 => x"00000000",    44 => x"00000000",
       45 => x"00000000",    46 => x"00000000",    47 => x"00000000",
       48 => x"5b9d0000",    49 => x"f800001e",    50 => x"34010002",
       51 => x"f8003e5b",    52 => x"e000002e",    53 => x"34000000",
       54 => x"34000000",    55 => x"34000000",    56 => x"00000000",
       57 => x"00000000",    58 => x"00000000",    59 => x"00000000",
       60 => x"00000000",    61 => x"00000000",    62 => x"00000000",
       63 => x"00000000",    64 => x"98000000",    65 => x"781c0001",
       66 => x"3b9cfffc",    67 => x"78010001",    68 => x"38214e68",
       69 => x"34020000",    70 => x"78030001",    71 => x"38636dd8",
       72 => x"c8611800",    73 => x"f8004481",    74 => x"34010000",
       75 => x"34020000",    76 => x"34030000",    77 => x"f800004d",
       78 => x"e0000000",    79 => x"379cffc4",    80 => x"5b810004",
       81 => x"5b820008",    82 => x"5b83000c",    83 => x"5b840010",
       84 => x"5b850014",    85 => x"5b860018",    86 => x"5b87001c",
       87 => x"5b880020",    88 => x"5b890024",    89 => x"5b8a0028",
       90 => x"5b9e0034",    91 => x"5b9f0038",    92 => x"2b81003c",
       93 => x"5b810030",    94 => x"bb800800",    95 => x"3421003c",
       96 => x"5b81002c",    97 => x"c3a00000",    98 => x"2b810004",
       99 => x"2b820008",   100 => x"2b83000c",   101 => x"2b840010",
      102 => x"2b850014",   103 => x"2b860018",   104 => x"2b87001c",
      105 => x"2b880020",   106 => x"2b890024",   107 => x"2b8a0028",
      108 => x"2b9d0030",   109 => x"2b9e0034",   110 => x"2b9f0038",
      111 => x"2b9c002c",   112 => x"34000000",   113 => x"c3c00000",
      114 => x"90001000",   115 => x"3401fffe",   116 => x"a0410800",
      117 => x"d0010000",   118 => x"90201000",   119 => x"3401fffe",
      120 => x"a0410800",   121 => x"d0210000",   122 => x"c3a00000",
      123 => x"90001000",   124 => x"3401fffe",   125 => x"a0410800",
      126 => x"d0010000",   127 => x"90201000",   128 => x"38420001",
      129 => x"d0220000",   130 => x"38210001",   131 => x"d0010000",
      132 => x"c3a00000",   133 => x"379cffe0",   134 => x"5b9d0004",
      135 => x"5b83000c",   136 => x"78030001",   137 => x"5b820008",
      138 => x"5b840010",   139 => x"5b850014",   140 => x"5b860018",
      141 => x"5b87001c",   142 => x"5b880020",   143 => x"38634e68",
      144 => x"28630000",   145 => x"5c600006",   146 => x"20210020",
      147 => x"44230004",   148 => x"b8400800",   149 => x"3782000c",
      150 => x"f8002abc",   151 => x"2b9d0004",   152 => x"379c0020",
      153 => x"c3a00000",   154 => x"379cffbc",   155 => x"5b8b003c",
      156 => x"5b8c0038",   157 => x"5b8d0034",   158 => x"5b8e0030",
      159 => x"5b8f002c",   160 => x"5b900028",   161 => x"5b910024",
      162 => x"5b920020",   163 => x"5b93001c",   164 => x"5b940018",
      165 => x"5b950014",   166 => x"5b960010",   167 => x"5b97000c",
      168 => x"5b980008",   169 => x"5b9d0004",   170 => x"f80041c1",
      171 => x"78030001",   172 => x"38633cc0",   173 => x"78010001",
      174 => x"28620000",   175 => x"38214e68",   176 => x"58200000",
      177 => x"78010001",   178 => x"3821f800",   179 => x"58220000",
      180 => x"f800317f",   181 => x"f800392c",   182 => x"f8003922",
      183 => x"78010001",   184 => x"382117fc",   185 => x"f8002abb",
      186 => x"34010001",   187 => x"f80030d9",   188 => x"f8003709",
      189 => x"78010001",   190 => x"38216d18",   191 => x"58200000",
      192 => x"f800362f",   193 => x"f80032be",   194 => x"34010000",
      195 => x"f8002dfd",   196 => x"34010000",   197 => x"34020050",
      198 => x"f800337c",   199 => x"37820040",   200 => x"34010000",
      201 => x"f80035c0",   202 => x"3402ffff",   203 => x"5c220010",
      204 => x"78010001",   205 => x"38211818",   206 => x"f8002aa6",
      207 => x"34010022",   208 => x"33810040",   209 => x"34010033",
      210 => x"33810041",   211 => x"34010044",   212 => x"33810042",
      213 => x"34010055",   214 => x"33810043",   215 => x"34010066",
      216 => x"33810044",   217 => x"34010077",   218 => x"33810045",
      219 => x"43830041",   220 => x"43840042",   221 => x"43850043",
      222 => x"43860044",   223 => x"43870045",   224 => x"43820040",
      225 => x"78010001",   226 => x"3821183c",   227 => x"f8002a91",
      228 => x"37810040",   229 => x"f8002c5e",   230 => x"34020001",
      231 => x"34010001",   232 => x"f8002bad",   233 => x"f8002e76",
      234 => x"f8002ffc",   235 => x"f8000550",   236 => x"78020001",
      237 => x"384243d8",   238 => x"34010002",   239 => x"f800325f",
      240 => x"f8003e62",   241 => x"f80028ea",   242 => x"f80027fe",
      243 => x"f80025d5",   244 => x"f8001fa8",   245 => x"34010003",
      246 => x"f800059b",   247 => x"f8000556",   248 => x"780f0001",
      249 => x"78130001",   250 => x"780b0001",   251 => x"78110001",
      252 => x"78100001",   253 => x"780c0001",   254 => x"780e0001",
      255 => x"780d0001",   256 => x"f800207f",   257 => x"39ef43dc",
      258 => x"34180004",   259 => x"3a73187c",   260 => x"396b6db8",
      261 => x"34120002",   262 => x"3a311870",   263 => x"34160001",
      264 => x"34150003",   265 => x"3a105d6c",   266 => x"398c4e68",
      267 => x"3417001b",   268 => x"39ce43cc",   269 => x"39ad6dac",
      270 => x"34010000",   271 => x"f8002bb8",   272 => x"29e40000",
      273 => x"7c230000",   274 => x"b820a000",   275 => x"64810000",
      276 => x"a0610800",   277 => x"44200008",   278 => x"34010000",
      279 => x"ba201000",   280 => x"fbffff6d",   281 => x"29610000",
      282 => x"34030001",   283 => x"58320004",   284 => x"e000000d",
      285 => x"66820000",   286 => x"7c840000",   287 => x"a0441000",
      288 => x"fc621800",   289 => x"cb031800",   290 => x"44410007",
      291 => x"34010000",   292 => x"ba601000",   293 => x"fbffff60",
      294 => x"29610000",   295 => x"34030002",   296 => x"58320008",
      297 => x"59f40000",   298 => x"44720009",   299 => x"44750004",
      300 => x"5c76000f",   301 => x"5a000000",   302 => x"e000000d",
      303 => x"f8002738",   304 => x"f80028c5",   305 => x"f80027d8",
      306 => x"e0000009",   307 => x"f8000516",   308 => x"5c350007",
      309 => x"34010002",   310 => x"34020000",   311 => x"34030001",
      312 => x"f8003e25",   313 => x"34010000",   314 => x"f800304e",
      315 => x"29810000",   316 => x"5c360009",   317 => x"f8000066",
      318 => x"f80038c9",   319 => x"44370003",   320 => x"29c10000",
      321 => x"5c200005",   322 => x"f8001f5a",   323 => x"59800000",
      324 => x"e0000002",   325 => x"f8001f61",   326 => x"29a10000",
      327 => x"44200002",   328 => x"f8000213",   329 => x"f80005c3",
      330 => x"f8004024",   331 => x"f8004107",   332 => x"e3ffffc2",
      333 => x"78010001",   334 => x"382143e0",   335 => x"28220000",
      336 => x"78010001",   337 => x"3821488c",   338 => x"e0000004",
      339 => x"28440000",   340 => x"44640004",   341 => x"3421000c",
      342 => x"28230000",   343 => x"5c60fffc",   344 => x"28210004",
      345 => x"c3a00000",   346 => x"379cfff4",   347 => x"5b9d0004",
      348 => x"5b810008",   349 => x"5b82000c",   350 => x"b8401800",
      351 => x"5c20000b",   352 => x"78020001",   353 => x"38423cc4",
      354 => x"28410000",   355 => x"54610007",   356 => x"78010001",
      357 => x"78020001",   358 => x"38421888",   359 => x"38214e7c",
      360 => x"f80029fe",   361 => x"e000000d",   362 => x"78030001",
      363 => x"38633cc8",   364 => x"28620000",   365 => x"37810008",
      366 => x"f80007f7",   367 => x"2b83000c",   368 => x"b8202000",
      369 => x"78020001",   370 => x"78010001",   371 => x"38214e7c",
      372 => x"3842188c",   373 => x"f80029f1",   374 => x"78010001",
      375 => x"38214e7c",   376 => x"2b9d0004",   377 => x"379c000c",
      378 => x"c3a00000",   379 => x"379cfff4",   380 => x"5b8b000c",
      381 => x"5b8c0008",   382 => x"5b9d0004",   383 => x"780b0001",
      384 => x"396b43e0",   385 => x"29610000",   386 => x"78020001",
      387 => x"38421894",   388 => x"282c0014",   389 => x"34010004",
      390 => x"f80024ce",   391 => x"fbffffc6",   392 => x"78020001",
      393 => x"b8201800",   394 => x"384218a4",   395 => x"34010007",
      396 => x"f80024c8",   397 => x"29810010",   398 => x"44200005",
      399 => x"29610000",   400 => x"28220000",   401 => x"34010009",
      402 => x"44410007",   403 => x"78020001",   404 => x"34010001",
      405 => x"384218a8",   406 => x"f80024be",   407 => x"34010000",
      408 => x"e0000006",   409 => x"78020001",   410 => x"34010004",
      411 => x"384218c0",   412 => x"f80024b8",   413 => x"34010001",
      414 => x"2b9d0004",   415 => x"2b8b000c",   416 => x"2b8c0008",
      417 => x"379c000c",   418 => x"c3a00000",   419 => x"379cff08",
      420 => x"5b8b0018",   421 => x"5b8c0014",   422 => x"5b8d0010",
      423 => x"5b8e000c",   424 => x"5b8f0008",   425 => x"5b9d0004",
      426 => x"78010001",   427 => x"382143e0",   428 => x"28210000",
      429 => x"780c0001",   430 => x"398c4e98",   431 => x"282b0014",
      432 => x"29810000",   433 => x"5c200008",   434 => x"f8002ff4",
      435 => x"78020001",   436 => x"384243cc",   437 => x"28420000",
      438 => x"a4401000",   439 => x"b4410800",   440 => x"59810000",
      441 => x"f8002fed",   442 => x"78030001",   443 => x"78020001",
      444 => x"386343cc",   445 => x"38424e98",   446 => x"28630000",
      447 => x"28420000",   448 => x"b4621000",   449 => x"c8220800",
      450 => x"4c200006",   451 => x"78010001",   452 => x"38214e94",
      453 => x"28210000",   454 => x"296200b8",   455 => x"4422018c",
      456 => x"f8002fde",   457 => x"78020001",   458 => x"38424e98",
      459 => x"58410000",   460 => x"296200b8",   461 => x"78010001",
      462 => x"38214e94",   463 => x"58220000",   464 => x"f80024ca",
      465 => x"78040001",   466 => x"34010001",   467 => x"34020001",
      468 => x"34030004",   469 => x"388418dc",   470 => x"f800249d",
      471 => x"78040001",   472 => x"388418fc",   473 => x"34030087",
      474 => x"34010002",   475 => x"34020001",   476 => x"f8002497",
      477 => x"378100e4",   478 => x"378200f0",   479 => x"f8002f79",
      480 => x"78020001",   481 => x"34010004",   482 => x"38421908",
      483 => x"f8002471",   484 => x"2b8200e8",   485 => x"2b8100e4",
      486 => x"f80023e3",   487 => x"78020001",   488 => x"b8201800",
      489 => x"384218a4",   490 => x"34010007",   491 => x"f8002469",
      492 => x"34020000",   493 => x"3781001c",   494 => x"f800024a",
      495 => x"78040001",   496 => x"34010004",   497 => x"34020001",
      498 => x"34030004",   499 => x"38841928",   500 => x"f800247f",
      501 => x"78040001",   502 => x"78050001",   503 => x"34010006",
      504 => x"34020001",   505 => x"34030007",   506 => x"38841938",
      507 => x"38a51940",   508 => x"f8002477",   509 => x"2b810048",
      510 => x"44200005",   511 => x"78020001",   512 => x"34010002",
      513 => x"38421948",   514 => x"e0000004",   515 => x"78020001",
      516 => x"34010001",   517 => x"38421954",   518 => x"f800244e",
      519 => x"2b810048",   520 => x"44200148",   521 => x"378100f8",
      522 => x"378200f4",   523 => x"f8002ecd",   524 => x"2b8300f4",
      525 => x"2b8400f8",   526 => x"78020001",   527 => x"34010087",
      528 => x"38421960",   529 => x"780c0001",   530 => x"f8002442",
      531 => x"398c43e0",   532 => x"29810000",   533 => x"282102c8",
      534 => x"28210010",   535 => x"282d0008",   536 => x"5da00038",
      537 => x"78020001",   538 => x"34010001",   539 => x"3842197c",
      540 => x"f8002438",   541 => x"fbffff5e",   542 => x"442d0135",
      543 => x"78020001",   544 => x"34010087",   545 => x"38421984",
      546 => x"f8002432",   547 => x"29810000",   548 => x"28210020",
      549 => x"28240010",   550 => x"28830004",   551 => x"4460000b",
      552 => x"78020001",   553 => x"384219a4",   554 => x"28840008",
      555 => x"4c030003",   556 => x"34010007",   557 => x"e0000003",
      558 => x"34010007",   559 => x"c8042000",   560 => x"f8002424",
      561 => x"e0000122",   562 => x"28830008",   563 => x"780b0001",
      564 => x"396b19b0",   565 => x"b9601000",   566 => x"34010007",
      567 => x"f800241d",   568 => x"78020001",   569 => x"34010087",
      570 => x"384219b8",   571 => x"f8002419",   572 => x"29810000",
      573 => x"b9601000",   574 => x"28210020",   575 => x"28230010",
      576 => x"34010007",   577 => x"2863001c",   578 => x"f8002412",
      579 => x"78020001",   580 => x"34010087",   581 => x"384219d8",
      582 => x"f800240e",   583 => x"29810000",   584 => x"b9601000",
      585 => x"28210020",   586 => x"28240004",   587 => x"34010007",
      588 => x"28830028",   589 => x"2884002c",   590 => x"f8002406",
      591 => x"e0000104",   592 => x"78010001",   593 => x"38214f24",
      594 => x"28210000",   595 => x"34020001",   596 => x"4841000e",
      597 => x"34020002",   598 => x"4c410004",   599 => x"34020003",
      600 => x"5c22000a",   601 => x"e0000005",   602 => x"78020001",
      603 => x"34010007",   604 => x"384219f8",   605 => x"e0000008",
      606 => x"78020001",   607 => x"34010007",   608 => x"38421a04",
      609 => x"e0000004",   610 => x"78020001",   611 => x"34010001",
      612 => x"38421a10",   613 => x"f80023ef",   614 => x"2b810050",
      615 => x"44200005",   616 => x"78020001",   617 => x"34010002",
      618 => x"38421a20",   619 => x"e0000004",   620 => x"78020001",
      621 => x"34010001",   622 => x"38421a2c",   623 => x"f80023e5",
      624 => x"2b81006c",   625 => x"44200007",   626 => x"2b810070",
      627 => x"44200005",   628 => x"78020001",   629 => x"34010002",
      630 => x"38421a38",   631 => x"e0000004",   632 => x"78020001",
      633 => x"34010001",   634 => x"38421a48",   635 => x"f80023d9",
      636 => x"78020001",   637 => x"34010007",   638 => x"38421a58",
      639 => x"f80023d5",   640 => x"378100ec",   641 => x"f80027d0",
      642 => x"78010001",   643 => x"38215d6c",   644 => x"28210000",
      645 => x"44200006",   646 => x"78020001",   647 => x"34010001",
      648 => x"38421a60",   649 => x"f80023cb",   650 => x"e0000009",
      651 => x"438300ec",   652 => x"438400ed",   653 => x"438500ee",
      654 => x"438600ef",   655 => x"78020001",   656 => x"34010002",
      657 => x"38421a70",   658 => x"f80023c2",   659 => x"fbfffee8",
      660 => x"442000bf",   661 => x"78020001",   662 => x"34010087",
      663 => x"38421a7c",   664 => x"f80023bc",   665 => x"78020001",
      666 => x"34010007",   667 => x"38422e58",   668 => x"356300c0",
      669 => x"f80023b7",   670 => x"78020001",   671 => x"34010087",
      672 => x"38421a98",   673 => x"f80023b3",   674 => x"296100bc",
      675 => x"44200005",   676 => x"78020001",   677 => x"34010002",
      678 => x"38421ab4",   679 => x"e0000004",   680 => x"78020001",
      681 => x"34010001",   682 => x"38421ab8",   683 => x"f80023a9",
      684 => x"78020001",   685 => x"34010087",   686 => x"38421ac0",
      687 => x"f80023a5",   688 => x"34010000",   689 => x"f8003e8a",
      690 => x"b8206000",   691 => x"20210001",   692 => x"44200005",
      693 => x"78020001",   694 => x"34010002",   695 => x"38421adc",
      696 => x"f800239c",   697 => x"218c0002",   698 => x"45800005",
      699 => x"78020001",   700 => x"34010002",   701 => x"38421ae4",
      702 => x"f8002396",   703 => x"78010001",   704 => x"38211b04",
      705 => x"f80028b3",   706 => x"78020001",   707 => x"34010004",
      708 => x"38421af0",   709 => x"f800238f",   710 => x"78020001",
      711 => x"34010087",   712 => x"38421b08",   713 => x"f800238b",
      714 => x"296200a4",   715 => x"296100a0",   716 => x"780d0001",
      717 => x"39ad1b24",   718 => x"fbfffe8c",   719 => x"b8201800",
      720 => x"b9a01000",   721 => x"34010007",   722 => x"f8002382",
      723 => x"78020001",   724 => x"34010087",   725 => x"38421b2c",
      726 => x"f800237e",   727 => x"296200b4",   728 => x"296100b0",
      729 => x"780c0001",   730 => x"398c1b64",   731 => x"fbfffe7f",
      732 => x"b8201800",   733 => x"b9a01000",   734 => x"34010007",
      735 => x"f8002375",   736 => x"78020001",   737 => x"34010087",
      738 => x"38421b48",   739 => x"f8002371",   740 => x"29630018",
      741 => x"2964001c",   742 => x"b9801000",   743 => x"34010007",
      744 => x"f800236c",   745 => x"78020001",   746 => x"34010087",
      747 => x"38421b7c",   748 => x"f8002368",   749 => x"29640024",
      750 => x"29630020",   751 => x"b9801000",   752 => x"34010007",
      753 => x"f8002363",   754 => x"296e00b4",   755 => x"296100a4",
      756 => x"78020001",   757 => x"3dce0001",   758 => x"38421b98",
      759 => x"c82e7000",   760 => x"780c0001",   761 => x"34010087",
      762 => x"398c1bb4",   763 => x"f8002359",   764 => x"b9c01800",
      765 => x"34010007",   766 => x"b9801000",   767 => x"f8002355",
      768 => x"29610018",   769 => x"296200a4",   770 => x"296f00a0",
      771 => x"1423001f",   772 => x"c8410800",   773 => x"f4221000",
      774 => x"c9e37800",   775 => x"c9e27800",   776 => x"2962001c",
      777 => x"296e0024",   778 => x"1443001f",   779 => x"c8221000",
      780 => x"f4410800",   781 => x"c9e37800",   782 => x"c9e17800",
      783 => x"29610020",   784 => x"1423001f",   785 => x"c8410800",
      786 => x"f4221000",   787 => x"c9e37800",   788 => x"15c3001f",
      789 => x"c82e7000",   790 => x"c9e27800",   791 => x"f5c10800",
      792 => x"c9e37800",   793 => x"78020001",   794 => x"c9e17800",
      795 => x"38421bbc",   796 => x"34010087",   797 => x"f8002337",
      798 => x"b9c01000",   799 => x"b9e00800",   800 => x"fbfffe3a",
      801 => x"b8201800",   802 => x"b9a01000",   803 => x"34010007",
      804 => x"f8002330",   805 => x"78020001",   806 => x"34010087",
      807 => x"38421bd8",   808 => x"f800232c",   809 => x"296300ec",
      810 => x"34010007",   811 => x"b9801000",   812 => x"f8002328",
      813 => x"78020001",   814 => x"34010087",   815 => x"38421bf4",
      816 => x"f8002324",   817 => x"296300a8",   818 => x"34010007",
      819 => x"b9801000",   820 => x"f8002320",   821 => x"78020001",
      822 => x"34010087",   823 => x"38421c10",   824 => x"f800231c",
      825 => x"296300e4",   826 => x"34010007",   827 => x"b9801000",
      828 => x"f8002318",   829 => x"78020001",   830 => x"34010087",
      831 => x"38421c2c",   832 => x"f8002314",   833 => x"78030001",
      834 => x"38634e74",   835 => x"28630000",   836 => x"34010007",
      837 => x"b9801000",   838 => x"f800230e",   839 => x"78020001",
      840 => x"34010087",   841 => x"38421c48",   842 => x"f800230a",
      843 => x"296300b8",   844 => x"78020001",   845 => x"34010007",
      846 => x"38421c64",   847 => x"f8002305",   848 => x"78010001",
      849 => x"38211c6c",   850 => x"f8002822",   851 => x"2b9d0004",
      852 => x"2b8b0018",   853 => x"2b8c0014",   854 => x"2b8d0010",
      855 => x"2b8e000c",   856 => x"2b8f0008",   857 => x"379c00f8",
      858 => x"c3a00000",   859 => x"379cff18",   860 => x"5b8b000c",
      861 => x"5b8c0008",   862 => x"5b9d0004",   863 => x"78010001",
      864 => x"382143e0",   865 => x"28210000",   866 => x"780c0001",
      867 => x"398c4e78",   868 => x"282b0014",   869 => x"29810000",
      870 => x"5c200008",   871 => x"f8002e3f",   872 => x"78020001",
      873 => x"384243cc",   874 => x"28420000",   875 => x"a4401000",
      876 => x"b4410800",   877 => x"59810000",   878 => x"78010001",
      879 => x"38216d04",   880 => x"28210000",   881 => x"296200b8",
      882 => x"5c220006",   883 => x"78010001",   884 => x"38214f24",
      885 => x"28220000",   886 => x"34010003",   887 => x"444100bb",
      888 => x"f8002e2e",   889 => x"78030001",   890 => x"78020001",
      891 => x"386343cc",   892 => x"38424e78",   893 => x"28630000",
      894 => x"28420000",   895 => x"b4621000",   896 => x"c8220800",
      897 => x"4c200006",   898 => x"78010001",   899 => x"38214f24",
      900 => x"28220000",   901 => x"34010003",   902 => x"5c4100ac",
      903 => x"f8002e1f",   904 => x"78020001",   905 => x"38424e78",
      906 => x"58410000",   907 => x"296200b8",   908 => x"78010001",
      909 => x"38216d04",   910 => x"58220000",   911 => x"378100d8",
      912 => x"378200e0",   913 => x"f8002dc7",   914 => x"34020000",
      915 => x"37810010",   916 => x"f80000a4",   917 => x"378100e8",
      918 => x"378200e4",   919 => x"f8002d41",   920 => x"2b8300e4",
      921 => x"2b8400e8",   922 => x"2b82003c",   923 => x"78010001",
      924 => x"38211c70",   925 => x"f80027d7",   926 => x"2b820044",
      927 => x"78010001",   928 => x"38211c84",   929 => x"7c420000",
      930 => x"f80027d2",   931 => x"fbfffdaa",   932 => x"b8201000",
      933 => x"78010001",   934 => x"38211c90",   935 => x"f80027cd",
      936 => x"78010001",   937 => x"38214f24",   938 => x"28220000",
      939 => x"34010003",   940 => x"5c41000a",   941 => x"29620010",
      942 => x"78010001",   943 => x"38211c98",   944 => x"20420001",
      945 => x"f80027c3",   946 => x"78010001",   947 => x"38211ca0",
      948 => x"356200c0",   949 => x"f80027bf",   950 => x"34010000",
      951 => x"f8003d84",   952 => x"b8201000",   953 => x"78010001",
      954 => x"38211cac",   955 => x"f80027b9",   956 => x"2b8200dc",
      957 => x"2b8300e0",   958 => x"78010001",   959 => x"38211cb4",
      960 => x"f80027b4",   961 => x"78010001",   962 => x"38214f24",
      963 => x"28220000",   964 => x"34010003",   965 => x"5c41004b",
      966 => x"296200a4",   967 => x"296100a0",   968 => x"fbfffd92",
      969 => x"b8201000",   970 => x"78010001",   971 => x"38211cc4",
      972 => x"f80027a8",   973 => x"296200b4",   974 => x"296100b0",
      975 => x"fbfffd8b",   976 => x"b8201000",   977 => x"78010001",
      978 => x"38211ccc",   979 => x"f80027a1",   980 => x"29620018",
      981 => x"2963001c",   982 => x"78010001",   983 => x"38211cd4",
      984 => x"f800279c",   985 => x"29620020",   986 => x"29630024",
      987 => x"78010001",   988 => x"38211ce8",   989 => x"f8002797",
      990 => x"296200b4",   991 => x"296300a4",   992 => x"78010001",
      993 => x"3c420001",   994 => x"38211cfc",   995 => x"c8621000",
      996 => x"f8002790",   997 => x"29620018",   998 => x"296100a4",
      999 => x"296300a0",  1000 => x"1444001f",  1001 => x"c8221000",
     1002 => x"f4410800",  1003 => x"c8641800",  1004 => x"c8611800",
     1005 => x"2961001c",  1006 => x"1424001f",  1007 => x"c8410800",
     1008 => x"f4221000",  1009 => x"c8641800",  1010 => x"c8621000",
     1011 => x"29630020",  1012 => x"1464001f",  1013 => x"c8231800",
     1014 => x"f4610800",  1015 => x"c8441000",  1016 => x"c8410800",
     1017 => x"29620024",  1018 => x"1444001f",  1019 => x"c8621000",
     1020 => x"f4431800",  1021 => x"c8240800",  1022 => x"c8230800",
     1023 => x"fbfffd5b",  1024 => x"b8201000",  1025 => x"78010001",
     1026 => x"38211d08",  1027 => x"f8002771",  1028 => x"296200ec",
     1029 => x"78010001",  1030 => x"38211d14",  1031 => x"f800276d",
     1032 => x"296200a8",  1033 => x"78010001",  1034 => x"38211d1c",
     1035 => x"f8002769",  1036 => x"296200b8",  1037 => x"78010001",
     1038 => x"38211d28",  1039 => x"f8002765",  1040 => x"3401ffff",
     1041 => x"f8003d35",  1042 => x"b8206000",  1043 => x"34010000",
     1044 => x"f8003d32",  1045 => x"b8205800",  1046 => x"34010001",
     1047 => x"f8003d2f",  1048 => x"78050001",  1049 => x"b8202000",
     1050 => x"b8a00800",  1051 => x"b9601800",  1052 => x"b9801000",
     1053 => x"38211d34",  1054 => x"780b0001",  1055 => x"f8002755",
     1056 => x"396b6d18",  1057 => x"34020002",  1058 => x"b9600800",
     1059 => x"f80034a8",  1060 => x"b8206000",  1061 => x"34020001",
     1062 => x"b9600800",  1063 => x"f80034a4",  1064 => x"2183ffff",
     1065 => x"08632710",  1066 => x"78010001",  1067 => x"15820010",
     1068 => x"14630010",  1069 => x"38211d48",  1070 => x"f8002746",
     1071 => x"78010001",  1072 => x"38211b04",  1073 => x"f8002743",
     1074 => x"34010000",  1075 => x"2b9d0004",  1076 => x"2b8b000c",
     1077 => x"2b8c0008",  1078 => x"379c00e8",  1079 => x"c3a00000",
     1080 => x"379cfff4",  1081 => x"5b8b0008",  1082 => x"5b9d0004",
     1083 => x"b8205800",  1084 => x"f800020d",  1085 => x"34020003",
     1086 => x"5c220003",  1087 => x"34010002",  1088 => x"e0000002",
     1089 => x"34010001",  1090 => x"59610028",  1091 => x"3562004c",
     1092 => x"35610048",  1093 => x"f80028aa",  1094 => x"34010000",
     1095 => x"59600040",  1096 => x"59600044",  1097 => x"59600088",
     1098 => x"5960008c",  1099 => x"3782000c",  1100 => x"34030000",
     1101 => x"f8003c5a",  1102 => x"44200006",  1103 => x"2b81000c",
     1104 => x"596100a0",  1105 => x"34010001",  1106 => x"596100a4",
     1107 => x"e0000003",  1108 => x"596000a0",  1109 => x"596000a4",
     1110 => x"34010000",  1111 => x"f8002870",  1112 => x"5961002c",
     1113 => x"34010001",  1114 => x"59610054",  1115 => x"59610050",
     1116 => x"34010000",  1117 => x"f8003be5",  1118 => x"59610034",
     1119 => x"34011f40",  1120 => x"596100b4",  1121 => x"78010001",
     1122 => x"382143d8",  1123 => x"28210000",  1124 => x"596100b8",
     1125 => x"596100bc",  1126 => x"35610014",  1127 => x"f8002815",
     1128 => x"34010000",  1129 => x"5960001c",  1130 => x"2b9d0004",
     1131 => x"2b8b0008",  1132 => x"379c000c",  1133 => x"c3a00000",
     1134 => x"c3a00000",  1135 => x"379cffbc",  1136 => x"5b8b0014",
     1137 => x"5b8c0010",  1138 => x"5b8d000c",  1139 => x"5b8e0008",
     1140 => x"5b9d0004",  1141 => x"5b830030",  1142 => x"78030001",
     1143 => x"38634e9c",  1144 => x"5b82002c",  1145 => x"5b840034",
     1146 => x"5b850038",  1147 => x"5b86003c",  1148 => x"5b870040",
     1149 => x"5b880044",  1150 => x"286d0000",  1151 => x"b8205800",
     1152 => x"b8407000",  1153 => x"34030000",  1154 => x"44200002",
     1155 => x"28230018",  1156 => x"b86d1800",  1157 => x"0063001c",
     1158 => x"4460001b",  1159 => x"780c0001",  1160 => x"398c4e9c",
     1161 => x"39a10001",  1162 => x"59810000",  1163 => x"29610028",
     1164 => x"37820018",  1165 => x"28230000",  1166 => x"b9600800",
     1167 => x"d8600000",  1168 => x"78030001",  1169 => x"38633ccc",
     1170 => x"28620000",  1171 => x"2b81001c",  1172 => x"598d0000",
     1173 => x"296b0334",  1174 => x"f8003f08",  1175 => x"780c0001",
     1176 => x"2b830018",  1177 => x"398c1d60",  1178 => x"b8202000",
     1179 => x"b9601000",  1180 => x"b9800800",  1181 => x"f80026d7",
     1182 => x"b9c00800",  1183 => x"37820030",  1184 => x"f80026b2",
     1185 => x"2b9d0004",  1186 => x"2b8b0014",  1187 => x"2b8c0010",
     1188 => x"2b8d000c",  1189 => x"2b8e0008",  1190 => x"379c0044",
     1191 => x"c3a00000",  1192 => x"379cfffc",  1193 => x"5b9d0004",
     1194 => x"b8402800",  1195 => x"5c600005",  1196 => x"78020001",
     1197 => x"38421d7c",  1198 => x"b8a01800",  1199 => x"e000000c",
     1200 => x"34020001",  1201 => x"5c620006",  1202 => x"78020001",
     1203 => x"38421d98",  1204 => x"b8a01800",  1205 => x"28240008",
     1206 => x"e0000005",  1207 => x"28240004",  1208 => x"78020001",
     1209 => x"38421db0",  1210 => x"b8a01800",  1211 => x"fbffffb4",
     1212 => x"2b9d0004",  1213 => x"379c0004",  1214 => x"c3a00000",
     1215 => x"379cffe8",  1216 => x"5b8b0018",  1217 => x"5b8c0014",
     1218 => x"5b8d0010",  1219 => x"5b8e000c",  1220 => x"5b9d0008",
     1221 => x"b8205800",  1222 => x"b8407000",  1223 => x"b8606800",
     1224 => x"4460001a",  1225 => x"40480000",  1226 => x"78020001",
     1227 => x"384249fc",  1228 => x"2108000f",  1229 => x"3d030002",
     1230 => x"282600e4",  1231 => x"b4431000",  1232 => x"28420000",
     1233 => x"282700e8",  1234 => x"78040001",  1235 => x"5b820004",
     1236 => x"34030001",  1237 => x"34020005",  1238 => x"38841dc8",
     1239 => x"b9a02800",  1240 => x"f8000048",  1241 => x"34010021",
     1242 => x"4c2d0006",  1243 => x"b9600800",  1244 => x"b9c01000",
     1245 => x"b9a01800",  1246 => x"f80015f5",  1247 => x"44200003",
     1248 => x"340d0000",  1249 => x"340e0000",  1250 => x"780c0001",
     1251 => x"29610000",  1252 => x"398c488c",  1253 => x"e000002d",
     1254 => x"44410003",  1255 => x"358c000c",  1256 => x"e000002a",
     1257 => x"59610004",  1258 => x"2961000c",  1259 => x"59600008",
     1260 => x"44200006",  1261 => x"29820004",  1262 => x"b9600800",
     1263 => x"34030000",  1264 => x"b9a02000",  1265 => x"fbffffb7",
     1266 => x"29840008",  1267 => x"b9a01800",  1268 => x"b9600800",
     1269 => x"b9c01000",  1270 => x"d8800000",  1271 => x"b8201800",
     1272 => x"44200006",  1273 => x"29620334",  1274 => x"29840004",
     1275 => x"78010001",  1276 => x"38211df4",  1277 => x"f8002677",
     1278 => x"29610004",  1279 => x"29630000",  1280 => x"29820004",
     1281 => x"4461000a",  1282 => x"59610000",  1283 => x"34010001",
     1284 => x"5961000c",  1285 => x"34030002",  1286 => x"b9600800",
     1287 => x"34040000",  1288 => x"fbffffa0",  1289 => x"34010000",
     1290 => x"e000000f",  1291 => x"b9600800",  1292 => x"5960000c",
     1293 => x"34030001",  1294 => x"34040000",  1295 => x"fbffff99",
     1296 => x"29610008",  1297 => x"e0000008",  1298 => x"29820000",
     1299 => x"5c40ffd3",  1300 => x"29620334",  1301 => x"78010001",
     1302 => x"38211e10",  1303 => x"f800265d",  1304 => x"34012710",
     1305 => x"2b9d0008",  1306 => x"2b8b0018",  1307 => x"2b8c0014",
     1308 => x"2b8d0010",  1309 => x"2b8e000c",  1310 => x"379c0018",
     1311 => x"c3a00000",  1312 => x"379cffe0",  1313 => x"5b8b000c",
     1314 => x"5b8c0008",  1315 => x"5b9d0004",  1316 => x"5b850014",
     1317 => x"5b840010",  1318 => x"78050001",  1319 => x"5b860018",
     1320 => x"5b87001c",  1321 => x"5b880020",  1322 => x"b8604800",
     1323 => x"b8806000",  1324 => x"38a51e30",  1325 => x"34030000",
     1326 => x"44200003",  1327 => x"28250334",  1328 => x"28230018",
     1329 => x"78060001",  1330 => x"38c64e9c",  1331 => x"28c10000",
     1332 => x"b8610800",  1333 => x"3c430002",  1334 => x"80230800",
     1335 => x"2021000f",  1336 => x"55210015",  1337 => x"78010001",
     1338 => x"38213d88",  1339 => x"b4231800",  1340 => x"78060001",
     1341 => x"28630000",  1342 => x"780b0001",  1343 => x"396b4ea0",
     1344 => x"b8c01000",  1345 => x"38421e38",  1346 => x"b9202000",
     1347 => x"b9600800",  1348 => x"f8002622",  1349 => x"b9600800",
     1350 => x"f80034af",  1351 => x"b9600800",  1352 => x"b9801000",
     1353 => x"37830014",  1354 => x"f8002639",  1355 => x"b9600800",
     1356 => x"f80034a9",  1357 => x"2b9d0004",  1358 => x"2b8b000c",
     1359 => x"2b8c0008",  1360 => x"379c0020",  1361 => x"c3a00000",
     1362 => x"379cfff8",  1363 => x"5b8b0008",  1364 => x"5b9d0004",
     1365 => x"3402001c",  1366 => x"b8201800",  1367 => x"340b0000",
     1368 => x"3405fffc",  1369 => x"34040003",  1370 => x"e0000009",
     1371 => x"3421ffd0",  1372 => x"202600ff",  1373 => x"50860002",
     1374 => x"e0000008",  1375 => x"bc220800",  1376 => x"34630001",
     1377 => x"b9615800",  1378 => x"3442fffc",  1379 => x"40610000",
     1380 => x"44200007",  1381 => x"5c45fff6",  1382 => x"78010001",
     1383 => x"78020001",  1384 => x"38211e44",  1385 => x"38423d78",
     1386 => x"f800260a",  1387 => x"b9600800",  1388 => x"2b9d0004",
     1389 => x"2b8b0008",  1390 => x"379c0008",  1391 => x"c3a00000",
     1392 => x"379cfffc",  1393 => x"5b9d0004",  1394 => x"34030001",
     1395 => x"34010003",  1396 => x"34020000",  1397 => x"f80039e8",
     1398 => x"34010000",  1399 => x"34020001",  1400 => x"f8003b95",
     1401 => x"34010000",  1402 => x"2b9d0004",  1403 => x"379c0004",
     1404 => x"c3a00000",  1405 => x"379cfff4",  1406 => x"5b8b000c",
     1407 => x"5b8c0008",  1408 => x"5b9d0004",  1409 => x"34010000",
     1410 => x"b8406000",  1411 => x"f8003abf",  1412 => x"45800005",
     1413 => x"642c0000",  1414 => x"c80c6000",  1415 => x"398c0001",
     1416 => x"e000000f",  1417 => x"780b0001",  1418 => x"396b4f20",
     1419 => x"5c2c0004",  1420 => x"59600000",  1421 => x"340cffff",
     1422 => x"e0000009",  1423 => x"29610000",  1424 => x"340c0001",
     1425 => x"5c200006",  1426 => x"78020001",  1427 => x"34010003",
     1428 => x"384243d8",  1429 => x"f8002db9",  1430 => x"596c0000",
     1431 => x"b9800800",  1432 => x"2b9d0004",  1433 => x"2b8b000c",
     1434 => x"2b8c0008",  1435 => x"379c000c",  1436 => x"c3a00000",
     1437 => x"34010000",  1438 => x"c3a00000",  1439 => x"379cfffc",
     1440 => x"5b9d0004",  1441 => x"34010000",  1442 => x"34020001",
     1443 => x"f8003b6a",  1444 => x"34010000",  1445 => x"2b9d0004",
     1446 => x"379c0004",  1447 => x"c3a00000",  1448 => x"379cfffc",
     1449 => x"5b9d0004",  1450 => x"282102c8",  1451 => x"28210010",
     1452 => x"2823000c",  1453 => x"44430004",  1454 => x"5822000c",
     1455 => x"b8400800",  1456 => x"f8002bd8",  1457 => x"34010000",
     1458 => x"2b9d0004",  1459 => x"379c0004",  1460 => x"c3a00000",
     1461 => x"379cfffc",  1462 => x"5b9d0004",  1463 => x"f8002bca",
     1464 => x"34020001",  1465 => x"5c200003",  1466 => x"f8003b43",
     1467 => x"7c220000",  1468 => x"b8400800",  1469 => x"2b9d0004",
     1470 => x"379c0004",  1471 => x"c3a00000",  1472 => x"379cfff8",
     1473 => x"5b8b0008",  1474 => x"5b9d0004",  1475 => x"b8202800",
     1476 => x"b8220800",  1477 => x"b8402000",  1478 => x"b8605800",
     1479 => x"44200005",  1480 => x"34010001",  1481 => x"b8a01000",
     1482 => x"b8801800",  1483 => x"f8002b2c",  1484 => x"45600005",
     1485 => x"1562001f",  1486 => x"34010002",  1487 => x"b9601800",
     1488 => x"f8002b27",  1489 => x"34010000",  1490 => x"2b9d0004",
     1491 => x"2b8b0008",  1492 => x"379c0008",  1493 => x"c3a00000",
     1494 => x"379cfffc",  1495 => x"5b9d0004",  1496 => x"b8201000",
     1497 => x"3401ffff",  1498 => x"f8003a79",  1499 => x"34010000",
     1500 => x"2b9d0004",  1501 => x"379c0004",  1502 => x"c3a00000",
     1503 => x"379cff24",  1504 => x"5b8b0014",  1505 => x"5b8c0010",
     1506 => x"5b8d000c",  1507 => x"5b8e0008",  1508 => x"5b9d0004",
     1509 => x"b8406000",  1510 => x"28220330",  1511 => x"b8807000",
     1512 => x"37810018",  1513 => x"b8605800",  1514 => x"b8a06800",
     1515 => x"fbfffe4d",  1516 => x"45c00005",  1517 => x"78010001",
     1518 => x"382143d4",  1519 => x"28210000",  1520 => x"59c10000",
     1521 => x"45a00003",  1522 => x"2b8100cc",  1523 => x"59a10000",
     1524 => x"2b82006c",  1525 => x"3401fffd",  1526 => x"44400013",
     1527 => x"45800007",  1528 => x"2b820060",  1529 => x"2b810058",
     1530 => x"b4410800",  1531 => x"2b8200a0",  1532 => x"b4220800",
     1533 => x"59810000",  1534 => x"2b820068",  1535 => x"3401fffd",
     1536 => x"44400009",  1537 => x"34010000",  1538 => x"45600007",
     1539 => x"2b830064",  1540 => x"2b82005c",  1541 => x"b4621000",
     1542 => x"2b8300a4",  1543 => x"b4431000",  1544 => x"59620000",
     1545 => x"2b9d0004",  1546 => x"2b8b0014",  1547 => x"2b8c0010",
     1548 => x"2b8d000c",  1549 => x"2b8e0008",  1550 => x"379c00dc",
     1551 => x"c3a00000",  1552 => x"34010000",  1553 => x"c3a00000",
     1554 => x"34010000",  1555 => x"c3a00000",  1556 => x"379cffec",
     1557 => x"5b8b000c",  1558 => x"5b8c0008",  1559 => x"5b9d0004",
     1560 => x"34040000",  1561 => x"b8406000",  1562 => x"b8605800",
     1563 => x"37820010",  1564 => x"37830014",  1565 => x"34050000",
     1566 => x"5b800014",  1567 => x"5b800010",  1568 => x"fbffffbf",
     1569 => x"34010001",  1570 => x"5d810003",  1571 => x"2b810010",
     1572 => x"e0000002",  1573 => x"2b810014",  1574 => x"59610000",
     1575 => x"34010001",  1576 => x"2b9d0004",  1577 => x"2b8b000c",
     1578 => x"2b8c0008",  1579 => x"379c0014",  1580 => x"c3a00000",
     1581 => x"379cfffc",  1582 => x"5b9d0004",  1583 => x"f80026d9",
     1584 => x"34010000",  1585 => x"2b9d0004",  1586 => x"379c0004",
     1587 => x"c3a00000",  1588 => x"379cfffc",  1589 => x"5b9d0004",
     1590 => x"f80026dd",  1591 => x"34010000",  1592 => x"2b9d0004",
     1593 => x"379c0004",  1594 => x"c3a00000",  1595 => x"379cfffc",
     1596 => x"5b9d0004",  1597 => x"f8002bf6",  1598 => x"f800339a",
     1599 => x"f80033a2",  1600 => x"78010001",  1601 => x"78020001",
     1602 => x"38421ee4",  1603 => x"38211eb4",  1604 => x"f8002530",
     1605 => x"34010000",  1606 => x"2b9d0004",  1607 => x"379c0004",
     1608 => x"c3a00000",  1609 => x"78010001",  1610 => x"38214f24",
     1611 => x"28210000",  1612 => x"c3a00000",  1613 => x"379cfff8",
     1614 => x"5b8b0008",  1615 => x"5b9d0004",  1616 => x"78010001",
     1617 => x"78020001",  1618 => x"38424a5c",  1619 => x"38214758",
     1620 => x"780b0001",  1621 => x"f8001981",  1622 => x"396b43e4",
     1623 => x"34030000",  1624 => x"b9600800",  1625 => x"34020000",
     1626 => x"fbfffe65",  1627 => x"78020001",  1628 => x"3842479c",
     1629 => x"58410000",  1630 => x"f8002b48",  1631 => x"78020001",
     1632 => x"38424f30",  1633 => x"58410000",  1634 => x"296102c8",
     1635 => x"28210010",  1636 => x"58200068",  1637 => x"f8000ae8",
     1638 => x"78010001",  1639 => x"38214f2c",  1640 => x"34020001",
     1641 => x"58220000",  1642 => x"34010000",  1643 => x"2b9d0004",
     1644 => x"2b8b0008",  1645 => x"379c0008",  1646 => x"c3a00000",
     1647 => x"379cfff4",  1648 => x"5b8b000c",  1649 => x"5b8c0008",
     1650 => x"5b9d0004",  1651 => x"780b0001",  1652 => x"396b43e4",
     1653 => x"296102c8",  1654 => x"34020000",  1655 => x"282c0010",
     1656 => x"29810000",  1657 => x"28230034",  1658 => x"b9600800",
     1659 => x"d8600000",  1660 => x"78010001",  1661 => x"34020000",
     1662 => x"340301b8",  1663 => x"59800040",  1664 => x"31800035",
     1665 => x"382144f4",  1666 => x"f8003e48",  1667 => x"78010001",
     1668 => x"38214f2c",  1669 => x"58200000",  1670 => x"0d60010c",
     1671 => x"f8000ac6",  1672 => x"78010001",  1673 => x"38214758",
     1674 => x"f8001995",  1675 => x"34010000",  1676 => x"2b9d0004",
     1677 => x"2b8b000c",  1678 => x"2b8c0008",  1679 => x"379c000c",
     1680 => x"c3a00000",  1681 => x"379cffec",  1682 => x"5b8b0014",
     1683 => x"5b8c0010",  1684 => x"5b8d000c",  1685 => x"5b8e0008",
     1686 => x"5b9d0004",  1687 => x"780b0001",  1688 => x"396b43e4",
     1689 => x"b8206000",  1690 => x"296102c8",  1691 => x"282d0010",
     1692 => x"78010001",  1693 => x"38214f24",  1694 => x"58200000",
     1695 => x"fbffffd0",  1696 => x"34010002",  1697 => x"45810016",
     1698 => x"34020003",  1699 => x"45820026",  1700 => x"34010001",
     1701 => x"5d81002e",  1702 => x"78010001",  1703 => x"31ac0004",
     1704 => x"38214a5c",  1705 => x"340e0006",  1706 => x"316c001d",
     1707 => x"302e0000",  1708 => x"34020000",  1709 => x"34010001",
     1710 => x"34030001",  1711 => x"f80038ae",  1712 => x"29610020",
     1713 => x"2821000c",  1714 => x"302e000e",  1715 => x"b9600800",
     1716 => x"f8001295",  1717 => x"380bea60",  1718 => x"e000001e",
     1719 => x"34010001",  1720 => x"31a10004",  1721 => x"3161001d",
     1722 => x"78010001",  1723 => x"38214a5c",  1724 => x"340effbb",
     1725 => x"302e0000",  1726 => x"34020000",  1727 => x"34010002",
     1728 => x"34030001",  1729 => x"f800389c",  1730 => x"29610020",
     1731 => x"2821000c",  1732 => x"302e000e",  1733 => x"b9600800",
     1734 => x"f8001283",  1735 => x"340b0fa0",  1736 => x"e000000c",
     1737 => x"31a10004",  1738 => x"3161001d",  1739 => x"78010001",
     1740 => x"38214a5c",  1741 => x"3402ffff",  1742 => x"30220000",
     1743 => x"34030001",  1744 => x"34010003",  1745 => x"34020000",
     1746 => x"f800388b",  1747 => x"340b0000",  1748 => x"f8002ad2",
     1749 => x"78020001",  1750 => x"b8207000",  1751 => x"b8400800",
     1752 => x"38211f00",  1753 => x"f800249b",  1754 => x"29a20000",
     1755 => x"780d0001",  1756 => x"39ad1f1c",  1757 => x"28430034",
     1758 => x"78020001",  1759 => x"b8400800",  1760 => x"382143e4",
     1761 => x"34020000",  1762 => x"d8600000",  1763 => x"e000000e",
     1764 => x"f8003a8a",  1765 => x"340103e8",  1766 => x"f8002ac5",
     1767 => x"f8002abf",  1768 => x"c82e1000",  1769 => x"51620006",
     1770 => x"78010001",  1771 => x"38211f0c",  1772 => x"f8002488",
     1773 => x"340bff8c",  1774 => x"e0000008",  1775 => x"b9a00800",
     1776 => x"f8002484",  1777 => x"34010000",  1778 => x"f8003950",
     1779 => x"5c200002",  1780 => x"5d61fff0",  1781 => x"340b0000",
     1782 => x"78010001",  1783 => x"38211b04",  1784 => x"f800247c",
     1785 => x"7d620000",  1786 => x"65810001",  1787 => x"a0410800",
     1788 => x"44200005",  1789 => x"78010001",  1790 => x"38214a5c",
     1791 => x"34020034",  1792 => x"30220000",  1793 => x"78010001",
     1794 => x"38214f24",  1795 => x"582c0000",  1796 => x"b9600800",
     1797 => x"2b9d0004",  1798 => x"2b8b0014",  1799 => x"2b8c0010",
     1800 => x"2b8d000c",  1801 => x"2b8e0008",  1802 => x"379c0014",
     1803 => x"c3a00000",  1804 => x"379cfff0",  1805 => x"5b8b0010",
     1806 => x"5b8c000c",  1807 => x"5b8d0008",  1808 => x"5b9d0004",
     1809 => x"34010000",  1810 => x"f80025b5",  1811 => x"78020001",
     1812 => x"38424f28",  1813 => x"b8205800",  1814 => x"28410000",
     1815 => x"442b0018",  1816 => x"78010001",  1817 => x"38214f2c",
     1818 => x"28210000",  1819 => x"584b0000",  1820 => x"65620000",
     1821 => x"7c210000",  1822 => x"a0410800",  1823 => x"44200005",
     1824 => x"fbffff4f",  1825 => x"78010001",  1826 => x"38211f20",
     1827 => x"f8002451",  1828 => x"78010001",  1829 => x"38214f2c",
     1830 => x"28210000",  1831 => x"7d6b0000",  1832 => x"64210000",
     1833 => x"a1615800",  1834 => x"45600005",  1835 => x"78010001",
     1836 => x"38211f38",  1837 => x"f8002447",  1838 => x"fbffff1f",
     1839 => x"78010001",  1840 => x"38214f2c",  1841 => x"28210000",
     1842 => x"44200022",  1843 => x"780b0001",  1844 => x"396b43e4",
     1845 => x"29610024",  1846 => x"29620038",  1847 => x"78040001",
     1848 => x"28250008",  1849 => x"3403007c",  1850 => x"b9600800",
     1851 => x"388444c8",  1852 => x"d8a00000",  1853 => x"b8201800",
     1854 => x"4801000f",  1855 => x"29610370",  1856 => x"34210001",
     1857 => x"59610370",  1858 => x"5c60000b",  1859 => x"780d0001",
     1860 => x"f8002a62",  1861 => x"39ad4f30",  1862 => x"29a20000",
     1863 => x"780c0001",  1864 => x"398c479c",  1865 => x"c8220800",
     1866 => x"29820000",  1867 => x"54410009",  1868 => x"e000000f",
     1869 => x"78010001",  1870 => x"382143e4",  1871 => x"28220040",
     1872 => x"fbfffd6f",  1873 => x"78020001",  1874 => x"3842479c",
     1875 => x"58410000",  1876 => x"34010000",  1877 => x"2b9d0004",
     1878 => x"2b8b0010",  1879 => x"2b8c000c",  1880 => x"2b8d0008",
     1881 => x"379c0010",  1882 => x"c3a00000",  1883 => x"f8002a4b",
     1884 => x"59a10000",  1885 => x"34020000",  1886 => x"b9600800",
     1887 => x"34030000",  1888 => x"fbfffd5f",  1889 => x"59810000",
     1890 => x"e3fffff2",  1891 => x"379cffe8",  1892 => x"5b9d0018",
     1893 => x"b8205000",  1894 => x"40610005",  1895 => x"40640000",
     1896 => x"40650001",  1897 => x"40660002",  1898 => x"40670003",
     1899 => x"40680004",  1900 => x"5b810004",  1901 => x"40610006",
     1902 => x"b8404800",  1903 => x"b9401000",  1904 => x"5b810008",
     1905 => x"40610007",  1906 => x"5b81000c",  1907 => x"40610008",
     1908 => x"5b810010",  1909 => x"40610009",  1910 => x"b9201800",
     1911 => x"5b810014",  1912 => x"78010001",  1913 => x"38211f50",
     1914 => x"f80023fa",  1915 => x"2b9d0018",  1916 => x"379c0018",
     1917 => x"c3a00000",  1918 => x"379cffd0",  1919 => x"5b8b0030",
     1920 => x"5b8c002c",  1921 => x"5b8d0028",  1922 => x"5b8e0024",
     1923 => x"5b8f0020",  1924 => x"5b90001c",  1925 => x"5b910018",
     1926 => x"5b920014",  1927 => x"5b930010",  1928 => x"5b94000c",
     1929 => x"5b950008",  1930 => x"5b9d0004",  1931 => x"b8603000",
     1932 => x"b8209800",  1933 => x"b8409000",  1934 => x"78010001",
     1935 => x"b880a800",  1936 => x"38211f88",  1937 => x"ba601000",
     1938 => x"ba401800",  1939 => x"b8c02000",  1940 => x"b8a0a000",
     1941 => x"78110001",  1942 => x"f80023de",  1943 => x"78100001",
     1944 => x"780f0001",  1945 => x"780e0001",  1946 => x"780d0001",
     1947 => x"b8205800",  1948 => x"340c0000",  1949 => x"3a311f9c",
     1950 => x"3a101fa4",  1951 => x"39ef1c28",  1952 => x"39ce1b04",
     1953 => x"39ad19a0",  1954 => x"e0000017",  1955 => x"5cc00006",
     1956 => x"ba200800",  1957 => x"ba601000",  1958 => x"ba401800",
     1959 => x"f80023cd",  1960 => x"b5615800",  1961 => x"b6ac1000",
     1962 => x"40420000",  1963 => x"ba000800",  1964 => x"358c0001",
     1965 => x"f80023c7",  1966 => x"21820003",  1967 => x"b42b5800",
     1968 => x"b9e03000",  1969 => x"5c400005",  1970 => x"2181000f",
     1971 => x"b9c03000",  1972 => x"44220002",  1973 => x"b9a03000",
     1974 => x"b8c00800",  1975 => x"f80023bd",  1976 => x"b5615800",
     1977 => x"2186000f",  1978 => x"4a8cffe9",  1979 => x"44c00005",
     1980 => x"78010001",  1981 => x"38211b04",  1982 => x"f80023b6",
     1983 => x"b42b5800",  1984 => x"b9600800",  1985 => x"2b9d0004",
     1986 => x"2b8b0030",  1987 => x"2b8c002c",  1988 => x"2b8d0028",
     1989 => x"2b8e0024",  1990 => x"2b8f0020",  1991 => x"2b90001c",
     1992 => x"2b910018",  1993 => x"2b920014",  1994 => x"2b930010",
     1995 => x"2b94000c",  1996 => x"2b950008",  1997 => x"379c0030",
     1998 => x"c3a00000",  1999 => x"379cffb8",  2000 => x"5b8b0048",
     2001 => x"5b8c0044",  2002 => x"5b8d0040",  2003 => x"5b8e003c",
     2004 => x"5b8f0038",  2005 => x"5b900034",  2006 => x"5b910030",
     2007 => x"5b92002c",  2008 => x"5b930028",  2009 => x"5b940024",
     2010 => x"5b950020",  2011 => x"5b96001c",  2012 => x"5b970018",
     2013 => x"5b980014",  2014 => x"5b9d0010",  2015 => x"b8608000",
     2016 => x"40430001",  2017 => x"b8206000",  2018 => x"34010002",
     2019 => x"2063000f",  2020 => x"b8406800",  2021 => x"404e0000",
     2022 => x"44610006",  2023 => x"78010001",  2024 => x"b9801000",
     2025 => x"38211fac",  2026 => x"f800238a",  2027 => x"e000013f",
     2028 => x"40450002",  2029 => x"40460003",  2030 => x"21ce000f",
     2031 => x"3ca50008",  2032 => x"78010001",  2033 => x"b8c52800",
     2034 => x"41a60004",  2035 => x"34030002",  2036 => x"b9c02000",
     2037 => x"344b0022",  2038 => x"38211fcc",  2039 => x"b9801000",
     2040 => x"f800237c",  2041 => x"41a2000c",  2042 => x"41a1000d",
     2043 => x"41a4000e",  2044 => x"41a30006",  2045 => x"3c420018",
     2046 => x"3c210010",  2047 => x"41a60007",  2048 => x"41a5000f",
     2049 => x"3c840008",  2050 => x"b8220800",  2051 => x"3c630008",
     2052 => x"b8812000",  2053 => x"78010001",  2054 => x"b8c31800",
     2055 => x"b8a42000",  2056 => x"b9801000",  2057 => x"38211ff8",
     2058 => x"f800236a",  2059 => x"78020001",  2060 => x"b9800800",
     2061 => x"3842201c",  2062 => x"35a30014",  2063 => x"fbffff54",
     2064 => x"41a3001e",  2065 => x"41a4001f",  2066 => x"41a50021",
     2067 => x"3c630008",  2068 => x"78010001",  2069 => x"b8831800",
     2070 => x"41a40020",  2071 => x"38212024",  2072 => x"b9801000",
     2073 => x"f800235b",  2074 => x"3401000c",  2075 => x"55c100d1",
     2076 => x"78010001",  2077 => x"3dce0002",  2078 => x"38213da8",
     2079 => x"b42e0800",  2080 => x"28210000",  2081 => x"c0200000",
     2082 => x"78010001",  2083 => x"b9801000",  2084 => x"38212050",
     2085 => x"f800234f",  2086 => x"41620002",  2087 => x"41610003",
     2088 => x"41640004",  2089 => x"3c420018",  2090 => x"3c210010",
     2091 => x"3c840008",  2092 => x"b8220800",  2093 => x"b8812000",
     2094 => x"41620006",  2095 => x"41610007",  2096 => x"41650008",
     2097 => x"3c420018",  2098 => x"3c210010",  2099 => x"3ca50008",
     2100 => x"b8220800",  2101 => x"b8a12800",  2102 => x"78030001",
     2103 => x"78010001",  2104 => x"41670005",  2105 => x"41660009",
     2106 => x"38212068",  2107 => x"b9801000",  2108 => x"38632078",
     2109 => x"e000001c",  2110 => x"78010001",  2111 => x"b9801000",
     2112 => x"38212084",  2113 => x"f8002333",  2114 => x"41620002",
     2115 => x"41610003",  2116 => x"41640004",  2117 => x"3c420018",
     2118 => x"3c210010",  2119 => x"3c840008",  2120 => x"b8220800",
     2121 => x"b8812000",  2122 => x"41620006",  2123 => x"41610007",
     2124 => x"41650008",  2125 => x"3c420018",  2126 => x"3c210010",
     2127 => x"3ca50008",  2128 => x"b8220800",  2129 => x"41670005",
     2130 => x"41660009",  2131 => x"b8a12800",  2132 => x"78030001",
     2133 => x"78010001",  2134 => x"38212068",  2135 => x"b9801000",
     2136 => x"386320a0",  2137 => x"b8e42000",  2138 => x"b8c52800",
     2139 => x"f8002319",  2140 => x"e000008e",  2141 => x"78010001",
     2142 => x"b9801000",  2143 => x"382120b0",  2144 => x"f8002314",
     2145 => x"41620002",  2146 => x"41610003",  2147 => x"41640004",
     2148 => x"3c420018",  2149 => x"3c210010",  2150 => x"3c840008",
     2151 => x"b8220800",  2152 => x"b8812000",  2153 => x"41620006",
     2154 => x"41610007",  2155 => x"41650008",  2156 => x"3c420018",
     2157 => x"3c210010",  2158 => x"3ca50008",  2159 => x"b8220800",
     2160 => x"b8a12800",  2161 => x"78030001",  2162 => x"78010001",
     2163 => x"41670005",  2164 => x"41660009",  2165 => x"38212068",
     2166 => x"b9801000",  2167 => x"386320cc",  2168 => x"e3ffffe1",
     2169 => x"78010001",  2170 => x"b9801000",  2171 => x"382120dc",
     2172 => x"f80022f8",  2173 => x"41620002",  2174 => x"41610003",
     2175 => x"41640004",  2176 => x"3c420018",  2177 => x"3c210010",
     2178 => x"3c840008",  2179 => x"b8220800",  2180 => x"b8812000",
     2181 => x"41620006",  2182 => x"41610007",  2183 => x"41650008",
     2184 => x"3c420018",  2185 => x"3c210010",  2186 => x"41670005",
     2187 => x"41660009",  2188 => x"3ca50008",  2189 => x"b8220800",
     2190 => x"780e0001",  2191 => x"39ce20f8",  2192 => x"b8a12800",
     2193 => x"78010001",  2194 => x"b9801000",  2195 => x"b9c01800",
     2196 => x"b8e42000",  2197 => x"b8c52800",  2198 => x"38212068",
     2199 => x"f80022dd",  2200 => x"3563000a",  2201 => x"b9800800",
     2202 => x"b9c01000",  2203 => x"fbfffec8",  2204 => x"340b0036",
     2205 => x"e0000080",  2206 => x"78010001",  2207 => x"b9801000",
     2208 => x"3821210c",  2209 => x"f80022d3",  2210 => x"41620002",
     2211 => x"41610003",  2212 => x"41640004",  2213 => x"3c420018",
     2214 => x"3c210010",  2215 => x"3c840008",  2216 => x"b8220800",
     2217 => x"b8812000",  2218 => x"41620006",  2219 => x"41610007",
     2220 => x"41650008",  2221 => x"3c420018",  2222 => x"3c210010",
     2223 => x"41670005",  2224 => x"41660009",  2225 => x"3ca50008",
     2226 => x"b8220800",  2227 => x"b8a12800",  2228 => x"78030001",
     2229 => x"78010001",  2230 => x"b8e42000",  2231 => x"b8c52800",
     2232 => x"b9801000",  2233 => x"38632128",  2234 => x"38212068",
     2235 => x"f80022b9",  2236 => x"41660010",  2237 => x"41670011",
     2238 => x"4165000f",  2239 => x"4164000e",  2240 => x"3cc60008",
     2241 => x"78010001",  2242 => x"78030001",  2243 => x"b8e63000",
     2244 => x"b9801000",  2245 => x"38632154",  2246 => x"38212140",
     2247 => x"f80022ad",  2248 => x"4163000d",  2249 => x"41640012",
     2250 => x"78010001",  2251 => x"b9801000",  2252 => x"38212178",
     2253 => x"f80022a7",  2254 => x"41610018",  2255 => x"41640013",
     2256 => x"41650014",  2257 => x"41660015",  2258 => x"41670016",
     2259 => x"41680017",  2260 => x"5b810004",  2261 => x"41610019",
     2262 => x"78030001",  2263 => x"b9801000",  2264 => x"5b810008",
     2265 => x"4161001a",  2266 => x"386321d0",  2267 => x"340b0040",
     2268 => x"5b81000c",  2269 => x"78010001",  2270 => x"382121a0",
     2271 => x"f8002295",  2272 => x"e000003d",  2273 => x"78010001",
     2274 => x"b9801000",  2275 => x"382121f0",  2276 => x"f8002290",
     2277 => x"78020001",  2278 => x"b9800800",  2279 => x"3842220c",
     2280 => x"b9601800",  2281 => x"fbfffe7a",  2282 => x"340b002c",
     2283 => x"e0000032",  2284 => x"340b0022",  2285 => x"e0000030",
     2286 => x"55f70009",  2287 => x"78010001",  2288 => x"b9801000",
     2289 => x"ba001800",  2290 => x"b9602000",  2291 => x"b9e02800",
     2292 => x"38212228",  2293 => x"f800227f",  2294 => x"e0000034",
     2295 => x"b5ab7000",  2296 => x"41d60002",  2297 => x"41c10003",
     2298 => x"41c30000",  2299 => x"3ed60008",  2300 => x"41c40001",
     2301 => x"b836b000",  2302 => x"41c10008",  2303 => x"41c50004",
     2304 => x"41c60005",  2305 => x"41c70006",  2306 => x"41c80007",
     2307 => x"5b810004",  2308 => x"41c10009",  2309 => x"3c630008",
     2310 => x"36d10004",  2311 => x"5b810008",  2312 => x"b8831800",
     2313 => x"baa00800",  2314 => x"b9801000",  2315 => x"ba202000",
     2316 => x"f8002268",  2317 => x"4df10007",  2318 => x"ba400800",
     2319 => x"b9801000",  2320 => x"ba201800",  2321 => x"b9e02000",
     2322 => x"f8002262",  2323 => x"e0000008",  2324 => x"b9800800",
     2325 => x"ba801000",  2326 => x"ba601800",  2327 => x"35c4000a",
     2328 => x"36c5fffa",  2329 => x"fbfffe65",  2330 => x"ba207800",
     2331 => x"b56f5800",  2332 => x"e000000b",  2333 => x"78150001",
     2334 => x"78140001",  2335 => x"78130001",  2336 => x"78120001",
     2337 => x"34180002",  2338 => x"34170009",  2339 => x"3ab5224c",
     2340 => x"3a9422b8",  2341 => x"3a7322c0",  2342 => x"3a52228c",
     2343 => x"4d700003",  2344 => x"ca0b7800",  2345 => x"49f8ffc5",
     2346 => x"78020001",  2347 => x"78030001",  2348 => x"b9800800",
     2349 => x"384222cc",  2350 => x"386322d4",  2351 => x"b9a02000",
     2352 => x"ba002800",  2353 => x"fbfffe4d",  2354 => x"2b9d0010",
     2355 => x"2b8b0048",  2356 => x"2b8c0044",  2357 => x"2b8d0040",
     2358 => x"2b8e003c",  2359 => x"2b8f0038",  2360 => x"2b900034",
     2361 => x"2b910030",  2362 => x"2b92002c",  2363 => x"2b930028",
     2364 => x"2b940024",  2365 => x"2b950020",  2366 => x"2b96001c",
     2367 => x"2b970018",  2368 => x"2b980014",  2369 => x"379c0048",
     2370 => x"c3a00000",  2371 => x"379cfff0",  2372 => x"5b8b0010",
     2373 => x"5b8c000c",  2374 => x"5b8d0008",  2375 => x"5b9d0004",
     2376 => x"b8205800",  2377 => x"b8406800",  2378 => x"b8606000",
     2379 => x"4480000f",  2380 => x"2881000c",  2381 => x"78070001",
     2382 => x"28850000",  2383 => x"28860004",  2384 => x"38e73cbc",
     2385 => x"5c200003",  2386 => x"78070001",  2387 => x"38e722dc",
     2388 => x"78010001",  2389 => x"382122e8",  2390 => x"b9601000",
     2391 => x"b8a01800",  2392 => x"b8a02000",  2393 => x"f800221b",
     2394 => x"b9600800",  2395 => x"b9a01000",  2396 => x"b9801800",
     2397 => x"fbfffe72",  2398 => x"34010000",  2399 => x"2b9d0004",
     2400 => x"2b8b0010",  2401 => x"2b8c000c",  2402 => x"2b8d0008",
     2403 => x"379c0010",  2404 => x"c3a00000",  2405 => x"379cffe8",
     2406 => x"5b8b0018",  2407 => x"5b8c0014",  2408 => x"5b8d0010",
     2409 => x"5b8e000c",  2410 => x"5b8f0008",  2411 => x"5b9d0004",
     2412 => x"282d0000",  2413 => x"b8207800",  2414 => x"282e0004",
     2415 => x"b8406000",  2416 => x"340b0000",  2417 => x"34010000",
     2418 => x"34040000",  2419 => x"544d0006",  2420 => x"b9a00800",
     2421 => x"f8003a76",  2422 => x"882c1000",  2423 => x"b9602000",
     2424 => x"c9a26800",  2425 => x"34030000",  2426 => x"34020001",
     2427 => x"e000000b",  2428 => x"3d850001",  2429 => x"3d6b0001",
     2430 => x"f5856000",  2431 => x"3c630001",  2432 => x"b58b5800",
     2433 => x"b8a06000",  2434 => x"3c450001",  2435 => x"f4451000",
     2436 => x"b4431800",  2437 => x"b8a01000",  2438 => x"1565001f",
     2439 => x"c8ac3000",  2440 => x"f4c53000",  2441 => x"c8ab2800",
     2442 => x"c8a62800",  2443 => x"00a5001f",  2444 => x"34060001",
     2445 => x"55ab0004",  2446 => x"5dab0002",  2447 => x"55cc0002",
     2448 => x"34060000",  2449 => x"a0a63000",  2450 => x"5cc0ffea",
     2451 => x"556d000d",  2452 => x"5d6d0002",  2453 => x"558e000b",
     2454 => x"c9cc2800",  2455 => x"f4ae7000",  2456 => x"c9ab6800",
     2457 => x"c9ae6800",  2458 => x"b8a07000",  2459 => x"b4822800",
     2460 => x"f4852000",  2461 => x"b4230800",  2462 => x"b4810800",
     2463 => x"b8a02000",  2464 => x"3c65001f",  2465 => x"00420001",
     2466 => x"00630001",  2467 => x"b8a21000",  2468 => x"b8622800",
     2469 => x"44a00006",  2470 => x"3d65001f",  2471 => x"018c0001",
     2472 => x"016b0001",  2473 => x"b8ac6000",  2474 => x"e3ffffe9",
     2475 => x"59e10000",  2476 => x"b9c00800",  2477 => x"59e40004",
     2478 => x"2b9d0004",  2479 => x"2b8b0018",  2480 => x"2b8c0014",
     2481 => x"2b8d0010",  2482 => x"2b8e000c",  2483 => x"2b8f0008",
     2484 => x"379c0018",  2485 => x"c3a00000",  2486 => x"379cfff8",
     2487 => x"5b8b0008",  2488 => x"5b9d0004",  2489 => x"b8405800",
     2490 => x"f80027ec",  2491 => x"b42b0800",  2492 => x"5c200002",
     2493 => x"34010001",  2494 => x"2b9d0004",  2495 => x"2b8b0008",
     2496 => x"379c0008",  2497 => x"c3a00000",  2498 => x"379cfff8",
     2499 => x"5b8b0008",  2500 => x"5b9d0004",  2501 => x"78040001",
     2502 => x"b8405800",  2503 => x"78050001",  2504 => x"34020006",
     2505 => x"34030001",  2506 => x"388423b4",  2507 => x"38a53ddc",
     2508 => x"b9603000",  2509 => x"fbfffb53",  2510 => x"45600005",
     2511 => x"1562001f",  2512 => x"34010002",  2513 => x"b9601800",
     2514 => x"f8002725",  2515 => x"34010000",  2516 => x"2b9d0004",
     2517 => x"2b8b0008",  2518 => x"379c0008",  2519 => x"c3a00000",
     2520 => x"379cfff4",  2521 => x"5b8b000c",  2522 => x"5b8c0008",
     2523 => x"5b9d0004",  2524 => x"b8206000",  2525 => x"b8405800",
     2526 => x"b8603000",  2527 => x"44600008",  2528 => x"78040001",
     2529 => x"78050001",  2530 => x"34020006",  2531 => x"34030001",
     2532 => x"388423c0",  2533 => x"38a53df4",  2534 => x"fbfffb3a",
     2535 => x"b9800800",  2536 => x"b9601000",  2537 => x"fbffffd9",
     2538 => x"2b9d0004",  2539 => x"2b8b000c",  2540 => x"2b8c0008",
     2541 => x"379c000c",  2542 => x"c3a00000",  2543 => x"379cfff0",
     2544 => x"5b8b0010",  2545 => x"5b8c000c",  2546 => x"5b8d0008",
     2547 => x"5b9d0004",  2548 => x"b8206800",  2549 => x"44400012",
     2550 => x"284b0000",  2551 => x"284c0004",  2552 => x"34040003",
     2553 => x"1561001f",  2554 => x"b9601000",  2555 => x"b9801800",
     2556 => x"f800273c",  2557 => x"78040001",  2558 => x"78050001",
     2559 => x"b9a00800",  2560 => x"34020006",  2561 => x"34030001",
     2562 => x"388423ec",  2563 => x"38a53e08",  2564 => x"b9603000",
     2565 => x"b9803800",  2566 => x"fbfffb1a",  2567 => x"34010000",
     2568 => x"2b9d0004",  2569 => x"2b8b0010",  2570 => x"2b8c000c",
     2571 => x"2b8d0008",  2572 => x"379c0010",  2573 => x"c3a00000",
     2574 => x"379cffe8",  2575 => x"5b8b000c",  2576 => x"5b8c0008",
     2577 => x"5b9d0004",  2578 => x"b8405800",  2579 => x"b8206000",
     2580 => x"37820018",  2581 => x"37810010",  2582 => x"f8002742",
     2583 => x"78020001",  2584 => x"38424e9c",  2585 => x"2b860014",
     2586 => x"2b870018",  2587 => x"28410000",  2588 => x"59660000",
     2589 => x"59670004",  2590 => x"20210001",  2591 => x"5c200009",
     2592 => x"78040001",  2593 => x"78050001",  2594 => x"b9800800",
     2595 => x"34020006",  2596 => x"34030002",  2597 => x"388423ec",
     2598 => x"38a53e18",  2599 => x"fbfffaf9",  2600 => x"34010000",
     2601 => x"2b9d0004",  2602 => x"2b8b000c",  2603 => x"2b8c0008",
     2604 => x"379c0018",  2605 => x"c3a00000",  2606 => x"379cffb4",
     2607 => x"5b8b001c",  2608 => x"5b8c0018",  2609 => x"5b8d0014",
     2610 => x"5b8e0010",  2611 => x"5b8f000c",  2612 => x"5b900008",
     2613 => x"5b9d0004",  2614 => x"28300058",  2615 => x"378c0040",
     2616 => x"b8407800",  2617 => x"b8206800",  2618 => x"78020001",
     2619 => x"340188f7",  2620 => x"b8607000",  2621 => x"0f81004c",
     2622 => x"38423d70",  2623 => x"b9800800",  2624 => x"34030006",
     2625 => x"b8805800",  2626 => x"f8003a0a",  2627 => x"b9801000",
     2628 => x"ba000800",  2629 => x"b9e01800",  2630 => x"b9c02000",
     2631 => x"37850020",  2632 => x"f8001df0",  2633 => x"b8206000",
     2634 => x"45600011",  2635 => x"2b81003c",  2636 => x"2b870024",
     2637 => x"2b880028",  2638 => x"78040001",  2639 => x"78050001",
     2640 => x"5961000c",  2641 => x"59670000",  2642 => x"59680004",
     2643 => x"59600008",  2644 => x"b9a00800",  2645 => x"34020005",
     2646 => x"34030002",  2647 => x"388423fc",  2648 => x"38a53e28",
     2649 => x"b9803000",  2650 => x"fbfffac6",  2651 => x"4c0c0010",
     2652 => x"78010001",  2653 => x"38214e9c",  2654 => x"28220000",
     2655 => x"29a10018",  2656 => x"b8410800",  2657 => x"00210014",
     2658 => x"34020001",  2659 => x"2021000f",  2660 => x"50410007",
     2661 => x"78010001",  2662 => x"3821241c",  2663 => x"b9e01000",
     2664 => x"b9c01800",  2665 => x"b9602000",  2666 => x"fbfffed9",
     2667 => x"b9800800",  2668 => x"2b9d0004",  2669 => x"2b8b001c",
     2670 => x"2b8c0018",  2671 => x"2b8d0014",  2672 => x"2b8e0010",
     2673 => x"2b8f000c",  2674 => x"2b900008",  2675 => x"379c004c",
     2676 => x"c3a00000",  2677 => x"379cffbc",  2678 => x"5b8b0014",
     2679 => x"5b8c0010",  2680 => x"5b8d000c",  2681 => x"5b8e0008",
     2682 => x"5b9d0004",  2683 => x"b8207000",  2684 => x"28210058",
     2685 => x"b8602800",  2686 => x"b8406800",  2687 => x"b8805800",
     2688 => x"37820038",  2689 => x"b8a02000",  2690 => x"b9a01800",
     2691 => x"37850018",  2692 => x"f8001d1c",  2693 => x"b8206000",
     2694 => x"4560000b",  2695 => x"2b81001c",  2696 => x"59610000",
     2697 => x"2b810020",  2698 => x"59610004",  2699 => x"2b810024",
     2700 => x"59610008",  2701 => x"2b810034",  2702 => x"5961000c",
     2703 => x"2b810030",  2704 => x"59610010",  2705 => x"4c0c0010",
     2706 => x"78040001",  2707 => x"38844e9c",  2708 => x"28820000",
     2709 => x"29c10018",  2710 => x"b8410800",  2711 => x"00210014",
     2712 => x"34020001",  2713 => x"2021000f",  2714 => x"50410007",
     2715 => x"78010001",  2716 => x"38212424",  2717 => x"b9a01000",
     2718 => x"b9801800",  2719 => x"b9602000",  2720 => x"fbfffea3",
     2721 => x"b9800800",  2722 => x"2b9d0004",  2723 => x"2b8b0014",
     2724 => x"2b8c0010",  2725 => x"2b8d000c",  2726 => x"2b8e0008",
     2727 => x"379c0044",  2728 => x"c3a00000",  2729 => x"379cfffc",
     2730 => x"5b9d0004",  2731 => x"28210058",  2732 => x"f8001ca1",
     2733 => x"34010000",  2734 => x"2b9d0004",  2735 => x"379c0004",
     2736 => x"c3a00000",  2737 => x"379cffd8",  2738 => x"5b8b0010",
     2739 => x"5b8c000c",  2740 => x"5b8d0008",  2741 => x"5b9d0004",
     2742 => x"b8205800",  2743 => x"28210058",  2744 => x"44200002",
     2745 => x"f8001c94",  2746 => x"b9600800",  2747 => x"f8000cfb",
     2748 => x"378c0014",  2749 => x"340188f7",  2750 => x"78020001",
     2751 => x"0f810020",  2752 => x"38423d70",  2753 => x"b9800800",
     2754 => x"34030006",  2755 => x"f8003989",  2756 => x"b9801800",
     2757 => x"34010001",  2758 => x"34020000",  2759 => x"f8001c4e",
     2760 => x"b8206000",  2761 => x"4420000e",  2762 => x"378d0024",
     2763 => x"b9a01000",  2764 => x"f8001c3a",  2765 => x"b9a01000",
     2766 => x"34030006",  2767 => x"35610060",  2768 => x"f800397c",
     2769 => x"3561004c",  2770 => x"596c0058",  2771 => x"b9a01000",
     2772 => x"34030006",  2773 => x"f8003977",  2774 => x"596c0044",
     2775 => x"34010000",  2776 => x"2b9d0004",  2777 => x"2b8b0010",
     2778 => x"2b8c000c",  2779 => x"2b8d0008",  2780 => x"379c0028",
     2781 => x"c3a00000",  2782 => x"379cfff8",  2783 => x"5b8b0008",
     2784 => x"5b9d0004",  2785 => x"78040001",  2786 => x"78050001",
     2787 => x"34020002",  2788 => x"34030002",  2789 => x"38842510",
     2790 => x"38a53e88",  2791 => x"b8205800",  2792 => x"fbfffa38",
     2793 => x"296302c8",  2794 => x"28610010",  2795 => x"28220064",
     2796 => x"34010000",  2797 => x"44400010",  2798 => x"34010001",
     2799 => x"59610004",  2800 => x"1061000b",  2801 => x"4062000c",
     2802 => x"29640028",  2803 => x"bc411000",  2804 => x"28830018",
     2805 => x"084203e8",  2806 => x"b9600800",  2807 => x"d8600000",
     2808 => x"596102d4",  2809 => x"296102c8",  2810 => x"28210010",
     2811 => x"58200064",  2812 => x"34010001",  2813 => x"2b9d0004",
     2814 => x"2b8b0008",  2815 => x"379c0008",  2816 => x"c3a00000",
     2817 => x"379cfff4",  2818 => x"5b8b000c",  2819 => x"5b8c0008",
     2820 => x"5b9d0004",  2821 => x"78040001",  2822 => x"78050001",
     2823 => x"b8606000",  2824 => x"34020002",  2825 => x"34030002",
     2826 => x"38842510",  2827 => x"38a53e9c",  2828 => x"b8205800",
     2829 => x"fbfffa13",  2830 => x"29820024",  2831 => x"296102c8",
     2832 => x"20430003",  2833 => x"28210010",  2834 => x"7c640000",
     2835 => x"58240038",  2836 => x"20440008",  2837 => x"20420004",
     2838 => x"7c840000",  2839 => x"7c420000",  2840 => x"30230035",
     2841 => x"58220044",  2842 => x"58240040",  2843 => x"29610020",
     2844 => x"28220010",  2845 => x"296102c8",  2846 => x"2c210008",
     2847 => x"0c41002c",  2848 => x"2b9d0004",  2849 => x"2b8b000c",
     2850 => x"2b8c0008",  2851 => x"379c000c",  2852 => x"c3a00000",
     2853 => x"379cfff8",  2854 => x"5b8b0008",  2855 => x"5b9d0004",
     2856 => x"282202c8",  2857 => x"78040001",  2858 => x"78050001",
     2859 => x"284b0010",  2860 => x"34030002",  2861 => x"34020002",
     2862 => x"38842510",  2863 => x"38a53ed4",  2864 => x"fbfff9f0",
     2865 => x"34010000",  2866 => x"31600005",  2867 => x"2b9d0004",
     2868 => x"2b8b0008",  2869 => x"379c0008",  2870 => x"c3a00000",
     2871 => x"379cfff8",  2872 => x"5b8b0008",  2873 => x"5b9d0004",
     2874 => x"78040001",  2875 => x"78050001",  2876 => x"b8205800",
     2877 => x"34020002",  2878 => x"34010000",  2879 => x"34030002",
     2880 => x"38842510",  2881 => x"38a53ee4",  2882 => x"fbfff9de",
     2883 => x"29610024",  2884 => x"44200006",  2885 => x"34020000",
     2886 => x"34030001",  2887 => x"34040002",  2888 => x"34060003",
     2889 => x"e000001f",  2890 => x"29610000",  2891 => x"29620040",
     2892 => x"58220014",  2893 => x"e000001d",  2894 => x"29650000",
     2895 => x"08410374",  2896 => x"b4a10800",  2897 => x"29650040",
     2898 => x"58250014",  2899 => x"28250368",  2900 => x"5ca30010",
     2901 => x"4025001d",  2902 => x"44a30004",  2903 => x"282102c8",
     2904 => x"5ca40009",  2905 => x"e0000005",  2906 => x"282102c8",
     2907 => x"28210010",  2908 => x"30230004",  2909 => x"e000000a",
     2910 => x"28210010",  2911 => x"30240004",  2912 => x"e0000007",
     2913 => x"28210010",  2914 => x"30260004",  2915 => x"e0000004",
     2916 => x"282102c8",  2917 => x"28210010",  2918 => x"30200004",
     2919 => x"34420001",  2920 => x"29610024",  2921 => x"4822ffe5",
     2922 => x"34010000",  2923 => x"2b9d0004",  2924 => x"2b8b0008",
     2925 => x"379c0008",  2926 => x"c3a00000",  2927 => x"379cfff4",
     2928 => x"5b8b000c",  2929 => x"5b8c0008",  2930 => x"5b9d0004",
     2931 => x"282202c8",  2932 => x"78040001",  2933 => x"78050001",
     2934 => x"284b0010",  2935 => x"34030002",  2936 => x"34020002",
     2937 => x"38842510",  2938 => x"38a53eec",  2939 => x"b8206000",
     2940 => x"fbfff9a4",  2941 => x"41630004",  2942 => x"3401012c",
     2943 => x"59610028",  2944 => x"34020001",  2945 => x"34010bb8",
     2946 => x"59610030",  2947 => x"59600008",  2948 => x"31600035",
     2949 => x"59600040",  2950 => x"59620014",  2951 => x"20630003",
     2952 => x"29610000",  2953 => x"5c620004",  2954 => x"28230034",
     2955 => x"b9800800",  2956 => x"e0000004",  2957 => x"28230034",
     2958 => x"34020000",  2959 => x"b9800800",  2960 => x"d8600000",
     2961 => x"34010000",  2962 => x"2b9d0004",  2963 => x"2b8b000c",
     2964 => x"2b8c0008",  2965 => x"379c000c",  2966 => x"c3a00000",
     2967 => x"379cfff0",  2968 => x"5b8b0010",  2969 => x"5b8c000c",
     2970 => x"5b8d0008",  2971 => x"5b9d0004",  2972 => x"78040001",
     2973 => x"78050001",  2974 => x"2c2d0002",  2975 => x"b8205800",
     2976 => x"b8406000",  2977 => x"34010000",  2978 => x"34020002",
     2979 => x"34030002",  2980 => x"38842510",  2981 => x"38a53e38",
     2982 => x"fbfff97a",  2983 => x"34010040",  2984 => x"4c2d0004",
     2985 => x"b9600800",  2986 => x"b9801000",  2987 => x"f8000466",
     2988 => x"2b9d0004",  2989 => x"2b8b0010",  2990 => x"2b8c000c",
     2991 => x"2b8d0008",  2992 => x"379c0010",  2993 => x"c3a00000",
     2994 => x"379cfff8",  2995 => x"5b8b0008",  2996 => x"5b9d0004",
     2997 => x"78040001",  2998 => x"78050001",  2999 => x"34020002",
     3000 => x"34030002",  3001 => x"38842510",  3002 => x"38a53e4c",
     3003 => x"b8205800",  3004 => x"fbfff964",  3005 => x"296102c8",
     3006 => x"34020040",  3007 => x"28210010",  3008 => x"40210004",
     3009 => x"44200006",  3010 => x"34030002",  3011 => x"44230004",
     3012 => x"b9600800",  3013 => x"f8000409",  3014 => x"3402004e",
     3015 => x"b8400800",  3016 => x"2b9d0004",  3017 => x"2b8b0008",
     3018 => x"379c0008",  3019 => x"c3a00000",  3020 => x"379cfff4",
     3021 => x"5b8b000c",  3022 => x"5b8c0008",  3023 => x"5b9d0004",
     3024 => x"78040001",  3025 => x"78050001",  3026 => x"34030002",
     3027 => x"b8406000",  3028 => x"38842510",  3029 => x"34020002",
     3030 => x"38a53e60",  3031 => x"b8205800",  3032 => x"fbfff948",
     3033 => x"296102c8",  3034 => x"34030000",  3035 => x"28210010",
     3036 => x"28210008",  3037 => x"44200007",  3038 => x"35630094",
     3039 => x"59800008",  3040 => x"b9600800",  3041 => x"b9801000",
     3042 => x"f80005c9",  3043 => x"34030001",  3044 => x"b8600800",
     3045 => x"2b9d0004",  3046 => x"2b8b000c",  3047 => x"2b8c0008",
     3048 => x"379c000c",  3049 => x"c3a00000",  3050 => x"379cfff8",
     3051 => x"5b8b0008",  3052 => x"5b9d0004",  3053 => x"78040001",
     3054 => x"78050001",  3055 => x"34020002",  3056 => x"34030002",
     3057 => x"38842510",  3058 => x"38a53e74",  3059 => x"b8205800",
     3060 => x"fbfff92c",  3061 => x"296102c8",  3062 => x"28220010",
     3063 => x"40410004",  3064 => x"20210002",  3065 => x"4420000b",
     3066 => x"40410035",  3067 => x"20210001",  3068 => x"44200008",
     3069 => x"28410008",  3070 => x"44200003",  3071 => x"28410040",
     3072 => x"5c200004",  3073 => x"b9600800",  3074 => x"34020009",
     3075 => x"f80000a1",  3076 => x"2b9d0004",  3077 => x"2b8b0008",
     3078 => x"379c0008",  3079 => x"c3a00000",  3080 => x"379cffdc",
     3081 => x"5b8b0010",  3082 => x"5b8c000c",  3083 => x"5b8d0008",
     3084 => x"5b9d0004",  3085 => x"28220020",  3086 => x"78040001",
     3087 => x"78050001",  3088 => x"284d0010",  3089 => x"282202c8",
     3090 => x"34030002",  3091 => x"38842510",  3092 => x"284c0010",
     3093 => x"38a53ea4",  3094 => x"34020002",  3095 => x"b8205800",
     3096 => x"fbfff908",  3097 => x"29620318",  3098 => x"2963031c",
     3099 => x"37810014",  3100 => x"f80010b2",  3101 => x"29810008",
     3102 => x"5c200019",  3103 => x"296200a0",  3104 => x"44410003",
     3105 => x"296100b4",  3106 => x"5c200008",  3107 => x"78040001",
     3108 => x"b9600800",  3109 => x"34020004",  3110 => x"34030001",
     3111 => x"3884251c",  3112 => x"fbfff8f8",  3113 => x"e0000013",
     3114 => x"b9600800",  3115 => x"f80011a4",  3116 => x"29a20004",
     3117 => x"29810000",  3118 => x"44400005",  3119 => x"28230034",
     3120 => x"34020000",  3121 => x"b9600800",  3122 => x"e0000004",
     3123 => x"28230034",  3124 => x"34020001",  3125 => x"b9600800",
     3126 => x"d8600000",  3127 => x"29620318",  3128 => x"b9600800",
     3129 => x"f800058c",  3130 => x"b9600800",  3131 => x"f80005b4",
     3132 => x"34010000",  3133 => x"2b9d0004",  3134 => x"2b8b0010",
     3135 => x"2b8c000c",  3136 => x"2b8d0008",  3137 => x"379c0024",
     3138 => x"c3a00000",  3139 => x"379cfff8",  3140 => x"5b8b0008",
     3141 => x"5b9d0004",  3142 => x"78040001",  3143 => x"78050001",
     3144 => x"34020002",  3145 => x"34030002",  3146 => x"38842510",
     3147 => x"38a53eb4",  3148 => x"b8205800",  3149 => x"fbfff8d3",
     3150 => x"b9600800",  3151 => x"f8000504",  3152 => x"34010000",
     3153 => x"2b9d0004",  3154 => x"2b8b0008",  3155 => x"379c0008",
     3156 => x"c3a00000",  3157 => x"379cffd8",  3158 => x"5b8b0010",
     3159 => x"5b8c000c",  3160 => x"5b8d0008",  3161 => x"5b9d0004",
     3162 => x"78050001",  3163 => x"b8806000",  3164 => x"78040001",
     3165 => x"b8406800",  3166 => x"34030002",  3167 => x"34020002",
     3168 => x"38842510",  3169 => x"38a53ec4",  3170 => x"b8205800",
     3171 => x"fbfff8bd",  3172 => x"34010001",  3173 => x"45810004",
     3174 => x"3401000c",  3175 => x"5d810036",  3176 => x"e0000022",
     3177 => x"296200ec",  3178 => x"5960031c",  3179 => x"37810024",
     3180 => x"4802000c",  3181 => x"1443001f",  3182 => x"00440010",
     3183 => x"3c630010",  3184 => x"3c420010",  3185 => x"b8641800",
     3186 => x"5b820028",  3187 => x"340203e8",  3188 => x"5b830024",
     3189 => x"fbfffcf0",  3190 => x"2b810028",  3191 => x"e000000d",
     3192 => x"c8021000",  3193 => x"1443001f",  3194 => x"00440010",
     3195 => x"3c630010",  3196 => x"3c420010",  3197 => x"b8641800",
     3198 => x"5b820028",  3199 => x"340203e8",  3200 => x"5b830024",
     3201 => x"fbfffce4",  3202 => x"2b810028",  3203 => x"c8010800",
     3204 => x"59610318",  3205 => x"356200e4",  3206 => x"b9600800",
     3207 => x"f8000fe6",  3208 => x"340c0100",  3209 => x"e0000014",
     3210 => x"296102c8",  3211 => x"b9a01000",  3212 => x"37830014",
     3213 => x"28240010",  3214 => x"b9600800",  3215 => x"340c0100",
     3216 => x"3484003c",  3217 => x"f8000416",  3218 => x"296102c8",
     3219 => x"34021000",  3220 => x"28210010",  3221 => x"2c23003c",
     3222 => x"5c620007",  3223 => x"40210004",  3224 => x"20210001",
     3225 => x"44200004",  3226 => x"b9600800",  3227 => x"34020006",
     3228 => x"f8000008",  3229 => x"b9800800",  3230 => x"2b9d0004",
     3231 => x"2b8b0010",  3232 => x"2b8c000c",  3233 => x"2b8d0008",
     3234 => x"379c0028",  3235 => x"c3a00000",  3236 => x"282302c8",
     3237 => x"34040006",  3238 => x"28630010",  3239 => x"44440004",
     3240 => x"34040009",  3241 => x"5c440008",  3242 => x"e0000004",
     3243 => x"34020001",  3244 => x"30620005",  3245 => x"e0000007",
     3246 => x"34020002",  3247 => x"30620005",  3248 => x"e0000006",
     3249 => x"40630005",  3250 => x"34020001",  3251 => x"5c620003",
     3252 => x"34020066",  3253 => x"e0000002",  3254 => x"34020064",
     3255 => x"58220004",  3256 => x"c3a00000",  3257 => x"379cfff4",
     3258 => x"5b8b000c",  3259 => x"5b8c0008",  3260 => x"5b9d0004",
     3261 => x"b8205800",  3262 => x"282102c8",  3263 => x"78050001",
     3264 => x"38a5246c",  3265 => x"282c0010",  3266 => x"34010001",
     3267 => x"41820005",  3268 => x"5c410003",  3269 => x"78050001",
     3270 => x"38a52954",  3271 => x"78040001",  3272 => x"b9600800",
     3273 => x"34020002",  3274 => x"34030001",  3275 => x"38842544",
     3276 => x"fbfff854",  3277 => x"41820005",  3278 => x"34010001",
     3279 => x"5c410003",  3280 => x"34010006",  3281 => x"e0000002",
     3282 => x"34010009",  3283 => x"59610004",  3284 => x"31800005",
     3285 => x"2b9d0004",  3286 => x"2b8b000c",  3287 => x"2b8c0008",
     3288 => x"379c000c",  3289 => x"c3a00000",  3290 => x"379cfffc",
     3291 => x"5b9d0004",  3292 => x"282202c8",  3293 => x"28420010",
     3294 => x"4043002c",  3295 => x"4460000a",  3296 => x"3463ffff",
     3297 => x"78040001",  3298 => x"3043002c",  3299 => x"38842568",
     3300 => x"34020002",  3301 => x"34030001",  3302 => x"fbfff83a",
     3303 => x"34010001",  3304 => x"e0000003",  3305 => x"fbffffd0",
     3306 => x"34010000",  3307 => x"2b9d0004",  3308 => x"379c0004",
     3309 => x"c3a00000",  3310 => x"379cffd8",  3311 => x"5b8b0018",
     3312 => x"5b8c0014",  3313 => x"5b8d0010",  3314 => x"5b8e000c",
     3315 => x"5b8f0008",  3316 => x"5b9d0004",  3317 => x"b8407000",
     3318 => x"2824000c",  3319 => x"282202c8",  3320 => x"b8205800",
     3321 => x"b8607800",  3322 => x"284d0010",  3323 => x"44800004",
     3324 => x"34010003",  3325 => x"31a1002c",  3326 => x"e000000c",
     3327 => x"282202e0",  3328 => x"44440008",  3329 => x"28220028",
     3330 => x"28440018",  3331 => x"34020000",  3332 => x"d8800000",
     3333 => x"296202e0",  3334 => x"c8220800",  3335 => x"4c20003c",
     3336 => x"340c0000",  3337 => x"e0000015",  3338 => x"29610028",
     3339 => x"340203e8",  3340 => x"28240018",  3341 => x"b9600800",
     3342 => x"d8800000",  3343 => x"596102e0",  3344 => x"296102c8",
     3345 => x"29620028",  3346 => x"4025000c",  3347 => x"1021000b",
     3348 => x"28440018",  3349 => x"bca12800",  3350 => x"b9600800",
     3351 => x"08a203e8",  3352 => x"d8800000",  3353 => x"596102d4",
     3354 => x"34021000",  3355 => x"b9600800",  3356 => x"f80003fb",
     3357 => x"b8206000",  3358 => x"45e0000e",  3359 => x"4162030d",
     3360 => x"3401000c",  3361 => x"5c41000b",  3362 => x"b9600800",
     3363 => x"b9c01000",  3364 => x"3783001c",  3365 => x"35a4003c",
     3366 => x"f8000381",  3367 => x"2da2003c",  3368 => x"34011001",
     3369 => x"5c410003",  3370 => x"34010065",  3371 => x"59610004",
     3372 => x"5d800004",  3373 => x"b9600800",  3374 => x"f8000aae",
     3375 => x"e0000003",  3376 => x"34010002",  3377 => x"59610004",
     3378 => x"29620004",  3379 => x"29610000",  3380 => x"44410002",
     3381 => x"596002d4",  3382 => x"296102c8",  3383 => x"28210010",
     3384 => x"28210028",  3385 => x"59610008",  3386 => x"b9800800",
     3387 => x"2b9d0004",  3388 => x"2b8b0018",  3389 => x"2b8c0014",
     3390 => x"2b8d0010",  3391 => x"2b8e000c",  3392 => x"2b8f0008",
     3393 => x"379c0028",  3394 => x"c3a00000",  3395 => x"b9600800",
     3396 => x"34020005",  3397 => x"f800124e",  3398 => x"b9600800",
     3399 => x"596002e0",  3400 => x"fbffff92",  3401 => x"340c0000",
     3402 => x"5c20ffc0",  3403 => x"e3ffffef",  3404 => x"379cffd8",
     3405 => x"5b8b0018",  3406 => x"5b8c0014",  3407 => x"5b8d0010",
     3408 => x"5b8e000c",  3409 => x"5b8f0008",  3410 => x"5b9d0004",
     3411 => x"b8407000",  3412 => x"2824000c",  3413 => x"282202c8",
     3414 => x"b8205800",  3415 => x"b8607800",  3416 => x"284c0010",
     3417 => x"44800004",  3418 => x"34010003",  3419 => x"3181002c",
     3420 => x"e000000c",  3421 => x"282202e0",  3422 => x"44440008",
     3423 => x"28220028",  3424 => x"28440018",  3425 => x"34020000",
     3426 => x"d8800000",  3427 => x"296202e0",  3428 => x"c8220800",
     3429 => x"4c200029",  3430 => x"340d0000",  3431 => x"e000000b",
     3432 => x"34021001",  3433 => x"b9600800",  3434 => x"f80003ad",
     3435 => x"b8206800",  3436 => x"29610028",  3437 => x"34023a98",
     3438 => x"28240018",  3439 => x"b9600800",  3440 => x"d8800000",
     3441 => x"596102e0",  3442 => x"45e0000e",  3443 => x"4162030d",
     3444 => x"3401000c",  3445 => x"5c41000b",  3446 => x"b9600800",
     3447 => x"b9c01000",  3448 => x"3783001c",  3449 => x"3584003c",
     3450 => x"f800032d",  3451 => x"2d82003c",  3452 => x"34011002",
     3453 => x"5c410003",  3454 => x"34010068",  3455 => x"59610004",
     3456 => x"45a00003",  3457 => x"34010002",  3458 => x"59610004",
     3459 => x"29810028",  3460 => x"59610008",  3461 => x"b9a00800",
     3462 => x"2b9d0004",  3463 => x"2b8b0018",  3464 => x"2b8c0014",
     3465 => x"2b8d0010",  3466 => x"2b8e000c",  3467 => x"2b8f0008",
     3468 => x"379c0028",  3469 => x"c3a00000",  3470 => x"b9600800",
     3471 => x"34020005",  3472 => x"f8001203",  3473 => x"b9600800",
     3474 => x"596002e0",  3475 => x"fbffff47",  3476 => x"340d0000",
     3477 => x"5c20ffd3",  3478 => x"e3ffffef",  3479 => x"379cfff4",
     3480 => x"5b8b000c",  3481 => x"5b8c0008",  3482 => x"5b9d0004",
     3483 => x"282202c8",  3484 => x"b8205800",  3485 => x"284c0010",
     3486 => x"2822000c",  3487 => x"44400004",  3488 => x"34010003",
     3489 => x"3181002c",  3490 => x"e000000b",  3491 => x"282302e0",
     3492 => x"44620013",  3493 => x"28220028",  3494 => x"28430018",
     3495 => x"34020000",  3496 => x"d8600000",  3497 => x"296202e0",
     3498 => x"c8220800",  3499 => x"4c200021",  3500 => x"e000000b",
     3501 => x"29810000",  3502 => x"28220000",  3503 => x"b9600800",
     3504 => x"d8400000",  3505 => x"29610028",  3506 => x"34023a98",
     3507 => x"28230018",  3508 => x"b9600800",  3509 => x"d8600000",
     3510 => x"596102e0",  3511 => x"29810000",  3512 => x"34020000",
     3513 => x"28230004",  3514 => x"b9600800",  3515 => x"d8600000",
     3516 => x"34020001",  3517 => x"5c220007",  3518 => x"34010067",
     3519 => x"59610004",  3520 => x"29810000",  3521 => x"28220008",
     3522 => x"b9600800",  3523 => x"d8400000",  3524 => x"29810028",
     3525 => x"59610008",  3526 => x"34010000",  3527 => x"2b9d0004",
     3528 => x"2b8b000c",  3529 => x"2b8c0008",  3530 => x"379c000c",
     3531 => x"c3a00000",  3532 => x"b9600800",  3533 => x"34020005",
     3534 => x"f80011c5",  3535 => x"29810000",  3536 => x"596002e0",
     3537 => x"28220008",  3538 => x"b9600800",  3539 => x"d8400000",
     3540 => x"b9600800",  3541 => x"fbffff05",  3542 => x"5c20ffd7",
     3543 => x"e3ffffef",  3544 => x"379cffd8",  3545 => x"5b8b0018",
     3546 => x"5b8c0014",  3547 => x"5b8d0010",  3548 => x"5b8e000c",
     3549 => x"5b8f0008",  3550 => x"5b9d0004",  3551 => x"b8407000",
     3552 => x"2824000c",  3553 => x"282202c8",  3554 => x"b8205800",
     3555 => x"b8607800",  3556 => x"284c0010",  3557 => x"44800004",
     3558 => x"34010003",  3559 => x"3181002c",  3560 => x"e000000c",
     3561 => x"282202e0",  3562 => x"44440008",  3563 => x"28220028",
     3564 => x"28440018",  3565 => x"34020000",  3566 => x"d8800000",
     3567 => x"296202e0",  3568 => x"c8220800",  3569 => x"4c200029",
     3570 => x"340d0000",  3571 => x"e000000b",  3572 => x"29610028",
     3573 => x"29820028",  3574 => x"28240018",  3575 => x"b9600800",
     3576 => x"d8800000",  3577 => x"596102e0",  3578 => x"34021002",
     3579 => x"b9600800",  3580 => x"f800031b",  3581 => x"b8206800",
     3582 => x"45e0000e",  3583 => x"4162030d",  3584 => x"3401000c",
     3585 => x"5c41000b",  3586 => x"b9600800",  3587 => x"b9c01000",
     3588 => x"3783001c",  3589 => x"3584003c",  3590 => x"f80002a1",
     3591 => x"2d82003c",  3592 => x"34011003",  3593 => x"5c410003",
     3594 => x"3401006a",  3595 => x"59610004",  3596 => x"45a00003",
     3597 => x"34010002",  3598 => x"59610004",  3599 => x"29810028",
     3600 => x"59610008",  3601 => x"b9a00800",  3602 => x"2b9d0004",
     3603 => x"2b8b0018",  3604 => x"2b8c0014",  3605 => x"2b8d0010",
     3606 => x"2b8e000c",  3607 => x"2b8f0008",  3608 => x"379c0028",
     3609 => x"c3a00000",  3610 => x"b9600800",  3611 => x"34020005",
     3612 => x"f8001177",  3613 => x"b9600800",  3614 => x"596002e0",
     3615 => x"fbfffebb",  3616 => x"340d0000",  3617 => x"5c20ffd3",
     3618 => x"e3ffffef",  3619 => x"379cffec",  3620 => x"5b8b0010",
     3621 => x"5b8c000c",  3622 => x"5b8d0008",  3623 => x"5b9d0004",
     3624 => x"282202c8",  3625 => x"b8206000",  3626 => x"284b0010",
     3627 => x"2822000c",  3628 => x"44400004",  3629 => x"34010003",
     3630 => x"3161002c",  3631 => x"e000000c",  3632 => x"282302e0",
     3633 => x"44620008",  3634 => x"28220028",  3635 => x"28430018",
     3636 => x"34020000",  3637 => x"d8600000",  3638 => x"298202e0",
     3639 => x"c8220800",  3640 => x"4c2000a9",  3641 => x"340d0000",
     3642 => x"e0000011",  3643 => x"29810028",  3644 => x"29620030",
     3645 => x"28230018",  3646 => x"b9800800",  3647 => x"d8600000",
     3648 => x"598102e0",  3649 => x"34021003",  3650 => x"b9800800",
     3651 => x"f80002d4",  3652 => x"b8206800",  3653 => x"3401006c",
     3654 => x"31610010",  3655 => x"29610014",  3656 => x"44200003",
     3657 => x"3401006e",  3658 => x"31610010",  3659 => x"41660010",
     3660 => x"78040001",  3661 => x"78050001",  3662 => x"b9800800",
     3663 => x"34020002",  3664 => x"34030001",  3665 => x"3884257c",
     3666 => x"38a53f18",  3667 => x"34c6ff94",  3668 => x"fbfff6cc",
     3669 => x"41620010",  3670 => x"34010008",  3671 => x"3442ff94",
     3672 => x"204200ff",  3673 => x"5441007f",  3674 => x"78010001",
     3675 => x"3c420002",  3676 => x"38213ef4",  3677 => x"b4220800",
     3678 => x"28210000",  3679 => x"c0200000",  3680 => x"29610000",
     3681 => x"34020000",  3682 => x"34030000",  3683 => x"2825002c",
     3684 => x"34040000",  3685 => x"b9800800",  3686 => x"d8a00000",
     3687 => x"5c200071",  3688 => x"3401006d",  3689 => x"31610010",
     3690 => x"29610000",  3691 => x"34020001",  3692 => x"28230024",
     3693 => x"b9800800",  3694 => x"d8600000",  3695 => x"5c200069",
     3696 => x"3401006e",  3697 => x"31610010",  3698 => x"29610000",
     3699 => x"34020001",  3700 => x"37830014",  3701 => x"28240028",
     3702 => x"b9800800",  3703 => x"d8800000",  3704 => x"34020001",
     3705 => x"5c22005f",  3706 => x"2b810014",  3707 => x"78040001",
     3708 => x"34020002",  3709 => x"00250010",  3710 => x"3c210010",
     3711 => x"5965001c",  3712 => x"59610018",  3713 => x"34030001",
     3714 => x"b9800800",  3715 => x"38842590",  3716 => x"fbfff69c",
     3717 => x"29650018",  3718 => x"78040001",  3719 => x"b9800800",
     3720 => x"34020002",  3721 => x"34030001",  3722 => x"388425b4",
     3723 => x"fbfff695",  3724 => x"3401006f",  3725 => x"31610010",
     3726 => x"29610000",  3727 => x"34020001",  3728 => x"28230020",
     3729 => x"b9800800",  3730 => x"d8600000",  3731 => x"5c200045",
     3732 => x"34010070",  3733 => x"31610010",  3734 => x"29610000",
     3735 => x"28220030",  3736 => x"b9800800",  3737 => x"d8400000",
     3738 => x"5c20003e",  3739 => x"34010071",  3740 => x"31610010",
     3741 => x"29610000",  3742 => x"34020002",  3743 => x"28230024",
     3744 => x"b9800800",  3745 => x"d8600000",  3746 => x"5c200036",
     3747 => x"34010072",  3748 => x"31610010",  3749 => x"29610000",
     3750 => x"34020002",  3751 => x"37830014",  3752 => x"28240028",
     3753 => x"b9800800",  3754 => x"d8800000",  3755 => x"34020001",
     3756 => x"5c22002c",  3757 => x"2b850014",  3758 => x"78040001",
     3759 => x"b9800800",  3760 => x"34020002",  3761 => x"34030001",
     3762 => x"388425d8",  3763 => x"fbfff66d",  3764 => x"2b810014",
     3765 => x"78040001",  3766 => x"34020002",  3767 => x"00250010",
     3768 => x"3c210010",  3769 => x"59650024",  3770 => x"59610020",
     3771 => x"34030001",  3772 => x"b9800800",  3773 => x"388425f0",
     3774 => x"fbfff662",  3775 => x"29650020",  3776 => x"78040001",
     3777 => x"b9800800",  3778 => x"34020002",  3779 => x"34030001",
     3780 => x"38842614",  3781 => x"fbfff65b",  3782 => x"34010073",
     3783 => x"31610010",  3784 => x"29610000",  3785 => x"34020002",
     3786 => x"28230020",  3787 => x"b9800800",  3788 => x"d8600000",
     3789 => x"5c20000b",  3790 => x"34010074",  3791 => x"31610010",
     3792 => x"b9800800",  3793 => x"34021004",  3794 => x"f8000245",
     3795 => x"b8206800",  3796 => x"34010069",  3797 => x"59810004",
     3798 => x"34010001",  3799 => x"59610014",  3800 => x"29610028",
     3801 => x"59810008",  3802 => x"b9a00800",  3803 => x"2b9d0004",
     3804 => x"2b8b0010",  3805 => x"2b8c000c",  3806 => x"2b8d0008",
     3807 => x"379c0014",  3808 => x"c3a00000",  3809 => x"b9800800",
     3810 => x"34020005",  3811 => x"f80010b0",  3812 => x"b9800800",
     3813 => x"598002e0",  3814 => x"fbfffdf4",  3815 => x"340d0000",
     3816 => x"5c20ff53",  3817 => x"e3fffff1",  3818 => x"379cffdc",
     3819 => x"5b8b0014",  3820 => x"5b8c0010",  3821 => x"5b8d000c",
     3822 => x"5b8e0008",  3823 => x"5b9d0004",  3824 => x"b8406800",
     3825 => x"282202c8",  3826 => x"b8205800",  3827 => x"b8607000",
     3828 => x"284c0010",  3829 => x"2822000c",  3830 => x"44400006",
     3831 => x"28220028",  3832 => x"28440018",  3833 => x"29820028",
     3834 => x"d8800000",  3835 => x"596102e0",  3836 => x"296102e0",
     3837 => x"44200009",  3838 => x"29610028",  3839 => x"34020000",
     3840 => x"28240018",  3841 => x"b9600800",  3842 => x"d8800000",
     3843 => x"296202e0",  3844 => x"c8220800",  3845 => x"4c200023",
     3846 => x"45c00018",  3847 => x"4162030d",  3848 => x"3401000c",
     3849 => x"5c410015",  3850 => x"b9600800",  3851 => x"b9a01000",
     3852 => x"37830018",  3853 => x"3584003c",  3854 => x"f8000199",
     3855 => x"2d81003c",  3856 => x"34021003",  3857 => x"5c220006",
     3858 => x"41820005",  3859 => x"34010001",  3860 => x"5c41000a",
     3861 => x"3401006a",  3862 => x"e0000007",  3863 => x"34021005",
     3864 => x"5c220006",  3865 => x"41820005",  3866 => x"34010002",
     3867 => x"5c410003",  3868 => x"3401006b",  3869 => x"59610004",
     3870 => x"29810028",  3871 => x"59610008",  3872 => x"34010000",
     3873 => x"2b9d0004",  3874 => x"2b8b0014",  3875 => x"2b8c0010",
     3876 => x"2b8d000c",  3877 => x"2b8e0008",  3878 => x"379c0024",
     3879 => x"c3a00000",  3880 => x"b9600800",  3881 => x"34020005",
     3882 => x"f8001069",  3883 => x"b9600800",  3884 => x"596002e0",
     3885 => x"fbfffd8c",  3886 => x"e3fffff2",  3887 => x"379cffd4",
     3888 => x"5b8b001c",  3889 => x"5b8c0018",  3890 => x"5b8d0014",
     3891 => x"5b8e0010",  3892 => x"5b8f000c",  3893 => x"5b900008",
     3894 => x"5b9d0004",  3895 => x"b8407000",  3896 => x"282202c8",
     3897 => x"2824000c",  3898 => x"b8205800",  3899 => x"284c0010",
     3900 => x"b8607800",  3901 => x"2d8d0048",  3902 => x"7dad0000",
     3903 => x"44800004",  3904 => x"34010003",  3905 => x"3181002c",
     3906 => x"e0000012",  3907 => x"282202e0",  3908 => x"44440022",
     3909 => x"28220028",  3910 => x"28440018",  3911 => x"34020000",
     3912 => x"d8800000",  3913 => x"296202e0",  3914 => x"c8220800",
     3915 => x"4c20003f",  3916 => x"e000001a",  3917 => x"29810000",
     3918 => x"28240030",  3919 => x"b9600800",  3920 => x"d8800000",
     3921 => x"b9600800",  3922 => x"fbfffd88",  3923 => x"4420002d",
     3924 => x"45a00008",  3925 => x"29810000",  3926 => x"34020000",
     3927 => x"34030000",  3928 => x"2825002c",  3929 => x"34040000",
     3930 => x"b9600800",  3931 => x"d8a00000",  3932 => x"2981004c",
     3933 => x"29700028",  3934 => x"340203e8",  3935 => x"f800348c",
     3936 => x"2a050018",  3937 => x"b8202000",  3938 => x"b8801000",
     3939 => x"b9600800",  3940 => x"d8a00000",  3941 => x"596102e0",
     3942 => x"45e00018",  3943 => x"4162030d",  3944 => x"3401000c",
     3945 => x"5c410015",  3946 => x"b9600800",  3947 => x"b9c01000",
     3948 => x"37830020",  3949 => x"3584003c",  3950 => x"f8000139",
     3951 => x"2d82003c",  3952 => x"34011004",  3953 => x"5c41000d",
     3954 => x"45a00005",  3955 => x"29810000",  3956 => x"28220030",
     3957 => x"b9600800",  3958 => x"d8400000",  3959 => x"41820005",
     3960 => x"34010001",  3961 => x"5c410003",  3962 => x"3401006b",
     3963 => x"e0000002",  3964 => x"34010068",  3965 => x"59610004",
     3966 => x"29810028",  3967 => x"59610008",  3968 => x"34010000",
     3969 => x"2b9d0004",  3970 => x"2b8b001c",  3971 => x"2b8c0018",
     3972 => x"2b8d0014",  3973 => x"2b8e0010",  3974 => x"2b8f000c",
     3975 => x"2b900008",  3976 => x"379c002c",  3977 => x"c3a00000",
     3978 => x"b9600800",  3979 => x"34020005",  3980 => x"f8001007",
     3981 => x"596002e0",  3982 => x"45a0ffc3",  3983 => x"e3ffffbe",
     3984 => x"379cfff0",  3985 => x"5b8b0010",  3986 => x"5b8c000c",
     3987 => x"5b8d0008",  3988 => x"5b9d0004",  3989 => x"282202c8",
     3990 => x"340d0001",  3991 => x"b8206000",  3992 => x"284b0010",
     3993 => x"29620000",  3994 => x"596d0008",  3995 => x"2842000c",
     3996 => x"d8400000",  3997 => x"41610005",  3998 => x"34020000",
     3999 => x"5c2d0005",  4000 => x"34021005",  4001 => x"b9800800",
     4002 => x"f8000175",  4003 => x"b8201000",  4004 => x"34010001",
     4005 => x"59610040",  4006 => x"3401ffff",  4007 => x"5c400009",
     4008 => x"41620005",  4009 => x"34010002",  4010 => x"5c410003",
     4011 => x"34010009",  4012 => x"e0000002",  4013 => x"34010006",
     4014 => x"59810004",  4015 => x"34010000",  4016 => x"2b9d0004",
     4017 => x"2b8b0010",  4018 => x"2b8c000c",  4019 => x"2b8d0008",
     4020 => x"379c0010",  4021 => x"c3a00000",  4022 => x"00430018",
     4023 => x"30220003",  4024 => x"30230000",  4025 => x"00430010",
     4026 => x"30230001",  4027 => x"00430008",  4028 => x"30230002",
     4029 => x"c3a00000",  4030 => x"40220000",  4031 => x"40230003",
     4032 => x"3c420018",  4033 => x"b8621000",  4034 => x"40230001",
     4035 => x"40210002",  4036 => x"3c630010",  4037 => x"3c210008",
     4038 => x"b8431000",  4039 => x"b8410800",  4040 => x"c3a00000",
     4041 => x"40220000",  4042 => x"40210001",  4043 => x"3c420008",
     4044 => x"b8410800",  4045 => x"c3a00000",  4046 => x"379cfff0",
     4047 => x"5b8b0010",  4048 => x"5b8c000c",  4049 => x"5b8d0008",
     4050 => x"5b9d0004",  4051 => x"28230020",  4052 => x"282202c8",
     4053 => x"b8205800",  4054 => x"2863000c",  4055 => x"28420010",
     4056 => x"282c003c",  4057 => x"4064000e",  4058 => x"340300ba",
     4059 => x"48830018",  4060 => x"28420000",  4061 => x"28430004",
     4062 => x"34020001",  4063 => x"d8600000",  4064 => x"ec016800",
     4065 => x"b9600800",  4066 => x"f8000967",  4067 => x"29610020",
     4068 => x"c80d6800",  4069 => x"21ad002e",  4070 => x"2821000c",
     4071 => x"35ad0006",  4072 => x"4021000e",  4073 => x"45a1000a",
     4074 => x"78010001",  4075 => x"b9a01000",  4076 => x"38212638",
     4077 => x"f8001b87",  4078 => x"29610020",  4079 => x"21ad00ff",
     4080 => x"2821000c",  4081 => x"302d000e",  4082 => x"318d0030",
     4083 => x"3401004e",  4084 => x"0d810002",  4085 => x"34010003",
     4086 => x"0d810040",  4087 => x"3401000a",  4088 => x"0d810042",
     4089 => x"34010800",  4090 => x"0d810044",  4091 => x"340130de",
     4092 => x"0d810046",  4093 => x"3401ad01",  4094 => x"0d810048",
     4095 => x"34012000",  4096 => x"0d81004a",  4097 => x"296102c8",
     4098 => x"28220010",  4099 => x"28430014",  4100 => x"40410004",
     4101 => x"44600002",  4102 => x"38210004",  4103 => x"28420008",
     4104 => x"44400002",  4105 => x"38210008",  4106 => x"0d81004c",
     4107 => x"2b9d0004",  4108 => x"2b8b0010",  4109 => x"2b8c000c",
     4110 => x"2b8d0008",  4111 => x"379c0010",  4112 => x"c3a00000",
     4113 => x"379cfff4",  4114 => x"5b8b000c",  4115 => x"5b8c0008",
     4116 => x"5b9d0004",  4117 => x"b8205800",  4118 => x"34210040",
     4119 => x"b8406000",  4120 => x"fbffffb1",  4121 => x"2d650044",
     4122 => x"2d640046",  4123 => x"78070001",  4124 => x"3ca50008",
     4125 => x"00860008",  4126 => x"38e73cd0",  4127 => x"b8a62800",
     4128 => x"28e60000",  4129 => x"64210003",  4130 => x"2d630048",
     4131 => x"e4a62800",  4132 => x"2d62004a",  4133 => x"a0250800",
     4134 => x"44200010",  4135 => x"3c840008",  4136 => x"00610008",
     4137 => x"2084ffff",  4138 => x"b8812000",  4139 => x"206300ff",
     4140 => x"3801dead",  4141 => x"e4812000",  4142 => x"64630001",
     4143 => x"a0831800",  4144 => x"44600006",  4145 => x"34012000",
     4146 => x"5c410004",  4147 => x"3561004c",  4148 => x"fbffff95",
     4149 => x"59810024",  4150 => x"2b9d0004",  4151 => x"2b8b000c",
     4152 => x"2b8c0008",  4153 => x"379c000c",  4154 => x"c3a00000",
     4155 => x"379cfff0",  4156 => x"5b8b0010",  4157 => x"5b8c000c",
     4158 => x"5b8d0008",  4159 => x"5b9d0004",  4160 => x"b8206000",
     4161 => x"282102c8",  4162 => x"204dffff",  4163 => x"28210010",
     4164 => x"40250005",  4165 => x"44a00003",  4166 => x"34012000",
     4167 => x"5da1000a",  4168 => x"78040001",  4169 => x"b9800800",
     4170 => x"34020005",  4171 => x"34030001",  4172 => x"38842650",
     4173 => x"b9a03000",  4174 => x"fbfff4d2",  4175 => x"34010000",
     4176 => x"e0000051",  4177 => x"298b003c",  4178 => x"34030008",
     4179 => x"41610000",  4180 => x"202100f0",  4181 => x"3821000c",
     4182 => x"31610000",  4183 => x"34010005",  4184 => x"31610020",
     4185 => x"29820020",  4186 => x"35610022",  4187 => x"28420014",
     4188 => x"f80033f0",  4189 => x"29810020",  4190 => x"28210014",
     4191 => x"2c210008",  4192 => x"0d6d0036",  4193 => x"00220008",
     4194 => x"3161002b",  4195 => x"34010003",  4196 => x"0d61002c",
     4197 => x"34010800",  4198 => x"0d610030",  4199 => x"340130de",
     4200 => x"0d610032",  4201 => x"3401ad01",  4202 => x"0d610034",
     4203 => x"3162002a",  4204 => x"34011003",  4205 => x"45a10005",
     4206 => x"34011004",  4207 => x"34020008",  4208 => x"5da1002d",
     4209 => x"e0000017",  4210 => x"298102c8",  4211 => x"35620038",
     4212 => x"28210010",  4213 => x"28230014",  4214 => x"44600005",
     4215 => x"40210034",  4216 => x"31610038",  4217 => x"30400001",
     4218 => x"e0000007",  4219 => x"40210034",  4220 => x"3c210008",
     4221 => x"38210001",  4222 => x"00230008",  4223 => x"31630038",
     4224 => x"30410001",  4225 => x"298102c8",  4226 => x"28220010",
     4227 => x"3561003a",  4228 => x"28420030",  4229 => x"fbffff31",
     4230 => x"34020014",  4231 => x"e0000016",  4232 => x"298102c8",
     4233 => x"28220010",  4234 => x"35610038",  4235 => x"2842001c",
     4236 => x"fbffff2a",  4237 => x"298102c8",  4238 => x"28220010",
     4239 => x"3561003c",  4240 => x"28420018",  4241 => x"fbffff25",
     4242 => x"298102c8",  4243 => x"28220010",  4244 => x"35610040",
     4245 => x"28420024",  4246 => x"fbffff20",  4247 => x"298102c8",
     4248 => x"28220010",  4249 => x"35610044",  4250 => x"28420020",
     4251 => x"fbffff1b",  4252 => x"34020018",  4253 => x"34410030",
     4254 => x"31600002",  4255 => x"31610003",  4256 => x"0d62002e",
     4257 => x"2b9d0004",  4258 => x"2b8b0010",  4259 => x"2b8c000c",
     4260 => x"2b8d0008",  4261 => x"379c0010",  4262 => x"c3a00000",
     4263 => x"379cffec",  4264 => x"5b8b0014",  4265 => x"5b8c0010",
     4266 => x"5b8d000c",  4267 => x"5b8e0008",  4268 => x"5b9d0004",
     4269 => x"b8405800",  4270 => x"b8607000",  4271 => x"34420022",
     4272 => x"b8206000",  4273 => x"b8600800",  4274 => x"34030008",
     4275 => x"b8806800",  4276 => x"f8003398",  4277 => x"3561002a",
     4278 => x"fbffff13",  4279 => x"0dc10008",  4280 => x"3561002c",
     4281 => x"fbffff10",  4282 => x"b8202800",  4283 => x"34040003",
     4284 => x"2d630030",  4285 => x"2d620032",  4286 => x"2d610034",
     4287 => x"44a40007",  4288 => x"78040001",  4289 => x"b9800800",
     4290 => x"34020005",  4291 => x"34030001",  4292 => x"38842684",
     4293 => x"e0000022",  4294 => x"3c650008",  4295 => x"78040001",
     4296 => x"00430008",  4297 => x"38843cd0",  4298 => x"b8a32800",
     4299 => x"28830000",  4300 => x"44a30007",  4301 => x"78040001",
     4302 => x"b9800800",  4303 => x"34020005",  4304 => x"34030001",
     4305 => x"388426d4",  4306 => x"e0000015",  4307 => x"3c450008",
     4308 => x"00230008",  4309 => x"20a5ffff",  4310 => x"b8a32800",
     4311 => x"3802dead",  4312 => x"44a20007",  4313 => x"78040001",
     4314 => x"b9800800",  4315 => x"34020005",  4316 => x"34030001",
     4317 => x"3884270c",  4318 => x"e0000009",  4319 => x"202500ff",
     4320 => x"34010001",  4321 => x"44a10008",  4322 => x"78040001",
     4323 => x"b9800800",  4324 => x"34020005",  4325 => x"34030001",
     4326 => x"38842750",  4327 => x"fbfff439",  4328 => x"e0000028",
     4329 => x"2d610036",  4330 => x"45a00002",  4331 => x"0da10000",
     4332 => x"34021003",  4333 => x"44220004",  4334 => x"34021004",
     4335 => x"5c220021",  4336 => x"e0000012",  4337 => x"298102c8",
     4338 => x"356e0038",  4339 => x"282d0010",  4340 => x"b9c00800",
     4341 => x"fbfffed4",  4342 => x"202100ff",  4343 => x"0da10048",
     4344 => x"b9c00800",  4345 => x"fbfffed0",  4346 => x"00210008",
     4347 => x"31a10050",  4348 => x"3561003a",  4349 => x"fbfffec1",
     4350 => x"298202c8",  4351 => x"28420010",  4352 => x"5841004c",
     4353 => x"e000000f",  4354 => x"298102c8",  4355 => x"282c0010",
     4356 => x"35610038",  4357 => x"fbfffeb9",  4358 => x"59810058",
     4359 => x"3561003c",  4360 => x"fbfffeb6",  4361 => x"59810054",
     4362 => x"35610040",  4363 => x"fbfffeb3",  4364 => x"59810060",
     4365 => x"35610044",  4366 => x"fbfffeb0",  4367 => x"5981005c",
     4368 => x"2b9d0004",  4369 => x"2b8b0014",  4370 => x"2b8c0010",
     4371 => x"2b8d000c",  4372 => x"2b8e0008",  4373 => x"379c0014",
     4374 => x"c3a00000",  4375 => x"379cfff4",  4376 => x"5b8b000c",
     4377 => x"5b8c0008",  4378 => x"5b9d0004",  4379 => x"2042ffff",
     4380 => x"b8205800",  4381 => x"fbffff1e",  4382 => x"b8206000",
     4383 => x"29610024",  4384 => x"29630070",  4385 => x"29620034",
     4386 => x"2827000c",  4387 => x"b5831800",  4388 => x"b9600800",
     4389 => x"356400f8",  4390 => x"34050000",  4391 => x"34060000",
     4392 => x"d8e00000",  4393 => x"78080001",  4394 => x"390849fc",
     4395 => x"4c2c000b",  4396 => x"29050030",  4397 => x"78040001",
     4398 => x"b9600800",  4399 => x"34020005",  4400 => x"34030001",
     4401 => x"38842794",  4402 => x"3406000c",  4403 => x"fbfff3ed",
     4404 => x"3401ffff",  4405 => x"e000000f",  4406 => x"296600f8",
     4407 => x"296700fc",  4408 => x"29080030",  4409 => x"78040001",
     4410 => x"b9600800",  4411 => x"34020005",  4412 => x"34030001",
     4413 => x"388427b4",  4414 => x"b9802800",  4415 => x"fbfff3e1",
     4416 => x"2961036c",  4417 => x"34210001",  4418 => x"5961036c",
     4419 => x"34010000",  4420 => x"2b9d0004",  4421 => x"2b8b000c",
     4422 => x"2b8c0008",  4423 => x"379c000c",  4424 => x"c3a00000",
     4425 => x"78020001",  4426 => x"384249f8",  4427 => x"58410000",
     4428 => x"c3a00000",  4429 => x"78010001",  4430 => x"38215210",
     4431 => x"28210000",  4432 => x"44200002",  4433 => x"58200010",
     4434 => x"c3a00000",  4435 => x"379cffec",  4436 => x"5b8b0014",
     4437 => x"5b8c0010",  4438 => x"5b8d000c",  4439 => x"5b8e0008",
     4440 => x"5b9d0004",  4441 => x"b8206800",  4442 => x"282102c8",
     4443 => x"780e0001",  4444 => x"39ce6db4",  4445 => x"282c0010",
     4446 => x"29c10000",  4447 => x"34020001",  4448 => x"29ab0014",
     4449 => x"fbfff30d",  4450 => x"29810000",  4451 => x"34020000",
     4452 => x"34030000",  4453 => x"2826001c",  4454 => x"35640028",
     4455 => x"b9a00800",  4456 => x"3565002c",  4457 => x"d8c00000",
     4458 => x"3402ffff",  4459 => x"5c200038",  4460 => x"29810000",
     4461 => x"34020000",  4462 => x"28230034",  4463 => x"b9a00800",
     4464 => x"d8600000",  4465 => x"34030010",  4466 => x"35a20358",
     4467 => x"b9600800",  4468 => x"f8003458",  4469 => x"29810000",
     4470 => x"596000a8",  4471 => x"28220018",  4472 => x"34010000",
     4473 => x"d8400000",  4474 => x"34010002",  4475 => x"59610014",
     4476 => x"29810058",  4477 => x"2d820054",  4478 => x"59600088",
     4479 => x"3c210010",  4480 => x"b8220800",  4481 => x"59610018",
     4482 => x"29810060",  4483 => x"2d82005c",  4484 => x"3c210010",
     4485 => x"b8220800",  4486 => x"5961001c",  4487 => x"2981001c",
     4488 => x"2d820018",  4489 => x"3c210010",  4490 => x"b8220800",
     4491 => x"59610020",  4492 => x"29810024",  4493 => x"2d820020",
     4494 => x"3c210010",  4495 => x"b8220800",  4496 => x"78020001",
     4497 => x"59610024",  4498 => x"384227d8",  4499 => x"356100c0",
     4500 => x"f8003398",  4501 => x"78010001",  4502 => x"38215210",
     4503 => x"582b0000",  4504 => x"29610010",  4505 => x"34020000",
     4506 => x"596000b8",  4507 => x"38210001",  4508 => x"59610010",
     4509 => x"78010001",  4510 => x"38215208",  4511 => x"58200000",
     4512 => x"29c10000",  4513 => x"fbfff2cd",  4514 => x"34020000",
     4515 => x"b8400800",  4516 => x"2b9d0004",  4517 => x"2b8b0014",
     4518 => x"2b8c0010",  4519 => x"2b8d000c",  4520 => x"2b8e0008",
     4521 => x"379c0014",  4522 => x"c3a00000",  4523 => x"28460000",
     4524 => x"28450004",  4525 => x"28440008",  4526 => x"28210014",
     4527 => x"28420010",  4528 => x"58260030",  4529 => x"58220040",
     4530 => x"34020001",  4531 => x"58250034",  4532 => x"58240038",
     4533 => x"5822003c",  4534 => x"28670000",  4535 => x"28660004",
     4536 => x"28650008",  4537 => x"2864000c",  4538 => x"28630010",
     4539 => x"58270044",  4540 => x"58260048",  4541 => x"5825004c",
     4542 => x"58240050",  4543 => x"58230054",  4544 => x"78010001",
     4545 => x"38215208",  4546 => x"58220000",  4547 => x"34010000",
     4548 => x"c3a00000",  4549 => x"379cfff8",  4550 => x"5b8b0008",
     4551 => x"5b9d0004",  4552 => x"282500b0",  4553 => x"282400b4",
     4554 => x"282300b8",  4555 => x"282b0014",  4556 => x"282700a8",
     4557 => x"282600ac",  4558 => x"59650060",  4559 => x"59640064",
     4560 => x"282500bc",  4561 => x"282400c0",  4562 => x"59630068",
     4563 => x"282300c4",  4564 => x"282100cc",  4565 => x"59670058",
     4566 => x"59640070",  4567 => x"5961007c",  4568 => x"34010001",
     4569 => x"59610078",  4570 => x"1441001f",  4571 => x"59630074",
     4572 => x"5966005c",  4573 => x"5965006c",  4574 => x"34030000",
     4575 => x"340403e8",  4576 => x"f8003197",  4577 => x"1423001f",
     4578 => x"2063ffff",  4579 => x"b4621000",  4580 => x"f4621800",
     4581 => x"00420010",  4582 => x"b4610800",  4583 => x"3c210010",
     4584 => x"b8221000",  4585 => x"34010000",  4586 => x"59620074",
     4587 => x"2b9d0004",  4588 => x"2b8b0008",  4589 => x"379c0008",
     4590 => x"c3a00000",  4591 => x"379cffbc",  4592 => x"5b8b003c",
     4593 => x"5b8c0038",  4594 => x"5b8d0034",  4595 => x"5b8e0030",
     4596 => x"5b8f002c",  4597 => x"5b900028",  4598 => x"5b910024",
     4599 => x"5b920020",  4600 => x"5b93001c",  4601 => x"5b940018",
     4602 => x"5b950014",  4603 => x"5b960010",  4604 => x"5b97000c",
     4605 => x"5b980008",  4606 => x"5b9d0004",  4607 => x"b8206000",
     4608 => x"282102c8",  4609 => x"298b0014",  4610 => x"282e0010",
     4611 => x"78010001",  4612 => x"38215208",  4613 => x"28210000",
     4614 => x"44200276",  4615 => x"2963003c",  4616 => x"44600007",
     4617 => x"29610050",  4618 => x"44200005",  4619 => x"29610064",
     4620 => x"44200003",  4621 => x"29610078",  4622 => x"5c200011",
     4623 => x"78010001",  4624 => x"3821520c",  4625 => x"28220000",
     4626 => x"34420001",  4627 => x"58220000",  4628 => x"34010005",
     4629 => x"4c220267",  4630 => x"29640050",  4631 => x"29650064",
     4632 => x"29660078",  4633 => x"78010001",  4634 => x"78020001",
     4635 => x"38423f54",  4636 => x"382127f8",  4637 => x"f8001957",
     4638 => x"e000025e",  4639 => x"29c10000",  4640 => x"28230038",
     4641 => x"44600004",  4642 => x"b9600800",  4643 => x"34020000",
     4644 => x"d8600000",  4645 => x"78010001",  4646 => x"38216db4",
     4647 => x"28210000",  4648 => x"34020001",  4649 => x"fbfff245",
     4650 => x"78010001",  4651 => x"3821520c",  4652 => x"58200000",
     4653 => x"296100b8",  4654 => x"29660030",  4655 => x"29670034",
     4656 => x"34210001",  4657 => x"596100b8",  4658 => x"78010001",
     4659 => x"38215208",  4660 => x"58200000",  4661 => x"29680038",
     4662 => x"2965006c",  4663 => x"29640074",  4664 => x"29610070",
     4665 => x"c8a62800",  4666 => x"c8882000",  4667 => x"c8270800",
     4668 => x"e0000002",  4669 => x"348403e8",  4670 => x"b8201800",
     4671 => x"3421ffff",  4672 => x"4804fffd",  4673 => x"b8a00800",
     4674 => x"78050001",  4675 => x"38a53cc8",  4676 => x"28a20000",
     4677 => x"e0000002",  4678 => x"b4621800",  4679 => x"b8205000",
     4680 => x"3421ffff",  4681 => x"4803fffd",  4682 => x"29610044",
     4683 => x"29650058",  4684 => x"29620060",  4685 => x"2969005c",
     4686 => x"c8a12800",  4687 => x"2961004c",  4688 => x"c8410800",
     4689 => x"29620048",  4690 => x"c9224800",  4691 => x"e0000002",
     4692 => x"342103e8",  4693 => x"b9201000",  4694 => x"3529ffff",
     4695 => x"4801fffd",  4696 => x"78090001",  4697 => x"39293cc8",
     4698 => x"292d0000",  4699 => x"e0000002",  4700 => x"b44d1000",
     4701 => x"b8a04800",  4702 => x"34a5ffff",  4703 => x"4802fffd",
     4704 => x"c8810800",  4705 => x"c9495000",  4706 => x"c8622000",
     4707 => x"e0000002",  4708 => x"342103e8",  4709 => x"b8801000",
     4710 => x"3484ffff",  4711 => x"4801fffd",  4712 => x"78040001",
     4713 => x"38843cc8",  4714 => x"b9401800",  4715 => x"28850000",
     4716 => x"e0000002",  4717 => x"b4451000",  4718 => x"b8602000",
     4719 => x"3463ffff",  4720 => x"4802fffd",  4721 => x"59610094",
     4722 => x"78010001",  4723 => x"38214e9c",  4724 => x"59620090",
     4725 => x"28210000",  4726 => x"29820018",  4727 => x"5964008c",
     4728 => x"b8220800",  4729 => x"00210010",  4730 => x"2021000f",
     4731 => x"44200032",  4732 => x"780d0001",  4733 => x"39ad2828",
     4734 => x"78050001",  4735 => x"b9800800",  4736 => x"34020004",
     4737 => x"34030002",  4738 => x"b9a02000",  4739 => x"38a52838",
     4740 => x"fbfff29c",  4741 => x"29660044",  4742 => x"29670048",
     4743 => x"2968004c",  4744 => x"78050001",  4745 => x"b9800800",
     4746 => x"34020004",  4747 => x"34030002",  4748 => x"b9a02000",
     4749 => x"38a52844",  4750 => x"fbfff292",  4751 => x"29660058",
     4752 => x"2967005c",  4753 => x"29680060",  4754 => x"78050001",
     4755 => x"b9800800",  4756 => x"34020004",  4757 => x"34030002",
     4758 => x"b9a02000",  4759 => x"38a52850",  4760 => x"fbfff288",
     4761 => x"2966006c",  4762 => x"29670070",  4763 => x"29680074",
     4764 => x"78050001",  4765 => x"b9800800",  4766 => x"34020004",
     4767 => x"34030002",  4768 => x"b9a02000",  4769 => x"38a5285c",
     4770 => x"fbfff27e",  4771 => x"2966008c",  4772 => x"29670090",
     4773 => x"29680094",  4774 => x"78050001",  4775 => x"b9800800",
     4776 => x"34020004",  4777 => x"34030002",  4778 => x"b9a02000",
     4779 => x"38a52868",  4780 => x"fbfff274",  4781 => x"2962008c",
     4782 => x"78050001",  4783 => x"38a53cd4",  4784 => x"28a40000",
     4785 => x"1441001f",  4786 => x"340300e8",  4787 => x"f80030c4",
     4788 => x"b8406800",  4789 => x"29620090",  4790 => x"b8207800",
     4791 => x"34030000",  4792 => x"1441001f",  4793 => x"340403e8",
     4794 => x"f80030bd",  4795 => x"29650094",  4796 => x"b5a21800",
     4797 => x"f5a36800",  4798 => x"14a2001f",  4799 => x"b5e10800",
     4800 => x"b4652800",  4801 => x"b5a10800",  4802 => x"f4651800",
     4803 => x"b4220800",  4804 => x"29640018",  4805 => x"29620020",
     4806 => x"b4611800",  4807 => x"2961001c",  4808 => x"297600a0",
     4809 => x"596300a0",  4810 => x"29630024",  4811 => x"b4821000",
     4812 => x"b4411000",  4813 => x"297400a4",  4814 => x"b4431000",
     4815 => x"596500a4",  4816 => x"1446001f",  4817 => x"4ca20003",
     4818 => x"596600a0",  4819 => x"596200a4",  4820 => x"296500a4",
     4821 => x"296100a0",  4822 => x"1477001f",  4823 => x"c8a21000",
     4824 => x"f4452800",  4825 => x"c8260800",  4826 => x"c8250800",
     4827 => x"1485001f",  4828 => x"b4642000",  4829 => x"f4641800",
     4830 => x"b6e5b800",  4831 => x"b477b800",  4832 => x"004d0001",
     4833 => x"3c23001f",  4834 => x"00250001",  4835 => x"b86d6800",
     4836 => x"b48d6800",  4837 => x"f48d2000",  4838 => x"b6e5b800",
     4839 => x"b497b800",  4840 => x"29640028",  4841 => x"1483001f",
     4842 => x"f800308d",  4843 => x"14350008",  4844 => x"1421001f",
     4845 => x"b5b5a800",  4846 => x"f5b56800",  4847 => x"b6e10800",
     4848 => x"b5a1b800",  4849 => x"29620030",  4850 => x"29610044",
     4851 => x"29720038",  4852 => x"29630034",  4853 => x"c8411000",
     4854 => x"2961004c",  4855 => x"ca419000",  4856 => x"29610048",
     4857 => x"c8611800",  4858 => x"e0000002",  4859 => x"365203e8",
     4860 => x"b8606800",  4861 => x"3463ffff",  4862 => x"4812fffd",
     4863 => x"78090001",  4864 => x"39293cc8",  4865 => x"29210000",
     4866 => x"e0000002",  4867 => x"b5a16800",  4868 => x"b8408800",
     4869 => x"3442ffff",  4870 => x"480dfffd",  4871 => x"378f0040",
     4872 => x"340203e8",  4873 => x"b9e00800",  4874 => x"5b970040",
     4875 => x"5b950044",  4876 => x"fbfff659",  4877 => x"78030001",
     4878 => x"38633cc8",  4879 => x"28620000",  4880 => x"b8208000",
     4881 => x"b9e00800",  4882 => x"fbfff653",  4883 => x"2b820044",
     4884 => x"b42d6800",  4885 => x"b6509000",  4886 => x"b6221000",
     4887 => x"340103e7",  4888 => x"e0000002",  4889 => x"3652fc18",
     4890 => x"b9a08800",  4891 => x"ba408000",  4892 => x"35ad0001",
     4893 => x"4a41fffc",  4894 => x"78040001",  4895 => x"78050001",
     4896 => x"38843cc4",  4897 => x"38a53cd8",  4898 => x"b8400800",
     4899 => x"28830000",  4900 => x"28a20000",  4901 => x"e0000002",
     4902 => x"b6228800",  4903 => x"b8207800",  4904 => x"ba206800",
     4905 => x"34210001",  4906 => x"4a23fffc",  4907 => x"2961002c",
     4908 => x"340203e8",  4909 => x"b9e0c000",  4910 => x"342103e7",
     4911 => x"f800306f",  4912 => x"b8209800",  4913 => x"4c110008",
     4914 => x"ba200800",  4915 => x"ba601000",  4916 => x"f8003097",
     4917 => x"4420000a",  4918 => x"083003e8",  4919 => x"ca216800",
     4920 => x"b6128000",  4921 => x"4da00006",  4922 => x"78090001",
     4923 => x"39293cc8",  4924 => x"29210000",  4925 => x"35efffff",
     4926 => x"b5a16800",  4927 => x"3401ffff",  4928 => x"5de10007",
     4929 => x"4c0d0006",  4930 => x"78020001",  4931 => x"38423cd8",
     4932 => x"28410000",  4933 => x"340f0000",  4934 => x"b5a16800",
     4935 => x"4da00007",  4936 => x"c8130800",  4937 => x"482d0005",
     4938 => x"5de00004",  4939 => x"b5b36800",  4940 => x"0a73fc18",
     4941 => x"b6138000",  4942 => x"78050001",  4943 => x"38a53cd4",
     4944 => x"28a40000",  4945 => x"1701001f",  4946 => x"bb001000",
     4947 => x"340300e8",  4948 => x"f8003023",  4949 => x"b820c000",
     4950 => x"1621001f",  4951 => x"b8409800",  4952 => x"34030000",
     4953 => x"340403e8",  4954 => x"ba201000",  4955 => x"f800301c",
     4956 => x"b6621800",  4957 => x"f6639800",  4958 => x"1642001f",
     4959 => x"b7010800",  4960 => x"b4729000",  4961 => x"b6610800",
     4962 => x"b4220800",  4963 => x"f4721800",  4964 => x"78020001",
     4965 => x"384249f8",  4966 => x"b4611800",  4967 => x"28410000",
     4968 => x"596300e8",  4969 => x"34020000",  4970 => x"596100bc",
     4971 => x"29c10000",  4972 => x"597200ec",  4973 => x"597700b0",
     4974 => x"28230004",  4975 => x"597500b4",  4976 => x"b9800800",
     4977 => x"d8600000",  4978 => x"34020001",  4979 => x"4422000c",
     4980 => x"78040001",  4981 => x"b9800800",  4982 => x"34020004",
     4983 => x"34030001",  4984 => x"38842874",  4985 => x"fbfff1a7",
     4986 => x"29c10000",  4987 => x"34020000",  4988 => x"28230034",
     4989 => x"b9800800",  4990 => x"d8600000",  4991 => x"29c10000",
     4992 => x"28210010",  4993 => x"d8200000",  4994 => x"5c200007",
     4995 => x"29630010",  4996 => x"3402fffd",  4997 => x"a0621000",
     4998 => x"59620010",  4999 => x"5de10009",  5000 => x"e000000a",
     5001 => x"78040001",  5002 => x"b9800800",  5003 => x"34020004",
     5004 => x"34030001",  5005 => x"38842898",  5006 => x"fbfff192",
     5007 => x"e00000e2",  5008 => x"34010002",  5009 => x"e0000003",
     5010 => x"45af0003",  5011 => x"34010001",  5012 => x"59610014",
     5013 => x"78040001",  5014 => x"b9800800",  5015 => x"34020004",
     5016 => x"b9e02800",  5017 => x"b9a03000",  5018 => x"34030002",
     5019 => x"388428a4",  5020 => x"ba003800",  5021 => x"fbfff183",
     5022 => x"29620014",  5023 => x"78010001",  5024 => x"38213f3c",
     5025 => x"3c420002",  5026 => x"78060001",  5027 => x"b4220800",
     5028 => x"28250000",  5029 => x"29610010",  5030 => x"38c63cbc",
     5031 => x"20210002",  5032 => x"44200003",  5033 => x"78060001",
     5034 => x"38c627e8",  5035 => x"78040001",  5036 => x"b9800800",
     5037 => x"34020004",  5038 => x"34030001",  5039 => x"388428c4",
     5040 => x"fbfff170",  5041 => x"29620014",  5042 => x"78010001",
     5043 => x"38213f3c",  5044 => x"3c420002",  5045 => x"b4221000",
     5046 => x"28420000",  5047 => x"356100c0",  5048 => x"f8003174",
     5049 => x"29620014",  5050 => x"34010004",  5051 => x"3442ffff",
     5052 => x"5441007e",  5053 => x"78010001",  5054 => x"3c420002",
     5055 => x"38213f28",  5056 => x"b4220800",  5057 => x"28210000",
     5058 => x"c0200000",  5059 => x"29c10000",  5060 => x"b9e01000",
     5061 => x"34030000",  5062 => x"28240014",  5063 => x"15e1001f",
     5064 => x"e0000006",  5065 => x"29c10000",  5066 => x"34020000",
     5067 => x"b9a01800",  5068 => x"28240014",  5069 => x"34010000",
     5070 => x"d8800000",  5071 => x"29610010",  5072 => x"38210002",
     5073 => x"59610010",  5074 => x"e0000043",  5075 => x"296500a8",
     5076 => x"78040001",  5077 => x"b9800800",  5078 => x"34020004",
     5079 => x"34030002",  5080 => x"388428dc",  5081 => x"b9a03000",
     5082 => x"ba003800",  5083 => x"fbfff145",  5084 => x"29c20000",
     5085 => x"296100a8",  5086 => x"28420018",  5087 => x"b6010800",
     5088 => x"596100a8",  5089 => x"d8400000",  5090 => x"29610010",
     5091 => x"38210002",  5092 => x"59610010",  5093 => x"34010005",
     5094 => x"59610014",  5095 => x"e0000053",  5096 => x"78090001",
     5097 => x"39293cd4",  5098 => x"29240000",  5099 => x"15e1001f",
     5100 => x"b9e01000",  5101 => x"340300e8",  5102 => x"f8002f89",
     5103 => x"b6027800",  5104 => x"1611001f",  5105 => x"f60f8000",
     5106 => x"b6210800",  5107 => x"b6018000",  5108 => x"15a1001f",
     5109 => x"34030000",  5110 => x"b9a01000",  5111 => x"340403e8",
     5112 => x"f8002f7f",  5113 => x"b5e21800",  5114 => x"f5e37800",
     5115 => x"b6010800",  5116 => x"b5e10800",  5117 => x"c8031000",
     5118 => x"48010002",  5119 => x"b8601000",  5120 => x"3401003b",
     5121 => x"4841000d",  5122 => x"29c10000",  5123 => x"34020001",
     5124 => x"28230034",  5125 => x"b9800800",  5126 => x"d8600000",
     5127 => x"296100b0",  5128 => x"59610080",  5129 => x"296100b4",
     5130 => x"59610084",  5131 => x"34010004",  5132 => x"59610014",
     5133 => x"e0000004",  5134 => x"29610088",  5135 => x"34210001",
     5136 => x"59610088",  5137 => x"29620088",  5138 => x"34010009",
     5139 => x"4c220027",  5140 => x"59600088",  5141 => x"34010003",
     5142 => x"e3ffffd0",  5143 => x"296300b4",  5144 => x"29610084",
     5145 => x"296400b0",  5146 => x"29620080",  5147 => x"c8610800",
     5148 => x"f4231800",  5149 => x"596100e4",  5150 => x"78010001",
     5151 => x"382149f8",  5152 => x"c8821000",  5153 => x"28210000",
     5154 => x"c8431000",  5155 => x"596200e0",  5156 => x"44200016",
     5157 => x"1601001f",  5158 => x"29c20000",  5159 => x"0021001e",
     5160 => x"b4308000",  5161 => x"296100a8",  5162 => x"16100002",
     5163 => x"28420018",  5164 => x"b6010800",  5165 => x"596100a8",
     5166 => x"d8400000",  5167 => x"296500a8",  5168 => x"78040001",
     5169 => x"b9800800",  5170 => x"34020006",  5171 => x"34030001",
     5172 => x"388428f8",  5173 => x"fbfff0eb",  5174 => x"296100b0",
     5175 => x"59610080",  5176 => x"296100b4",  5177 => x"59610084",
     5178 => x"29620014",  5179 => x"34010004",  5180 => x"44410004",
     5181 => x"296100f0",  5182 => x"34210001",  5183 => x"596100f0",
     5184 => x"296400e8",  5185 => x"296300ec",  5186 => x"1481001f",
     5187 => x"98611800",  5188 => x"c8611000",  5189 => x"98812000",
     5190 => x"f4431800",  5191 => x"c8810800",  5192 => x"c8230800",
     5193 => x"48200005",  5194 => x"5c200007",  5195 => x"340101f4",
     5196 => x"54410002",  5197 => x"e0000004",  5198 => x"296100f4",
     5199 => x"34210001",  5200 => x"596100f4",  5201 => x"296500a4",
     5202 => x"296400a0",  5203 => x"ca851800",  5204 => x"f4740800",
     5205 => x"cac41000",  5206 => x"c8411000",  5207 => x"48020007",
     5208 => x"34010001",  5209 => x"48400013",  5210 => x"5c400011",
     5211 => x"340203e8",  5212 => x"54620010",  5213 => x"e000000e",
     5214 => x"c8140800",  5215 => x"7c220000",  5216 => x"c8161800",
     5217 => x"c8621800",  5218 => x"c8251000",  5219 => x"f4410800",
     5220 => x"c8641800",  5221 => x"c8611800",  5222 => x"34010001",
     5223 => x"48600005",  5224 => x"5c600003",  5225 => x"340303e8",
     5226 => x"54430002",  5227 => x"34010000",  5228 => x"202100ff",
     5229 => x"44200004",  5230 => x"296100f8",  5231 => x"34210001",
     5232 => x"596100f8",  5233 => x"78010001",  5234 => x"38216db4",
     5235 => x"28210000",  5236 => x"34020000",  5237 => x"fbffeff9",
     5238 => x"29c10000",  5239 => x"28230038",  5240 => x"44600004",
     5241 => x"b9600800",  5242 => x"34020001",  5243 => x"d8600000",
     5244 => x"34010000",  5245 => x"2b9d0004",  5246 => x"2b8b003c",
     5247 => x"2b8c0038",  5248 => x"2b8d0034",  5249 => x"2b8e0030",
     5250 => x"2b8f002c",  5251 => x"2b900028",  5252 => x"2b910024",
     5253 => x"2b920020",  5254 => x"2b93001c",  5255 => x"2b940018",
     5256 => x"2b950014",  5257 => x"2b960010",  5258 => x"2b97000c",
     5259 => x"2b980008",  5260 => x"379c0044",  5261 => x"c3a00000",
     5262 => x"379cffe8",  5263 => x"5b8b0018",  5264 => x"5b8c0014",
     5265 => x"5b8d0010",  5266 => x"5b8e000c",  5267 => x"5b8f0008",
     5268 => x"5b9d0004",  5269 => x"b8407800",  5270 => x"28220020",
     5271 => x"b8205800",  5272 => x"b8607000",  5273 => x"284d0008",
     5274 => x"28220024",  5275 => x"282c02c8",  5276 => x"28440000",
     5277 => x"d8800000",  5278 => x"48010058",  5279 => x"29610020",
     5280 => x"34030008",  5281 => x"2824000c",  5282 => x"4161004c",
     5283 => x"30810004",  5284 => x"4161004d",  5285 => x"30810005",
     5286 => x"4161004e",  5287 => x"30810006",  5288 => x"3401ffff",
     5289 => x"30810007",  5290 => x"3401fffe",  5291 => x"30810008",
     5292 => x"4161004f",  5293 => x"30810009",  5294 => x"41610050",
     5295 => x"3081000a",  5296 => x"41610051",  5297 => x"3081000b",
     5298 => x"29610020",  5299 => x"2824000c",  5300 => x"b9800800",
     5301 => x"34820004",  5302 => x"f8002f96",  5303 => x"29610020",
     5304 => x"35620374",  5305 => x"28210000",  5306 => x"3180000a",
     5307 => x"c8410800",  5308 => x"14210002",  5309 => x"0821d775",
     5310 => x"0d810008",  5311 => x"41a10042",  5312 => x"3181000b",
     5313 => x"34010014",  5314 => x"3181000c",  5315 => x"41a10043",
     5316 => x"3181000d",  5317 => x"34010002",  5318 => x"3181000e",
     5319 => x"78010001",  5320 => x"382149c4",  5321 => x"28240000",
     5322 => x"4480000f",  5323 => x"b9600800",  5324 => x"b9e01000",
     5325 => x"b9c01800",  5326 => x"d8800000",  5327 => x"4420000a",
     5328 => x"78040001",  5329 => x"78050001",  5330 => x"b9600800",
     5331 => x"34020002",  5332 => x"34030001",  5333 => x"38842964",
     5334 => x"38a53f64",  5335 => x"fbfff049",  5336 => x"e000001e",
     5337 => x"29610020",  5338 => x"78040001",  5339 => x"34020003",
     5340 => x"2825000c",  5341 => x"34030001",  5342 => x"b9600800",
     5343 => x"40a5000e",  5344 => x"38842980",  5345 => x"fbfff03f",
     5346 => x"29610020",  5347 => x"78040001",  5348 => x"34020003",
     5349 => x"2825000c",  5350 => x"34030001",  5351 => x"b9600800",
     5352 => x"40a5000f",  5353 => x"38842994",  5354 => x"fbfff036",
     5355 => x"2962003c",  5356 => x"b9600800",  5357 => x"f8000634",
     5358 => x"4162001d",  5359 => x"34010001",  5360 => x"44410003",
     5361 => x"34010004",  5362 => x"e0000002",  5363 => x"34010006",
     5364 => x"59610004",  5365 => x"e0000003",  5366 => x"340103e8",
     5367 => x"59610008",  5368 => x"34010000",  5369 => x"2b9d0004",
     5370 => x"2b8b0018",  5371 => x"2b8c0014",  5372 => x"2b8d0010",
     5373 => x"2b8e000c",  5374 => x"2b8f0008",  5375 => x"379c0018",
     5376 => x"c3a00000",  5377 => x"379cfff4",  5378 => x"5b8b000c",
     5379 => x"5b8c0008",  5380 => x"5b9d0004",  5381 => x"2822000c",
     5382 => x"b8205800",  5383 => x"44400006",  5384 => x"28220028",
     5385 => x"28430018",  5386 => x"34020fa0",  5387 => x"d8600000",
     5388 => x"596102dc",  5389 => x"296102dc",  5390 => x"44200009",
     5391 => x"29610028",  5392 => x"34020000",  5393 => x"28230018",
     5394 => x"b9600800",  5395 => x"d8600000",  5396 => x"296202dc",
     5397 => x"c8220800",  5398 => x"4c200014",  5399 => x"296c02dc",
     5400 => x"34010000",  5401 => x"4580000a",  5402 => x"29610028",
     5403 => x"34020000",  5404 => x"28230018",  5405 => x"b9600800",
     5406 => x"d8600000",  5407 => x"c9810800",  5408 => x"a4201000",
     5409 => x"1442001f",  5410 => x"a0220800",  5411 => x"59610008",
     5412 => x"34010000",  5413 => x"2b9d0004",  5414 => x"2b8b000c",
     5415 => x"2b8c0008",  5416 => x"379c000c",  5417 => x"c3a00000",
     5418 => x"b9600800",  5419 => x"34020004",  5420 => x"f8000a67",
     5421 => x"34010001",  5422 => x"59610004",  5423 => x"e3fffff5",
     5424 => x"340203e8",  5425 => x"58220008",  5426 => x"34010000",
     5427 => x"c3a00000",  5428 => x"379cfff0",  5429 => x"5b8b0010",
     5430 => x"5b8c000c",  5431 => x"5b8d0008",  5432 => x"5b9d0004",
     5433 => x"78040001",  5434 => x"388449c4",  5435 => x"2884000c",
     5436 => x"b8205800",  5437 => x"b8406800",  5438 => x"b8606000",
     5439 => x"44800003",  5440 => x"d8800000",  5441 => x"5c20001f",
     5442 => x"2961000c",  5443 => x"4420000b",  5444 => x"296102c8",
     5445 => x"29630028",  5446 => x"4022000c",  5447 => x"1021000b",
     5448 => x"28630018",  5449 => x"bc411000",  5450 => x"b9600800",
     5451 => x"084203e8",  5452 => x"d8600000",  5453 => x"596102d4",
     5454 => x"4580000f",  5455 => x"4161030d",  5456 => x"44200008",
     5457 => x"3402000b",  5458 => x"5c22000b",  5459 => x"b9600800",
     5460 => x"b9a01000",  5461 => x"b9801800",  5462 => x"f8000352",
     5463 => x"e0000005",  5464 => x"b9600800",  5465 => x"b9a01000",
     5466 => x"b9801800",  5467 => x"f8000370",  5468 => x"5c200004",
     5469 => x"b9600800",  5470 => x"f800027e",  5471 => x"44200003",
     5472 => x"34010002",  5473 => x"59610004",  5474 => x"29620004",
     5475 => x"29610000",  5476 => x"44410002",  5477 => x"596002d4",
     5478 => x"296c02d4",  5479 => x"34010000",  5480 => x"4580000a",
     5481 => x"29610028",  5482 => x"34020000",  5483 => x"28230018",
     5484 => x"b9600800",  5485 => x"d8600000",  5486 => x"c9810800",
     5487 => x"a4201000",  5488 => x"1442001f",  5489 => x"a0220800",
     5490 => x"59610008",  5491 => x"34010000",  5492 => x"2b9d0004",
     5493 => x"2b8b0010",  5494 => x"2b8c000c",  5495 => x"2b8d0008",
     5496 => x"379c0010",  5497 => x"c3a00000",  5498 => x"34010000",
     5499 => x"c3a00000",  5500 => x"379cffec",  5501 => x"5b8b0014",
     5502 => x"5b8c0010",  5503 => x"5b8d000c",  5504 => x"5b8e0008",
     5505 => x"5b9d0004",  5506 => x"344b00b2",  5507 => x"3d6b0002",
     5508 => x"b8407000",  5509 => x"b42b5800",  5510 => x"29620004",
     5511 => x"b8206000",  5512 => x"340d0000",  5513 => x"44400008",
     5514 => x"28220028",  5515 => x"28430018",  5516 => x"34020000",
     5517 => x"d8600000",  5518 => x"29620004",  5519 => x"c8220800",
     5520 => x"4c200009",  5521 => x"b9a00800",  5522 => x"2b9d0004",
     5523 => x"2b8b0014",  5524 => x"2b8c0010",  5525 => x"2b8d000c",
     5526 => x"2b8e0008",  5527 => x"379c0014",  5528 => x"c3a00000",
     5529 => x"b9800800",  5530 => x"b9c01000",  5531 => x"f80009f8",
     5532 => x"340d0001",  5533 => x"59600004",  5534 => x"e3fffff3",
     5535 => x"379cffec",  5536 => x"5b8b0014",  5537 => x"5b8c0010",
     5538 => x"5b8d000c",  5539 => x"5b8e0008",  5540 => x"5b9d0004",
     5541 => x"b8407000",  5542 => x"2822000c",  5543 => x"b8205800",
     5544 => x"b8606800",  5545 => x"340c0000",  5546 => x"44400014",
     5547 => x"282302c8",  5548 => x"34020001",  5549 => x"1063000d",
     5550 => x"f80009f4",  5551 => x"296302c8",  5552 => x"b9600800",
     5553 => x"34020003",  5554 => x"1063000b",  5555 => x"f80009ef",
     5556 => x"29630344",  5557 => x"34020001",  5558 => x"34010000",
     5559 => x"5c620002",  5560 => x"29610340",  5561 => x"0d61007e",
     5562 => x"b9600800",  5563 => x"f80005d9",  5564 => x"b8206000",
     5565 => x"48010047",  5566 => x"b9600800",  5567 => x"34020001",
     5568 => x"fbffffbc",  5569 => x"44200010",  5570 => x"296302c8",
     5571 => x"b9600800",  5572 => x"34020001",  5573 => x"1063000d",
     5574 => x"f80009dc",  5575 => x"29630344",  5576 => x"34020001",
     5577 => x"34010000",  5578 => x"5c620002",  5579 => x"29610340",
     5580 => x"0d61007e",  5581 => x"b9600800",  5582 => x"f8000613",
     5583 => x"48010046",  5584 => x"340c0000",  5585 => x"b9600800",
     5586 => x"34020003",  5587 => x"fbffffa9",  5588 => x"44200010",
     5589 => x"29630344",  5590 => x"34020001",  5591 => x"34010000",
     5592 => x"5c620002",  5593 => x"29610340",  5594 => x"0d61007e",
     5595 => x"b9600800",  5596 => x"f80005b8",  5597 => x"48010038",
     5598 => x"296302c8",  5599 => x"b9600800",  5600 => x"34020003",
     5601 => x"1063000b",  5602 => x"340c0000",  5603 => x"f80009bf",
     5604 => x"45a00020",  5605 => x"78010001",  5606 => x"382149c4",
     5607 => x"28250010",  5608 => x"4164030d",  5609 => x"44a00007",
     5610 => x"b9600800",  5611 => x"b9c01000",  5612 => x"b9a01800",
     5613 => x"d8a00000",  5614 => x"b8202000",  5615 => x"48010042",
     5616 => x"34010001",  5617 => x"44810010",  5618 => x"3401000b",
     5619 => x"44810003",  5620 => x"5c800010",  5621 => x"e0000006",
     5622 => x"b9600800",  5623 => x"b9c01000",  5624 => x"b9a01800",
     5625 => x"f80002af",  5626 => x"e0000005",  5627 => x"b9600800",
     5628 => x"b9c01000",  5629 => x"b9a01800",  5630 => x"f80002cd",
     5631 => x"b8206000",  5632 => x"e0000004",  5633 => x"b9600800",
     5634 => x"356200e4",  5635 => x"f800066a",  5636 => x"45800006",
     5637 => x"34010001",  5638 => x"4581000f",  5639 => x"3401ffff",
     5640 => x"5d81000e",  5641 => x"e0000029",  5642 => x"29610020",
     5643 => x"2821000c",  5644 => x"4022000e",  5645 => x"340100ff",
     5646 => x"44410004",  5647 => x"4162001d",  5648 => x"34010002",
     5649 => x"5c410005",  5650 => x"34010004",  5651 => x"59610004",
     5652 => x"e0000002",  5653 => x"340c0000",  5654 => x"296e02d8",
     5655 => x"340d0000",  5656 => x"45c0000a",  5657 => x"29610028",
     5658 => x"34020000",  5659 => x"28230018",  5660 => x"b9600800",
     5661 => x"d8600000",  5662 => x"c9c16800",  5663 => x"a5a00800",
     5664 => x"1421001f",  5665 => x"a1a16800",  5666 => x"296e02d0",
     5667 => x"34010000",  5668 => x"45c0000a",  5669 => x"29610028",
     5670 => x"34020000",  5671 => x"28230018",  5672 => x"b9600800",
     5673 => x"d8600000",  5674 => x"c9c10800",  5675 => x"a4201000",
     5676 => x"1442001f",  5677 => x"a0220800",  5678 => x"4da10007",
     5679 => x"b9a00800",  5680 => x"e0000005",  5681 => x"b8206000",
     5682 => x"34010002",  5683 => x"59610004",  5684 => x"340101f4",
     5685 => x"59610008",  5686 => x"b9800800",  5687 => x"2b9d0004",
     5688 => x"2b8b0014",  5689 => x"2b8c0010",  5690 => x"2b8d000c",
     5691 => x"2b8e0008",  5692 => x"379c0014",  5693 => x"c3a00000",
     5694 => x"379cfff0",  5695 => x"5b8b000c",  5696 => x"5b8c0008",
     5697 => x"5b9d0004",  5698 => x"b8406000",  5699 => x"2822000c",
     5700 => x"b8205800",  5701 => x"4440000c",  5702 => x"282202c8",
     5703 => x"28250028",  5704 => x"4044000c",  5705 => x"1042000b",
     5706 => x"bc821000",  5707 => x"28a40018",  5708 => x"084203e8",
     5709 => x"5b830010",  5710 => x"d8800000",  5711 => x"2b830010",
     5712 => x"596102d4",  5713 => x"4460000d",  5714 => x"4161030d",
     5715 => x"44200007",  5716 => x"3402000b",  5717 => x"5c220009",
     5718 => x"b9600800",  5719 => x"b9801000",  5720 => x"f8000250",
     5721 => x"e0000004",  5722 => x"b9600800",  5723 => x"b9801000",
     5724 => x"f800026f",  5725 => x"5c200004",  5726 => x"b9600800",
     5727 => x"f800017d",  5728 => x"44200003",  5729 => x"34010002",
     5730 => x"59610004",  5731 => x"29620004",  5732 => x"29610000",
     5733 => x"44410002",  5734 => x"596002d4",  5735 => x"340103e8",
     5736 => x"59610008",  5737 => x"34010000",  5738 => x"2b9d0004",
     5739 => x"2b8b000c",  5740 => x"2b8c0008",  5741 => x"379c0010",
     5742 => x"c3a00000",  5743 => x"379cfff8",  5744 => x"5b8b0008",
     5745 => x"5b9d0004",  5746 => x"b8205800",  5747 => x"4460000d",
     5748 => x"4024030d",  5749 => x"44800007",  5750 => x"34050008",
     5751 => x"44850007",  5752 => x"3405000b",  5753 => x"5c850007",
     5754 => x"f8000198",  5755 => x"e0000004",  5756 => x"f80001b1",
     5757 => x"e0000002",  5758 => x"f80001e9",  5759 => x"5c200004",
     5760 => x"b9600800",  5761 => x"f800015b",  5762 => x"44200003",
     5763 => x"34010002",  5764 => x"59610004",  5765 => x"340103e8",
     5766 => x"59610008",  5767 => x"34010000",  5768 => x"2b9d0004",
     5769 => x"2b8b0008",  5770 => x"379c0008",  5771 => x"c3a00000",
     5772 => x"379cffd4",  5773 => x"5b8b0014",  5774 => x"5b8c0010",
     5775 => x"5b8d000c",  5776 => x"5b8e0008",  5777 => x"5b9d0004",
     5778 => x"b8205800",  5779 => x"2821000c",  5780 => x"b8407000",
     5781 => x"b8606800",  5782 => x"44200023",  5783 => x"34020000",
     5784 => x"34030014",  5785 => x"35610080",  5786 => x"f8002e30",
     5787 => x"b9600800",  5788 => x"f80006da",  5789 => x"78010001",
     5790 => x"382149c4",  5791 => x"28240014",  5792 => x"44800007",
     5793 => x"b9600800",  5794 => x"b9c01000",  5795 => x"b9a01800",
     5796 => x"d8800000",  5797 => x"b8206000",  5798 => x"5c20005f",
     5799 => x"4161001c",  5800 => x"29630028",  5801 => x"202100fd",
     5802 => x"3161001c",  5803 => x"296102c8",  5804 => x"28630018",
     5805 => x"4022000c",  5806 => x"1021000b",  5807 => x"bc411000",
     5808 => x"b9600800",  5809 => x"084203e8",  5810 => x"d8600000",
     5811 => x"296302c8",  5812 => x"596102d4",  5813 => x"34020000",
     5814 => x"1063000a",  5815 => x"b9600800",  5816 => x"f80008ea",
     5817 => x"45a00049",  5818 => x"4161030d",  5819 => x"34020008",
     5820 => x"44220012",  5821 => x"54220003",  5822 => x"5c200044",
     5823 => x"e000000a",  5824 => x"34020009",  5825 => x"44220014",
     5826 => x"3402000b",  5827 => x"5c22003f",  5828 => x"b9600800",
     5829 => x"b9c01000",  5830 => x"b9a01800",  5831 => x"f800014b",
     5832 => x"e000000a",  5833 => x"b9600800",  5834 => x"b9c01000",
     5835 => x"b9a01800",  5836 => x"f8000161",  5837 => x"e0000005",
     5838 => x"b9600800",  5839 => x"b9c01000",  5840 => x"b9a01800",
     5841 => x"f8000196",  5842 => x"b8206000",  5843 => x"5c200032",
     5844 => x"e000002e",  5845 => x"34010035",  5846 => x"340c0001",
     5847 => x"4c2d002e",  5848 => x"378c0018",  5849 => x"b9c00800",
     5850 => x"b9801000",  5851 => x"f80004a2",  5852 => x"296102c8",
     5853 => x"37820024",  5854 => x"34030008",  5855 => x"f8002d4c",
     5856 => x"5c20001c",  5857 => x"2d6202f2",  5858 => x"2d61032a",
     5859 => x"5c410019",  5860 => x"296102c8",  5861 => x"2c220008",
     5862 => x"2f81002c",  5863 => x"5c410015",  5864 => x"4161001c",
     5865 => x"20210001",  5866 => x"44200012",  5867 => x"b9801000",
     5868 => x"356100bc",  5869 => x"f8000619",  5870 => x"78010001",
     5871 => x"382149c4",  5872 => x"28220018",  5873 => x"44400006",
     5874 => x"b9600800",  5875 => x"d8400000",  5876 => x"b8206000",
     5877 => x"5c200010",  5878 => x"e0000003",  5879 => x"b9600800",
     5880 => x"f80006d7",  5881 => x"4161032d",  5882 => x"316102ee",
     5883 => x"e0000007",  5884 => x"78040001",  5885 => x"b9600800",
     5886 => x"34020005",  5887 => x"34030002",  5888 => x"388429ac",
     5889 => x"fbffee1f",  5890 => x"b9600800",  5891 => x"f80000d9",
     5892 => x"b8206000",  5893 => x"296102cc",  5894 => x"44200009",
     5895 => x"29610028",  5896 => x"34020000",  5897 => x"28230018",
     5898 => x"b9600800",  5899 => x"d8600000",  5900 => x"296202cc",
     5901 => x"c8220800",  5902 => x"4c200033",  5903 => x"3401ffff",
     5904 => x"45810005",  5905 => x"7d810001",  5906 => x"c8010800",
     5907 => x"a1816000",  5908 => x"e0000003",  5909 => x"34010002",
     5910 => x"59610004",  5911 => x"29620004",  5912 => x"29610000",
     5913 => x"44410005",  5914 => x"596002d4",  5915 => x"596002cc",
     5916 => x"b9600800",  5917 => x"f8000659",  5918 => x"296e02d4",
     5919 => x"340d0000",  5920 => x"45c0000a",  5921 => x"29610028",
     5922 => x"34020000",  5923 => x"28230018",  5924 => x"b9600800",
     5925 => x"d8600000",  5926 => x"c9c16800",  5927 => x"a5a00800",
     5928 => x"1421001f",  5929 => x"a1a16800",  5930 => x"296e02cc",
     5931 => x"b9a00800",  5932 => x"45c0000a",  5933 => x"29610028",
     5934 => x"34020000",  5935 => x"28230018",  5936 => x"b9600800",
     5937 => x"d8600000",  5938 => x"c9c10800",  5939 => x"a4201000",
     5940 => x"1442001f",  5941 => x"a0220800",  5942 => x"4da10002",
     5943 => x"b9a00800",  5944 => x"59610008",  5945 => x"b9800800",
     5946 => x"2b9d0004",  5947 => x"2b8b0014",  5948 => x"2b8c0010",
     5949 => x"2b8d000c",  5950 => x"2b8e0008",  5951 => x"379c002c",
     5952 => x"c3a00000",  5953 => x"b9600800",  5954 => x"34020000",
     5955 => x"f8000850",  5956 => x"b9600800",  5957 => x"596002cc",
     5958 => x"f80004f6",  5959 => x"29630100",  5960 => x"29620104",
     5961 => x"296500f8",  5962 => x"296400fc",  5963 => x"b8206000",
     5964 => x"29610108",  5965 => x"596300b0",  5966 => x"296302c8",
     5967 => x"596200b4",  5968 => x"596100b8",  5969 => x"596500a8",
     5970 => x"596400ac",  5971 => x"1063000a",  5972 => x"b9600800",
     5973 => x"34020000",  5974 => x"f800084c",  5975 => x"29620020",
     5976 => x"356100a8",  5977 => x"28430008",  5978 => x"b8201000",
     5979 => x"34630018",  5980 => x"f80005bd",  5981 => x"e3ffffb2",
     5982 => x"379cfff8",  5983 => x"5b8b0008",  5984 => x"5b9d0004",
     5985 => x"282202c8",  5986 => x"28240028",  5987 => x"b8205800",
     5988 => x"4043000c",  5989 => x"1042000b",  5990 => x"bc621000",
     5991 => x"28830018",  5992 => x"084203e8",  5993 => x"d8600000",
     5994 => x"596102d4",  5995 => x"2b9d0004",  5996 => x"2b8b0008",
     5997 => x"379c0008",  5998 => x"c3a00000",  5999 => x"379cffe4",
     6000 => x"5b8b001c",  6001 => x"5b8c0018",  6002 => x"5b8d0014",
     6003 => x"5b8e0010",  6004 => x"5b8f000c",  6005 => x"5b900008",
     6006 => x"5b9d0004",  6007 => x"340c0000",  6008 => x"b8205800",
     6009 => x"b8407000",  6010 => x"342f030c",  6011 => x"34300320",
     6012 => x"e0000013",  6013 => x"098d0058",  6014 => x"ba000800",
     6015 => x"3403000a",  6016 => x"35a20110",  6017 => x"b5621000",
     6018 => x"f8002ca9",  6019 => x"5c20000b",  6020 => x"b56d0800",
     6021 => x"b9e01000",  6022 => x"34030024",  6023 => x"34210144",
     6024 => x"f8002cc4",  6025 => x"b56d5800",  6026 => x"b9c00800",
     6027 => x"3562011c",  6028 => x"f80003be",  6029 => x"e0000020",
     6030 => x"358c0001",  6031 => x"2d63010c",  6032 => x"486cffed",
     6033 => x"34010004",  6034 => x"54610003",  6035 => x"34630001",
     6036 => x"0d63010c",  6037 => x"2d6d010c",  6038 => x"35620320",
     6039 => x"3403000a",  6040 => x"35adffff",  6041 => x"09ac0058",
     6042 => x"35810110",  6043 => x"b5610800",  6044 => x"f8002cb0",
     6045 => x"b56c0800",  6046 => x"34030024",  6047 => x"b9e01000",
     6048 => x"34210144",  6049 => x"f8002cab",  6050 => x"b56c1000",
     6051 => x"b9c00800",  6052 => x"3442011c",  6053 => x"f80003a5",
     6054 => x"78040001",  6055 => x"b9600800",  6056 => x"34020003",
     6057 => x"34030001",  6058 => x"388429dc",  6059 => x"b9a02800",
     6060 => x"fbffed74",  6061 => x"2b9d0004",  6062 => x"2b8b001c",
     6063 => x"2b8c0018",  6064 => x"2b8d0014",  6065 => x"2b8e0010",
     6066 => x"2b8f000c",  6067 => x"2b900008",  6068 => x"379c001c",
     6069 => x"c3a00000",  6070 => x"4022001e",  6071 => x"34030001",
     6072 => x"44430009",  6073 => x"44400008",  6074 => x"34030002",
     6075 => x"5c430008",  6076 => x"34020012",  6077 => x"58220070",
     6078 => x"3402000e",  6079 => x"58220074",  6080 => x"e0000003",
     6081 => x"58200070",  6082 => x"58200074",  6083 => x"28240070",
     6084 => x"2825002c",  6085 => x"34020000",  6086 => x"b4a42800",
     6087 => x"20a30003",  6088 => x"44600003",  6089 => x"34020004",
     6090 => x"c8431000",  6091 => x"b4a22800",  6092 => x"28260030",
     6093 => x"28220074",  6094 => x"5825003c",  6095 => x"34030000",
     6096 => x"b4c23000",  6097 => x"20c70003",  6098 => x"44e00003",
     6099 => x"34030004",  6100 => x"c8671800",  6101 => x"b4c31800",
     6102 => x"c8a42000",  6103 => x"c8621000",  6104 => x"58230040",
     6105 => x"58240034",  6106 => x"58220038",  6107 => x"c3a00000",
     6108 => x"379cfff4",  6109 => x"5b8b000c",  6110 => x"5b8c0008",
     6111 => x"5b9d0004",  6112 => x"78020001",  6113 => x"384249c4",
     6114 => x"28420020",  6115 => x"b8205800",  6116 => x"44400006",
     6117 => x"d8400000",  6118 => x"b8206000",  6119 => x"34010001",
     6120 => x"45810018",  6121 => x"480c0018",  6122 => x"296102d4",
     6123 => x"340c0000",  6124 => x"44200015",  6125 => x"29610028",
     6126 => x"34020000",  6127 => x"28230018",  6128 => x"b9600800",
     6129 => x"d8600000",  6130 => x"296202d4",  6131 => x"c8220800",
     6132 => x"4c200013",  6133 => x"e000000c",  6134 => x"4162001d",
     6135 => x"34010002",  6136 => x"44410004",  6137 => x"34010006",
     6138 => x"59610004",  6139 => x"e0000006",  6140 => x"34010004",
     6141 => x"59610004",  6142 => x"b9600800",  6143 => x"fbffff5f",
     6144 => x"340c0000",  6145 => x"b9800800",  6146 => x"2b9d0004",
     6147 => x"2b8b000c",  6148 => x"2b8c0008",  6149 => x"379c000c",
     6150 => x"c3a00000",  6151 => x"b9600800",  6152 => x"34020002",
     6153 => x"f800078a",  6154 => x"29610020",  6155 => x"596002d4",
     6156 => x"0d60010c",  6157 => x"2821000c",  6158 => x"4022000e",
     6159 => x"340100ff",  6160 => x"5c41ffe6",  6161 => x"e3ffffeb",
     6162 => x"379cfff4",  6163 => x"5b8b000c",  6164 => x"5b8c0008",
     6165 => x"5b9d0004",  6166 => x"3404003f",  6167 => x"b8205800",
     6168 => x"340cffff",  6169 => x"4c83000e",  6170 => x"fbffff55",
     6171 => x"b9600800",  6172 => x"fbffff42",  6173 => x"b9600800",
     6174 => x"f800015a",  6175 => x"59610004",  6176 => x"78010001",
     6177 => x"382149c4",  6178 => x"28220024",  6179 => x"340c0000",
     6180 => x"44400003",  6181 => x"b9600800",  6182 => x"d8400000",
     6183 => x"b9800800",  6184 => x"2b9d0004",  6185 => x"2b8b000c",
     6186 => x"2b8c0008",  6187 => x"379c000c",  6188 => x"c3a00000",
     6189 => x"379cffe0",  6190 => x"5b8b0014",  6191 => x"5b8c0010",
     6192 => x"5b8d000c",  6193 => x"5b8e0008",  6194 => x"5b9d0004",
     6195 => x"b8205800",  6196 => x"3401002b",  6197 => x"b8407000",
     6198 => x"340cffff",  6199 => x"4c230028",  6200 => x"4161001c",
     6201 => x"340c0000",  6202 => x"20210001",  6203 => x"44200024",
     6204 => x"296300ec",  6205 => x"296200f0",  6206 => x"296100f4",
     6207 => x"296500e4",  6208 => x"296400e8",  6209 => x"5963009c",
     6210 => x"596200a0",  6211 => x"2963031c",  6212 => x"29620318",
     6213 => x"596100a4",  6214 => x"59650094",  6215 => x"356100d0",
     6216 => x"59640098",  6217 => x"f8000485",  6218 => x"41610313",
     6219 => x"20210002",  6220 => x"44200007",  6221 => x"4161001c",
     6222 => x"38210002",  6223 => x"3161001c",  6224 => x"2d61032a",
     6225 => x"0d6102ec",  6226 => x"e000000d",  6227 => x"378d0018",
     6228 => x"b9c00800",  6229 => x"b9a01000",  6230 => x"f80002ed",
     6231 => x"4161001c",  6232 => x"b9a01000",  6233 => x"202100fd",
     6234 => x"3161001c",  6235 => x"35610080",  6236 => x"f80004aa",
     6237 => x"b9600800",  6238 => x"f8000551",  6239 => x"b9800800",
     6240 => x"2b9d0004",  6241 => x"2b8b0014",  6242 => x"2b8c0010",
     6243 => x"2b8d000c",  6244 => x"2b8e0008",  6245 => x"379c0020",
     6246 => x"c3a00000",  6247 => x"379cffe4",  6248 => x"5b8b0010",
     6249 => x"5b8c000c",  6250 => x"5b8d0008",  6251 => x"5b9d0004",
     6252 => x"b8205800",  6253 => x"b8400800",  6254 => x"3402002b",
     6255 => x"3404ffff",  6256 => x"4c430031",  6257 => x"4162001c",
     6258 => x"20430001",  6259 => x"5c600004",  6260 => x"78010001",
     6261 => x"382129fc",  6262 => x"e0000005",  6263 => x"20420002",
     6264 => x"5c400007",  6265 => x"78010001",  6266 => x"38212a38",
     6267 => x"78020001",  6268 => x"38423f74",  6269 => x"f80012f7",
     6270 => x"e0000022",  6271 => x"2d6402ec",  6272 => x"2d63032a",
     6273 => x"44830007",  6274 => x"78010001",  6275 => x"78020001",
     6276 => x"38423f74",  6277 => x"38212a70",  6278 => x"f80012ee",
     6279 => x"e0000019",  6280 => x"378d0014",  6281 => x"b9a01000",
     6282 => x"f80002ec",  6283 => x"4161001c",  6284 => x"356c0080",
     6285 => x"b9a01000",  6286 => x"202100fd",  6287 => x"3161001c",
     6288 => x"b9800800",  6289 => x"f8000475",  6290 => x"78030001",
     6291 => x"386349c4",  6292 => x"28640028",  6293 => x"44800009",
     6294 => x"b9600800",  6295 => x"b9801000",  6296 => x"356300d0",
     6297 => x"d8800000",  6298 => x"b8202000",  6299 => x"34010001",
     6300 => x"44810004",  6301 => x"48040004",  6302 => x"b9600800",
     6303 => x"f8000510",  6304 => x"34040000",  6305 => x"b8800800",
     6306 => x"2b9d0004",  6307 => x"2b8b0010",  6308 => x"2b8c000c",
     6309 => x"2b8d0008",  6310 => x"379c001c",  6311 => x"c3a00000",
     6312 => x"379cfff0",  6313 => x"5b8b0010",  6314 => x"5b8c000c",
     6315 => x"5b8d0008",  6316 => x"5b9d0004",  6317 => x"b8406800",
     6318 => x"3402003f",  6319 => x"b8205800",  6320 => x"340cffff",
     6321 => x"4c430013",  6322 => x"78040001",  6323 => x"34030002",
     6324 => x"38842ab0",  6325 => x"34020003",  6326 => x"fbffec6a",
     6327 => x"b9a01000",  6328 => x"b9600800",  6329 => x"fbfffeb6",
     6330 => x"b9600800",  6331 => x"f80000bd",  6332 => x"59610004",
     6333 => x"78010001",  6334 => x"382149c4",  6335 => x"28220024",
     6336 => x"340c0000",  6337 => x"44400003",  6338 => x"b9600800",
     6339 => x"d8400000",  6340 => x"b9800800",  6341 => x"2b9d0004",
     6342 => x"2b8b0010",  6343 => x"2b8c000c",  6344 => x"2b8d0008",
     6345 => x"379c0010",  6346 => x"c3a00000",  6347 => x"34010000",
     6348 => x"c3a00000",  6349 => x"379cfffc",  6350 => x"5b9d0004",
     6351 => x"34030008",  6352 => x"f8002b5b",  6353 => x"2b9d0004",
     6354 => x"379c0004",  6355 => x"c3a00000",  6356 => x"379cffe0",
     6357 => x"5b8b0020",  6358 => x"5b8c001c",  6359 => x"5b8d0018",
     6360 => x"5b8e0014",  6361 => x"5b8f0010",  6362 => x"5b90000c",
     6363 => x"5b910008",  6364 => x"5b9d0004",  6365 => x"780e0001",
     6366 => x"39ce3f94",  6367 => x"78040001",  6368 => x"b8406800",
     6369 => x"b8606000",  6370 => x"34020003",  6371 => x"34030002",
     6372 => x"38842e58",  6373 => x"b9c02800",  6374 => x"b8207800",
     6375 => x"35b10021",  6376 => x"fbffec38",  6377 => x"35900021",
     6378 => x"ba200800",  6379 => x"ba001000",  6380 => x"fbffffe1",
     6381 => x"5c200033",  6382 => x"2d81002a",  6383 => x"2dab002a",
     6384 => x"c9615800",  6385 => x"35620001",  6386 => x"34010002",
     6387 => x"54410043",  6388 => x"29e20020",  6389 => x"34030001",
     6390 => x"35a10048",  6391 => x"28420014",  6392 => x"5d63000b",
     6393 => x"fbffffd4",  6394 => x"5c20003c",  6395 => x"78040001",
     6396 => x"b9e00800",  6397 => x"34020003",  6398 => x"34030001",
     6399 => x"38842ae0",  6400 => x"b9c02800",  6401 => x"3406008f",
     6402 => x"e000000e",  6403 => x"3403ffff",  6404 => x"358c0048",
     6405 => x"5d63000e",  6406 => x"b9800800",  6407 => x"fbffffc6",
     6408 => x"5c20002e",  6409 => x"78040001",  6410 => x"b9e00800",
     6411 => x"34020003",  6412 => x"34030001",  6413 => x"38842ae0",
     6414 => x"b9c02800",  6415 => x"34060098",  6416 => x"fbffec10",
     6417 => x"340b0000",  6418 => x"e0000024",  6419 => x"b9801000",
     6420 => x"fbffffb9",  6421 => x"b8205800",  6422 => x"5c200020",
     6423 => x"78040001",  6424 => x"b9e00800",  6425 => x"34020003",
     6426 => x"34030001",  6427 => x"38842af0",  6428 => x"b9c02800",
     6429 => x"340600a0",  6430 => x"fbffec02",  6431 => x"e0000017",
     6432 => x"41ab001a",  6433 => x"4181001a",  6434 => x"5d61000e",
     6435 => x"41ab001c",  6436 => x"4181001c",  6437 => x"5d61000b",
     6438 => x"41ab001d",  6439 => x"4181001d",  6440 => x"5d610008",
     6441 => x"2da2001e",  6442 => x"2d81001e",  6443 => x"340b0000",
     6444 => x"5c41000a",  6445 => x"41ab0020",  6446 => x"41810020",
     6447 => x"45610003",  6448 => x"c9615800",  6449 => x"e0000005",
     6450 => x"ba200800",  6451 => x"ba001000",  6452 => x"fbffff99",
     6453 => x"b8205800",  6454 => x"b9600800",  6455 => x"2b9d0004",
     6456 => x"2b8b0020",  6457 => x"2b8c001c",  6458 => x"2b8d0018",
     6459 => x"2b8e0014",  6460 => x"2b8f0010",  6461 => x"2b90000c",
     6462 => x"2b910008",  6463 => x"379c0020",  6464 => x"c3a00000",
     6465 => x"379cfffc",  6466 => x"5b9d0004",  6467 => x"34020000",
     6468 => x"34030014",  6469 => x"f8002b85",  6470 => x"2b9d0004",
     6471 => x"379c0004",  6472 => x"c3a00000",  6473 => x"379cfff0",
     6474 => x"5b8b0010",  6475 => x"5b8c000c",  6476 => x"5b8d0008",
     6477 => x"5b9d0004",  6478 => x"b8206800",  6479 => x"28210020",
     6480 => x"282c0014",  6481 => x"282b000c",  6482 => x"28210010",
     6483 => x"0c200000",  6484 => x"34210004",  6485 => x"fbffffec",
     6486 => x"29a10020",  6487 => x"28210010",  6488 => x"34210018",
     6489 => x"fbffffe8",  6490 => x"b9800800",  6491 => x"34020000",
     6492 => x"34030020",  6493 => x"f8002b6d",  6494 => x"29610004",
     6495 => x"3402ffa0",  6496 => x"59810000",  6497 => x"29610008",
     6498 => x"59810004",  6499 => x"29610004",  6500 => x"59810010",
     6501 => x"29610008",  6502 => x"59810014",  6503 => x"2d61000e",
     6504 => x"0d810018",  6505 => x"2d610010",  6506 => x"0d81001a",
     6507 => x"41610012",  6508 => x"3181001c",  6509 => x"41610013",
     6510 => x"3181001d",  6511 => x"29a10020",  6512 => x"28210018",
     6513 => x"3022001c",  6514 => x"2b9d0004",  6515 => x"2b8b0010",
     6516 => x"2b8c000c",  6517 => x"2b8d0008",  6518 => x"379c0010",
     6519 => x"c3a00000",  6520 => x"379cff8c",  6521 => x"5b8b0018",
     6522 => x"5b8c0014",  6523 => x"5b8d0010",  6524 => x"5b8e000c",
     6525 => x"5b8f0008",  6526 => x"5b9d0004",  6527 => x"2c22010c",
     6528 => x"b8205800",  6529 => x"340d0000",  6530 => x"340c0001",
     6531 => x"5c400014",  6532 => x"28230000",  6533 => x"b8406800",
     6534 => x"34020006",  6535 => x"5c620010",  6536 => x"fbffffc1",
     6537 => x"29610000",  6538 => x"e0000105",  6539 => x"09820058",
     6540 => x"09a30058",  6541 => x"b9600800",  6542 => x"34420110",
     6543 => x"34630110",  6544 => x"b5621000",  6545 => x"b5631800",
     6546 => x"fbffff42",  6547 => x"48010002",  6548 => x"e0000002",
     6549 => x"b9806800",  6550 => x"358c0001",  6551 => x"2d66010c",
     6552 => x"48ccfff3",  6553 => x"78040001",  6554 => x"b9600800",
     6555 => x"34020003",  6556 => x"34030001",  6557 => x"38842b00",
     6558 => x"b9a02800",  6559 => x"fbffeb81",  6560 => x"1d61010e",
     6561 => x"442d0022",  6562 => x"0d6d010e",  6563 => x"296c0020",
     6564 => x"340f0000",  6565 => x"340e0001",  6566 => x"e0000015",
     6567 => x"29820000",  6568 => x"09c10374",  6569 => x"b4410800",
     6570 => x"2c23010c",  6571 => x"4460000f",  6572 => x"09e40374",
     6573 => x"1c23010e",  6574 => x"b4442000",  6575 => x"1c82010e",
     6576 => x"08630058",  6577 => x"08420058",  6578 => x"34630110",
     6579 => x"b4231800",  6580 => x"34420110",  6581 => x"b4821000",
     6582 => x"fbffff1e",  6583 => x"48010002",  6584 => x"e0000002",
     6585 => x"b9c07800",  6586 => x"35ce0001",  6587 => x"2981000c",
     6588 => x"2c21000c",  6589 => x"482effea",  6590 => x"2981001c",
     6591 => x"442f0004",  6592 => x"34010001",  6593 => x"598f001c",
     6594 => x"59810020",  6595 => x"4162001d",  6596 => x"34010002",
     6597 => x"44410063",  6598 => x"2d61010c",  6599 => x"5c200004",
     6600 => x"29620000",  6601 => x"34010004",  6602 => x"444100c5",
     6603 => x"29610020",  6604 => x"09ac0058",  6605 => x"2821000c",
     6606 => x"4023000a",  6607 => x"4022000b",  6608 => x"40290004",
     6609 => x"40280005",  6610 => x"40270006",  6611 => x"40260007",
     6612 => x"40250008",  6613 => x"40240009",  6614 => x"33830047",
     6615 => x"33890041",  6616 => x"33880042",  6617 => x"33870043",
     6618 => x"33860044",  6619 => x"33850045",  6620 => x"33840046",
     6621 => x"33820048",  6622 => x"2c22000e",  6623 => x"35830110",
     6624 => x"b5631800",  6625 => x"0f82003c",  6626 => x"2c220010",
     6627 => x"0f82003e",  6628 => x"40220012",  6629 => x"3382003a",
     6630 => x"40220013",  6631 => x"0f80004a",  6632 => x"33820040",
     6633 => x"28220004",  6634 => x"5b820068",  6635 => x"28210008",
     6636 => x"37820020",  6637 => x"5b81006c",  6638 => x"b9600800",
     6639 => x"fbfffee5",  6640 => x"4162001d",  6641 => x"34030001",
     6642 => x"44430029",  6643 => x"29620020",  6644 => x"78050001",
     6645 => x"38a53fa4",  6646 => x"2844000c",  6647 => x"1086000e",
     6648 => x"48060004",  6649 => x"48010023",  6650 => x"5c200019",
     6651 => x"e0000006",  6652 => x"48010020",  6653 => x"44200004",
     6654 => x"2c81000c",  6655 => x"5c23000a",  6656 => x"e0000028",
     6657 => x"78040001",  6658 => x"b9600800",  6659 => x"34020003",
     6660 => x"34030001",  6661 => x"38842b20",  6662 => x"fbffeb1a",
     6663 => x"34010002",  6664 => x"e0000087",  6665 => x"29630338",
     6666 => x"2841001c",  6667 => x"4461001d",  6668 => x"b56c1000",
     6669 => x"37810041",  6670 => x"34420131",  6671 => x"5b85001c",
     6672 => x"fbfffebd",  6673 => x"2b85001c",  6674 => x"5c20000c",
     6675 => x"78040001",  6676 => x"b9600800",  6677 => x"34020003",
     6678 => x"34030001",  6679 => x"38842b2c",  6680 => x"fbffeb08",
     6681 => x"34010007",  6682 => x"e0000075",  6683 => x"4c200003",
     6684 => x"b9600800",  6685 => x"fbffff2c",  6686 => x"78040001",
     6687 => x"78050001",  6688 => x"b9600800",  6689 => x"34020003",
     6690 => x"34030001",  6691 => x"38842b3c",  6692 => x"38a53fa4",
     6693 => x"fbffeafb",  6694 => x"34010006",  6695 => x"e0000068",
     6696 => x"09a30058",  6697 => x"29620020",  6698 => x"b5631800",
     6699 => x"2c64013a",  6700 => x"284c0018",  6701 => x"28410014",
     6702 => x"28420010",  6703 => x"34840001",  6704 => x"0c440000",
     6705 => x"34620150",  6706 => x"28450008",  6707 => x"2844000c",
     6708 => x"58250000",  6709 => x"58240004",  6710 => x"2c420010",
     6711 => x"0c220008",  6712 => x"34620128",  6713 => x"404e0009",
     6714 => x"4045000f",  6715 => x"40440010",  6716 => x"404a000a",
     6717 => x"4049000b",  6718 => x"4048000c",  6719 => x"4047000d",
     6720 => x"4046000e",  6721 => x"302e0010",  6722 => x"30250016",
     6723 => x"302a0011",  6724 => x"30290012",  6725 => x"30280013",
     6726 => x"30270014",  6727 => x"30260015",  6728 => x"30240017",
     6729 => x"28440004",  6730 => x"346e0120",  6731 => x"58240018",
     6732 => x"41c4000a",  6733 => x"3024001c",  6734 => x"40420008",
     6735 => x"3022001d",  6736 => x"4061013c",  6737 => x"3181001c",
     6738 => x"1dc50008",  6739 => x"1d810000",  6740 => x"4425000e",
     6741 => x"78040001",  6742 => x"b9600800",  6743 => x"34020003",
     6744 => x"34030001",  6745 => x"38842b48",  6746 => x"fbffeac6",
     6747 => x"2dc10008",  6748 => x"34020000",  6749 => x"0d810000",
     6750 => x"29610028",  6751 => x"28230004",  6752 => x"b9600800",
     6753 => x"d8600000",  6754 => x"09ad0058",  6755 => x"b56d0800",
     6756 => x"34210141",  6757 => x"4022000b",  6758 => x"20420004",
     6759 => x"7c420000",  6760 => x"59820004",  6761 => x"4022000b",
     6762 => x"20420002",  6763 => x"7c420000",  6764 => x"59820008",
     6765 => x"4022000b",  6766 => x"20420001",  6767 => x"5982000c",
     6768 => x"4022000b",  6769 => x"20420010",  6770 => x"7c420000",
     6771 => x"59820010",  6772 => x"4022000b",  6773 => x"20420020",
     6774 => x"7c420000",  6775 => x"59820014",  6776 => x"4021000b",
     6777 => x"20210008",  6778 => x"7c210000",  6779 => x"59810018",
     6780 => x"78010001",  6781 => x"382149c4",  6782 => x"2824001c",
     6783 => x"44800007",  6784 => x"b56d1000",  6785 => x"b8406800",
     6786 => x"b9600800",  6787 => x"34420144",  6788 => x"35a3011c",
     6789 => x"d8800000",  6790 => x"78040001",  6791 => x"78050001",
     6792 => x"b9600800",  6793 => x"34020003",  6794 => x"34030001",
     6795 => x"38842b5c",  6796 => x"38a53fa4",  6797 => x"fbffea93",
     6798 => x"34010009",  6799 => x"2b9d0004",  6800 => x"2b8b0018",
     6801 => x"2b8c0014",  6802 => x"2b8d0010",  6803 => x"2b8e000c",
     6804 => x"2b8f0008",  6805 => x"379c0074",  6806 => x"c3a00000",
     6807 => x"379cffec",  6808 => x"5b8b0014",  6809 => x"5b8c0010",
     6810 => x"5b8d000c",  6811 => x"5b8e0008",  6812 => x"5b9d0004",
     6813 => x"b8406000",  6814 => x"28220024",  6815 => x"b8607000",
     6816 => x"28230070",  6817 => x"2847000c",  6818 => x"28220034",
     6819 => x"b8806800",  6820 => x"b5831800",  6821 => x"342400f8",
     6822 => x"b9a02800",  6823 => x"34060000",  6824 => x"b8205800",
     6825 => x"d8e00000",  6826 => x"78070001",  6827 => x"38e749fc",
     6828 => x"3dc20002",  6829 => x"4c2c000c",  6830 => x"b4e23800",
     6831 => x"28e50000",  6832 => x"78040001",  6833 => x"b9600800",
     6834 => x"34020005",  6835 => x"34030001",  6836 => x"38842794",
     6837 => x"b9c03000",  6838 => x"fbffea6a",  6839 => x"3401ffff",
     6840 => x"e0000014",  6841 => x"b4e24000",  6842 => x"296600f8",
     6843 => x"296700fc",  6844 => x"29080000",  6845 => x"78040001",
     6846 => x"b9600800",  6847 => x"34020005",  6848 => x"34030001",
     6849 => x"388427b4",  6850 => x"b9802800",  6851 => x"fbffea5d",
     6852 => x"34010001",  6853 => x"5da10003",  6854 => x"29620104",
     6855 => x"44400005",  6856 => x"2961036c",  6857 => x"34210001",
     6858 => x"5961036c",  6859 => x"34010000",  6860 => x"2b9d0004",
     6861 => x"2b8b0014",  6862 => x"2b8c0010",  6863 => x"2b8d000c",
     6864 => x"2b8e0008",  6865 => x"379c0014",  6866 => x"c3a00000",
     6867 => x"379cfff0",  6868 => x"5b8b0010",  6869 => x"5b8c000c",
     6870 => x"5b8d0008",  6871 => x"5b9d0004",  6872 => x"b8205800",
     6873 => x"40410000",  6874 => x"b8406000",  6875 => x"34030002",
     6876 => x"00210004",  6877 => x"356d0320",  6878 => x"3161030c",
     6879 => x"40410000",  6880 => x"2021000f",  6881 => x"3161030d",
     6882 => x"40410001",  6883 => x"2021000f",  6884 => x"3161030e",
     6885 => x"2c410002",  6886 => x"0d610310",  6887 => x"40410004",
     6888 => x"34420006",  6889 => x"31610312",  6890 => x"35610313",
     6891 => x"f8002961",  6892 => x"35820008",  6893 => x"34030004",
     6894 => x"3561031c",  6895 => x"f800295d",  6896 => x"3582000c",
     6897 => x"34030004",  6898 => x"35610318",  6899 => x"f8002959",
     6900 => x"35820014",  6901 => x"34030008",  6902 => x"b9a00800",
     6903 => x"f8002955",  6904 => x"2d81001c",  6905 => x"296202c8",
     6906 => x"34030008",  6907 => x"0d610328",  6908 => x"2d81001e",
     6909 => x"0d61032a",  6910 => x"41810020",  6911 => x"3161032c",
     6912 => x"41810021",  6913 => x"3161032d",  6914 => x"b9a00800",
     6915 => x"f8002928",  6916 => x"3403ffff",  6917 => x"44200015",
     6918 => x"29610020",  6919 => x"28210014",  6920 => x"2c220008",
     6921 => x"4440000a",  6922 => x"b9a01000",  6923 => x"34030008",
     6924 => x"f800291f",  6925 => x"5c200009",  6926 => x"29610020",
     6927 => x"28210014",  6928 => x"2c220008",  6929 => x"2d610328",
     6930 => x"5c410004",  6931 => x"4161001c",  6932 => x"38210001",
     6933 => x"e0000003",  6934 => x"4161001c",  6935 => x"202100fe",
     6936 => x"3161001c",  6937 => x"34030000",  6938 => x"b8600800",
     6939 => x"2b9d0004",  6940 => x"2b8b0010",  6941 => x"2b8c000c",
     6942 => x"2b8d0008",  6943 => x"379c0010",  6944 => x"c3a00000",
     6945 => x"379cfff4",  6946 => x"5b8b000c",  6947 => x"5b8c0008",
     6948 => x"5b9d0004",  6949 => x"30400000",  6950 => x"b8206000",
     6951 => x"282102c8",  6952 => x"b8405800",  6953 => x"34030008",
     6954 => x"4021000e",  6955 => x"30410001",  6956 => x"29810020",
     6957 => x"2821000c",  6958 => x"40210014",  6959 => x"30410004",
     6960 => x"34010002",  6961 => x"30410006",  6962 => x"34410008",
     6963 => x"34020000",  6964 => x"f8002996",  6965 => x"298202c8",
     6966 => x"35610014",  6967 => x"34030008",  6968 => x"f8002914",
     6969 => x"298102c8",  6970 => x"2c210008",  6971 => x"0d61001c",
     6972 => x"3401007f",  6973 => x"31610021",  6974 => x"2b9d0004",
     6975 => x"2b8b000c",  6976 => x"2b8c0008",  6977 => x"379c000c",
     6978 => x"c3a00000",  6979 => x"2c230022",  6980 => x"0c430004",
     6981 => x"28230024",  6982 => x"58430000",  6983 => x"28210028",
     6984 => x"58410008",  6985 => x"c3a00000",  6986 => x"379cfff4",
     6987 => x"5b8b000c",  6988 => x"5b8c0008",  6989 => x"5b9d0004",
     6990 => x"b8205800",  6991 => x"2c210022",  6992 => x"b8406000",
     6993 => x"34030008",  6994 => x"0c410004",  6995 => x"29610024",
     6996 => x"58410000",  6997 => x"29610028",  6998 => x"58410008",
     6999 => x"2d61002c",  7000 => x"0c41000c",  7001 => x"4161002f",
     7002 => x"3041000e",  7003 => x"41610030",  7004 => x"30410010",
     7005 => x"41610031",  7006 => x"30410011",  7007 => x"2d610032",
     7008 => x"0c410012",  7009 => x"41610034",  7010 => x"30410014",
     7011 => x"34410015",  7012 => x"35620035",  7013 => x"f80028e7",
     7014 => x"2d61003d",  7015 => x"0d81001e",  7016 => x"4161003f",
     7017 => x"31810020",  7018 => x"78010001",  7019 => x"382149c4",
     7020 => x"28230030",  7021 => x"44600004",  7022 => x"b9600800",
     7023 => x"b9801000",  7024 => x"d8600000",  7025 => x"2b9d0004",
     7026 => x"2b8b000c",  7027 => x"2b8c0008",  7028 => x"379c000c",
     7029 => x"c3a00000",  7030 => x"2c230022",  7031 => x"0c430004",
     7032 => x"28230024",  7033 => x"58430000",  7034 => x"28210028",
     7035 => x"58410008",  7036 => x"c3a00000",  7037 => x"379cfff4",
     7038 => x"5b8b000c",  7039 => x"5b8c0008",  7040 => x"5b9d0004",
     7041 => x"b8205800",  7042 => x"2c210022",  7043 => x"b8406000",
     7044 => x"34030008",  7045 => x"0c410004",  7046 => x"29610024",
     7047 => x"58410000",  7048 => x"29610028",  7049 => x"58410008",
     7050 => x"3441000c",  7051 => x"3562002c",  7052 => x"f80028c0",
     7053 => x"2d610034",  7054 => x"0d810014",  7055 => x"2b9d0004",
     7056 => x"2b8b000c",  7057 => x"2b8c0008",  7058 => x"379c000c",
     7059 => x"c3a00000",  7060 => x"379cfff4",  7061 => x"5b8b000c",
     7062 => x"5b8c0008",  7063 => x"5b9d0004",  7064 => x"282b003c",
     7065 => x"b8206000",  7066 => x"34020000",  7067 => x"41610000",
     7068 => x"3403000a",  7069 => x"202100f0",  7070 => x"3821000b",
     7071 => x"31610000",  7072 => x"34010040",  7073 => x"0d610002",
     7074 => x"2d810306",  7075 => x"34210001",  7076 => x"2021ffff",
     7077 => x"0d810306",  7078 => x"0d61001e",  7079 => x"34010005",
     7080 => x"31610020",  7081 => x"298102c8",  7082 => x"4021000b",
     7083 => x"31610021",  7084 => x"35610022",  7085 => x"f800291d",
     7086 => x"29810020",  7087 => x"34030008",  7088 => x"28220018",
     7089 => x"28210014",  7090 => x"2c420000",  7091 => x"0d62002c",
     7092 => x"4021001c",  7093 => x"3161002f",  7094 => x"29810020",
     7095 => x"28210014",  7096 => x"40210018",  7097 => x"31610030",
     7098 => x"29810020",  7099 => x"28210014",  7100 => x"40210019",
     7101 => x"31610031",  7102 => x"29810020",  7103 => x"28210014",
     7104 => x"2c22001a",  7105 => x"0d620032",  7106 => x"4021001d",
     7107 => x"31610034",  7108 => x"29810020",  7109 => x"28220014",
     7110 => x"35610035",  7111 => x"34420010",  7112 => x"f8002884",
     7113 => x"29810020",  7114 => x"28220010",  7115 => x"28210018",
     7116 => x"2c420000",  7117 => x"0d62003d",  7118 => x"4021001c",
     7119 => x"34020040",  7120 => x"3161003f",  7121 => x"78010001",
     7122 => x"382149c4",  7123 => x"2823002c",  7124 => x"44600004",
     7125 => x"b9800800",  7126 => x"d8600000",  7127 => x"b8201000",
     7128 => x"b9800800",  7129 => x"3403000b",  7130 => x"34040000",
     7131 => x"fbfffebc",  7132 => x"2b9d0004",  7133 => x"2b8b000c",
     7134 => x"2b8c0008",  7135 => x"379c000c",  7136 => x"c3a00000",
     7137 => x"379cffc8",  7138 => x"5b8b0018",  7139 => x"5b8c0014",
     7140 => x"5b8d0010",  7141 => x"5b8e000c",  7142 => x"5b8f0008",
     7143 => x"5b9d0004",  7144 => x"28220028",  7145 => x"378c001c",
     7146 => x"b8205800",  7147 => x"28430000",  7148 => x"b9801000",
     7149 => x"378f0030",  7150 => x"d8600000",  7151 => x"b9800800",
     7152 => x"b9e01000",  7153 => x"f8000103",  7154 => x"296c003c",
     7155 => x"340efff0",  7156 => x"340d002c",  7157 => x"41810000",
     7158 => x"0d8d0002",  7159 => x"34020000",  7160 => x"a02e0800",
     7161 => x"31810000",  7162 => x"2d6102f0",  7163 => x"34030008",
     7164 => x"34210001",  7165 => x"2021ffff",  7166 => x"0d6102f0",
     7167 => x"31800020",  7168 => x"0d81001e",  7169 => x"296102c8",
     7170 => x"4021000d",  7171 => x"31810021",  7172 => x"35810008",
     7173 => x"f80028c5",  7174 => x"2f810034",  7175 => x"3402002c",
     7176 => x"34030000",  7177 => x"0d810022",  7178 => x"2b810030",
     7179 => x"34040001",  7180 => x"59810024",  7181 => x"2b810038",
     7182 => x"59810028",  7183 => x"b9600800",  7184 => x"fbfffe87",
     7185 => x"5c200023",  7186 => x"29610020",  7187 => x"356c00f8",
     7188 => x"b9801000",  7189 => x"28230008",  7190 => x"b9800800",
     7191 => x"34630018",  7192 => x"f8000101",  7193 => x"b9e01000",
     7194 => x"b9800800",  7195 => x"f80000d9",  7196 => x"2961003c",
     7197 => x"34030008",  7198 => x"34040000",  7199 => x"40220000",
     7200 => x"0c2d0002",  7201 => x"a04e7000",  7202 => x"39ce0008",
     7203 => x"302e0000",  7204 => x"2d6202f0",  7205 => x"0c22001e",
     7206 => x"34020002",  7207 => x"30220020",  7208 => x"296202c8",
     7209 => x"4042000d",  7210 => x"30220021",  7211 => x"2f820034",
     7212 => x"0c220022",  7213 => x"2b820030",  7214 => x"58220024",
     7215 => x"2b820038",  7216 => x"58220028",  7217 => x"b9600800",
     7218 => x"3402002c",  7219 => x"fbfffe64",  7220 => x"2b9d0004",
     7221 => x"2b8b0018",  7222 => x"2b8c0014",  7223 => x"2b8d0010",
     7224 => x"2b8e000c",  7225 => x"2b8f0008",  7226 => x"379c0038",
     7227 => x"c3a00000",  7228 => x"379cffd4",  7229 => x"5b8b000c",
     7230 => x"5b8c0008",  7231 => x"5b9d0004",  7232 => x"28220028",
     7233 => x"378b0010",  7234 => x"b8206000",  7235 => x"28430000",
     7236 => x"b9601000",  7237 => x"d8600000",  7238 => x"37820024",
     7239 => x"b9600800",  7240 => x"f80000ac",  7241 => x"298b003c",
     7242 => x"34020000",  7243 => x"34030008",  7244 => x"41610000",
     7245 => x"202100f0",  7246 => x"38210001",  7247 => x"31610000",
     7248 => x"3401002c",  7249 => x"0d610002",  7250 => x"2d8102f2",
     7251 => x"34210001",  7252 => x"2021ffff",  7253 => x"0d8102f2",
     7254 => x"0d61001e",  7255 => x"34010001",  7256 => x"31610020",
     7257 => x"3401007f",  7258 => x"31610021",  7259 => x"35610008",
     7260 => x"f800286e",  7261 => x"2f810028",  7262 => x"3402002c",
     7263 => x"34030001",  7264 => x"0d610022",  7265 => x"2b810024",
     7266 => x"34040001",  7267 => x"59610024",  7268 => x"2b81002c",
     7269 => x"59610028",  7270 => x"b9800800",  7271 => x"fbfffe30",
     7272 => x"2b9d0004",  7273 => x"2b8b000c",  7274 => x"2b8c0008",
     7275 => x"379c002c",  7276 => x"c3a00000",  7277 => x"379cffe8",
     7278 => x"5b8b000c",  7279 => x"5b8c0008",  7280 => x"5b9d0004",
     7281 => x"b8206000",  7282 => x"b8400800",  7283 => x"37820010",
     7284 => x"f8000080",  7285 => x"298b003c",  7286 => x"34020000",
     7287 => x"34030008",  7288 => x"41610000",  7289 => x"202100f0",
     7290 => x"38210009",  7291 => x"31610000",  7292 => x"34010036",
     7293 => x"0d610002",  7294 => x"41810312",  7295 => x"31610004",
     7296 => x"35610008",  7297 => x"f8002849",  7298 => x"2981031c",
     7299 => x"35820320",  7300 => x"34030008",  7301 => x"59610008",
     7302 => x"29810318",  7303 => x"5961000c",  7304 => x"2d81032a",
     7305 => x"0d61001e",  7306 => x"34010003",  7307 => x"31610020",
     7308 => x"298102c8",  7309 => x"4021000a",  7310 => x"31610021",
     7311 => x"2f810014",  7312 => x"0d610022",  7313 => x"2b810010",
     7314 => x"59610024",  7315 => x"2b810018",  7316 => x"59610028",
     7317 => x"3561002c",  7318 => x"f80027b6",  7319 => x"2d810328",
     7320 => x"34020036",  7321 => x"34030009",  7322 => x"0d610034",
     7323 => x"34040000",  7324 => x"b9800800",  7325 => x"fbfffdfa",
     7326 => x"2b9d0004",  7327 => x"2b8b000c",  7328 => x"2b8c0008",
     7329 => x"379c0018",  7330 => x"c3a00000",  7331 => x"379cfff0",
     7332 => x"5b8b0010",  7333 => x"5b8c000c",  7334 => x"5b8d0008",
     7335 => x"5b9d0004",  7336 => x"78030001",  7337 => x"282d0004",
     7338 => x"38633cc8",  7339 => x"28620000",  7340 => x"b8205800",
     7341 => x"b9a00800",  7342 => x"f80026f0",  7343 => x"78030001",
     7344 => x"296c0000",  7345 => x"38633cc8",  7346 => x"28620000",
     7347 => x"b42c6000",  7348 => x"596c0000",  7349 => x"b9a00800",
     7350 => x"f8002715",  7351 => x"59610004",  7352 => x"4c0c0007",
     7353 => x"4c20000f",  7354 => x"358cffff",  7355 => x"78030001",
     7356 => x"596c0000",  7357 => x"38633cc8",  7358 => x"e0000007",
     7359 => x"45800009",  7360 => x"4c010008",  7361 => x"358c0001",
     7362 => x"78030001",  7363 => x"596c0000",  7364 => x"38633cd8",
     7365 => x"28620000",  7366 => x"b4220800",  7367 => x"59610004",
     7368 => x"2b9d0004",  7369 => x"2b8b0010",  7370 => x"2b8c000c",
     7371 => x"2b8d0008",  7372 => x"379c0010",  7373 => x"c3a00000",
     7374 => x"379cffe8",  7375 => x"5b8b0008",  7376 => x"5b9d0004",
     7377 => x"5b82000c",  7378 => x"5b830010",  7379 => x"5b830014",
     7380 => x"5b820018",  7381 => x"b8205800",  7382 => x"4c600006",
     7383 => x"78010001",  7384 => x"78020001",  7385 => x"38212bdc",
     7386 => x"38423fb8",  7387 => x"f8000e99",  7388 => x"2b810018",
     7389 => x"38028000",  7390 => x"2b830014",  7391 => x"b4221000",
     7392 => x"f4220800",  7393 => x"00420010",  7394 => x"b4230800",
     7395 => x"3c230010",  7396 => x"00210010",  7397 => x"b8431000",
     7398 => x"78030001",  7399 => x"38633cc8",  7400 => x"5b820018",
     7401 => x"28620000",  7402 => x"5b810014",  7403 => x"37810014",
     7404 => x"fbffec79",  7405 => x"59610004",  7406 => x"2b810018",
     7407 => x"59610000",  7408 => x"2b9d0004",  7409 => x"2b8b0008",
     7410 => x"379c0018",  7411 => x"c3a00000",  7412 => x"379cfffc",
     7413 => x"5b9d0004",  7414 => x"28230000",  7415 => x"48030003",
     7416 => x"28210004",  7417 => x"4c200006",  7418 => x"78010001",
     7419 => x"38212c08",  7420 => x"f8000e78",  7421 => x"3401ffff",
     7422 => x"e0000005",  7423 => x"58410008",  7424 => x"58430000",
     7425 => x"0c400004",  7426 => x"34010000",  7427 => x"2b9d0004",
     7428 => x"379c0004",  7429 => x"c3a00000",  7430 => x"379cfffc",
     7431 => x"5b9d0004",  7432 => x"78050001",  7433 => x"38a53cdc",
     7434 => x"28430000",  7435 => x"28a40000",  7436 => x"54640006",
     7437 => x"28420008",  7438 => x"58230000",  7439 => x"58220004",
     7440 => x"34010000",  7441 => x"e0000005",  7442 => x"78010001",
     7443 => x"38212c44",  7444 => x"f8000e60",  7445 => x"3401ffff",
     7446 => x"2b9d0004",  7447 => x"379c0004",  7448 => x"c3a00000",
     7449 => x"379cfffc",  7450 => x"5b9d0004",  7451 => x"28660000",
     7452 => x"28450000",  7453 => x"28630004",  7454 => x"28420004",
     7455 => x"b4c52800",  7456 => x"58250000",  7457 => x"b4621000",
     7458 => x"58220004",  7459 => x"fbffff80",  7460 => x"2b9d0004",
     7461 => x"379c0004",  7462 => x"c3a00000",  7463 => x"379cfffc",
     7464 => x"5b9d0004",  7465 => x"28460000",  7466 => x"28650000",
     7467 => x"c8c52800",  7468 => x"58250000",  7469 => x"28450004",
     7470 => x"28620004",  7471 => x"c8a21000",  7472 => x"58220004",
     7473 => x"fbffff72",  7474 => x"2b9d0004",  7475 => x"379c0004",
     7476 => x"c3a00000",  7477 => x"379cfffc",  7478 => x"5b9d0004",
     7479 => x"78040001",  7480 => x"38843ce0",  7481 => x"28230000",
     7482 => x"28820000",  7483 => x"a0621000",  7484 => x"4c400005",
     7485 => x"3442ffff",  7486 => x"3404fffe",  7487 => x"b8441000",
     7488 => x"34420001",  7489 => x"78050001",  7490 => x"38a53cc8",
     7491 => x"28a40000",  7492 => x"88441000",  7493 => x"28240004",
     7494 => x"b4441000",  7495 => x"0064001f",  7496 => x"b4831800",
     7497 => x"14630001",  7498 => x"58230000",  7499 => x"0043001f",
     7500 => x"b4621000",  7501 => x"14420001",  7502 => x"58220004",
     7503 => x"fbffff54",  7504 => x"2b9d0004",  7505 => x"379c0004",
     7506 => x"c3a00000",  7507 => x"379cfff8",  7508 => x"5b8b0008",
     7509 => x"5b9d0004",  7510 => x"28250000",  7511 => x"78030001",
     7512 => x"b8201000",  7513 => x"38632c94",  7514 => x"4805000a",
     7515 => x"78030001",  7516 => x"38631c28",  7517 => x"5ca00007",
     7518 => x"28210004",  7519 => x"78030001",  7520 => x"38632c94",
     7521 => x"48a10003",  7522 => x"78030001",  7523 => x"38631c28",
     7524 => x"28410004",  7525 => x"14a4001f",  7526 => x"780b0001",
     7527 => x"1426001f",  7528 => x"98853800",  7529 => x"396b5214",
     7530 => x"98c12800",  7531 => x"78020001",  7532 => x"b9600800",
     7533 => x"38422c98",  7534 => x"c8e42000",  7535 => x"c8a62800",
     7536 => x"f8000df6",  7537 => x"b9600800",  7538 => x"2b9d0004",
     7539 => x"2b8b0008",  7540 => x"379c0008",  7541 => x"c3a00000",
     7542 => x"379cfff8",  7543 => x"5b8b0008",  7544 => x"5b9d0004",
     7545 => x"28220020",  7546 => x"28240028",  7547 => x"b8205800",
     7548 => x"28430004",  7549 => x"58600038",  7550 => x"28430014",
     7551 => x"0c20010c",  7552 => x"0c600008",  7553 => x"28830014",
     7554 => x"44600013",  7555 => x"d8600000",  7556 => x"3402ffff",
     7557 => x"5c220008",  7558 => x"78040001",  7559 => x"b9600800",
     7560 => x"34020004",  7561 => x"34030001",  7562 => x"38842ca4",
     7563 => x"fbffe795",  7564 => x"34010000",  7565 => x"29620020",
     7566 => x"c8010800",  7567 => x"3c21000a",  7568 => x"28420004",
     7569 => x"1423001f",  7570 => x"5841002c",  7571 => x"58430028",
     7572 => x"e000000d",  7573 => x"28420008",  7574 => x"28420038",
     7575 => x"20420001",  7576 => x"5c430005",  7577 => x"28840008",
     7578 => x"34020000",  7579 => x"34030000",  7580 => x"d8800000",
     7581 => x"29610020",  7582 => x"28210004",  7583 => x"58200028",
     7584 => x"5820002c",  7585 => x"29610020",  7586 => x"78040001",
     7587 => x"34020004",  7588 => x"28260004",  7589 => x"34030001",
     7590 => x"b9600800",  7591 => x"28c50028",  7592 => x"28c6002c",
     7593 => x"38842cc0",  7594 => x"fbffe776",  7595 => x"2b9d0004",
     7596 => x"2b8b0008",  7597 => x"379c0008",  7598 => x"c3a00000",
     7599 => x"379cfff0",  7600 => x"5b8b0010",  7601 => x"5b8c000c",
     7602 => x"5b8d0008",  7603 => x"5b9d0004",  7604 => x"b8205800",
     7605 => x"28210020",  7606 => x"35620094",  7607 => x"35630080",
     7608 => x"282d0004",  7609 => x"356c00d0",  7610 => x"b9a00800",
     7611 => x"fbffff6c",  7612 => x"b9a01000",  7613 => x"b9801800",
     7614 => x"b9a00800",  7615 => x"fbffff68",  7616 => x"b9800800",
     7617 => x"fbffff92",  7618 => x"78040001",  7619 => x"b8202800",
     7620 => x"34020004",  7621 => x"b9600800",  7622 => x"34030003",
     7623 => x"38842ce0",  7624 => x"fbffe758",  7625 => x"2b9d0004",
     7626 => x"2b8b0010",  7627 => x"2b8c000c",  7628 => x"2b8d0008",
     7629 => x"379c0010",  7630 => x"c3a00000",  7631 => x"379cffb8",
     7632 => x"5b8b0024",  7633 => x"5b8c0020",  7634 => x"5b8d001c",
     7635 => x"5b8e0018",  7636 => x"5b8f0014",  7637 => x"5b900010",
     7638 => x"5b91000c",  7639 => x"5b920008",  7640 => x"5b9d0004",
     7641 => x"28220020",  7642 => x"b8205800",  7643 => x"284d0004",
     7644 => x"284c0010",  7645 => x"28220080",  7646 => x"5c400008",
     7647 => x"28230084",  7648 => x"5c620006",  7649 => x"78040001",
     7650 => x"34020004",  7651 => x"34030002",  7652 => x"38842cf8",
     7653 => x"e000006e",  7654 => x"35af0014",  7655 => x"357000bc",
     7656 => x"357100a8",  7657 => x"b9e00800",  7658 => x"ba001000",
     7659 => x"ba201800",  7660 => x"fbffff3b",  7661 => x"357200d0",
     7662 => x"b9e01000",  7663 => x"ba401800",  7664 => x"b9e00800",
     7665 => x"fbffff36",  7666 => x"ba400800",  7667 => x"fbffff60",
     7668 => x"78040001",  7669 => x"b8202800",  7670 => x"34020004",
     7671 => x"34030003",  7672 => x"38842d18",  7673 => x"b9600800",
     7674 => x"fbffe726",  7675 => x"35610080",  7676 => x"fbffff57",
     7677 => x"78040001",  7678 => x"b8202800",  7679 => x"34020004",
     7680 => x"34030002",  7681 => x"38842d30",  7682 => x"b9600800",
     7683 => x"fbffe71d",  7684 => x"35610094",  7685 => x"fbffff4e",
     7686 => x"78040001",  7687 => x"b8202800",  7688 => x"34020004",
     7689 => x"34030002",  7690 => x"38842d38",  7691 => x"b9600800",
     7692 => x"fbffe714",  7693 => x"ba200800",  7694 => x"fbffff45",
     7695 => x"78040001",  7696 => x"b8202800",  7697 => x"34020004",
     7698 => x"34030002",  7699 => x"38842d40",  7700 => x"b9600800",
     7701 => x"fbffe70b",  7702 => x"ba000800",  7703 => x"fbffff3c",
     7704 => x"78040001",  7705 => x"b8202800",  7706 => x"34020004",
     7707 => x"34030002",  7708 => x"38842d48",  7709 => x"b9600800",
     7710 => x"fbffe702",  7711 => x"b9a00800",  7712 => x"fbffff33",
     7713 => x"78040001",  7714 => x"b8202800",  7715 => x"34020004",
     7716 => x"34030001",  7717 => x"38842d50",  7718 => x"b9600800",
     7719 => x"fbffe6f9",  7720 => x"b9e00800",  7721 => x"fbffff2a",
     7722 => x"78040001",  7723 => x"b8202800",  7724 => x"38842d68",
     7725 => x"b9600800",  7726 => x"34020004",  7727 => x"34030001",
     7728 => x"fbffe6f0",  7729 => x"29610020",  7730 => x"358e0018",
     7731 => x"28220004",  7732 => x"b9c00800",  7733 => x"34430014",
     7734 => x"fbfffee3",  7735 => x"b9c00800",  7736 => x"fbfffefd",
     7737 => x"b9c00800",  7738 => x"fbffff19",  7739 => x"78040001",
     7740 => x"b8202800",  7741 => x"34020004",  7742 => x"b9600800",
     7743 => x"34030001",  7744 => x"38842d80",  7745 => x"fbffe6df",
     7746 => x"29610020",  7747 => x"28220010",  7748 => x"28260004",
     7749 => x"28420018",  7750 => x"5c400142",  7751 => x"28210008",
     7752 => x"28270030",  7753 => x"44e2013c",  7754 => x"28c20000",
     7755 => x"5c400003",  7756 => x"28c30014",  7757 => x"44620008",
     7758 => x"78040001",  7759 => x"b9600800",  7760 => x"34020004",
     7761 => x"34030001",  7762 => x"38842d94",  7763 => x"fbffe6cd",
     7764 => x"e0000134",  7765 => x"28c50004",  7766 => x"48a70003",
     7767 => x"28c20018",  7768 => x"4ce2012d",  7769 => x"28c60018",
     7770 => x"78040001",  7771 => x"b9600800",  7772 => x"34020004",
     7773 => x"34030001",  7774 => x"38842dc0",  7775 => x"fbffe6c1",
     7776 => x"e0000128",  7777 => x"2982001c",  7778 => x"59a20034",
     7779 => x"1c220040",  7780 => x"29a10034",  7781 => x"3444ffff",
     7782 => x"1423001f",  7783 => x"98612800",  7784 => x"c8a32800",
     7785 => x"3403001f",  7786 => x"c8621800",  7787 => x"94a33800",
     7788 => x"34820001",  7789 => x"34630001",  7790 => x"3484ffff",
     7791 => x"5ce0fffc",  7792 => x"34030001",  7793 => x"bc621000",
     7794 => x"4c460002",  7795 => x"59a20038",  7796 => x"29a30038",
     7797 => x"4c620003",  7798 => x"34630001",  7799 => x"59a30038",
     7800 => x"2982001c",  7801 => x"4c400002",  7802 => x"5981001c",
     7803 => x"2982001c",  7804 => x"4c400002",  7805 => x"5980001c",
     7806 => x"2985001c",  7807 => x"08210003",  7808 => x"4c25000d",
     7809 => x"78040001",  7810 => x"b9600800",  7811 => x"34020004",
     7812 => x"34030001",  7813 => x"38842e04",  7814 => x"fbffe69a",
     7815 => x"29a10034",  7816 => x"29a20038",  7817 => x"3c210001",
     7818 => x"34420001",  7819 => x"b4410800",  7820 => x"5981001c",
     7821 => x"29af0038",  7822 => x"29a20034",  7823 => x"35900004",
     7824 => x"35e1ffff",  7825 => x"88220800",  7826 => x"2982001c",
     7827 => x"b4220800",  7828 => x"b9e01000",  7829 => x"f8002509",
     7830 => x"59a10034",  7831 => x"78040001",  7832 => x"b8203000",
     7833 => x"b9e02800",  7834 => x"38842e1c",  7835 => x"5981001c",
     7836 => x"34020004",  7837 => x"b9600800",  7838 => x"34030001",
     7839 => x"fbffe681",  7840 => x"b9a01000",  7841 => x"b9c01800",
     7842 => x"ba000800",  7843 => x"fbfffe84",  7844 => x"ba000800",
     7845 => x"fbfffeae",  7846 => x"78040001",  7847 => x"b8202800",
     7848 => x"34020004",  7849 => x"b9600800",  7850 => x"34030001",
     7851 => x"38842e40",  7852 => x"fbffe674",  7853 => x"296f0020",
     7854 => x"29e10008",  7855 => x"2825002c",  7856 => x"44a00011",
     7857 => x"29820004",  7858 => x"44400007",  7859 => x"78040001",
     7860 => x"b9600800",  7861 => x"34020004",  7862 => x"34030001",
     7863 => x"38842e5c",  7864 => x"e3ffff9b",  7865 => x"29820008",
     7866 => x"4ca20007",  7867 => x"78040001",  7868 => x"b9600800",
     7869 => x"34020004",  7870 => x"34030001",  7871 => x"38842e8c",
     7872 => x"e00000c3",  7873 => x"29820004",  7874 => x"44400031",
     7875 => x"28220038",  7876 => x"20410001",  7877 => x"5c2000c3",
     7878 => x"20420002",  7879 => x"5c410019",  7880 => x"296300c4",
     7881 => x"296200c8",  7882 => x"296100cc",  7883 => x"5b830030",
     7884 => x"29e30010",  7885 => x"296500bc",  7886 => x"296400c0",
     7887 => x"378c0028",  7888 => x"5b820034",  7889 => x"5b810038",
     7890 => x"b9801000",  7891 => x"b9800800",  7892 => x"34630018",
     7893 => x"5b850028",  7894 => x"5b84002c",  7895 => x"fbfffe42",
     7896 => x"29610028",  7897 => x"b9801000",  7898 => x"28230004",
     7899 => x"b9600800",  7900 => x"d8600000",  7901 => x"b9600800",
     7902 => x"fbfffe98",  7903 => x"e00000a9",  7904 => x"29820008",
     7905 => x"78030001",  7906 => x"38633ce4",  7907 => x"28610000",
     7908 => x"ec021000",  7909 => x"78050001",  7910 => x"c8021000",
     7911 => x"38a53ce8",  7912 => x"a0411000",  7913 => x"28a10000",
     7914 => x"b4411000",  7915 => x"29610028",  7916 => x"c8021000",
     7917 => x"28230010",  7918 => x"5c600002",  7919 => x"2823000c",
     7920 => x"b9600800",  7921 => x"d8600000",  7922 => x"e0000096",
     7923 => x"29830008",  7924 => x"29ed0004",  7925 => x"78050001",
     7926 => x"1462001f",  7927 => x"29b0002c",  7928 => x"00640016",
     7929 => x"3c63000a",  7930 => x"29ae0028",  7931 => x"3c42000a",
     7932 => x"b4708000",  7933 => x"b8821000",  7934 => x"f4701800",
     7935 => x"b44e1000",  7936 => x"b4627000",  7937 => x"1c22003e",
     7938 => x"38a53ce8",  7939 => x"28a40000",  7940 => x"1441001f",
     7941 => x"34030000",  7942 => x"59ae0028",  7943 => x"59b0002c",
     7944 => x"f800246f",  7945 => x"00430016",  7946 => x"3c21000a",
     7947 => x"3c42000a",  7948 => x"b8610800",  7949 => x"49c1000b",
     7950 => x"5dc10002",  7951 => x"56020009",  7952 => x"c8021000",
     7953 => x"7c430000",  7954 => x"c8010800",  7955 => x"c8230800",
     7956 => x"482e0004",  7957 => x"5c2e0005",  7958 => x"54500002",
     7959 => x"e0000003",  7960 => x"59a10028",  7961 => x"59a2002c",
     7962 => x"29a10028",  7963 => x"29a2002c",  7964 => x"48200003",
     7965 => x"5c200004",  7966 => x"44410003",  7967 => x"340d0000",
     7968 => x"e0000002",  7969 => x"340dffff",  7970 => x"5b810044",
     7971 => x"5b820048",  7972 => x"45a00007",  7973 => x"c8021000",
     7974 => x"7c430000",  7975 => x"c8010800",  7976 => x"c8230800",
     7977 => x"5b810044",  7978 => x"5b820048",  7979 => x"29e20008",
     7980 => x"37810044",  7981 => x"1c42003e",  7982 => x"fbffea37",
     7983 => x"45a00009",  7984 => x"2b810048",  7985 => x"2b820044",
     7986 => x"c8010800",  7987 => x"7c230000",  7988 => x"c8021000",
     7989 => x"c8431000",  7990 => x"5b820044",  7991 => x"5b810048",
     7992 => x"29820008",  7993 => x"1441001f",  7994 => x"00430016",
     7995 => x"3c21000a",  7996 => x"ec026000",  7997 => x"3c42000a",
     7998 => x"b8610800",  7999 => x"c80c6000",  8000 => x"5b81003c",
     8001 => x"5b820040",  8002 => x"45800007",  8003 => x"c8021000",
     8004 => x"7c430000",  8005 => x"c8010800",  8006 => x"c8230800",
     8007 => x"5b81003c",  8008 => x"5b820040",  8009 => x"29610020",
     8010 => x"28220008",  8011 => x"3781003c",  8012 => x"1c42003c",
     8013 => x"fbffea18",  8014 => x"45800009",  8015 => x"2b810040",
     8016 => x"2b82003c",  8017 => x"c8010800",  8018 => x"7c230000",
     8019 => x"c8021000",  8020 => x"c8431000",  8021 => x"5b82003c",
     8022 => x"5b810040",  8023 => x"2b830048",  8024 => x"2b820040",
     8025 => x"2b81003c",  8026 => x"2b840044",  8027 => x"b4621000",
     8028 => x"f4621800",  8029 => x"b4810800",  8030 => x"b4610800",
     8031 => x"48200003",  8032 => x"5c200006",  8033 => x"44410005",
     8034 => x"3c210016",  8035 => x"0042000a",  8036 => x"b8221000",
     8037 => x"e0000009",  8038 => x"c8021000",  8039 => x"7c430000",
     8040 => x"c8010800",  8041 => x"c8230800",  8042 => x"3c210016",
     8043 => x"0042000a",  8044 => x"b8221000",  8045 => x"c8021000",
     8046 => x"29610020",  8047 => x"28210008",  8048 => x"28250038",
     8049 => x"20a50001",  8050 => x"5ca00008",  8051 => x"29640028",
     8052 => x"c8021000",  8053 => x"28830010",  8054 => x"5c650002",
     8055 => x"2883000c",  8056 => x"b9600800",  8057 => x"d8600000",
     8058 => x"29610020",  8059 => x"78040001",  8060 => x"34020004",
     8061 => x"28210004",  8062 => x"34030002",  8063 => x"38842ec8",
     8064 => x"2825002c",  8065 => x"b9600800",  8066 => x"14a5000a",
     8067 => x"fbffe59d",  8068 => x"e0000004",  8069 => x"29a60038",
     8070 => x"4c06fedb",  8071 => x"e3fffedc",  8072 => x"2b9d0004",
     8073 => x"2b8b0024",  8074 => x"2b8c0020",  8075 => x"2b8d001c",
     8076 => x"2b8e0018",  8077 => x"2b8f0014",  8078 => x"2b900010",
     8079 => x"2b91000c",  8080 => x"2b920008",  8081 => x"379c0048",
     8082 => x"c3a00000",  8083 => x"379cfffc",  8084 => x"5b9d0004",
     8085 => x"78030001",  8086 => x"3c420002",  8087 => x"38634a3c",
     8088 => x"b4622800",  8089 => x"28a50000",  8090 => x"78040001",
     8091 => x"34020006",  8092 => x"34030001",  8093 => x"38842ee0",
     8094 => x"fbffe582",  8095 => x"2b9d0004",  8096 => x"379c0004",
     8097 => x"c3a00000",  8098 => x"379cfff0",  8099 => x"5b8b0010",
     8100 => x"5b8c000c",  8101 => x"5b8d0008",  8102 => x"5b9d0004",
     8103 => x"b8205800",  8104 => x"78010001",  8105 => x"3821522c",
     8106 => x"b8406800",  8107 => x"28220000",  8108 => x"5c400005",
     8109 => x"29620020",  8110 => x"2844000c",  8111 => x"28820008",
     8112 => x"58220000",  8113 => x"78040001",  8114 => x"78010001",
     8115 => x"3884522c",  8116 => x"38213cec",  8117 => x"28260000",
     8118 => x"28850000",  8119 => x"340c0190",  8120 => x"bd836000",
     8121 => x"88a62800",  8122 => x"b9801000",  8123 => x"34a53039",
     8124 => x"00a10010",  8125 => x"88a62800",  8126 => x"202107ff",
     8127 => x"34a53039",  8128 => x"58850000",  8129 => x"00a50010",
     8130 => x"3c24000a",  8131 => x"20a103ff",  8132 => x"b8240800",
     8133 => x"f8002436",  8134 => x"3d820001",  8135 => x"b4221000",
     8136 => x"29610028",  8137 => x"28230018",  8138 => x"b9600800",
     8139 => x"d8600000",  8140 => x"35a200b2",  8141 => x"3c420002",
     8142 => x"b5625800",  8143 => x"59610004",  8144 => x"2b9d0004",
     8145 => x"2b8b0010",  8146 => x"2b8c000c",  8147 => x"2b8d0008",
     8148 => x"379c0010",  8149 => x"c3a00000",  8150 => x"379cfff0",
     8151 => x"5b8b0010",  8152 => x"5b8c000c",  8153 => x"5b8d0008",
     8154 => x"5b9d0004",  8155 => x"282b000c",  8156 => x"b8206000",
     8157 => x"34010001",  8158 => x"59610000",  8159 => x"29810024",
     8160 => x"48200002",  8161 => x"34010001",  8162 => x"0d61000c",
     8163 => x"29810008",  8164 => x"5c200002",  8165 => x"59820008",
     8166 => x"298d0008",  8167 => x"3561000e",  8168 => x"34030004",
     8169 => x"b9a01000",  8170 => x"f8002462",  8171 => x"2d62000c",
     8172 => x"34010001",  8173 => x"5c410004",  8174 => x"29810000",
     8175 => x"4021001d",  8176 => x"64210002",  8177 => x"59610018",
     8178 => x"41a10044",  8179 => x"2d67000c",  8180 => x"34060002",
     8181 => x"31610012",  8182 => x"41a10045",  8183 => x"34050001",
     8184 => x"3404ffff",  8185 => x"31610013",  8186 => x"41a10046",
     8187 => x"31610014",  8188 => x"34010000",  8189 => x"e000000c",
     8190 => x"08220374",  8191 => x"29880000",  8192 => x"b5021000",
     8193 => x"44600004",  8194 => x"4043001d",  8195 => x"44660002",
     8196 => x"59600018",  8197 => x"58410338",  8198 => x"58450000",
     8199 => x"0c44010e",  8200 => x"34210001",  8201 => x"29630018",
     8202 => x"48e1fff4",  8203 => x"44600006",  8204 => x"78010001",
     8205 => x"38212f70",  8206 => x"f8000b66",  8207 => x"3401ffff",
     8208 => x"3161000e",  8209 => x"78010001",  8210 => x"382149c4",
     8211 => x"28230004",  8212 => x"34010000",  8213 => x"44600004",
     8214 => x"b9800800",  8215 => x"b9a01000",  8216 => x"d8600000",
     8217 => x"2b9d0004",  8218 => x"2b8b0010",  8219 => x"2b8c000c",
     8220 => x"2b8d0008",  8221 => x"379c0010",  8222 => x"c3a00000",
     8223 => x"379cfffc",  8224 => x"5b9d0004",  8225 => x"78020001",
     8226 => x"384249c4",  8227 => x"28430008",  8228 => x"34020000",
     8229 => x"44600003",  8230 => x"d8600000",  8231 => x"b8201000",
     8232 => x"b8400800",  8233 => x"2b9d0004",  8234 => x"379c0004",
     8235 => x"c3a00000",  8236 => x"379cfffc",  8237 => x"5b9d0004",
     8238 => x"b8201000",  8239 => x"78010001",  8240 => x"38212f94",
     8241 => x"f8000b43",  8242 => x"2b9d0004",  8243 => x"379c0004",
     8244 => x"c3a00000",  8245 => x"379cffcc",  8246 => x"5b8b0010",
     8247 => x"5b8c000c",  8248 => x"5b8d0008",  8249 => x"5b9d0004",
     8250 => x"378b0014",  8251 => x"34020000",  8252 => x"34030024",
     8253 => x"b9600800",  8254 => x"f800248c",  8255 => x"78030001",
     8256 => x"b9600800",  8257 => x"34040000",  8258 => x"34020000",
     8259 => x"38635230",  8260 => x"34080020",  8261 => x"34070008",
     8262 => x"e0000004",  8263 => x"34840001",  8264 => x"34210004",
     8265 => x"44870017",  8266 => x"b4432800",  8267 => x"e0000004",
     8268 => x"30a00000",  8269 => x"34420001",  8270 => x"34a50001",
     8271 => x"40a60000",  8272 => x"44c8fffc",  8273 => x"44c0000d",
     8274 => x"b4432800",  8275 => x"58250000",  8276 => x"e0000002",
     8277 => x"34420001",  8278 => x"b4432800",  8279 => x"40a50000",
     8280 => x"7ca90000",  8281 => x"7ca60020",  8282 => x"a1263000",
     8283 => x"5cc0fffa",  8284 => x"5ca6ffeb",  8285 => x"e0000003",
     8286 => x"340c0000",  8287 => x"448c0021",  8288 => x"2b810014",
     8289 => x"340c0000",  8290 => x"40220000",  8291 => x"34010023",
     8292 => x"4441001c",  8293 => x"780b0001",  8294 => x"780c0001",
     8295 => x"396b4dc8",  8296 => x"398c4e68",  8297 => x"e0000011",
     8298 => x"29610000",  8299 => x"f80024a0",  8300 => x"b8206800",
     8301 => x"5c20000c",  8302 => x"29620004",  8303 => x"37810018",
     8304 => x"d8400000",  8305 => x"b8206000",  8306 => x"4c2d000e",
     8307 => x"29620000",  8308 => x"78010001",  8309 => x"b9801800",
     8310 => x"38212f9c",  8311 => x"f8000afd",  8312 => x"e0000008",
     8313 => x"356b0008",  8314 => x"2b820014",  8315 => x"558bffef",
     8316 => x"78010001",  8317 => x"38212fb4",  8318 => x"f8000af6",
     8319 => x"340cffea",  8320 => x"b9800800",  8321 => x"2b9d0004",
     8322 => x"2b8b0010",  8323 => x"2b8c000c",  8324 => x"2b8d0008",
     8325 => x"379c0034",  8326 => x"c3a00000",  8327 => x"379cfff8",
     8328 => x"5b8b0008",  8329 => x"5b9d0004",  8330 => x"780b0001",
     8331 => x"396b5284",  8332 => x"29650000",  8333 => x"78020001",
     8334 => x"34240001",  8335 => x"b8201800",  8336 => x"38425230",
     8337 => x"b4220800",  8338 => x"c8a31800",  8339 => x"b4821000",
     8340 => x"f80023f1",  8341 => x"29610000",  8342 => x"3421ffff",
     8343 => x"59610000",  8344 => x"2b9d0004",  8345 => x"2b8b0008",
     8346 => x"379c0008",  8347 => x"c3a00000",  8348 => x"78010001",
     8349 => x"3821528c",  8350 => x"58200000",  8351 => x"78010001",
     8352 => x"38215284",  8353 => x"58200000",  8354 => x"78010001",
     8355 => x"38215288",  8356 => x"58200000",  8357 => x"c3a00000",
     8358 => x"379cfff4",  8359 => x"5b8b000c",  8360 => x"5b8c0008",
     8361 => x"5b9d0004",  8362 => x"780b0001",  8363 => x"396b5288",
     8364 => x"29610000",  8365 => x"340c0001",  8366 => x"442c000f",
     8367 => x"34020002",  8368 => x"44220099",  8369 => x"5c2000a1",
     8370 => x"78010001",  8371 => x"38212fd0",  8372 => x"f8000ac0",
     8373 => x"78010001",  8374 => x"3821528c",  8375 => x"58200000",
     8376 => x"78010001",  8377 => x"38215284",  8378 => x"58200000",
     8379 => x"596c0000",  8380 => x"e0000096",  8381 => x"f800194a",
     8382 => x"48010094",  8383 => x"3402001b",  8384 => x"44220008",
     8385 => x"78020001",  8386 => x"38425290",  8387 => x"28430000",
     8388 => x"6424005b",  8389 => x"00650010",  8390 => x"a0a42000",
     8391 => x"44800006",  8392 => x"78010001",  8393 => x"38215290",
     8394 => x"78020001",  8395 => x"58220000",  8396 => x"e0000003",
     8397 => x"b8230800",  8398 => x"58410000",  8399 => x"78010001",
     8400 => x"38215290",  8401 => x"282b0000",  8402 => x"216100ff",
     8403 => x"4420007f",  8404 => x"3401007e",  8405 => x"4561002e",
     8406 => x"49610006",  8407 => x"34010009",  8408 => x"4561006d",
     8409 => x"3401000d",  8410 => x"5d610042",  8411 => x"e0000020",
     8412 => x"78020001",  8413 => x"38423cf0",  8414 => x"28410000",
     8415 => x"45610010",  8416 => x"78020001",  8417 => x"38423cf4",
     8418 => x"28410000",  8419 => x"45610004",  8420 => x"3401007f",
     8421 => x"5d610037",  8422 => x"e0000027",  8423 => x"78010001",
     8424 => x"3821528c",  8425 => x"28220000",  8426 => x"4c02005b",
     8427 => x"3442ffff",  8428 => x"58220000",  8429 => x"34010044",
     8430 => x"e000000b",  8431 => x"78010001",  8432 => x"78020001",
     8433 => x"3821528c",  8434 => x"38425284",  8435 => x"28230000",
     8436 => x"28420000",  8437 => x"4c620050",  8438 => x"34630001",
     8439 => x"58230000",  8440 => x"34010043",  8441 => x"fbffff33",
     8442 => x"e000004b",  8443 => x"78010001",  8444 => x"38211b04",
     8445 => x"f8000a77",  8446 => x"78010001",  8447 => x"38215288",
     8448 => x"34020002",  8449 => x"58220000",  8450 => x"e0000043",
     8451 => x"78010001",  8452 => x"78020001",  8453 => x"3821528c",
     8454 => x"38425284",  8455 => x"28210000",  8456 => x"28420000",
     8457 => x"4422003c",  8458 => x"fbffff7d",  8459 => x"34010050",
     8460 => x"e3ffffed",  8461 => x"780b0001",  8462 => x"396b528c",
     8463 => x"29610000",  8464 => x"4c010035",  8465 => x"34010044",
     8466 => x"fbffff1a",  8467 => x"34010050",  8468 => x"fbffff18",
     8469 => x"29610000",  8470 => x"3421ffff",  8471 => x"fbffff70",
     8472 => x"29610000",  8473 => x"3421ffff",  8474 => x"59610000",
     8475 => x"e000002a",  8476 => x"78010001",  8477 => x"a1610800",
     8478 => x"5c200027",  8479 => x"78010001",  8480 => x"38215284",
     8481 => x"28240000",  8482 => x"3401004f",  8483 => x"48810022",
     8484 => x"78010001",  8485 => x"3821528c",  8486 => x"28230000",
     8487 => x"44640008",  8488 => x"78020001",  8489 => x"34610001",
     8490 => x"38425230",  8491 => x"b4220800",  8492 => x"b4621000",
     8493 => x"c8831800",  8494 => x"f8002357",  8495 => x"78010001",
     8496 => x"3821528c",  8497 => x"28230000",  8498 => x"78020001",
     8499 => x"38425230",  8500 => x"b4431000",  8501 => x"304b0000",
     8502 => x"34620001",  8503 => x"58220000",  8504 => x"78010001",
     8505 => x"38215284",  8506 => x"28220000",  8507 => x"34420001",
     8508 => x"58220000",  8509 => x"34010040",  8510 => x"fbfffeee",
     8511 => x"78020001",  8512 => x"38425290",  8513 => x"28420000",
     8514 => x"78010001",  8515 => x"38212fd8",  8516 => x"f8000a30",
     8517 => x"78010001",  8518 => x"38215290",  8519 => x"58200000",
     8520 => x"e000000a",  8521 => x"78020001",  8522 => x"38425284",
     8523 => x"28420000",  8524 => x"78010001",  8525 => x"38215230",
     8526 => x"b4220800",  8527 => x"30200000",  8528 => x"fbfffee5",
     8529 => x"59600000",  8530 => x"2b9d0004",  8531 => x"2b8b000c",
     8532 => x"2b8c0008",  8533 => x"379c000c",  8534 => x"c3a00000",
     8535 => x"34030000",  8536 => x"34070009",  8537 => x"34050005",
     8538 => x"e0000014",  8539 => x"3486ffd0",  8540 => x"20c800ff",
     8541 => x"55070004",  8542 => x"3c630004",  8543 => x"b4c31800",
     8544 => x"e000000d",  8545 => x"3486ffbf",  8546 => x"20c600ff",
     8547 => x"54c50004",  8548 => x"3c630004",  8549 => x"3484ffc9",
     8550 => x"e0000006",  8551 => x"3486ff9f",  8552 => x"20c600ff",
     8553 => x"54c50007",  8554 => x"3c630004",  8555 => x"3484ffa9",
     8556 => x"b4831800",  8557 => x"34210001",  8558 => x"40240000",
     8559 => x"5c80ffec",  8560 => x"58430000",  8561 => x"c3a00000",
     8562 => x"34030000",  8563 => x"34050009",  8564 => x"e0000007",
     8565 => x"3484ffd0",  8566 => x"208600ff",  8567 => x"54c50006",
     8568 => x"0863000a",  8569 => x"34210001",  8570 => x"b4831800",
     8571 => x"40240000",  8572 => x"5c80fff9",  8573 => x"58430000",
     8574 => x"c3a00000",  8575 => x"379cffec",  8576 => x"5b8b0014",
     8577 => x"5b8c0010",  8578 => x"5b8d000c",  8579 => x"5b8e0008",
     8580 => x"5b9d0004",  8581 => x"78010001",  8582 => x"38216a58",
     8583 => x"40210000",  8584 => x"340bffff",  8585 => x"4420001c",
     8586 => x"780b0001",  8587 => x"780e0001",  8588 => x"780d0001",
     8589 => x"340c0000",  8590 => x"396b5230",  8591 => x"39ce5284",
     8592 => x"39ad2ff4",  8593 => x"b9600800",  8594 => x"34020050",
     8595 => x"b9801800",  8596 => x"f800149a",  8597 => x"59c10000",
     8598 => x"48200007",  8599 => x"340b0000",  8600 => x"5d80000d",
     8601 => x"78010001",  8602 => x"38212fdc",  8603 => x"f80009d9",
     8604 => x"e0000009",  8605 => x"b5610800",  8606 => x"3020ffff",
     8607 => x"b9601000",  8608 => x"b9a00800",  8609 => x"f80009d3",
     8610 => x"fbfffe93",  8611 => x"340c0001",  8612 => x"e3ffffed",
     8613 => x"b9600800",  8614 => x"2b9d0004",  8615 => x"2b8b0014",
     8616 => x"2b8c0010",  8617 => x"2b8d000c",  8618 => x"2b8e0008",
     8619 => x"379c0014",  8620 => x"c3a00000",  8621 => x"379cfff8",
     8622 => x"5b8b0008",  8623 => x"5b9d0004",  8624 => x"78010001",
     8625 => x"38216db8",  8626 => x"28210000",  8627 => x"78030001",
     8628 => x"386343c0",  8629 => x"28620000",  8630 => x"282b000c",
     8631 => x"78030001",  8632 => x"78010001",  8633 => x"3863301c",
     8634 => x"38213004",  8635 => x"f80009b9",  8636 => x"78040001",
     8637 => x"78030001",  8638 => x"388443c4",  8639 => x"386343c8",
     8640 => x"28820000",  8641 => x"28630000",  8642 => x"78010001",
     8643 => x"3821303c",  8644 => x"f80009b0",  8645 => x"216b000f",
     8646 => x"356b0001",  8647 => x"78010001",  8648 => x"34020080",
     8649 => x"3d6b0004",  8650 => x"3821304c",  8651 => x"34030800",
     8652 => x"f80009a8",  8653 => x"3561ff80",  8654 => x"3402000f",
     8655 => x"50410006",  8656 => x"78010001",  8657 => x"38213074",
     8658 => x"b9601000",  8659 => x"35630010",  8660 => x"f80009a0",
     8661 => x"34010000",  8662 => x"2b9d0004",  8663 => x"2b8b0008",
     8664 => x"379c0008",  8665 => x"c3a00000",  8666 => x"379cffe8",
     8667 => x"5b8b0010",  8668 => x"5b8c000c",  8669 => x"5b8d0008",
     8670 => x"5b9d0004",  8671 => x"b8205800",  8672 => x"28210000",
     8673 => x"78020001",  8674 => x"384230a4",  8675 => x"f8002328",
     8676 => x"5c200011",  8677 => x"2963000c",  8678 => x"3402ffea",
     8679 => x"44610086",  8680 => x"29610004",  8681 => x"f80004b9",
     8682 => x"b8206800",  8683 => x"29610008",  8684 => x"f80004b6",
     8685 => x"b8206000",  8686 => x"2961000c",  8687 => x"f80004b3",
     8688 => x"b8201800",  8689 => x"b9801000",  8690 => x"b9a00800",
     8691 => x"f8001d6a",  8692 => x"e0000078",  8693 => x"29610000",
     8694 => x"78020001",  8695 => x"384230ac",  8696 => x"f8002313",
     8697 => x"b8201800",  8698 => x"5c200007",  8699 => x"29610004",
     8700 => x"3402ffea",  8701 => x"44230070",  8702 => x"f80004a4",
     8703 => x"f8001e43",  8704 => x"e0000060",  8705 => x"29610000",
     8706 => x"78020001",  8707 => x"384230b0",  8708 => x"f8002307",
     8709 => x"5c200003",  8710 => x"f8001ed5",  8711 => x"e0000065",
     8712 => x"29610000",  8713 => x"78020001",  8714 => x"384230b8",
     8715 => x"f8002300",  8716 => x"5c20000d",  8717 => x"29630008",
     8718 => x"3402ffea",  8719 => x"4461005e",  8720 => x"29610004",
     8721 => x"f8000491",  8722 => x"b8206000",  8723 => x"29610008",
     8724 => x"f800048e",  8725 => x"b8201000",  8726 => x"b9800800",
     8727 => x"f8001e3c",  8728 => x"e0000054",  8729 => x"29610000",
     8730 => x"78020001",  8731 => x"384230bc",  8732 => x"f80022ef",
     8733 => x"b8201800",  8734 => x"5c20000e",  8735 => x"29610004",
     8736 => x"3402ffea",  8737 => x"4423004c",  8738 => x"f8000480",
     8739 => x"37820018",  8740 => x"37830014",  8741 => x"f8001e56",
     8742 => x"2b820018",  8743 => x"2b830014",  8744 => x"78010001",
     8745 => x"382130c0",  8746 => x"f800094a",  8747 => x"e0000041",
     8748 => x"29610000",  8749 => x"78020001",  8750 => x"384230c8",
     8751 => x"f80022dc",  8752 => x"b8201800",  8753 => x"5c200007",
     8754 => x"29610004",  8755 => x"3402ffea",  8756 => x"44230039",
     8757 => x"f800046d",  8758 => x"f8001de8",  8759 => x"e0000035",
     8760 => x"29610000",  8761 => x"78020001",  8762 => x"384230d0",
     8763 => x"f80022d0",  8764 => x"b8201800",  8765 => x"5c200007",
     8766 => x"29610004",  8767 => x"3402ffea",  8768 => x"4423002d",
     8769 => x"f8000461",  8770 => x"f8001df3",  8771 => x"e0000029",
     8772 => x"29610000",  8773 => x"78020001",  8774 => x"384230d8",
     8775 => x"f80022c4",  8776 => x"5c20000d",  8777 => x"29630008",
     8778 => x"3402ffea",  8779 => x"44610022",  8780 => x"29610004",
     8781 => x"f8000455",  8782 => x"b8206000",  8783 => x"29610008",
     8784 => x"f8000452",  8785 => x"b8201000",  8786 => x"b9800800",
     8787 => x"f8001f02",  8788 => x"e0000018",  8789 => x"29610000",
     8790 => x"78020001",  8791 => x"384230e0",  8792 => x"f80022b3",
     8793 => x"b8201800",  8794 => x"5c20000b",  8795 => x"29610004",
     8796 => x"3402ffea",  8797 => x"44230010",  8798 => x"f8000444",
     8799 => x"f8001ee7",  8800 => x"b8201000",  8801 => x"78010001",
     8802 => x"382138c0",  8803 => x"f8000911",  8804 => x"e0000008",
     8805 => x"29610000",  8806 => x"78020001",  8807 => x"384230e8",
     8808 => x"f80022a3",  8809 => x"3402ffea",  8810 => x"5c200003",
     8811 => x"f8001f9d",  8812 => x"34020000",  8813 => x"b8400800",
     8814 => x"2b9d0004",  8815 => x"2b8b0010",  8816 => x"2b8c000c",
     8817 => x"2b8d0008",  8818 => x"379c0018",  8819 => x"c3a00000",
     8820 => x"379cffb4",  8821 => x"5b8b002c",  8822 => x"5b8c0028",
     8823 => x"5b8d0024",  8824 => x"5b8e0020",  8825 => x"5b8f001c",
     8826 => x"5b900018",  8827 => x"5b910014",  8828 => x"5b920010",
     8829 => x"5b93000c",  8830 => x"5b940008",  8831 => x"5b9d0004",
     8832 => x"b8205800",  8833 => x"28210000",  8834 => x"44200015",
     8835 => x"78020001",  8836 => x"384230f8",  8837 => x"f8002286",
     8838 => x"b8206000",  8839 => x"5c200010",  8840 => x"f8000f2c",
     8841 => x"5c2c0005",  8842 => x"78010001",  8843 => x"38213100",
     8844 => x"f80008e8",  8845 => x"e0000004",  8846 => x"78010001",
     8847 => x"38214aa8",  8848 => x"f8000f2b",  8849 => x"78020001",
     8850 => x"38424aa8",  8851 => x"78010001",  8852 => x"30400010",
     8853 => x"38212e58",  8854 => x"e000004d",  8855 => x"29610000",
     8856 => x"78020001",  8857 => x"3842310c",  8858 => x"f8002271",
     8859 => x"5c200009",  8860 => x"f80011c7",  8861 => x"3402ffff",
     8862 => x"340c0000",  8863 => x"5c2200b3",  8864 => x"78010001",
     8865 => x"38213114",  8866 => x"f80008d2",  8867 => x"e00000af",
     8868 => x"29610010",  8869 => x"44200040",  8870 => x"29610000",
     8871 => x"78020001",  8872 => x"38423128",  8873 => x"f8002262",
     8874 => x"5c20003b",  8875 => x"29610004",  8876 => x"356c0004",
     8877 => x"f80022a3",  8878 => x"34020010",  8879 => x"54220005",
     8880 => x"29610004",  8881 => x"f800229f",  8882 => x"3c220018",
     8883 => x"14420018",  8884 => x"34030000",  8885 => x"37840030",
     8886 => x"e0000007",  8887 => x"29810000",  8888 => x"b4832800",
     8889 => x"b4230800",  8890 => x"40210000",  8891 => x"34630001",
     8892 => x"30a10000",  8893 => x"b0600800",  8894 => x"4841fff9",
     8895 => x"b4811000",  8896 => x"34030020",  8897 => x"3404000f",
     8898 => x"e0000005",  8899 => x"34210001",  8900 => x"30430000",
     8901 => x"b0200800",  8902 => x"34420001",  8903 => x"4c81fffc",
     8904 => x"29610008",  8905 => x"f80003d9",  8906 => x"5b810044",
     8907 => x"2961000c",  8908 => x"f80003d6",  8909 => x"5b810048",
     8910 => x"29610010",  8911 => x"f80003d3",  8912 => x"5b810040",
     8913 => x"34020001",  8914 => x"37810030",  8915 => x"34030000",
     8916 => x"f80011a4",  8917 => x"3c220018",  8918 => x"3401fffe",
     8919 => x"14420018",  8920 => x"5c410004",  8921 => x"78010001",
     8922 => x"3821312c",  8923 => x"e0000067",  8924 => x"3401ffff",
     8925 => x"5c410004",  8926 => x"78010001",  8927 => x"3821313c",
     8928 => x"e0000062",  8929 => x"78010001",  8930 => x"38213148",
     8931 => x"f8000891",  8932 => x"e000006d",  8933 => x"29610000",
     8934 => x"44200033",  8935 => x"78020001",  8936 => x"38423158",
     8937 => x"f8002222",  8938 => x"5c20002f",  8939 => x"78100001",
     8940 => x"780f0001",  8941 => x"780e0001",  8942 => x"340c0000",
     8943 => x"340b0000",  8944 => x"34120001",  8945 => x"37910030",
     8946 => x"3414ffff",  8947 => x"3a103194",  8948 => x"37930040",
     8949 => x"39ef2fd8",  8950 => x"39ce319c",  8951 => x"ba200800",
     8952 => x"34020000",  8953 => x"b9801800",  8954 => x"f800117e",
     8955 => x"5d60000b",  8956 => x"b0201000",  8957 => x"5c4b0004",
     8958 => x"78010001",  8959 => x"38213160",  8960 => x"e0000042",
     8961 => x"5c540004",  8962 => x"78010001",  8963 => x"38213178",
     8964 => x"e000003e",  8965 => x"b8409000",  8966 => x"358c0001",
     8967 => x"ba000800",  8968 => x"b9801000",  8969 => x"f800086b",
     8970 => x"ba206800",  8971 => x"41a20000",  8972 => x"b9e00800",
     8973 => x"35ad0001",  8974 => x"f8000866",  8975 => x"5db3fffc",
     8976 => x"2b820044",  8977 => x"2b830048",  8978 => x"2b840040",
     8979 => x"356b0001",  8980 => x"b9c00800",  8981 => x"b1605800",
     8982 => x"f800085e",  8983 => x"4a4bffe0",  8984 => x"e0000039",
     8985 => x"29610000",  8986 => x"4420002a",  8987 => x"78020001",
     8988 => x"384231bc",  8989 => x"f80021ee",  8990 => x"5c200026",
     8991 => x"78020001",  8992 => x"38424aa8",  8993 => x"40430000",
     8994 => x"5c610004",  8995 => x"78010001",  8996 => x"382131c4",
     8997 => x"e000001d",  8998 => x"378b0030",  8999 => x"b9600800",
     9000 => x"34030010",  9001 => x"f80022a3",  9002 => x"b9600800",
     9003 => x"f80011bd",  9004 => x"4c010014",  9005 => x"2b820044",
     9006 => x"2b830048",  9007 => x"2b840040",  9008 => x"78010001",
     9009 => x"382131dc",  9010 => x"f8000842",  9011 => x"2b820044",
     9012 => x"78010001",  9013 => x"38214e6c",  9014 => x"58220000",
     9015 => x"2b820048",  9016 => x"78010001",  9017 => x"38214e70",
     9018 => x"58220000",  9019 => x"2b820040",  9020 => x"78010001",
     9021 => x"382143d4",  9022 => x"58220000",  9023 => x"e0000012",
     9024 => x"78010001",  9025 => x"38213204",  9026 => x"f8000832",
     9027 => x"e000000e",  9028 => x"29610000",  9029 => x"340c0000",
     9030 => x"4420000c",  9031 => x"78020001",  9032 => x"3842321c",
     9033 => x"f80021c2",  9034 => x"b8201000",  9035 => x"5c200007",
     9036 => x"29610004",  9037 => x"340cffea",  9038 => x"44220004",
     9039 => x"f8000353",  9040 => x"f80009e2",  9041 => x"340c0000",
     9042 => x"b9800800",  9043 => x"2b9d0004",  9044 => x"2b8b002c",
     9045 => x"2b8c0028",  9046 => x"2b8d0024",  9047 => x"2b8e0020",
     9048 => x"2b8f001c",  9049 => x"2b900018",  9050 => x"2b910014",
     9051 => x"2b920010",  9052 => x"2b93000c",  9053 => x"2b940008",
     9054 => x"379c004c",  9055 => x"c3a00000",  9056 => x"379cfff8",
     9057 => x"5b8b0008",  9058 => x"5b9d0004",  9059 => x"b8205800",
     9060 => x"28210000",  9061 => x"5c200011",  9062 => x"78010001",
     9063 => x"38216dac",  9064 => x"28220000",  9065 => x"340b0000",
     9066 => x"64420000",  9067 => x"58220000",  9068 => x"78010001",
     9069 => x"38216d04",  9070 => x"28230000",  9071 => x"3463ffff",
     9072 => x"58230000",  9073 => x"5c4b002b",  9074 => x"78010001",
     9075 => x"38213224",  9076 => x"f8000800",  9077 => x"e0000027",
     9078 => x"78020001",  9079 => x"38423238",  9080 => x"f8002193",
     9081 => x"5c200007",  9082 => x"f800096b",  9083 => x"b8201000",
     9084 => x"78010001",  9085 => x"38213704",  9086 => x"f80007f6",
     9087 => x"e000001c",  9088 => x"29610000",  9089 => x"78020001",
     9090 => x"3842250c",  9091 => x"f8002188",  9092 => x"5c20000b",
     9093 => x"78010001",  9094 => x"38216dac",  9095 => x"34020001",
     9096 => x"58220000",  9097 => x"78010001",  9098 => x"38216d04",
     9099 => x"28220000",  9100 => x"3442ffff",  9101 => x"58220000",
     9102 => x"e000000d",  9103 => x"29610000",  9104 => x"78020001",
     9105 => x"3842323c",  9106 => x"f8002179",  9107 => x"340bffea",
     9108 => x"5c200008",  9109 => x"78010001",  9110 => x"38216dac",
     9111 => x"58200000",  9112 => x"78010001",  9113 => x"38213224",
     9114 => x"f80007da",  9115 => x"340b0000",  9116 => x"b9600800",
     9117 => x"2b9d0004",  9118 => x"2b8b0008",  9119 => x"379c0008",
     9120 => x"c3a00000",  9121 => x"379cfff8",  9122 => x"5b8b0008",
     9123 => x"5b9d0004",  9124 => x"b8205800",  9125 => x"28210000",
     9126 => x"78020001",  9127 => x"384230c8",  9128 => x"f8002163",
     9129 => x"5c200003",  9130 => x"fbffe2a3",  9131 => x"e0000008",
     9132 => x"29610000",  9133 => x"78020001",  9134 => x"384230d0",
     9135 => x"f800215c",  9136 => x"3402ffea",  9137 => x"5c200003",
     9138 => x"fbffe2bd",  9139 => x"b8201000",  9140 => x"b8400800",
     9141 => x"2b9d0004",  9142 => x"2b8b0008",  9143 => x"379c0008",
     9144 => x"c3a00000",  9145 => x"379cfff8",  9146 => x"5b8b0008",
     9147 => x"5b9d0004",  9148 => x"b8205800",  9149 => x"28210000",
     9150 => x"78020001",  9151 => x"38423244",  9152 => x"f800214b",
     9153 => x"34020001",  9154 => x"44200018",  9155 => x"29610000",
     9156 => x"78020001",  9157 => x"38422954",  9158 => x"f8002145",
     9159 => x"34020002",  9160 => x"44200012",  9161 => x"29610000",
     9162 => x"78020001",  9163 => x"3842246c",  9164 => x"f800213f",
     9165 => x"34020003",  9166 => x"4420000c",  9167 => x"fbffe27a",
     9168 => x"3c210002",  9169 => x"78020001",  9170 => x"38423fd0",
     9171 => x"b4411000",  9172 => x"28420000",  9173 => x"78010001",
     9174 => x"38212e58",  9175 => x"f800079d",  9176 => x"34010000",
     9177 => x"e0000003",  9178 => x"b8400800",  9179 => x"fbffe2b6",
     9180 => x"2b9d0004",  9181 => x"2b8b0008",  9182 => x"379c0008",
     9183 => x"c3a00000",  9184 => x"379cfff0",  9185 => x"5b8b000c",
     9186 => x"5b8c0008",  9187 => x"5b9d0004",  9188 => x"b8205800",
     9189 => x"28210000",  9190 => x"4420000b",  9191 => x"78020001",
     9192 => x"3842325c",  9193 => x"f8002122",  9194 => x"b8206000",
     9195 => x"5c200006",  9196 => x"37810010",  9197 => x"f8000f35",
     9198 => x"340bffff",  9199 => x"49810021",  9200 => x"e000001c",
     9201 => x"29610000",  9202 => x"340b0000",  9203 => x"5c20001d",
     9204 => x"37810010",  9205 => x"34020000",  9206 => x"f8001133",
     9207 => x"4d61000a",  9208 => x"2b820010",  9209 => x"78010001",
     9210 => x"38213264",  9211 => x"f8000779",  9212 => x"2b820010",
     9213 => x"78010001",  9214 => x"382143d8",  9215 => x"58220000",
     9216 => x"e0000010",  9217 => x"78010001",  9218 => x"3821328c",
     9219 => x"f8000771",  9220 => x"37810010",  9221 => x"f8000f1d",
     9222 => x"340bffff",  9223 => x"48010009",  9224 => x"2b820010",
     9225 => x"78010001",  9226 => x"382143d8",  9227 => x"58220000",
     9228 => x"37810010",  9229 => x"34020001",  9230 => x"f800111b",
     9231 => x"b8205800",  9232 => x"b9600800",  9233 => x"2b9d0004",
     9234 => x"2b8b000c",  9235 => x"2b8c0008",  9236 => x"379c0010",
     9237 => x"c3a00000",  9238 => x"379cffe8",  9239 => x"5b8b000c",
     9240 => x"5b8c0008",  9241 => x"5b9d0004",  9242 => x"b8205800",
     9243 => x"37820018",  9244 => x"37810010",  9245 => x"f8000d3b",
     9246 => x"29610008",  9247 => x"44200014",  9248 => x"29610000",
     9249 => x"78020001",  9250 => x"384232c0",  9251 => x"f80020e8",
     9252 => x"5c20000f",  9253 => x"fbffe224",  9254 => x"34030003",
     9255 => x"3402fff0",  9256 => x"4423003f",  9257 => x"29610004",
     9258 => x"f8000278",  9259 => x"b8206000",  9260 => x"29610008",
     9261 => x"f8000275",  9262 => x"b8201800",  9263 => x"b9801000",
     9264 => x"1581001f",  9265 => x"34040003",  9266 => x"e0000020",
     9267 => x"29610000",  9268 => x"4420000f",  9269 => x"78020001",
     9270 => x"384232c4",  9271 => x"f80020d4",  9272 => x"5c20000b",
     9273 => x"fbffe210",  9274 => x"34020003",  9275 => x"44220023",
     9276 => x"29610004",  9277 => x"f8000265",  9278 => x"b8201000",
     9279 => x"34030000",  9280 => x"1421001f",  9281 => x"34040001",
     9282 => x"e0000010",  9283 => x"29610000",  9284 => x"44200010",
     9285 => x"78020001",  9286 => x"384232cc",  9287 => x"f80020c4",
     9288 => x"5c20000c",  9289 => x"fbffe200",  9290 => x"34020003",
     9291 => x"44220013",  9292 => x"29610004",  9293 => x"f8000255",
     9294 => x"b8201800",  9295 => x"34020000",  9296 => x"34010000",
     9297 => x"34040002",  9298 => x"f8000ce6",  9299 => x"e0000013",
     9300 => x"29610000",  9301 => x"44200009",  9302 => x"78020001",
     9303 => x"384232d4",  9304 => x"f80020b3",  9305 => x"5c200005",
     9306 => x"78010001",  9307 => x"382130c0",  9308 => x"2b820014",
     9309 => x"e0000007",  9310 => x"2b820014",  9311 => x"2b810010",
     9312 => x"f8000169",  9313 => x"b8201000",  9314 => x"78010001",
     9315 => x"382132d8",  9316 => x"2b830018",  9317 => x"f800070f",
     9318 => x"34020000",  9319 => x"b8400800",  9320 => x"2b9d0004",
     9321 => x"2b8b000c",  9322 => x"2b8c0008",  9323 => x"379c0018",
     9324 => x"c3a00000",  9325 => x"78010001",  9326 => x"38214e68",
     9327 => x"34020001",  9328 => x"58220000",  9329 => x"34010000",
     9330 => x"c3a00000",  9331 => x"379cfffc",  9332 => x"5b9d0004",
     9333 => x"f8000d8c",  9334 => x"34010000",  9335 => x"2b9d0004",
     9336 => x"379c0004",  9337 => x"c3a00000",  9338 => x"379cffec",
     9339 => x"5b8b0010",  9340 => x"5b8c000c",  9341 => x"5b8d0008",
     9342 => x"5b9d0004",  9343 => x"340b0000",  9344 => x"b8406800",
     9345 => x"340c0006",  9346 => x"37820014",  9347 => x"fbfffcd4",
     9348 => x"2b830014",  9349 => x"b5ab1000",  9350 => x"356b0001",
     9351 => x"30430000",  9352 => x"40220000",  9353 => x"6442003a",
     9354 => x"b4220800",  9355 => x"5d6cfff7",  9356 => x"2b9d0004",
     9357 => x"2b8b0010",  9358 => x"2b8c000c",  9359 => x"2b8d0008",
     9360 => x"379c0014",  9361 => x"c3a00000",  9362 => x"379cfff0",
     9363 => x"5b8b0008",  9364 => x"5b9d0004",  9365 => x"b8205800",
     9366 => x"28210000",  9367 => x"44200005",  9368 => x"78020001",
     9369 => x"38423300",  9370 => x"f8002071",  9371 => x"5c200004",
     9372 => x"3781000c",  9373 => x"f80007df",  9374 => x"e000002b",
     9375 => x"29610000",  9376 => x"78020001",  9377 => x"38423304",
     9378 => x"f8002069",  9379 => x"5c200008",  9380 => x"378b000c",
     9381 => x"b9600800",  9382 => x"f80007d6",  9383 => x"b9601000",
     9384 => x"34010000",  9385 => x"f80011e0",  9386 => x"e000001f",
     9387 => x"29610000",  9388 => x"78020001",  9389 => x"384232c0",
     9390 => x"f800205d",  9391 => x"5c20000b",  9392 => x"29630004",
     9393 => x"44610009",  9394 => x"378b000c",  9395 => x"b8600800",
     9396 => x"b9601000",  9397 => x"fbffffc5",  9398 => x"b9600800",
     9399 => x"f80007b1",  9400 => x"f80008ac",  9401 => x"e0000010",
     9402 => x"29610000",  9403 => x"78020001",  9404 => x"3842330c",
     9405 => x"f800204e",  9406 => x"b8201800",  9407 => x"3402ffea",
     9408 => x"5c200013",  9409 => x"29610004",  9410 => x"44230011",
     9411 => x"378b000c",  9412 => x"b9601000",  9413 => x"fbffffb5",
     9414 => x"34010000",  9415 => x"b9601000",  9416 => x"f80011b8",
     9417 => x"4382000c",  9418 => x"4383000d",  9419 => x"4384000e",
     9420 => x"4385000f",  9421 => x"43860010",  9422 => x"43870011",
     9423 => x"78010001",  9424 => x"38213314",  9425 => x"f80006a3",
     9426 => x"34020000",  9427 => x"b8400800",  9428 => x"2b9d0004",
     9429 => x"2b8b0008",  9430 => x"379c0010",  9431 => x"c3a00000",
     9432 => x"379cfff4",  9433 => x"5b8b000c",  9434 => x"5b8c0008",
     9435 => x"5b9d0004",  9436 => x"34020050",  9437 => x"b8205800",
     9438 => x"34010000",  9439 => x"f80009f5",  9440 => x"5c200006",
     9441 => x"78010001",  9442 => x"38213344",  9443 => x"f8000691",
     9444 => x"340bffff",  9445 => x"e0000031",  9446 => x"29610000",
     9447 => x"4420000c",  9448 => x"78020001",  9449 => x"3842310c",
     9450 => x"f8002021",  9451 => x"5c200008",  9452 => x"f8001072",
     9453 => x"340b0000",  9454 => x"4c2b0028",  9455 => x"78010001",
     9456 => x"38213358",  9457 => x"f8000683",  9458 => x"e0000024",
     9459 => x"29610004",  9460 => x"44200012",  9461 => x"29610000",
     9462 => x"78020001",  9463 => x"38423128",  9464 => x"f8002013",
     9465 => x"b8206000",  9466 => x"5c20000c",  9467 => x"b9600800",
     9468 => x"f8001077",  9469 => x"4c2c0004",  9470 => x"78010001",
     9471 => x"38213378",  9472 => x"e0000003",  9473 => x"78010001",
     9474 => x"38213394",  9475 => x"f8000671",  9476 => x"340b0000",
     9477 => x"e0000011",  9478 => x"29610000",  9479 => x"44200007",
     9480 => x"78020001",  9481 => x"38423158",  9482 => x"f8002001",
     9483 => x"5c200003",  9484 => x"f80010e1",  9485 => x"e3fffff7",
     9486 => x"29610000",  9487 => x"340b0000",  9488 => x"44200006",
     9489 => x"78020001",  9490 => x"3842339c",  9491 => x"f8001ff8",
     9492 => x"5c200002",  9493 => x"fbfffc6a",  9494 => x"b9600800",
     9495 => x"2b9d0004",  9496 => x"2b8b000c",  9497 => x"2b8c0008",
     9498 => x"379c000c",  9499 => x"c3a00000",  9500 => x"379cfff8",
     9501 => x"5b8b0008",  9502 => x"5b9d0004",  9503 => x"b8205800",
     9504 => x"28210000",  9505 => x"4420000c",  9506 => x"78020001",
     9507 => x"384233ac",  9508 => x"f8001fe7",  9509 => x"5c200008",
     9510 => x"34010001",  9511 => x"fbffec22",  9512 => x"78010001",
     9513 => x"382143d0",  9514 => x"34020001",  9515 => x"58220000",
     9516 => x"e000000b",  9517 => x"29610000",  9518 => x"44200009",
     9519 => x"78020001",  9520 => x"384233b4",  9521 => x"f8001fda",
     9522 => x"5c200005",  9523 => x"fbffec16",  9524 => x"78010001",
     9525 => x"382143d0",  9526 => x"58200000",  9527 => x"78010001",
     9528 => x"382143d0",  9529 => x"28210000",  9530 => x"78020001",
     9531 => x"384233a8",  9532 => x"44200003",  9533 => x"78020001",
     9534 => x"384233a4",  9535 => x"78010001",  9536 => x"382133bc",
     9537 => x"f8000633",  9538 => x"34010000",  9539 => x"2b9d0004",
     9540 => x"2b8b0008",  9541 => x"379c0008",  9542 => x"c3a00000",
     9543 => x"379cfff0",  9544 => x"5b8b0010",  9545 => x"5b8c000c",
     9546 => x"5b8d0008",  9547 => x"5b9d0004",  9548 => x"78010001",
     9549 => x"382133d8",  9550 => x"780b0001",  9551 => x"780d0001",
     9552 => x"780c0001",  9553 => x"f8000623",  9554 => x"396b4dc8",
     9555 => x"39ad4e68",  9556 => x"398c33f0",  9557 => x"e0000005",
     9558 => x"29620000",  9559 => x"b9800800",  9560 => x"356b0008",
     9561 => x"f800061b",  9562 => x"55abfffc",  9563 => x"34010000",
     9564 => x"2b9d0004",  9565 => x"2b8b0010",  9566 => x"2b8c000c",
     9567 => x"2b8d0008",  9568 => x"379c0010",  9569 => x"c3a00000",
     9570 => x"379cfff8",  9571 => x"5b9d0004",  9572 => x"b8201000",
     9573 => x"28210000",  9574 => x"4420000d",  9575 => x"28420004",
     9576 => x"5c40000b",  9577 => x"37820008",  9578 => x"fbfffc08",
     9579 => x"2b820008",  9580 => x"78010001",  9581 => x"382143cc",
     9582 => x"084203e8",  9583 => x"58220000",  9584 => x"78010001",
     9585 => x"38211b04",  9586 => x"e0000003",  9587 => x"78010001",
     9588 => x"38213400",  9589 => x"f80005ff",  9590 => x"34010000",
     9591 => x"2b9d0004",  9592 => x"379c0008",  9593 => x"c3a00000",
     9594 => x"379cffe8",  9595 => x"5b8b0010",  9596 => x"5b8c000c",
     9597 => x"5b9b0008",  9598 => x"5b9d0004",  9599 => x"b820d800",
     9600 => x"28210000",  9601 => x"44200005",  9602 => x"78020001",
     9603 => x"38423300",  9604 => x"f8001f87",  9605 => x"5c200004",
     9606 => x"37810018",  9607 => x"f80004ca",  9608 => x"e0000018",
     9609 => x"2b610000",  9610 => x"78020001",  9611 => x"384232c0",
     9612 => x"f8001f7f",  9613 => x"b8201800",  9614 => x"3402ffea",
     9615 => x"5c200021",  9616 => x"2b610004",  9617 => x"4423001f",
     9618 => x"379b0018",  9619 => x"378c001c",  9620 => x"378b0014",
     9621 => x"b9601000",  9622 => x"fbfffbdc",  9623 => x"2b820014",
     9624 => x"33620000",  9625 => x"40220000",  9626 => x"377b0001",
     9627 => x"6442002e",  9628 => x"b4220800",  9629 => x"5f6cfff8",
     9630 => x"37810018",  9631 => x"f80004bb",  9632 => x"78010001",
     9633 => x"38215d6c",  9634 => x"28210000",  9635 => x"44200005",
     9636 => x"78010001",  9637 => x"38213424",  9638 => x"f80005ce",
     9639 => x"e0000008",  9640 => x"43820018",  9641 => x"43830019",
     9642 => x"4384001a",  9643 => x"4385001b",  9644 => x"78010001",
     9645 => x"38213440",  9646 => x"f80005c6",  9647 => x"34020000",
     9648 => x"b8400800",  9649 => x"2b9d0004",  9650 => x"2b8b0010",
     9651 => x"2b8c000c",  9652 => x"2b9b0008",  9653 => x"379c0018",
     9654 => x"c3a00000",  9655 => x"379cfffc",  9656 => x"5b9d0004",
     9657 => x"28210000",  9658 => x"44200005",  9659 => x"fbffdf97",
     9660 => x"78020001",  9661 => x"38424e9c",  9662 => x"58410000",
     9663 => x"78020001",  9664 => x"38424e9c",  9665 => x"28420000",
     9666 => x"78010001",  9667 => x"38213460",  9668 => x"f80005b0",
     9669 => x"34010000",  9670 => x"2b9d0004",  9671 => x"379c0004",
     9672 => x"c3a00000",  9673 => x"379cffd8",  9674 => x"5b8b0028",
     9675 => x"5b8c0024",  9676 => x"5b8d0020",  9677 => x"5b8e001c",
     9678 => x"5b8f0018",  9679 => x"5b900014",  9680 => x"5b910010",
     9681 => x"5b92000c",  9682 => x"5b9d0008",  9683 => x"78030001",
     9684 => x"38633cf8",  9685 => x"b8406000",  9686 => x"b8400800",
     9687 => x"28620000",  9688 => x"f8001e23",  9689 => x"78030001",
     9690 => x"38633cf8",  9691 => x"28620000",  9692 => x"b8205800",
     9693 => x"b9800800",  9694 => x"f8001e0d",  9695 => x"b8206000",
     9696 => x"3402003c",  9697 => x"b9600800",  9698 => x"f8001e19",
     9699 => x"34020e10",  9700 => x"b8208800",  9701 => x"b9600800",
     9702 => x"f8001e15",  9703 => x"3402003c",  9704 => x"f8001e03",
     9705 => x"34020e10",  9706 => x"b8207800",  9707 => x"b9600800",
     9708 => x"f8001dff",  9709 => x"b8208000",  9710 => x"34020007",
     9711 => x"35810004",  9712 => x"f8001e0b",  9713 => x"b8209000",
     9714 => x"340b07b2",  9715 => x"e000000f",  9716 => x"3402016d",
     9717 => x"5da0000b",  9718 => x"34020064",  9719 => x"b9600800",
     9720 => x"f8001dd3",  9721 => x"3402016e",  9722 => x"5c2d0006",
     9723 => x"34020190",  9724 => x"b9600800",  9725 => x"f8001dce",
     9726 => x"64220000",  9727 => x"3442016d",  9728 => x"c9826000",
     9729 => x"356b0001",  9730 => x"216d0003",  9731 => x"3402016d",
     9732 => x"5da0000b",  9733 => x"34020064",  9734 => x"b9600800",
     9735 => x"f8001dc4",  9736 => x"3402016e",  9737 => x"5c2d0006",
     9738 => x"34020190",  9739 => x"b9600800",  9740 => x"f8001dbf",
     9741 => x"64220000",  9742 => x"3442016d",  9743 => x"5182ffe5",
     9744 => x"34020064",  9745 => x"b9600800",  9746 => x"f8001db9",
     9747 => x"34020190",  9748 => x"b8207000",  9749 => x"b9600800",
     9750 => x"f8001db5",  9751 => x"78030001",  9752 => x"34020000",
     9753 => x"64250000",  9754 => x"38633fe0",  9755 => x"e000000d",
     9756 => x"34040000",  9757 => x"5da00004",  9758 => x"34040001",
     9759 => x"5dcd0002",  9760 => x"b8a02000",  9761 => x"0884000c",
     9762 => x"b4822000",  9763 => x"3c840002",  9764 => x"34420001",
     9765 => x"b4642000",  9766 => x"28810000",  9767 => x"c9816000",
     9768 => x"34040000",  9769 => x"5da00004",  9770 => x"34040001",
     9771 => x"5dcd0002",  9772 => x"b8a02000",  9773 => x"0884000c",
     9774 => x"b4822000",  9775 => x"3c840002",  9776 => x"b4642000",
     9777 => x"28810000",  9778 => x"5181ffea",  9779 => x"3e450002",
     9780 => x"78030001",  9781 => x"38634040",  9782 => x"b4652800",
     9783 => x"3c420002",  9784 => x"78030001",  9785 => x"3863405c",
     9786 => x"b4622000",  9787 => x"28840000",  9788 => x"28a30000",
     9789 => x"780d0001",  9790 => x"39ad5294",  9791 => x"78020001",
     9792 => x"b9a00800",  9793 => x"38423480",  9794 => x"35850001",
     9795 => x"b9603000",  9796 => x"ba003800",  9797 => x"b9e04000",
     9798 => x"5b910004",  9799 => x"f800051f",  9800 => x"b9a00800",
     9801 => x"2b9d0008",  9802 => x"2b8b0028",  9803 => x"2b8c0024",
     9804 => x"2b8d0020",  9805 => x"2b8e001c",  9806 => x"2b8f0018",
     9807 => x"2b900014",  9808 => x"2b910010",  9809 => x"2b92000c",
     9810 => x"379c0028",  9811 => x"c3a00000",  9812 => x"379cffdc",
     9813 => x"5b8b0008",  9814 => x"5b9d0004",  9815 => x"5b840014",
     9816 => x"20240080",  9817 => x"64840000",  9818 => x"5b830010",
     9819 => x"78030001",  9820 => x"b8204800",  9821 => x"b8600800",
     9822 => x"34030002",  9823 => x"5b82000c",  9824 => x"b8405800",
     9825 => x"382134a0",  9826 => x"c8641000",  9827 => x"2123007f",
     9828 => x"5b850018",  9829 => x"5b86001c",  9830 => x"5b870020",
     9831 => x"5b880024",  9832 => x"f800050c",  9833 => x"37820010",
     9834 => x"b9600800",  9835 => x"f80004e7",  9836 => x"78010001",
     9837 => x"382134ac",  9838 => x"f8000506",  9839 => x"2b9d0004",
     9840 => x"2b8b0008",  9841 => x"379c0024",  9842 => x"c3a00000",
     9843 => x"379cffe0",  9844 => x"5b8b000c",  9845 => x"5b8c0008",
     9846 => x"5b9d0004",  9847 => x"b8404800",  9848 => x"78020001",
     9849 => x"b8205000",  9850 => x"b8400800",  9851 => x"b8605800",
     9852 => x"b9401000",  9853 => x"b9201800",  9854 => x"382134b0",
     9855 => x"b8806000",  9856 => x"5b840010",  9857 => x"5b850014",
     9858 => x"5b860018",  9859 => x"5b87001c",  9860 => x"5b880020",
     9861 => x"f80004ef",  9862 => x"21620080",  9863 => x"78030001",
     9864 => x"64420000",  9865 => x"b8600800",  9866 => x"34030002",
     9867 => x"c8621000",  9868 => x"382134a0",  9869 => x"2163007f",
     9870 => x"f80004e6",  9871 => x"37820014",  9872 => x"b9800800",
     9873 => x"f80004c1",  9874 => x"78010001",  9875 => x"382134ac",
     9876 => x"f80004e0",  9877 => x"2b9d0004",  9878 => x"2b8b000c",
     9879 => x"2b8c0008",  9880 => x"379c0020",  9881 => x"c3a00000",
     9882 => x"379cfffc",  9883 => x"5b9d0004",  9884 => x"78010001",
     9885 => x"382134bc",  9886 => x"f80004d6",  9887 => x"2b9d0004",
     9888 => x"379c0004",  9889 => x"c3a00000",  9890 => x"40240000",
     9891 => x"3402002d",  9892 => x"34030001",  9893 => x"5c820003",
     9894 => x"34210001",  9895 => x"3403ffff",  9896 => x"34020000",
     9897 => x"34050009",  9898 => x"e0000004",  9899 => x"0842000a",
     9900 => x"34210001",  9901 => x"b4821000",  9902 => x"40240000",
     9903 => x"3484ffd0",  9904 => x"208600ff",  9905 => x"50a6fffa",
     9906 => x"88430800",  9907 => x"c3a00000",  9908 => x"379cfff4",
     9909 => x"5b8b000c",  9910 => x"5b8c0008",  9911 => x"5b9d0004",
     9912 => x"b8206000",  9913 => x"f8000aed",  9914 => x"342b0001",
     9915 => x"f8000aeb",  9916 => x"5c2bffff",  9917 => x"b9800800",
     9918 => x"e0000002",  9919 => x"3421ffff",  9920 => x"4820ffff",
     9921 => x"f8000ae5",  9922 => x"c82b0800",  9923 => x"2b9d0004",
     9924 => x"2b8b000c",  9925 => x"2b8c0008",  9926 => x"379c000c",
     9927 => x"c3a00000",  9928 => x"379cfff0",  9929 => x"5b8b0010",
     9930 => x"5b8c000c",  9931 => x"5b8d0008",  9932 => x"5b9d0004",
     9933 => x"340b0400",  9934 => x"340c0400",  9935 => x"e0000003",
     9936 => x"b58b6000",  9937 => x"3d6b0001",  9938 => x"b9800800",
     9939 => x"fbffffe1",  9940 => x"4420fffc",  9941 => x"158c0001",
     9942 => x"156b0002",  9943 => x"e0000009",  9944 => x"b56c6800",
     9945 => x"b9a00800",  9946 => x"fbffffda",  9947 => x"5c200002",
     9948 => x"b9a06000",  9949 => x"0161001f",  9950 => x"b42b5800",
     9951 => x"156b0001",  9952 => x"5d60fff8",  9953 => x"78010001",
     9954 => x"382152d4",  9955 => x"582c0000",  9956 => x"78010001",
     9957 => x"b9801000",  9958 => x"38213514",  9959 => x"f800048d",
     9960 => x"2b9d0004",  9961 => x"2b8b0010",  9962 => x"2b8c000c",
     9963 => x"2b8d0008",  9964 => x"379c0010",  9965 => x"c3a00000",
     9966 => x"379cfffc",  9967 => x"5b9d0004",  9968 => x"78020001",
     9969 => x"384252d4",  9970 => x"28430000",  9971 => x"34042710",
     9972 => x"0865000a",  9973 => x"e0000004",  9974 => x"3442ffff",
     9975 => x"4840ffff",  9976 => x"3421d8f0",  9977 => x"50810003",
     9978 => x"b8a01000",  9979 => x"e3fffffc",  9980 => x"88230800",
     9981 => x"340203e8",  9982 => x"f8001ced",  9983 => x"e0000002",
     9984 => x"3421ffff",  9985 => x"4820ffff",  9986 => x"34010000",
     9987 => x"2b9d0004",  9988 => x"379c0004",  9989 => x"c3a00000",
     9990 => x"379cfffc",  9991 => x"5b9d0004",  9992 => x"b8400800",
     9993 => x"f8000573",  9994 => x"34010000",  9995 => x"2b9d0004",
     9996 => x"379c0004",  9997 => x"c3a00000",  9998 => x"78020001",
     9999 => x"384252d8", 10000 => x"58410018", 10001 => x"58410240",
    10002 => x"58410468", 10003 => x"58410690", 10004 => x"c3a00000",
    10005 => x"379cff24", 10006 => x"5b8b0014", 10007 => x"5b8c0010",
    10008 => x"5b8d000c", 10009 => x"5b8e0008", 10010 => x"5b9d0004",
    10011 => x"78010001", 10012 => x"b8607000", 10013 => x"382152d8",
    10014 => x"340c0000", 10015 => x"34020004", 10016 => x"28230000",
    10017 => x"5c600009", 10018 => x"78040001", 10019 => x"b8801000",
    10020 => x"37810018", 10021 => x"3842352c", 10022 => x"fbffdd12",
    10023 => x"340b0000", 10024 => x"4961001d", 10025 => x"e0000006",
    10026 => x"358c0001", 10027 => x"34210228", 10028 => x"5d82fff4",
    10029 => x"340b0000", 10030 => x"e0000017", 10031 => x"098d0228",
    10032 => x"780c0001", 10033 => x"398c52d8", 10034 => x"b5ac5800",
    10035 => x"b9c01000", 10036 => x"3403000e", 10037 => x"35610004",
    10038 => x"f8001d16", 10039 => x"35610012", 10040 => x"f8000544",
    10041 => x"2b8100d0", 10042 => x"34020200", 10043 => x"0d600220",
    10044 => x"59610018", 10045 => x"2b8100b8", 10046 => x"5961001c",
    10047 => x"35610220", 10048 => x"0c200002", 10049 => x"0c220004",
    10050 => x"0c200006", 10051 => x"34010001", 10052 => x"59610000",
    10053 => x"b9600800", 10054 => x"2b9d0004", 10055 => x"2b8b0014",
    10056 => x"2b8c0010", 10057 => x"2b8d000c", 10058 => x"2b8e0008",
    10059 => x"379c00dc", 10060 => x"c3a00000", 10061 => x"44200002",
    10062 => x"58200000", 10063 => x"34010000", 10064 => x"c3a00000",
    10065 => x"379cffe8", 10066 => x"5b8b0018", 10067 => x"5b8c0014",
    10068 => x"5b8d0010", 10069 => x"5b8e000c", 10070 => x"5b8f0008",
    10071 => x"5b9d0004", 10072 => x"b8205800", 10073 => x"59620010",
    10074 => x"b8407000", 10075 => x"b8807800", 10076 => x"b8a06000",
    10077 => x"282d0008", 10078 => x"44600005", 10079 => x"b8a00800",
    10080 => x"3402fc18", 10081 => x"f8001c3d", 10082 => x"b42d6800",
    10083 => x"c9cf2000", 10084 => x"b8801800", 10085 => x"4c800002",
    10086 => x"b48c1800", 10087 => x"0181001f", 10088 => x"b42c0800",
    10089 => x"14210001", 10090 => x"b4242000", 10091 => x"4c800002",
    10092 => x"b48c2000", 10093 => x"49840002", 10094 => x"c88c2000",
    10095 => x"09820003", 10096 => x"1445001f", 10097 => x"00a5001e",
    10098 => x"b4a21000", 10099 => x"14420002", 10100 => x"48620006",
    10101 => x"1582001f", 10102 => x"0042001e", 10103 => x"b44c1000",
    10104 => x"14420002", 10105 => x"4c62000d", 10106 => x"b4812000",
    10107 => x"596d0008", 10108 => x"5964000c", 10109 => x"4984000a",
    10110 => x"c88c2000", 10111 => x"5964000c", 10112 => x"b9800800",
    10113 => x"340203e8", 10114 => x"f8001c1c", 10115 => x"b5a10800",
    10116 => x"59610008", 10117 => x"e0000002", 10118 => x"5963000c",
    10119 => x"78030001", 10120 => x"38633cc4", 10121 => x"29610008",
    10122 => x"28620000", 10123 => x"4c41000d", 10124 => x"78030001",
    10125 => x"38633cd8", 10126 => x"28620000", 10127 => x"29630000",
    10128 => x"b4220800", 10129 => x"29620004", 10130 => x"59610008",
    10131 => x"34410001", 10132 => x"f4411000", 10133 => x"59610004",
    10134 => x"b4431000", 10135 => x"59620000", 10136 => x"2b9d0004",
    10137 => x"2b8b0018", 10138 => x"2b8c0014", 10139 => x"2b8d0010",
    10140 => x"2b8e000c", 10141 => x"2b8f0008", 10142 => x"379c0018",
    10143 => x"c3a00000", 10144 => x"379cffb8", 10145 => x"5b8b0020",
    10146 => x"5b8c001c", 10147 => x"5b8d0018", 10148 => x"5b8e0014",
    10149 => x"5b8f0010", 10150 => x"5b90000c", 10151 => x"5b910008",
    10152 => x"5b9d0004", 10153 => x"b8407800", 10154 => x"2c220226",
    10155 => x"b8205800", 10156 => x"b8806800", 10157 => x"b8a06000",
    10158 => x"34010000", 10159 => x"4440007f", 10160 => x"2d610222",
    10161 => x"3442ffff", 10162 => x"0d620226", 10163 => x"b5612000",
    10164 => x"40840020", 10165 => x"34210001", 10166 => x"2021ffff",
    10167 => x"3384004a", 10168 => x"0d610222", 10169 => x"34040200",
    10170 => x"2d620224", 10171 => x"5c240002", 10172 => x"0d600222",
    10173 => x"2d610222", 10174 => x"b5612000", 10175 => x"40840020",
    10176 => x"34210001", 10177 => x"2021ffff", 10178 => x"3384004b",
    10179 => x"0d610222", 10180 => x"34040200", 10181 => x"5c240002",
    10182 => x"0d600222", 10183 => x"34420002", 10184 => x"2042ffff",
    10185 => x"0d620224", 10186 => x"3787004a", 10187 => x"3785003c",
    10188 => x"34060200", 10189 => x"e000000b", 10190 => x"2d610222",
    10191 => x"b5612000", 10192 => x"40840020", 10193 => x"34210001",
    10194 => x"2021ffff", 10195 => x"30a40000", 10196 => x"0d610222",
    10197 => x"34a50001", 10198 => x"5c260002", 10199 => x"0d600222",
    10200 => x"5ca7fff6", 10201 => x"3442000e", 10202 => x"2042ffff",
    10203 => x"0d620224", 10204 => x"3787003c", 10205 => x"37850024",
    10206 => x"34060200", 10207 => x"e000000b", 10208 => x"2d610222",
    10209 => x"b5612000", 10210 => x"40840020", 10211 => x"34210001",
    10212 => x"2021ffff", 10213 => x"30a40000", 10214 => x"0d610222",
    10215 => x"34a50001", 10216 => x"5c260002", 10217 => x"0d600222",
    10218 => x"5ca7fff6", 10219 => x"34420018", 10220 => x"2f8e004a",
    10221 => x"2042ffff", 10222 => x"0d620224", 10223 => x"b9a00800",
    10224 => x"51cd0002", 10225 => x"b9c00800", 10226 => x"b4613000",
    10227 => x"34050200", 10228 => x"e000000c", 10229 => x"2d640222",
    10230 => x"b5642000", 10231 => x"40840020", 10232 => x"30640000",
    10233 => x"2d640222", 10234 => x"34630001", 10235 => x"34840001",
    10236 => x"2084ffff", 10237 => x"0d640222", 10238 => x"5c850002",
    10239 => x"0d600222", 10240 => x"5c66fff5", 10241 => x"b4410800",
    10242 => x"0d610224", 10243 => x"2f810048", 10244 => x"37820042",
    10245 => x"34030006", 10246 => x"0de1000c", 10247 => x"b9e00800",
    10248 => x"f8001c44", 10249 => x"35e10006", 10250 => x"3782003c",
    10251 => x"34030006", 10252 => x"f8001c40", 10253 => x"4580001d",
    10254 => x"2b900034", 10255 => x"2b8f0028", 10256 => x"34010000",
    10257 => x"59900014", 10258 => x"598f0018", 10259 => x"f80018ea",
    10260 => x"b8208800", 10261 => x"35820010", 10262 => x"34030000",
    10263 => x"34010000", 10264 => x"f800188f", 10265 => x"2b81002c",
    10266 => x"43820024", 10267 => x"29640018", 10268 => x"59810000",
    10269 => x"2b810030", 10270 => x"59900008", 10271 => x"5980000c",
    10272 => x"59810004", 10273 => x"222100ff", 10274 => x"64210000",
    10275 => x"b9e01800", 10276 => x"a0220800", 10277 => x"29820010",
    10278 => x"5981001c", 10279 => x"34051f40", 10280 => x"b9800800",
    10281 => x"fbffff28", 10282 => x"35cefff2", 10283 => x"b9a00800",
    10284 => x"51cd0002", 10285 => x"b9c00800", 10286 => x"2b9d0004",
    10287 => x"2b8b0020", 10288 => x"2b8c001c", 10289 => x"2b8d0018",
    10290 => x"2b8e0014", 10291 => x"2b8f0010", 10292 => x"2b90000c",
    10293 => x"2b910008", 10294 => x"379c0048", 10295 => x"c3a00000",
    10296 => x"379cffbc", 10297 => x"5b8b001c", 10298 => x"5b8c0018",
    10299 => x"5b8d0014", 10300 => x"5b8e0010", 10301 => x"5b8f000c",
    10302 => x"5b900008", 10303 => x"5b9d0004", 10304 => x"378c0038",
    10305 => x"b8208000", 10306 => x"b8607800", 10307 => x"b9800800",
    10308 => x"34030006", 10309 => x"b8807000", 10310 => x"b8406800",
    10311 => x"b8a05800", 10312 => x"f8001c04", 10313 => x"36020012",
    10314 => x"34030006", 10315 => x"3781003e", 10316 => x"f8001c00",
    10317 => x"2da1000c", 10318 => x"b9e01000", 10319 => x"35c3000e",
    10320 => x"0f810044", 10321 => x"37840020", 10322 => x"b9800800",
    10323 => x"f80007de", 10324 => x"4560000a", 10325 => x"2b820028",
    10326 => x"5960000c", 10327 => x"59620000", 10328 => x"2b82002c",
    10329 => x"59620004", 10330 => x"2b820030", 10331 => x"59620008",
    10332 => x"43820020", 10333 => x"5962001c", 10334 => x"2b9d0004",
    10335 => x"2b8b001c", 10336 => x"2b8c0018", 10337 => x"2b8d0014",
    10338 => x"2b8e0010", 10339 => x"2b8f000c", 10340 => x"2b900008",
    10341 => x"379c0044", 10342 => x"c3a00000", 10343 => x"379cffc4",
    10344 => x"5b8b0020", 10345 => x"5b8c001c", 10346 => x"5b8d0018",
    10347 => x"5b8e0014", 10348 => x"5b8f0010", 10349 => x"5b90000c",
    10350 => x"5b9b0008", 10351 => x"5b9d0004", 10352 => x"780b0001",
    10353 => x"396b5d58", 10354 => x"78020001", 10355 => x"b9600800",
    10356 => x"38425b78", 10357 => x"340301e0", 10358 => x"37840024",
    10359 => x"f800070e", 10360 => x"b8207000", 10361 => x"4c01006d",
    10362 => x"780c0001", 10363 => x"398c52d8", 10364 => x"340d0000",
    10365 => x"b9808000", 10366 => x"b9607800", 10367 => x"341b0004",
    10368 => x"09ab0228", 10369 => x"29810000", 10370 => x"b5705800",
    10371 => x"44200009", 10372 => x"b9e00800", 10373 => x"35620004",
    10374 => x"34030006", 10375 => x"f8001ba4", 10376 => x"5c200004",
    10377 => x"2de2000c", 10378 => x"2d810010", 10379 => x"44410005",
    10380 => x"35ad0001", 10381 => x"358c0228", 10382 => x"5dbbfff2",
    10383 => x"e0000057", 10384 => x"2d630224", 10385 => x"35c10028",
    10386 => x"48230054", 10387 => x"2d620220", 10388 => x"21c1ffff",
    10389 => x"00250008", 10390 => x"b5622000", 10391 => x"34420001",
    10392 => x"0f81003e", 10393 => x"2042ffff", 10394 => x"30850020",
    10395 => x"0d620220", 10396 => x"34040200", 10397 => x"5c440002",
    10398 => x"0d600220", 10399 => x"2d620220", 10400 => x"4385003f",
    10401 => x"b5622000", 10402 => x"34420001", 10403 => x"2042ffff",
    10404 => x"30850020", 10405 => x"0d620220", 10406 => x"34040200",
    10407 => x"5c440002", 10408 => x"0d600220", 10409 => x"3463fffe",
    10410 => x"78020001", 10411 => x"2063ffff", 10412 => x"38425d58",
    10413 => x"0d630224", 10414 => x"3446000e", 10415 => x"34050200",
    10416 => x"e000000b", 10417 => x"2d640220", 10418 => x"40480000",
    10419 => x"34420001", 10420 => x"b5643800", 10421 => x"34840001",
    10422 => x"2084ffff", 10423 => x"30e80020", 10424 => x"0d640220",
    10425 => x"5c850002", 10426 => x"0d600220", 10427 => x"5c46fff6",
    10428 => x"3463fff2", 10429 => x"2063ffff", 10430 => x"0d630224",
    10431 => x"379b003c", 10432 => x"37820024", 10433 => x"34050200",
    10434 => x"e000000b", 10435 => x"2d640220", 10436 => x"40470000",
    10437 => x"34420001", 10438 => x"b5643000", 10439 => x"34840001",
    10440 => x"2084ffff", 10441 => x"30c70020", 10442 => x"0d640220",
    10443 => x"5c850002", 10444 => x"0d600220", 10445 => x"5c5bfff6",
    10446 => x"3463ffe8", 10447 => x"78020001", 10448 => x"2063ffff",
    10449 => x"38425b78", 10450 => x"0d630224", 10451 => x"b4223000",
    10452 => x"34050200", 10453 => x"e000000b", 10454 => x"2d640220",
    10455 => x"40480000", 10456 => x"34420001", 10457 => x"b5643800",
    10458 => x"34840001", 10459 => x"2084ffff", 10460 => x"30e80020",
    10461 => x"0d640220", 10462 => x"5c850002", 10463 => x"0d600220",
    10464 => x"5c46fff6", 10465 => x"c8610800", 10466 => x"0d610224",
    10467 => x"2d610226", 10468 => x"34210001", 10469 => x"0d610226",
    10470 => x"2b9d0004", 10471 => x"2b8b0020", 10472 => x"2b8c001c",
    10473 => x"2b8d0018", 10474 => x"2b8e0014", 10475 => x"2b8f0010",
    10476 => x"2b90000c", 10477 => x"2b9b0008", 10478 => x"379c003c",
    10479 => x"c3a00000", 10480 => x"379cffe8", 10481 => x"5b8b0008",
    10482 => x"5b9d0004", 10483 => x"378b000c", 10484 => x"b9600800",
    10485 => x"34020000", 10486 => x"3403000e", 10487 => x"f8001bd3",
    10488 => x"b9600800", 10489 => x"340200ff", 10490 => x"34030006",
    10491 => x"f8001bcf", 10492 => x"34010806", 10493 => x"0f810018",
    10494 => x"34020000", 10495 => x"b9601800", 10496 => x"34010000",
    10497 => x"fbfffe14", 10498 => x"78020001", 10499 => x"38425d68",
    10500 => x"58410000", 10501 => x"2b9d0004", 10502 => x"2b8b0008",
    10503 => x"379c0018", 10504 => x"c3a00000", 10505 => x"379cff38",
    10506 => x"5b8b0028", 10507 => x"5b8c0024", 10508 => x"5b8d0020",
    10509 => x"5b8e001c", 10510 => x"5b8f0018", 10511 => x"5b900014",
    10512 => x"5b910010", 10513 => x"5b92000c", 10514 => x"5b930008",
    10515 => x"5b9d0004", 10516 => x"78010001", 10517 => x"38215d6c",
    10518 => x"282c0000", 10519 => x"5d800047", 10520 => x"780b0001",
    10521 => x"396b5d68", 10522 => x"29610000", 10523 => x"378e00ac",
    10524 => x"378d002c", 10525 => x"b9c01000", 10526 => x"b9a01800",
    10527 => x"34040080", 10528 => x"34050000", 10529 => x"fbfffe7f",
    10530 => x"4d81003c", 10531 => x"3402001b", 10532 => x"4c41003a",
    10533 => x"378c00c4", 10534 => x"b9800800", 10535 => x"f800012a",
    10536 => x"43810032", 10537 => x"5c200035", 10538 => x"43930033",
    10539 => x"34010001", 10540 => x"5e610032", 10541 => x"378f0044",
    10542 => x"b9e00800", 10543 => x"b9801000", 10544 => x"34030004",
    10545 => x"f8001afa", 10546 => x"5c20002c", 10547 => x"379000bc",
    10548 => x"37920034", 10549 => x"ba401000", 10550 => x"34030006",
    10551 => x"ba000800", 10552 => x"f8001b14", 10553 => x"3791003a",
    10554 => x"ba201000", 10555 => x"34030004", 10556 => x"378100c8",
    10557 => x"f8001b0f", 10558 => x"34010008", 10559 => x"3381002e",
    10560 => x"34010006", 10561 => x"33810030", 10562 => x"34010004",
    10563 => x"33810031", 10564 => x"34010002", 10565 => x"33810033",
    10566 => x"ba400800", 10567 => x"3380002c", 10568 => x"3393002d",
    10569 => x"3380002f", 10570 => x"33800032", 10571 => x"f8000331",
    10572 => x"b9801000", 10573 => x"34030004", 10574 => x"ba200800",
    10575 => x"f8001afd", 10576 => x"ba001000", 10577 => x"34030006",
    10578 => x"3781003e", 10579 => x"f8001af9", 10580 => x"378200c8",
    10581 => x"34030004", 10582 => x"b9e00800", 10583 => x"f8001af5",
    10584 => x"29610000", 10585 => x"b9c01000", 10586 => x"b9a01800",
    10587 => x"3404001c", 10588 => x"34050000", 10589 => x"fbfffedb",
    10590 => x"2b9d0004", 10591 => x"2b8b0028", 10592 => x"2b8c0024",
    10593 => x"2b8d0020", 10594 => x"2b8e001c", 10595 => x"2b8f0018",
    10596 => x"2b900014", 10597 => x"2b910010", 10598 => x"2b92000c",
    10599 => x"2b930008", 10600 => x"379c00c8", 10601 => x"c3a00000",
    10602 => x"379cffe0", 10603 => x"5b8b0018", 10604 => x"5b8c0014",
    10605 => x"5b8d0010", 10606 => x"5b8e000c", 10607 => x"5b8f0008",
    10608 => x"5b9d0004", 10609 => x"378d001c", 10610 => x"b8205800",
    10611 => x"b9a00800", 10612 => x"f80000dd", 10613 => x"41620000",
    10614 => x"34010045", 10615 => x"340c0000", 10616 => x"5c41004a",
    10617 => x"356e0010", 10618 => x"b9a01000", 10619 => x"b9c00800",
    10620 => x"34030004", 10621 => x"f8001aae", 10622 => x"b8201000",
    10623 => x"5c200043", 10624 => x"41640009", 10625 => x"34030001",
    10626 => x"416d0002", 10627 => x"41610003", 10628 => x"b8406000",
    10629 => x"5c83003d", 10630 => x"41630014", 10631 => x"34020008",
    10632 => x"5c62003a", 10633 => x"3dad0008", 10634 => x"b9a16800",
    10635 => x"35adffe8", 10636 => x"34010040", 10637 => x"4c2d0002",
    10638 => x"340d0040", 10639 => x"356f000c", 10640 => x"b9e01000",
    10641 => x"34030004", 10642 => x"37810020", 10643 => x"f8001ab9",
    10644 => x"35ac0018", 10645 => x"34010045", 10646 => x"31610000",
    10647 => x"15810008", 10648 => x"3782001c", 10649 => x"31610002",
    10650 => x"3401003f", 10651 => x"31610008", 10652 => x"34010001",
    10653 => x"31610009", 10654 => x"34030004", 10655 => x"31600001",
    10656 => x"316c0003", 10657 => x"31600004", 10658 => x"31600005",
    10659 => x"31600006", 10660 => x"31600007", 10661 => x"3160000a",
    10662 => x"3160000b", 10663 => x"b9e00800", 10664 => x"f8001aa4",
    10665 => x"34030004", 10666 => x"37820020", 10667 => x"b9c00800",
    10668 => x"f8001aa0", 10669 => x"35ad0005", 10670 => x"01a1001f",
    10671 => x"31600014", 10672 => x"b42d6800", 10673 => x"15a20001",
    10674 => x"31600015", 10675 => x"31600016", 10676 => x"31600017",
    10677 => x"35610014", 10678 => x"f8000015", 10679 => x"2021ffff",
    10680 => x"00220008", 10681 => x"31610017", 10682 => x"31620016",
    10683 => x"b9600800", 10684 => x"3402000a", 10685 => x"f800000e",
    10686 => x"2021ffff", 10687 => x"00220008", 10688 => x"3161000b",
    10689 => x"3162000a", 10690 => x"b9800800", 10691 => x"2b9d0004",
    10692 => x"2b8b0018", 10693 => x"2b8c0014", 10694 => x"2b8d0010",
    10695 => x"2b8e000c", 10696 => x"2b8f0008", 10697 => x"379c0020",
    10698 => x"c3a00000", 10699 => x"34030000", 10700 => x"34040000",
    10701 => x"e0000005", 10702 => x"2c250000", 10703 => x"34840001",
    10704 => x"34210002", 10705 => x"b4651800", 10706 => x"4844fffc",
    10707 => x"00610010", 10708 => x"2063ffff", 10709 => x"b4611800",
    10710 => x"00610010", 10711 => x"b4231800", 10712 => x"a4600800",
    10713 => x"2021ffff", 10714 => x"c3a00000", 10715 => x"379cffe8",
    10716 => x"5b8b0008", 10717 => x"5b9d0004", 10718 => x"78010001",
    10719 => x"378b000c", 10720 => x"38215d6c", 10721 => x"34020000",
    10722 => x"3403000e", 10723 => x"58200000", 10724 => x"b9600800",
    10725 => x"f8001ae5", 10726 => x"b9600800", 10727 => x"f8000295",
    10728 => x"34010800", 10729 => x"0f810018", 10730 => x"34020000",
    10731 => x"b9601800", 10732 => x"34010000", 10733 => x"fbfffd28",
    10734 => x"78020001", 10735 => x"38425d74", 10736 => x"58410000",
    10737 => x"2b9d0004", 10738 => x"2b8b0008", 10739 => x"379c0018",
    10740 => x"c3a00000", 10741 => x"379cfe50", 10742 => x"5b8b0010",
    10743 => x"5b8c000c", 10744 => x"5b8d0008", 10745 => x"5b9d0004",
    10746 => x"78020001", 10747 => x"38425d74", 10748 => x"28410000",
    10749 => x"378c0014", 10750 => x"378201a4", 10751 => x"b9801800",
    10752 => x"34040190", 10753 => x"34050000", 10754 => x"fbfffd9e",
    10755 => x"b8205800", 10756 => x"4c010019", 10757 => x"78020001",
    10758 => x"38425d6c", 10759 => x"28410000", 10760 => x"44200004",
    10761 => x"b9800800", 10762 => x"b9601000", 10763 => x"f8000110",
    10764 => x"78010001", 10765 => x"38215d6c", 10766 => x"282d0000",
    10767 => x"5da0000e", 10768 => x"378c0014", 10769 => x"b9800800",
    10770 => x"b9601000", 10771 => x"fbffff57", 10772 => x"b8202000",
    10773 => x"4da10008", 10774 => x"78020001", 10775 => x"38425d74",
    10776 => x"28410000", 10777 => x"b9801800", 10778 => x"378201a4",
    10779 => x"34050000", 10780 => x"fbfffe1c", 10781 => x"78010001",
    10782 => x"38215d6c", 10783 => x"28210000", 10784 => x"4420001d",
    10785 => x"78010001", 10786 => x"38215d78", 10787 => x"28210000",
    10788 => x"5c200019", 10789 => x"78010001", 10790 => x"38215d7c",
    10791 => x"28220000", 10792 => x"378b0014", 10793 => x"378c01a4",
    10794 => x"34420001", 10795 => x"58220000", 10796 => x"b9600800",
    10797 => x"f8000058", 10798 => x"b8206800", 10799 => x"340200ff",
    10800 => x"34030006", 10801 => x"b9800800", 10802 => x"f8001a98",
    10803 => x"78050001", 10804 => x"34010800", 10805 => x"38a55d74",
    10806 => x"0f8101b0", 10807 => x"28a10000", 10808 => x"b9801000",
    10809 => x"b9601800", 10810 => x"b9a02000", 10811 => x"34050000",
    10812 => x"fbfffdfc", 10813 => x"78010001", 10814 => x"38215d6c",
    10815 => x"28210000", 10816 => x"4420000b", 10817 => x"78010001",
    10818 => x"38215d78", 10819 => x"28220000", 10820 => x"78040001",
    10821 => x"38843cfc", 10822 => x"28830000", 10823 => x"34420001",
    10824 => x"58220000", 10825 => x"5c430002", 10826 => x"58200000",
    10827 => x"2b9d0004", 10828 => x"2b8b0010", 10829 => x"2b8c000c",
    10830 => x"2b8d0008", 10831 => x"379c01b0", 10832 => x"c3a00000",
    10833 => x"379cfffc", 10834 => x"5b9d0004", 10835 => x"78020001",
    10836 => x"38425d70", 10837 => x"34030004", 10838 => x"f80019f6",
    10839 => x"2b9d0004", 10840 => x"379c0004", 10841 => x"c3a00000",
    10842 => x"379cffe4", 10843 => x"5b8b0014", 10844 => x"5b8c0010",
    10845 => x"5b8d000c", 10846 => x"5b8e0008", 10847 => x"5b9d0004",
    10848 => x"78030001", 10849 => x"780b0001", 10850 => x"396b5d70",
    10851 => x"b8206000", 10852 => x"38636dc8", 10853 => x"286d0000",
    10854 => x"b9801000", 10855 => x"34030004", 10856 => x"b9600800",
    10857 => x"f80019e3", 10858 => x"41610001", 10859 => x"416e0000",
    10860 => x"3c210010", 10861 => x"3dce0018", 10862 => x"b9c17000",
    10863 => x"41610003", 10864 => x"b9c17000", 10865 => x"41610002",
    10866 => x"378b0018", 10867 => x"3c210008", 10868 => x"b9c17000",
    10869 => x"b9600800", 10870 => x"f8000206", 10871 => x"b9800800",
    10872 => x"59ae0018", 10873 => x"b9601000", 10874 => x"f8000913",
    10875 => x"78010001", 10876 => x"38215d6c", 10877 => x"58200000",
    10878 => x"2b9d0004", 10879 => x"2b8b0014", 10880 => x"2b8c0010",
    10881 => x"2b8d000c", 10882 => x"2b8e0008", 10883 => x"379c001c",
    10884 => x"c3a00000", 10885 => x"379cffe8", 10886 => x"5b8b0018",
    10887 => x"5b8c0014", 10888 => x"5b8d0010", 10889 => x"5b8e000c",
    10890 => x"5b8f0008", 10891 => x"5b9d0004", 10892 => x"340c0001",
    10893 => x"b8205800", 10894 => x"302c001c", 10895 => x"302c001d",
    10896 => x"34010006", 10897 => x"3161001e", 10898 => x"3160001f",
    10899 => x"35610020", 10900 => x"b8406800", 10901 => x"f80001e7",
    10902 => x"41620024", 10903 => x"41610020", 10904 => x"34030002",
    10905 => x"356e0008", 10906 => x"98410800", 10907 => x"31610020",
    10908 => x"41620025", 10909 => x"41610021", 10910 => x"316d0025",
    10911 => x"356f0010", 10912 => x"98410800", 10913 => x"41620022",
    10914 => x"31610021", 10915 => x"15a10008", 10916 => x"98221000",
    10917 => x"31620022", 10918 => x"41620023", 10919 => x"31610024",
    10920 => x"35610026", 10921 => x"984d1000", 10922 => x"31620023",
    10923 => x"34020000", 10924 => x"f8001a1e", 10925 => x"34020000",
    10926 => x"34030004", 10927 => x"35610028", 10928 => x"f8001a1a",
    10929 => x"34020000", 10930 => x"34030004", 10931 => x"3561002c",
    10932 => x"f8001a16", 10933 => x"34020000", 10934 => x"34030004",
    10935 => x"35610030", 10936 => x"f8001a12", 10937 => x"34020000",
    10938 => x"34030004", 10939 => x"35610034", 10940 => x"f8001a0e",
    10941 => x"356d0038", 10942 => x"34020000", 10943 => x"34030010",
    10944 => x"b9a00800", 10945 => x"f8001a09", 10946 => x"b9a00800",
    10947 => x"f80001b9", 10948 => x"34020000", 10949 => x"34030040",
    10950 => x"35610048", 10951 => x"f8001a03", 10952 => x"34020000",
    10953 => x"34030080", 10954 => x"35610088", 10955 => x"f80019ff",
    10956 => x"34020000", 10957 => x"34030040", 10958 => x"35610108",
    10959 => x"f80019fb", 10960 => x"34020000", 10961 => x"34030004",
    10962 => x"b9c00800", 10963 => x"f80019f7", 10964 => x"356d000c",
    10965 => x"340200ff", 10966 => x"34030004", 10967 => x"b9a00800",
    10968 => x"f80019f2", 10969 => x"34010011", 10970 => x"31610011",
    10971 => x"34010044", 10972 => x"34020034", 10973 => x"31610015",
    10974 => x"34010043", 10975 => x"31620013", 10976 => x"31610017",
    10977 => x"31620019", 10978 => x"31600010", 10979 => x"340200a0",
    10980 => x"316c0012", 10981 => x"31600014", 10982 => x"31600016",
    10983 => x"316c0018", 10984 => x"3160001a", 10985 => x"3160001b",
    10986 => x"b9c00800", 10987 => x"fbfffee0", 10988 => x"2022ffff",
    10989 => x"5c400002", 10990 => x"3802ffff", 10991 => x"00410008",
    10992 => x"3162001b", 10993 => x"3161001a", 10994 => x"34010045",
    10995 => x"31610000", 10996 => x"34010001", 10997 => x"31610002",
    10998 => x"34010048", 10999 => x"31610003", 11000 => x"3401003f",
    11001 => x"31610008", 11002 => x"34010011", 11003 => x"31610009",
    11004 => x"31600001", 11005 => x"31600004", 11006 => x"31600005",
    11007 => x"31600006", 11008 => x"31600007", 11009 => x"3160000a",
    11010 => x"3160000b", 11011 => x"b9a00800", 11012 => x"34020000",
    11013 => x"34030004", 11014 => x"f80019c4", 11015 => x"34030004",
    11016 => x"b9e00800", 11017 => x"340200ff", 11018 => x"f80019c0",
    11019 => x"b9600800", 11020 => x"3402000a", 11021 => x"fbfffebe",
    11022 => x"2021ffff", 11023 => x"00220008", 11024 => x"3161000b",
    11025 => x"34010148", 11026 => x"3162000a", 11027 => x"2b9d0004",
    11028 => x"2b8b0018", 11029 => x"2b8c0014", 11030 => x"2b8d0010",
    11031 => x"2b8e000c", 11032 => x"2b8f0008", 11033 => x"379c0018",
    11034 => x"c3a00000", 11035 => x"379cffe0", 11036 => x"5b8b0014",
    11037 => x"5b8c0010", 11038 => x"5b8d000c", 11039 => x"5b8e0008",
    11040 => x"5b9d0004", 11041 => x"378d0018", 11042 => x"b8205800",
    11043 => x"b9a00800", 11044 => x"b8407000", 11045 => x"f8000157",
    11046 => x"34010148", 11047 => x"340c0000", 11048 => x"5dc10022",
    11049 => x"41620000", 11050 => x"34010045", 11051 => x"5c41001f",
    11052 => x"41620009", 11053 => x"34010011", 11054 => x"5c41001c",
    11055 => x"41610016", 11056 => x"5c20001a", 11057 => x"41620017",
    11058 => x"34010044", 11059 => x"5c410017", 11060 => x"41610014",
    11061 => x"5c200015", 11062 => x"41620015", 11063 => x"34010043",
    11064 => x"5c410012", 11065 => x"35610038", 11066 => x"b9a01000",
    11067 => x"34030006", 11068 => x"f80018ef", 11069 => x"5c20000d",
    11070 => x"3561002c", 11071 => x"fbffff1b", 11072 => x"37810020",
    11073 => x"fbffff10", 11074 => x"43820020", 11075 => x"43830021",
    11076 => x"43840022", 11077 => x"43850023", 11078 => x"78010001",
    11079 => x"38213530", 11080 => x"f800002c", 11081 => x"340c0001",
    11082 => x"b9800800", 11083 => x"2b9d0004", 11084 => x"2b8b0014",
    11085 => x"2b8c0010", 11086 => x"2b8d000c", 11087 => x"2b8e0008",
    11088 => x"379c0020", 11089 => x"c3a00000", 11090 => x"379cfff4",
    11091 => x"5b8b000c", 11092 => x"5b8c0008", 11093 => x"5b9d0004",
    11094 => x"780b0001", 11095 => x"b8202000", 11096 => x"396b5d80",
    11097 => x"b8401800", 11098 => x"b9600800", 11099 => x"b8801000",
    11100 => x"f8000027", 11101 => x"b8206000", 11102 => x"b9600800",
    11103 => x"f8000e96", 11104 => x"b9800800", 11105 => x"2b9d0004",
    11106 => x"2b8b000c", 11107 => x"2b8c0008", 11108 => x"379c000c",
    11109 => x"c3a00000", 11110 => x"379cffe0", 11111 => x"5b9d0004",
    11112 => x"5b83000c", 11113 => x"3783000c", 11114 => x"5b820008",
    11115 => x"5b840010", 11116 => x"5b850014", 11117 => x"5b860018",
    11118 => x"5b87001c", 11119 => x"5b880020", 11120 => x"f8000013",
    11121 => x"2b9d0004", 11122 => x"379c0020", 11123 => x"c3a00000",
    11124 => x"379cffdc", 11125 => x"5b9d0004", 11126 => x"5b82000c",
    11127 => x"3782000c", 11128 => x"5b810008", 11129 => x"5b830010",
    11130 => x"5b840014", 11131 => x"5b850018", 11132 => x"5b86001c",
    11133 => x"5b870020", 11134 => x"5b880024", 11135 => x"fbffffd3",
    11136 => x"2b9d0004", 11137 => x"379c0024", 11138 => x"c3a00000",
    11139 => x"379cff94", 11140 => x"5b8b0044", 11141 => x"5b8c0040",
    11142 => x"5b8d003c", 11143 => x"5b8e0038", 11144 => x"5b8f0034",
    11145 => x"5b900030", 11146 => x"5b91002c", 11147 => x"5b920028",
    11148 => x"5b930024", 11149 => x"5b940020", 11150 => x"5b95001c",
    11151 => x"5b960018", 11152 => x"5b970014", 11153 => x"5b980010",
    11154 => x"5b99000c", 11155 => x"5b9b0008", 11156 => x"5b9d0004",
    11157 => x"78160001", 11158 => x"b820c800", 11159 => x"b840a000",
    11160 => x"b8209800", 11161 => x"34180025", 11162 => x"34090069",
    11163 => x"34080070", 11164 => x"34070058", 11165 => x"34060063",
    11166 => x"34050064", 11167 => x"341b002a", 11168 => x"340a0030",
    11169 => x"34170010", 11170 => x"37950060", 11171 => x"3ad63558",
    11172 => x"e0000093", 11173 => x"34110001", 11174 => x"34100020",
    11175 => x"340e000a", 11176 => x"44380004", 11177 => x"32610000",
    11178 => x"e0000038", 11179 => x"34100030", 11180 => x"36940001",
    11181 => x"42810000", 11182 => x"4429003c", 11183 => x"5429000d",
    11184 => x"44270037", 11185 => x"54270008", 11186 => x"443b0018",
    11187 => x"543b0004", 11188 => x"44200085", 11189 => x"5c380017",
    11190 => x"e000002b", 11191 => x"5c2a0015", 11192 => x"e3fffff3",
    11193 => x"44260019", 11194 => x"5c250012", 11195 => x"e000002f",
    11196 => x"4428002b", 11197 => x"54280006", 11198 => x"3402006e",
    11199 => x"44220077", 11200 => x"3404006f", 11201 => x"5c24000b",
    11202 => x"e0000022", 11203 => x"34020075", 11204 => x"44220026",
    11205 => x"34040078", 11206 => x"44240021", 11207 => x"34020073",
    11208 => x"5c220004", 11209 => x"e000000e", 11210 => x"286e0000",
    11211 => x"34630004", 11212 => x"3422ffcf", 11213 => x"204200ff",
    11214 => x"34040008", 11215 => x"5444ffdd", 11216 => x"3431ffd0",
    11217 => x"e3ffffdb", 11218 => x"28610000", 11219 => x"34630004",
    11220 => x"32610000", 11221 => x"36730001", 11222 => x"e0000060",
    11223 => x"b8600800", 11224 => x"28210000", 11225 => x"34630004",
    11226 => x"e0000004", 11227 => x"32620000", 11228 => x"34210001",
    11229 => x"36730001", 11230 => x"40220000", 11231 => x"5c40fffc",
    11232 => x"e0000056", 11233 => x"32780000", 11234 => x"36730001",
    11235 => x"e0000053", 11236 => x"3401000a", 11237 => x"45c10004",
    11238 => x"e0000004", 11239 => x"340e0010", 11240 => x"e0000002",
    11241 => x"340e0008", 11242 => x"286d0000", 11243 => x"34720004",
    11244 => x"65c3000a", 11245 => x"01a4001f", 11246 => x"340f0000",
    11247 => x"a0831800", 11248 => x"44600003", 11249 => x"c80d6800",
    11250 => x"340f0001", 11251 => x"340c0010", 11252 => x"e0000019",
    11253 => x"b9a00800", 11254 => x"b9c01000", 11255 => x"5b85004c",
    11256 => x"5b860050", 11257 => x"5b870054", 11258 => x"5b880058",
    11259 => x"5b89005c", 11260 => x"5b8a0048", 11261 => x"f80017fe",
    11262 => x"b6c11800", 11263 => x"40630000", 11264 => x"358cffff",
    11265 => x"b6ac5800", 11266 => x"b9a00800", 11267 => x"31630000",
    11268 => x"b9c01000", 11269 => x"f80017e6", 11270 => x"2b8a0048",
    11271 => x"2b89005c", 11272 => x"2b880058", 11273 => x"2b870054",
    11274 => x"2b860050", 11275 => x"2b85004c", 11276 => x"b8206800",
    11277 => x"7d840000", 11278 => x"7da30000", 11279 => x"a0831800",
    11280 => x"5c60ffe5", 11281 => x"5d970004", 11282 => x"34020030",
    11283 => x"3382006f", 11284 => x"340c000f", 11285 => x"66020020",
    11286 => x"a1e21000", 11287 => x"4440000b", 11288 => x"358cffff",
    11289 => x"b6ac1000", 11290 => x"3403002d", 11291 => x"30430000",
    11292 => x"340f0000", 11293 => x"e0000005", 11294 => x"358cffff",
    11295 => x"b6ac1000", 11296 => x"30500000", 11297 => x"e0000003",
    11298 => x"caf10800", 11299 => x"b42f0800", 11300 => x"4981fffa",
    11301 => x"45e00005", 11302 => x"358cffff", 11303 => x"b6ac0800",
    11304 => x"3402002d", 11305 => x"30220000", 11306 => x"caec1800",
    11307 => x"ba600800", 11308 => x"3404000f", 11309 => x"e0000006",
    11310 => x"b6ac1000", 11311 => x"40420000", 11312 => x"358c0001",
    11313 => x"30220000", 11314 => x"34210001", 11315 => x"4c8cfffb",
    11316 => x"b6639800", 11317 => x"ba401800", 11318 => x"36940001",
    11319 => x"42810000", 11320 => x"5c20ff6d", 11321 => x"ca790800",
    11322 => x"32600000", 11323 => x"2b9d0004", 11324 => x"2b8b0044",
    11325 => x"2b8c0040", 11326 => x"2b8d003c", 11327 => x"2b8e0038",
    11328 => x"2b8f0034", 11329 => x"2b900030", 11330 => x"2b91002c",
    11331 => x"2b920028", 11332 => x"2b930024", 11333 => x"2b940020",
    11334 => x"2b95001c", 11335 => x"2b960018", 11336 => x"2b970014",
    11337 => x"2b980010", 11338 => x"2b99000c", 11339 => x"2b9b0008",
    11340 => x"379c006c", 11341 => x"c3a00000", 11342 => x"78020001",
    11343 => x"14210002", 11344 => x"38426dbc", 11345 => x"28420000",
    11346 => x"202100ff", 11347 => x"3c210010", 11348 => x"5841002c",
    11349 => x"28410030", 11350 => x"4c20ffff", 11351 => x"28410030",
    11352 => x"2021ffff", 11353 => x"c3a00000", 11354 => x"14210002",
    11355 => x"78030001", 11356 => x"38636dbc", 11357 => x"202100ff",
    11358 => x"28630000", 11359 => x"2042ffff", 11360 => x"78048000",
    11361 => x"3c210010", 11362 => x"b8441000", 11363 => x"b8411000",
    11364 => x"5862002c", 11365 => x"28610030", 11366 => x"4c20ffff",
    11367 => x"c3a00000", 11368 => x"40240002", 11369 => x"40230003",
    11370 => x"78020001", 11371 => x"3c840018", 11372 => x"3c630010",
    11373 => x"38426dbc", 11374 => x"b8831800", 11375 => x"40240005",
    11376 => x"28420000", 11377 => x"b8641800", 11378 => x"40240004",
    11379 => x"3c840008", 11380 => x"b8641800", 11381 => x"58430028",
    11382 => x"40230001", 11383 => x"40210000", 11384 => x"3c210008",
    11385 => x"b8610800", 11386 => x"58410024", 11387 => x"c3a00000",
    11388 => x"78020001", 11389 => x"38426dbc", 11390 => x"28430000",
    11391 => x"28630028", 11392 => x"30230005", 11393 => x"28430000",
    11394 => x"28630028", 11395 => x"00630008", 11396 => x"30230004",
    11397 => x"28430000", 11398 => x"28630028", 11399 => x"00630010",
    11400 => x"30230003", 11401 => x"28430000", 11402 => x"28630028",
    11403 => x"00630018", 11404 => x"30230002", 11405 => x"28430000",
    11406 => x"28630024", 11407 => x"30230001", 11408 => x"28420000",
    11409 => x"28420024", 11410 => x"00420008", 11411 => x"30220000",
    11412 => x"c3a00000", 11413 => x"379cfff4", 11414 => x"5b8b000c",
    11415 => x"5b8c0008", 11416 => x"5b9d0004", 11417 => x"780b0001",
    11418 => x"b8406000", 11419 => x"396b6dbc", 11420 => x"5c200004",
    11421 => x"29610000", 11422 => x"58200000", 11423 => x"e0000022",
    11424 => x"29610000", 11425 => x"58200000", 11426 => x"28220034",
    11427 => x"78010001", 11428 => x"3821356c", 11429 => x"fbfffecf",
    11430 => x"f80000be", 11431 => x"29610000", 11432 => x"340200e0",
    11433 => x"58220000", 11434 => x"78010001", 11435 => x"38215e00",
    11436 => x"34020800", 11437 => x"582c0000", 11438 => x"34010000",
    11439 => x"fbffffab", 11440 => x"340100c8", 11441 => x"f80004fa",
    11442 => x"34010000", 11443 => x"38028000", 11444 => x"fbffffa6",
    11445 => x"34010000", 11446 => x"34020000", 11447 => x"fbffffa3",
    11448 => x"34010010", 11449 => x"34020000", 11450 => x"fbffffa0",
    11451 => x"7d820000", 11452 => x"34010000", 11453 => x"c8021000",
    11454 => x"20421200", 11455 => x"34420140", 11456 => x"fbffff9a",
    11457 => x"34010000", 11458 => x"2b9d0004", 11459 => x"2b8b000c",
    11460 => x"2b8c0008", 11461 => x"379c000c", 11462 => x"c3a00000",
    11463 => x"379cfff0", 11464 => x"5b8b000c", 11465 => x"5b8c0008",
    11466 => x"5b9d0004", 11467 => x"78020001", 11468 => x"38425e00",
    11469 => x"284b0000", 11470 => x"b8206000", 11471 => x"34010004",
    11472 => x"fbffff7e", 11473 => x"7d6b0000", 11474 => x"0f810012",
    11475 => x"34010004", 11476 => x"c80b5800", 11477 => x"fbffff79",
    11478 => x"216b0020", 11479 => x"0f810012", 11480 => x"356b0004",
    11481 => x"45800004", 11482 => x"34010014", 11483 => x"fbffff73",
    11484 => x"0d810000", 11485 => x"2f810012", 11486 => x"a1610800",
    11487 => x"e42b0800", 11488 => x"2b9d0004", 11489 => x"2b8b000c",
    11490 => x"2b8c0008", 11491 => x"379c0010", 11492 => x"c3a00000",
    11493 => x"379cfffc", 11494 => x"5b9d0004", 11495 => x"34010040",
    11496 => x"fbffff66", 11497 => x"00210004", 11498 => x"2021001f",
    11499 => x"08210320", 11500 => x"2b9d0004", 11501 => x"379c0004",
    11502 => x"c3a00000", 11503 => x"379cfff4", 11504 => x"5b8b000c",
    11505 => x"5b8c0008", 11506 => x"5b9d0004", 11507 => x"78030001",
    11508 => x"38634e6c", 11509 => x"b8405800", 11510 => x"28620000",
    11511 => x"58220000", 11512 => x"78010001", 11513 => x"38214e70",
    11514 => x"282c0000", 11515 => x"34010040", 11516 => x"fbffff52",
    11517 => x"00210004", 11518 => x"2021001f", 11519 => x"08210320",
    11520 => x"b42c0800", 11521 => x"59610000", 11522 => x"34010000",
    11523 => x"2b9d0004", 11524 => x"2b8b000c", 11525 => x"2b8c0008",
    11526 => x"379c000c", 11527 => x"c3a00000", 11528 => x"379cfffc",
    11529 => x"5b9d0004", 11530 => x"34010040", 11531 => x"fbffff43",
    11532 => x"38220001", 11533 => x"34010040", 11534 => x"fbffff4c",
    11535 => x"34010000", 11536 => x"2b9d0004", 11537 => x"379c0004",
    11538 => x"c3a00000", 11539 => x"379cfffc", 11540 => x"5b9d0004",
    11541 => x"34010040", 11542 => x"fbffff38", 11543 => x"3402fffe",
    11544 => x"a0221000", 11545 => x"34010040", 11546 => x"fbffff40",
    11547 => x"34010000", 11548 => x"2b9d0004", 11549 => x"379c0004",
    11550 => x"c3a00000", 11551 => x"379cfff8", 11552 => x"5b8b0008",
    11553 => x"5b9d0004", 11554 => x"780b0001", 11555 => x"396b6dbc",
    11556 => x"29610000", 11557 => x"28220004", 11558 => x"38420010",
    11559 => x"58220004", 11560 => x"34010001", 11561 => x"f8000482",
    11562 => x"29610000", 11563 => x"28210004", 11564 => x"20210020",
    11565 => x"7c210000", 11566 => x"2b9d0004", 11567 => x"2b8b0008",
    11568 => x"379c0008", 11569 => x"c3a00000", 11570 => x"379cfff8",
    11571 => x"5b8b0008", 11572 => x"5b9d0004", 11573 => x"b8205800",
    11574 => x"34010044", 11575 => x"fbffff17", 11576 => x"38220020",
    11577 => x"45600003", 11578 => x"3402ffdf", 11579 => x"a0221000",
    11580 => x"34010044", 11581 => x"fbffff1d", 11582 => x"34010000",
    11583 => x"2b9d0004", 11584 => x"2b8b0008", 11585 => x"379c0008",
    11586 => x"c3a00000", 11587 => x"379cfff8", 11588 => x"5b8b0008",
    11589 => x"5b9d0004", 11590 => x"78020001", 11591 => x"38426d00",
    11592 => x"28420000", 11593 => x"780b0001", 11594 => x"396b6dbc",
    11595 => x"59620000", 11596 => x"fbffff1c", 11597 => x"34010001",
    11598 => x"fbffffe4", 11599 => x"78020001", 11600 => x"38423d00",
    11601 => x"28410000", 11602 => x"78040001", 11603 => x"38843d04",
    11604 => x"58200000", 11605 => x"29610000", 11606 => x"28830000",
    11607 => x"34020003", 11608 => x"58200000", 11609 => x"5822000c",
    11610 => x"58230008", 11611 => x"78030001", 11612 => x"38633d08",
    11613 => x"58220004", 11614 => x"28620000", 11615 => x"5822003c",
    11616 => x"2b9d0004", 11617 => x"2b8b0008", 11618 => x"379c0008",
    11619 => x"c3a00000", 11620 => x"379cfffc", 11621 => x"5b9d0004",
    11622 => x"78010001", 11623 => x"78040001", 11624 => x"38214abc",
    11625 => x"38843d0c", 11626 => x"28220000", 11627 => x"28830000",
    11628 => x"44430012", 11629 => x"78030001", 11630 => x"38634ba0",
    11631 => x"780500ff", 11632 => x"e000000d", 11633 => x"28240000",
    11634 => x"3c870018", 11635 => x"00860018", 11636 => x"b8e63000",
    11637 => x"a0853800", 11638 => x"00e70008", 11639 => x"2084ff00",
    11640 => x"3c840008", 11641 => x"b8c73000", 11642 => x"b8c42000",
    11643 => x"58240000", 11644 => x"34210004", 11645 => x"5461fff4",
    11646 => x"78010001", 11647 => x"78050001", 11648 => x"38214abc",
    11649 => x"38a53d0c", 11650 => x"28240000", 11651 => x"28a30000",
    11652 => x"44830005", 11653 => x"78010001", 11654 => x"38213574",
    11655 => x"fbfffded", 11656 => x"e000004f", 11657 => x"78020001",
    11658 => x"38425e04", 11659 => x"28430000", 11660 => x"5c600016",
    11661 => x"2824000c", 11662 => x"34031234", 11663 => x"0084000d",
    11664 => x"2084ffff", 11665 => x"5c83000b", 11666 => x"28240014",
    11667 => x"34035678", 11668 => x"0084000d", 11669 => x"2084ffff",
    11670 => x"5c830006", 11671 => x"2823001c", 11672 => x"38019abc",
    11673 => x"0063000d", 11674 => x"2063ffff", 11675 => x"44610005",
    11676 => x"78010001", 11677 => x"3821359c", 11678 => x"fbfffdd6",
    11679 => x"e0000038", 11680 => x"34010001", 11681 => x"58410000",
    11682 => x"78020001", 11683 => x"38423d10", 11684 => x"28430000",
    11685 => x"78020001", 11686 => x"38426dbc", 11687 => x"28420000",
    11688 => x"78010001", 11689 => x"38214abc", 11690 => x"28460024",
    11691 => x"28250014", 11692 => x"2824001c", 11693 => x"2827000c",
    11694 => x"20c6ffff", 11695 => x"3cc6000d", 11696 => x"a0832000",
    11697 => x"a0a32800", 11698 => x"a0e31800", 11699 => x"b8c31800",
    11700 => x"5823000c", 11701 => x"28430028", 11702 => x"00630010",
    11703 => x"3c63000d", 11704 => x"b8651800", 11705 => x"58230014",
    11706 => x"28430028", 11707 => x"2063ffff", 11708 => x"3c63000d",
    11709 => x"b8641800", 11710 => x"5823001c", 11711 => x"78010001",
    11712 => x"78030001", 11713 => x"58400014", 11714 => x"34040000",
    11715 => x"38214ac0", 11716 => x"38634ba0", 11717 => x"e000000f",
    11718 => x"28250000", 11719 => x"28270004", 11720 => x"34210008",
    11721 => x"20a60fff", 11722 => x"3ce70014", 11723 => x"00a5000c",
    11724 => x"58460018", 11725 => x"b8e52800", 11726 => x"3ca50008",
    11727 => x"2087003f", 11728 => x"38a50040", 11729 => x"b8a72800",
    11730 => x"58450014", 11731 => x"34840001", 11732 => x"5461fff2",
    11733 => x"34010080", 11734 => x"58410014", 11735 => x"2b9d0004",
    11736 => x"379c0004", 11737 => x"c3a00000", 11738 => x"78030001",
    11739 => x"38636db8", 11740 => x"44400004", 11741 => x"28620000",
    11742 => x"58410004", 11743 => x"c3a00000", 11744 => x"28620000",
    11745 => x"58410008", 11746 => x"c3a00000", 11747 => x"78030001",
    11748 => x"38636db8", 11749 => x"44400004", 11750 => x"28620000",
    11751 => x"58410004", 11752 => x"c3a00000", 11753 => x"28620000",
    11754 => x"58410008", 11755 => x"c3a00000", 11756 => x"3401012c",
    11757 => x"34000000", 11758 => x"3421ffff", 11759 => x"5c20fffe",
    11760 => x"c3a00000", 11761 => x"379cfff8", 11762 => x"5b8b0008",
    11763 => x"5b9d0004", 11764 => x"202100ff", 11765 => x"3c2b0003",
    11766 => x"78020001", 11767 => x"38424ba0", 11768 => x"b44b5800",
    11769 => x"29610004", 11770 => x"34020000", 11771 => x"fbffffdf",
    11772 => x"fbfffff0", 11773 => x"29610000", 11774 => x"34020000",
    11775 => x"fbffffdb", 11776 => x"fbffffec", 11777 => x"2b9d0004",
    11778 => x"2b8b0008", 11779 => x"379c0008", 11780 => x"c3a00000",
    11781 => x"379cfff8", 11782 => x"5b8b0008", 11783 => x"5b9d0004",
    11784 => x"202100ff", 11785 => x"3c2b0003", 11786 => x"78020001",
    11787 => x"38424ba0", 11788 => x"b44b5800", 11789 => x"29610004",
    11790 => x"34020001", 11791 => x"fbffffcb", 11792 => x"fbffffdc",
    11793 => x"29610000", 11794 => x"34020001", 11795 => x"fbffffc7",
    11796 => x"fbffffd8", 11797 => x"29610004", 11798 => x"34020000",
    11799 => x"fbffffc3", 11800 => x"fbffffd4", 11801 => x"29610000",
    11802 => x"34020000", 11803 => x"fbffffbf", 11804 => x"fbffffd0",
    11805 => x"2b9d0004", 11806 => x"2b8b0008", 11807 => x"379c0008",
    11808 => x"c3a00000", 11809 => x"379cfff8", 11810 => x"5b8b0008",
    11811 => x"5b9d0004", 11812 => x"202100ff", 11813 => x"3c2b0003",
    11814 => x"78020001", 11815 => x"38424ba0", 11816 => x"b44b5800",
    11817 => x"29610004", 11818 => x"34020000", 11819 => x"fbffffaf",
    11820 => x"fbffffc0", 11821 => x"29610000", 11822 => x"34020001",
    11823 => x"fbffffab", 11824 => x"fbffffbc", 11825 => x"29610004",
    11826 => x"34020001", 11827 => x"fbffffa7", 11828 => x"fbffffb8",
    11829 => x"2b9d0004", 11830 => x"2b8b0008", 11831 => x"379c0008",
    11832 => x"c3a00000", 11833 => x"379cffec", 11834 => x"5b8b0014",
    11835 => x"5b8c0010", 11836 => x"5b8d000c", 11837 => x"5b8e0008",
    11838 => x"5b9d0004", 11839 => x"202100ff", 11840 => x"78030001",
    11841 => x"3c2b0003", 11842 => x"38634ba0", 11843 => x"204e00ff",
    11844 => x"340d0008", 11845 => x"b46b5800", 11846 => x"29610004",
    11847 => x"21c20080", 11848 => x"35adffff", 11849 => x"fbffff91",
    11850 => x"fbffffa2", 11851 => x"29610000", 11852 => x"34020001",
    11853 => x"3dce0001", 11854 => x"fbffff8c", 11855 => x"fbffff9d",
    11856 => x"29610000", 11857 => x"34020000", 11858 => x"21ad00ff",
    11859 => x"fbffff87", 11860 => x"356c0004", 11861 => x"fbffff97",
    11862 => x"21ce00ff", 11863 => x"5da0ffef", 11864 => x"29810000",
    11865 => x"34020001", 11866 => x"fbffff80", 11867 => x"fbffff91",
    11868 => x"29610000", 11869 => x"34020001", 11870 => x"fbffff7c",
    11871 => x"fbffff8d", 11872 => x"78010001", 11873 => x"38216db8",
    11874 => x"28210000", 11875 => x"298d0000", 11876 => x"34020000",
    11877 => x"28210004", 11878 => x"a02d6800", 11879 => x"29610000",
    11880 => x"fbffff72", 11881 => x"fbffff83", 11882 => x"29810000",
    11883 => x"34020000", 11884 => x"fbffff6e", 11885 => x"fbffff7f",
    11886 => x"7da10000", 11887 => x"2b9d0004", 11888 => x"2b8b0014",
    11889 => x"2b8c0010", 11890 => x"2b8d000c", 11891 => x"2b8e0008",
    11892 => x"379c0014", 11893 => x"c3a00000", 11894 => x"379cffe0",
    11895 => x"5b8b0020", 11896 => x"5b8c001c", 11897 => x"5b8d0018",
    11898 => x"5b8e0014", 11899 => x"5b8f0010", 11900 => x"5b90000c",
    11901 => x"5b910008", 11902 => x"5b9d0004", 11903 => x"202100ff",
    11904 => x"3c2b0003", 11905 => x"78040001", 11906 => x"38844ba0",
    11907 => x"b48b5800", 11908 => x"29610004", 11909 => x"b8407800",
    11910 => x"34020001", 11911 => x"207000ff", 11912 => x"fbffff52",
    11913 => x"fbffff63", 11914 => x"29610000", 11915 => x"34020000",
    11916 => x"780d0001", 11917 => x"fbffff4d", 11918 => x"340c0000",
    11919 => x"fbffff5d", 11920 => x"340e0000", 11921 => x"39ad6db8",
    11922 => x"34110008", 11923 => x"29610000", 11924 => x"34020001",
    11925 => x"3d8c0001", 11926 => x"fbffff44", 11927 => x"fbffff55",
    11928 => x"29a10000", 11929 => x"29620004", 11930 => x"218c00ff",
    11931 => x"28210004", 11932 => x"a0220800", 11933 => x"44200002",
    11934 => x"398c0001", 11935 => x"29610000", 11936 => x"34020000",
    11937 => x"35ce0001", 11938 => x"fbffff38", 11939 => x"fbffff49",
    11940 => x"5dd1ffef", 11941 => x"46000004", 11942 => x"29610004",
    11943 => x"34020001", 11944 => x"e0000003", 11945 => x"29610004",
    11946 => x"34020000", 11947 => x"fbffff2f", 11948 => x"fbffff40",
    11949 => x"29610000", 11950 => x"34020001", 11951 => x"fbffff2b",
    11952 => x"fbffff3c", 11953 => x"29610000", 11954 => x"34020000",
    11955 => x"fbffff27", 11956 => x"fbffff38", 11957 => x"31ec0000",
    11958 => x"2b9d0004", 11959 => x"2b8b0020", 11960 => x"2b8c001c",
    11961 => x"2b8d0018", 11962 => x"2b8e0014", 11963 => x"2b8f0010",
    11964 => x"2b90000c", 11965 => x"2b910008", 11966 => x"379c0020",
    11967 => x"c3a00000", 11968 => x"379cfff8", 11969 => x"5b8b0008",
    11970 => x"5b9d0004", 11971 => x"202100ff", 11972 => x"3c2b0003",
    11973 => x"78020001", 11974 => x"38424ba0", 11975 => x"b44b5800",
    11976 => x"29610000", 11977 => x"34020001", 11978 => x"fbffff10",
    11979 => x"fbffff21", 11980 => x"29610004", 11981 => x"34020001",
    11982 => x"fbffff0c", 11983 => x"fbffff1d", 11984 => x"2b9d0004",
    11985 => x"2b8b0008", 11986 => x"379c0008", 11987 => x"c3a00000",
    11988 => x"379cfff4", 11989 => x"5b8b000c", 11990 => x"5b8c0008",
    11991 => x"5b9d0004", 11992 => x"202b00ff", 11993 => x"b9600800",
    11994 => x"204c00ff", 11995 => x"fbffff16", 11996 => x"3d820001",
    11997 => x"b9600800", 11998 => x"204200fe", 11999 => x"fbffff5a",
    12000 => x"b8206000", 12001 => x"b9600800", 12002 => x"fbffff3f",
    12003 => x"65810000", 12004 => x"2b9d0004", 12005 => x"2b8b000c",
    12006 => x"2b8c0008", 12007 => x"379c000c", 12008 => x"c3a00000",
    12009 => x"379cffe8", 12010 => x"5b8b0018", 12011 => x"5b8c0014",
    12012 => x"5b8d0010", 12013 => x"5b8e000c", 12014 => x"5b8f0008",
    12015 => x"5b9d0004", 12016 => x"780b0001", 12017 => x"396b5e08",
    12018 => x"296d000c", 12019 => x"296f0004", 12020 => x"b8206000",
    12021 => x"3dad0002", 12022 => x"c84f0800", 12023 => x"b9a01000",
    12024 => x"b8607000", 12025 => x"f8001502", 12026 => x"b42f1000",
    12027 => x"b5af6800", 12028 => x"b44e0800", 12029 => x"542d0006",
    12030 => x"b9800800", 12031 => x"b9c01800", 12032 => x"f800154c",
    12033 => x"b8206000", 12034 => x"e0000009", 12035 => x"c9a26800",
    12036 => x"b9a01800", 12037 => x"b9800800", 12038 => x"f8001546",
    12039 => x"29620004", 12040 => x"b58d0800", 12041 => x"c9cd1800",
    12042 => x"f8001542", 12043 => x"b9800800", 12044 => x"2b9d0004",
    12045 => x"2b8b0018", 12046 => x"2b8c0014", 12047 => x"2b8d0010",
    12048 => x"2b8e000c", 12049 => x"2b8f0008", 12050 => x"379c0018",
    12051 => x"c3a00000", 12052 => x"379cffe8", 12053 => x"5b8b0018",
    12054 => x"5b8c0014", 12055 => x"5b8d0010", 12056 => x"5b8e000c",
    12057 => x"5b8f0008", 12058 => x"5b9d0004", 12059 => x"780b0001",
    12060 => x"396b5e08", 12061 => x"296f000c", 12062 => x"296e0004",
    12063 => x"b8406800", 12064 => x"3def0002", 12065 => x"c82e0800",
    12066 => x"b9e01000", 12067 => x"f80014d8", 12068 => x"b42e6000",
    12069 => x"b58d0800", 12070 => x"b5ee7000", 12071 => x"542e0006",
    12072 => x"b9800800", 12073 => x"34020000", 12074 => x"b9a01800",
    12075 => x"f800159f", 12076 => x"e000000b", 12077 => x"c9cc7000",
    12078 => x"34020000", 12079 => x"b9c01800", 12080 => x"b9800800",
    12081 => x"f8001599", 12082 => x"29610004", 12083 => x"34020000",
    12084 => x"c9ae1800", 12085 => x"f8001595", 12086 => x"b9800800",
    12087 => x"2b9d0004", 12088 => x"2b8b0018", 12089 => x"2b8c0014",
    12090 => x"2b8d0010", 12091 => x"2b8e000c", 12092 => x"2b8f0008",
    12093 => x"379c0018", 12094 => x"c3a00000", 12095 => x"379cfff4",
    12096 => x"5b8b000c", 12097 => x"5b8c0008", 12098 => x"5b9d0004",
    12099 => x"780c0001", 12100 => x"398c6dcc", 12101 => x"29810000",
    12102 => x"780b0001", 12103 => x"396b5e08", 12104 => x"58200000",
    12105 => x"34020200", 12106 => x"78010001", 12107 => x"38216230",
    12108 => x"5962000c", 12109 => x"34020800", 12110 => x"59610004",
    12111 => x"59610000", 12112 => x"fbffffc4", 12113 => x"29620004",
    12114 => x"29810000", 12115 => x"58220008", 12116 => x"2962000c",
    12117 => x"5822000c", 12118 => x"34020002", 12119 => x"5822004c",
    12120 => x"34020400", 12121 => x"58220000", 12122 => x"2b9d0004",
    12123 => x"2b8b000c", 12124 => x"2b8c0008", 12125 => x"379c000c",
    12126 => x"c3a00000", 12127 => x"379cfff4", 12128 => x"5b8b000c",
    12129 => x"5b8c0008", 12130 => x"5b9d0004", 12131 => x"780b0001",
    12132 => x"396b6dcc", 12133 => x"29630000", 12134 => x"340c0002",
    12135 => x"78010001", 12136 => x"586c0040", 12137 => x"78020001",
    12138 => x"586c004c", 12139 => x"38215e08", 12140 => x"38426230",
    12141 => x"58220004", 12142 => x"00420002", 12143 => x"34040800",
    12144 => x"5824000c", 12145 => x"344401ff", 12146 => x"3c840010",
    12147 => x"2042ffff", 12148 => x"b8821000", 12149 => x"58620020",
    12150 => x"78020001", 12151 => x"38425e30", 12152 => x"58220014",
    12153 => x"34020100", 12154 => x"5822001c", 12155 => x"58200020",
    12156 => x"58200024", 12157 => x"fbffffc2", 12158 => x"29610000",
    12159 => x"582c0044", 12160 => x"2b9d0004", 12161 => x"2b8b000c",
    12162 => x"2b8c0008", 12163 => x"379c000c", 12164 => x"c3a00000",
    12165 => x"379cffc4", 12166 => x"5b8b0028", 12167 => x"5b8c0024",
    12168 => x"5b8d0020", 12169 => x"5b8e001c", 12170 => x"5b8f0018",
    12171 => x"5b900014", 12172 => x"5b910010", 12173 => x"5b92000c",
    12174 => x"5b930008", 12175 => x"5b9d0004", 12176 => x"b8805800",
    12177 => x"78040001", 12178 => x"38846dcc", 12179 => x"28840000",
    12180 => x"b8209000", 12181 => x"b8408800", 12182 => x"2881004c",
    12183 => x"b8608000", 12184 => x"340c0000", 12185 => x"20210002",
    12186 => x"4420008a", 12187 => x"780e0001", 12188 => x"39ce5e08",
    12189 => x"29c20000", 12190 => x"28430000", 12191 => x"48030009",
    12192 => x"28810000", 12193 => x"20210200", 12194 => x"5c200004",
    12195 => x"78010001", 12196 => x"382135c4", 12197 => x"fbfffbcf",
    12198 => x"fbffff99", 12199 => x"e000007d", 12200 => x"20610001",
    12201 => x"206d0ffe", 12202 => x"c9a16800", 12203 => x"35af0003",
    12204 => x"01ef0002", 12205 => x"78044000", 12206 => x"a0642000",
    12207 => x"35ef0001", 12208 => x"340cffff", 12209 => x"5c800054",
    12210 => x"7d610000", 12211 => x"0063001d", 12212 => x"a0611800",
    12213 => x"4464003e", 12214 => x"b44d1000", 12215 => x"34030004",
    12216 => x"37810038", 12217 => x"fbffff30", 12218 => x"29c30000",
    12219 => x"35b3fffa", 12220 => x"35adfffe", 12221 => x"b46d1000",
    12222 => x"3781003e", 12223 => x"34030002", 12224 => x"fbffff29",
    12225 => x"78010001", 12226 => x"38213d14", 12227 => x"282c0000",
    12228 => x"37820034", 12229 => x"3781002c", 12230 => x"2b8d0038",
    12231 => x"f8000191", 12232 => x"78020001", 12233 => x"38423d18",
    12234 => x"28410000", 12235 => x"a1ac6000", 12236 => x"01ad001c",
    12237 => x"502c000e", 12238 => x"78030001", 12239 => x"38633d1c",
    12240 => x"2b820034", 12241 => x"28610000", 12242 => x"54410009",
    12243 => x"2b820030", 12244 => x"2b81002c", 12245 => x"3444ffff",
    12246 => x"f4441000", 12247 => x"3421ffff", 12248 => x"b4410800",
    12249 => x"5b81002c", 12250 => x"5b840030", 12251 => x"78020001",
    12252 => x"38423d20", 12253 => x"28410000", 12254 => x"2b820030",
    12255 => x"2183000f", 12256 => x"c86d1800", 12257 => x"a0410800",
    12258 => x"5961000c", 12259 => x"6461fff1", 12260 => x"64630001",
    12261 => x"59600008", 12262 => x"b8231800", 12263 => x"44600004",
    12264 => x"34010001", 12265 => x"59610004", 12266 => x"e0000002",
    12267 => x"59600004", 12268 => x"2f81003e", 12269 => x"3d8c0003",
    12270 => x"ba606800", 12271 => x"20210800", 12272 => x"64210000",
    12273 => x"596c0010", 12274 => x"31610000", 12275 => x"b9a06000",
    12276 => x"520d0002", 12277 => x"ba006000", 12278 => x"780b0001",
    12279 => x"396b5e08", 12280 => x"29610024", 12281 => x"29620000",
    12282 => x"3403000e", 12283 => x"34210001", 12284 => x"59610024",
    12285 => x"34420004", 12286 => x"ba400800", 12287 => x"fbfffeea",
    12288 => x"29630000", 12289 => x"ba200800", 12290 => x"34620012",
    12291 => x"3583fff2", 12292 => x"fbfffee5", 12293 => x"780b0001",
    12294 => x"396b5e08", 12295 => x"3dee0002", 12296 => x"29610000",
    12297 => x"b9c01000", 12298 => x"fbffff0a", 12299 => x"78030001",
    12300 => x"38636dcc", 12301 => x"286d0000", 12302 => x"29610000",
    12303 => x"59af0010", 12304 => x"2962000c", 12305 => x"296f0004",
    12306 => x"3c420002", 12307 => x"c82f0800", 12308 => x"b42e0800",
    12309 => x"f80013e6", 12310 => x"b42f0800", 12311 => x"59610000",
    12312 => x"29a20010", 12313 => x"28210000", 12314 => x"4801000a",
    12315 => x"29a10000", 12316 => x"20210200", 12317 => x"44200002",
    12318 => x"fbffff21", 12319 => x"78010001", 12320 => x"38216dcc",
    12321 => x"28210000", 12322 => x"34020002", 12323 => x"5822004c",
    12324 => x"b9800800", 12325 => x"2b9d0004", 12326 => x"2b8b0028",
    12327 => x"2b8c0024", 12328 => x"2b8d0020", 12329 => x"2b8e001c",
    12330 => x"2b8f0018", 12331 => x"2b900014", 12332 => x"2b910010",
    12333 => x"2b92000c", 12334 => x"2b930008", 12335 => x"379c003c",
    12336 => x"c3a00000", 12337 => x"379cffd8", 12338 => x"5b8b001c",
    12339 => x"5b8c0018", 12340 => x"5b8d0014", 12341 => x"5b8e0010",
    12342 => x"5b8f000c", 12343 => x"5b900008", 12344 => x"5b9d0004",
    12345 => x"780d0001", 12346 => x"39ad5e08", 12347 => x"b8605800",
    12348 => x"34030100", 12349 => x"59a3001c", 12350 => x"59a30018",
    12351 => x"78030001", 12352 => x"38636dcc", 12353 => x"b8207800",
    12354 => x"b8407000", 12355 => x"78010001", 12356 => x"28620000",
    12357 => x"38215e30", 12358 => x"59a10014", 12359 => x"59a10010",
    12360 => x"58410004", 12361 => x"35630010", 12362 => x"34020000",
    12363 => x"b8806000", 12364 => x"f800147e", 12365 => x"29a10010",
    12366 => x"3402003c", 12367 => x"b9601800", 12368 => x"34210004",
    12369 => x"51620002", 12370 => x"3403003c", 12371 => x"34020000",
    12372 => x"780d0001", 12373 => x"f8001475", 12374 => x"39ad5e08",
    12375 => x"29a10010", 12376 => x"b9e01000", 12377 => x"3403000e",
    12378 => x"34210004", 12379 => x"f80013f1", 12380 => x"29a10010",
    12381 => x"b9c01000", 12382 => x"3563fff2", 12383 => x"34210012",
    12384 => x"f80013ec", 12385 => x"3401003b", 12386 => x"502b0002",
    12387 => x"e0000002", 12388 => x"340b003c", 12389 => x"35630001",
    12390 => x"7d810000", 12391 => x"00630001", 12392 => x"3c21001e",
    12393 => x"78048000", 12394 => x"b8642000", 12395 => x"b8812000",
    12396 => x"78010001", 12397 => x"38215e08", 12398 => x"28220010",
    12399 => x"3c630002", 12400 => x"78010001", 12401 => x"58440000",
    12402 => x"38216dcc", 12403 => x"b4431000", 12404 => x"58400000",
    12405 => x"28220000", 12406 => x"340d0000", 12407 => x"b8207800",
    12408 => x"28430000", 12409 => x"341003e8", 12410 => x"38630001",
    12411 => x"58430000", 12412 => x"29e10000", 12413 => x"282e0000",
    12414 => x"21c10002", 12415 => x"5c200009", 12416 => x"34010001",
    12417 => x"35ad0001", 12418 => x"f8000129", 12419 => x"5db0fff9",
    12420 => x"78010001", 12421 => x"382135e4", 12422 => x"b9c01000",
    12423 => x"fbfffaed", 12424 => x"45800046", 12425 => x"780d0001",
    12426 => x"340e0000", 12427 => x"39ad6dcc", 12428 => x"340f0064",
    12429 => x"29a10000", 12430 => x"28220000", 12431 => x"20420800",
    12432 => x"5c40000a", 12433 => x"34010001", 12434 => x"35ce0001",
    12435 => x"f8000118", 12436 => x"5dcffff9", 12437 => x"78010001",
    12438 => x"38213614", 12439 => x"fbfffadd", 12440 => x"340e0000",
    12441 => x"e0000003", 12442 => x"282e0014", 12443 => x"21ce0001",
    12444 => x"78010001", 12445 => x"38216dcc", 12446 => x"28210000",
    12447 => x"282d0018", 12448 => x"28230014", 12449 => x"00630006",
    12450 => x"2063ffff", 12451 => x"44600006", 12452 => x"78020001",
    12453 => x"34010000", 12454 => x"38423644", 12455 => x"34040000",
    12456 => x"fbffcfdd", 12457 => x"78020001", 12458 => x"38423d14",
    12459 => x"28410000", 12460 => x"37820028", 12461 => x"a1a16800",
    12462 => x"37810020", 12463 => x"f80000a9", 12464 => x"78030001",
    12465 => x"38633d18", 12466 => x"28610000", 12467 => x"502d000e",
    12468 => x"78030001", 12469 => x"38633d1c", 12470 => x"2b820028",
    12471 => x"28610000", 12472 => x"54410009", 12473 => x"2b830024",
    12474 => x"2b820020", 12475 => x"3461ffff", 12476 => x"f4611800",
    12477 => x"3442ffff", 12478 => x"b4621000", 12479 => x"5b820020",
    12480 => x"5b810024", 12481 => x"2b810020", 12482 => x"318e0000",
    12483 => x"3dad0003", 12484 => x"59810008", 12485 => x"2b810024",
    12486 => x"59800004", 12487 => x"598d0010", 12488 => x"5981000c",
    12489 => x"78010001", 12490 => x"38215e08", 12491 => x"28220020",
    12492 => x"34420001", 12493 => x"58220020", 12494 => x"b9600800",
    12495 => x"2b9d0004", 12496 => x"2b8b001c", 12497 => x"2b8c0018",
    12498 => x"2b8d0014", 12499 => x"2b8e0010", 12500 => x"2b8f000c",
    12501 => x"2b900008", 12502 => x"379c0028", 12503 => x"c3a00000",
    12504 => x"78030001", 12505 => x"38635e08", 12506 => x"28640020",
    12507 => x"58240000", 12508 => x"28610024", 12509 => x"58410000",
    12510 => x"c3a00000", 12511 => x"78010001", 12512 => x"38216d10",
    12513 => x"28210000", 12514 => x"28220008", 12515 => x"2821000c",
    12516 => x"202100ff", 12517 => x"c3a00000", 12518 => x"78010001",
    12519 => x"78030001", 12520 => x"38633d24", 12521 => x"38216d10",
    12522 => x"28210000", 12523 => x"28620000", 12524 => x"78040001",
    12525 => x"38843d28", 12526 => x"58220000", 12527 => x"58200014",
    12528 => x"28830000", 12529 => x"58200018", 12530 => x"58200010",
    12531 => x"58230000", 12532 => x"58220000", 12533 => x"5820001c",
    12534 => x"c3a00000", 12535 => x"379cffe8", 12536 => x"5b8b0018",
    12537 => x"5b8c0014", 12538 => x"5b8d0010", 12539 => x"5b8e000c",
    12540 => x"5b8f0008", 12541 => x"5b9d0004", 12542 => x"780b0001",
    12543 => x"b8207800", 12544 => x"34010001", 12545 => x"b8406800",
    12546 => x"b8607000", 12547 => x"396b366c", 12548 => x"5de10003",
    12549 => x"780b0001", 12550 => x"396b3670", 12551 => x"15ac001f",
    12552 => x"b9c00800", 12553 => x"f800131e", 12554 => x"218c0002",
    12555 => x"358c002b", 12556 => x"78020001", 12557 => x"b8202800",
    12558 => x"38423678", 12559 => x"34010000", 12560 => x"b9601800",
    12561 => x"b9802000", 12562 => x"fbffcf73", 12563 => x"78020001",
    12564 => x"34010002", 12565 => x"38426d10", 12566 => x"5de1000e",
    12567 => x"28410000", 12568 => x"15a2001f", 12569 => x"20420007",
    12570 => x"b44e7000", 12571 => x"f44e1000", 12572 => x"01ce0003",
    12573 => x"b44d6800", 12574 => x"3dad001d", 12575 => x"58200014",
    12576 => x"58200018", 12577 => x"b9ae7000", 12578 => x"582e0010",
    12579 => x"e0000006", 12580 => x"28420000", 12581 => x"21ad00ff",
    12582 => x"584e0014", 12583 => x"584d0018", 12584 => x"58400010",
    12585 => x"78010001", 12586 => x"38216d10", 12587 => x"28210000",
    12588 => x"28220000", 12589 => x"38420004", 12590 => x"58220000",
    12591 => x"34010000", 12592 => x"2b9d0004", 12593 => x"2b8b0018",
    12594 => x"2b8c0014", 12595 => x"2b8d0010", 12596 => x"2b8e000c",
    12597 => x"2b8f0008", 12598 => x"379c0018", 12599 => x"c3a00000",
    12600 => x"78050001", 12601 => x"38a56d10", 12602 => x"28a50000",
    12603 => x"202100ff", 12604 => x"00630003", 12605 => x"58a20014",
    12606 => x"58a10018", 12607 => x"58a30010", 12608 => x"34010003",
    12609 => x"5c810007", 12610 => x"28a20000", 12611 => x"3401fff3",
    12612 => x"a0410800", 12613 => x"38210008", 12614 => x"58a10000",
    12615 => x"c3a00000", 12616 => x"34010001", 12617 => x"5c810007",
    12618 => x"28a2001c", 12619 => x"3401ffe7", 12620 => x"a0410800",
    12621 => x"38210008", 12622 => x"58a1001c", 12623 => x"c3a00000",
    12624 => x"34010002", 12625 => x"5c810006", 12626 => x"28a2001c",
    12627 => x"3401ffe7", 12628 => x"a0410800", 12629 => x"38210010",
    12630 => x"58a1001c", 12631 => x"c3a00000", 12632 => x"379cffe0",
    12633 => x"5b8b0020", 12634 => x"5b8c001c", 12635 => x"5b8d0018",
    12636 => x"5b8e0014", 12637 => x"5b8f0010", 12638 => x"5b90000c",
    12639 => x"5b910008", 12640 => x"5b9d0004", 12641 => x"b8206000",
    12642 => x"78010001", 12643 => x"38213d14", 12644 => x"282f0000",
    12645 => x"780b0001", 12646 => x"b8406800", 12647 => x"396b6d10",
    12648 => x"fbffff77", 12649 => x"b8208800", 12650 => x"29610000",
    12651 => x"b8408000", 12652 => x"282e0004", 12653 => x"a1cf7000",
    12654 => x"fbffff71", 12655 => x"5c31fff9", 12656 => x"5c50fff8",
    12657 => x"45800003", 12658 => x"59810000", 12659 => x"59820004",
    12660 => x"45a00003", 12661 => x"3dc10003", 12662 => x"59a10000",
    12663 => x"2b9d0004", 12664 => x"2b8b0020", 12665 => x"2b8c001c",
    12666 => x"2b8d0018", 12667 => x"2b8e0014", 12668 => x"2b8f0010",
    12669 => x"2b90000c", 12670 => x"2b910008", 12671 => x"379c0020",
    12672 => x"c3a00000", 12673 => x"78010001", 12674 => x"38216d10",
    12675 => x"28210000", 12676 => x"28210000", 12677 => x"20210004",
    12678 => x"64210000", 12679 => x"c3a00000", 12680 => x"78020001",
    12681 => x"38426d10", 12682 => x"28420000", 12683 => x"2843001c",
    12684 => x"44200003", 12685 => x"38630006", 12686 => x"e0000003",
    12687 => x"3401fff9", 12688 => x"a0611800", 12689 => x"5843001c",
    12690 => x"34010000", 12691 => x"c3a00000", 12692 => x"78020001",
    12693 => x"38426dd0", 12694 => x"28420000", 12695 => x"78030001",
    12696 => x"38636db8", 12697 => x"58620000", 12698 => x"44200005",
    12699 => x"28430010", 12700 => x"78018000", 12701 => x"b8610800",
    12702 => x"e0000006", 12703 => x"78040001", 12704 => x"38843d20",
    12705 => x"28430010", 12706 => x"28810000", 12707 => x"a0610800",
    12708 => x"58410010", 12709 => x"c3a00000", 12710 => x"78010001",
    12711 => x"38216db8", 12712 => x"28210000", 12713 => x"28210014",
    12714 => x"c3a00000", 12715 => x"78020001", 12716 => x"38426db8",
    12717 => x"28420000", 12718 => x"28430014", 12719 => x"b4230800",
    12720 => x"28430014", 12721 => x"c8611800", 12722 => x"4803fffe",
    12723 => x"c3a00000", 12724 => x"78010001", 12725 => x"38216db8",
    12726 => x"28210000", 12727 => x"28210004", 12728 => x"20210080",
    12729 => x"64210000", 12730 => x"c3a00000", 12731 => x"379cffe0",
    12732 => x"5b8b001c", 12733 => x"5b8c0018", 12734 => x"5b8d0014",
    12735 => x"5b8e0010", 12736 => x"5b8f000c", 12737 => x"5b900008",
    12738 => x"5b9d0004", 12739 => x"b8208000", 12740 => x"34010001",
    12741 => x"fbfffcfb", 12742 => x"34010001", 12743 => x"fbfffc2a",
    12744 => x"340200a0", 12745 => x"34010001", 12746 => x"fbfffc6f",
    12747 => x"34020000", 12748 => x"34010001", 12749 => x"fbfffc6c",
    12750 => x"34010001", 12751 => x"fbfffc36", 12752 => x"340200a1",
    12753 => x"34010001", 12754 => x"fbfffc67", 12755 => x"378d0023",
    12756 => x"b9a01000", 12757 => x"34030001", 12758 => x"34010001",
    12759 => x"fbfffc9f", 12760 => x"34010001", 12761 => x"fbfffc48",
    12762 => x"34010001", 12763 => x"438c0023", 12764 => x"fbfffc15",
    12765 => x"34010001", 12766 => x"340200a1", 12767 => x"fbfffc5a",
    12768 => x"340bffd9", 12769 => x"340f000f", 12770 => x"340e0017",
    12771 => x"34030000", 12772 => x"34010001", 12773 => x"b9a01000",
    12774 => x"fbfffc90", 12775 => x"43830023", 12776 => x"b5836000",
    12777 => x"218c00ff", 12778 => x"556f0003", 12779 => x"b60b0800",
    12780 => x"30230000", 12781 => x"356b0001", 12782 => x"5d6efff5",
    12783 => x"37820023", 12784 => x"34030001", 12785 => x"34010001",
    12786 => x"fbfffc84", 12787 => x"34010001", 12788 => x"fbfffc2d",
    12789 => x"43810023", 12790 => x"fc2c6000", 12791 => x"c80c0800",
    12792 => x"2b9d0004", 12793 => x"2b8b001c", 12794 => x"2b8c0018",
    12795 => x"2b8d0014", 12796 => x"2b8e0010", 12797 => x"2b8f000c",
    12798 => x"2b900008", 12799 => x"379c0020", 12800 => x"c3a00000",
    12801 => x"379cffe0", 12802 => x"5b9b0008", 12803 => x"341b0020",
    12804 => x"b77cd800", 12805 => x"5b8b0020", 12806 => x"5b8c001c",
    12807 => x"5b8d0018", 12808 => x"5b8e0014", 12809 => x"5b8f0010",
    12810 => x"5b90000c", 12811 => x"5b9d0004", 12812 => x"780b0001",
    12813 => x"780c0001", 12814 => x"bb807800", 12815 => x"34020001",
    12816 => x"396b4c88", 12817 => x"398c3698", 12818 => x"e0000012",
    12819 => x"bb808000", 12820 => x"379cffe4", 12821 => x"378e000b",
    12822 => x"01ce0003", 12823 => x"35a2002c", 12824 => x"3dce0003",
    12825 => x"34030014", 12826 => x"b9c00800", 12827 => x"f8001231",
    12828 => x"31c00013", 12829 => x"29a20020", 12830 => x"29630074",
    12831 => x"b9800800", 12832 => x"b9c02000", 12833 => x"fbfff953",
    12834 => x"34020000", 12835 => x"ba00e000", 12836 => x"b9600800",
    12837 => x"f8001090", 12838 => x"b8206800", 12839 => x"5c20ffec",
    12840 => x"b9e0e000", 12841 => x"2b9d0004", 12842 => x"2b8b0020",
    12843 => x"2b8c001c", 12844 => x"2b8d0018", 12845 => x"2b8e0014",
    12846 => x"2b8f0010", 12847 => x"2b90000c", 12848 => x"2b9b0008",
    12849 => x"379c0020", 12850 => x"c3a00000", 12851 => x"379cffec",
    12852 => x"5b8b0014", 12853 => x"5b8c0010", 12854 => x"5b8d000c",
    12855 => x"5b8e0008", 12856 => x"5b9d0004", 12857 => x"780b0001",
    12858 => x"396b6a30", 12859 => x"29610000", 12860 => x"5c200007",
    12861 => x"78010001", 12862 => x"38214c88", 12863 => x"f8001054",
    12864 => x"29610000", 12865 => x"34210001", 12866 => x"59610000",
    12867 => x"780b0001", 12868 => x"396b4bb0", 12869 => x"780c0001",
    12870 => x"356d00d8", 12871 => x"398c4c88", 12872 => x"e0000009",
    12873 => x"29620008", 12874 => x"2963000c", 12875 => x"29640010",
    12876 => x"296e0000", 12877 => x"b9800800", 12878 => x"f8001119",
    12879 => x"59c10000", 12880 => x"356b0018", 12881 => x"5d6dfff8",
    12882 => x"2b9d0004", 12883 => x"2b8b0014", 12884 => x"2b8c0010",
    12885 => x"2b8d000c", 12886 => x"2b8e0008", 12887 => x"379c0014",
    12888 => x"c3a00000", 12889 => x"379cfff4", 12890 => x"5b8b000c",
    12891 => x"5b8c0008", 12892 => x"5b9d0004", 12893 => x"34020000",
    12894 => x"b8206000", 12895 => x"f80002ca", 12896 => x"b8205800",
    12897 => x"4c200005", 12898 => x"78010001", 12899 => x"382136c0",
    12900 => x"b9601000", 12901 => x"e0000004", 12902 => x"29820000",
    12903 => x"78010001", 12904 => x"382136ec", 12905 => x"fbfff90b",
    12906 => x"b9600800", 12907 => x"2b9d0004", 12908 => x"2b8b000c",
    12909 => x"2b8c0008", 12910 => x"379c000c", 12911 => x"c3a00000",
    12912 => x"379cfffc", 12913 => x"5b9d0004", 12914 => x"78010001",
    12915 => x"38216a34", 12916 => x"58200000", 12917 => x"78020001",
    12918 => x"78010001", 12919 => x"38216a48", 12920 => x"38426a38",
    12921 => x"3403ffff", 12922 => x"58230000", 12923 => x"58430000",
    12924 => x"58200008", 12925 => x"58400008", 12926 => x"58400004",
    12927 => x"58200004", 12928 => x"5840000c", 12929 => x"5820000c",
    12930 => x"34020000", 12931 => x"34010000", 12932 => x"f8000dcf",
    12933 => x"2b9d0004", 12934 => x"379c0004", 12935 => x"c3a00000",
    12936 => x"379cfff4", 12937 => x"5b8b000c", 12938 => x"5b8c0008",
    12939 => x"5b9d0004", 12940 => x"b8206000", 12941 => x"34010000",
    12942 => x"f8000e6f", 12943 => x"b8205800", 12944 => x"34020000",
    12945 => x"5c20008b", 12946 => x"fbfffa8d", 12947 => x"78030001",
    12948 => x"38636a38", 12949 => x"28650008", 12950 => x"78020001",
    12951 => x"38426a34", 12952 => x"b8202000", 12953 => x"28420000",
    12954 => x"44ab0004", 12955 => x"34010001", 12956 => x"5ca1001d",
    12957 => x"e0000010", 12958 => x"34010001", 12959 => x"44810005",
    12960 => x"28610004", 12961 => x"34210001", 12962 => x"58610004",
    12963 => x"e0000002", 12964 => x"58600004", 12965 => x"78030001",
    12966 => x"38636a38", 12967 => x"28650004", 12968 => x"34010004",
    12969 => x"4c250010", 12970 => x"34010001", 12971 => x"58610008",
    12972 => x"e0000002", 12973 => x"44850003", 12974 => x"58600004",
    12975 => x"e000000a", 12976 => x"28650004", 12977 => x"34010004",
    12978 => x"34a50001", 12979 => x"58650004", 12980 => x"4c250005",
    12981 => x"34010002", 12982 => x"58610008", 12983 => x"3441fe0c",
    12984 => x"5861000c", 12985 => x"78030001", 12986 => x"38636a48",
    12987 => x"28650008", 12988 => x"44a00004", 12989 => x"34010001",
    12990 => x"5ca1001c", 12991 => x"e000000f", 12992 => x"44850005",
    12993 => x"28610004", 12994 => x"34210001", 12995 => x"58610004",
    12996 => x"e0000002", 12997 => x"58600004", 12998 => x"78030001",
    12999 => x"38636a48", 13000 => x"28640004", 13001 => x"34010004",
    13002 => x"4c240010", 13003 => x"34010001", 13004 => x"58610008",
    13005 => x"e0000002", 13006 => x"44800003", 13007 => x"58600004",
    13008 => x"e000000a", 13009 => x"28640004", 13010 => x"34010004",
    13011 => x"34840001", 13012 => x"58640004", 13013 => x"4c240005",
    13014 => x"34010002", 13015 => x"58610008", 13016 => x"3441fe0c",
    13017 => x"5861000c", 13018 => x"3401251b", 13019 => x"4c22003a",
    13020 => x"78020001", 13021 => x"38426a38", 13022 => x"28430008",
    13023 => x"34010002", 13024 => x"5c610008", 13025 => x"78020001",
    13026 => x"38426a48", 13027 => x"28410008", 13028 => x"5c230004",
    13029 => x"2844000c", 13030 => x"34011f3f", 13031 => x"e0000008",
    13032 => x"78020001", 13033 => x"3842370c", 13034 => x"34010000",
    13035 => x"fbffcd9a", 13036 => x"3402ffff", 13037 => x"e000002f",
    13038 => x"3484e0c0", 13039 => x"4881ffff", 13040 => x"78020001",
    13041 => x"38426a48", 13042 => x"5844000c", 13043 => x"78020001",
    13044 => x"38426a38", 13045 => x"2843000c", 13046 => x"34011f3f",
    13047 => x"e0000002", 13048 => x"3463e0c0", 13049 => x"4861ffff",
    13050 => x"78020001", 13051 => x"38426a38", 13052 => x"5843000c",
    13053 => x"4c640003", 13054 => x"348bf060", 13055 => x"e0000004",
    13056 => x"340b0000", 13057 => x"4c830002", 13058 => x"348b0fa0",
    13059 => x"b5635800", 13060 => x"0161001f", 13061 => x"b42b5800",
    13062 => x"156b0001", 13063 => x"4d600003", 13064 => x"356b1f40",
    13065 => x"e0000004", 13066 => x"34011f3f", 13067 => x"4c2b0002",
    13068 => x"356be0c0", 13069 => x"78020001", 13070 => x"38423728",
    13071 => x"34010000", 13072 => x"b9602800", 13073 => x"fbffcd74",
    13074 => x"34020001", 13075 => x"598b0000", 13076 => x"e0000008",
    13077 => x"78010001", 13078 => x"34420064", 13079 => x"38216a34",
    13080 => x"58220000", 13081 => x"34010000", 13082 => x"f8000d39",
    13083 => x"34020000", 13084 => x"b8400800", 13085 => x"2b9d0004",
    13086 => x"2b8b000c", 13087 => x"2b8c0008", 13088 => x"379c000c",
    13089 => x"c3a00000", 13090 => x"379cfff8", 13091 => x"5b8b0008",
    13092 => x"5b9d0004", 13093 => x"78020001", 13094 => x"b8205800",
    13095 => x"b8400800", 13096 => x"3821375c", 13097 => x"fbfff84b",
    13098 => x"e0000003", 13099 => x"34010064", 13100 => x"fbfffe7f",
    13101 => x"34010000", 13102 => x"fbfff999", 13103 => x"4420fffc",
    13104 => x"34010003", 13105 => x"34020000", 13106 => x"34030001",
    13107 => x"f8000c2a", 13108 => x"78020001", 13109 => x"b8400800",
    13110 => x"38213774", 13111 => x"fbfff83d", 13112 => x"e0000003",
    13113 => x"34010064", 13114 => x"fbfffe71", 13115 => x"34010000",
    13116 => x"f8000d06", 13117 => x"4420fffc", 13118 => x"78020001",
    13119 => x"b8400800", 13120 => x"38211b04", 13121 => x"fbfff833",
    13122 => x"78020001", 13123 => x"b8400800", 13124 => x"38213784",
    13125 => x"fbfff82f", 13126 => x"fbffff2a", 13127 => x"b9600800",
    13128 => x"fbffff40", 13129 => x"4420fffe", 13130 => x"2b9d0004",
    13131 => x"2b8b0008", 13132 => x"379c0008", 13133 => x"c3a00000",
    13134 => x"379cfff0", 13135 => x"5b8b000c", 13136 => x"5b8c0008",
    13137 => x"5b9d0004", 13138 => x"b8405800", 13139 => x"34020003",
    13140 => x"5c220020", 13141 => x"fbffff1b", 13142 => x"b9600800",
    13143 => x"fbffff31", 13144 => x"4420fffe", 13145 => x"4c200002",
    13146 => x"e000001a", 13147 => x"37810010", 13148 => x"34020000",
    13149 => x"f80001cc", 13150 => x"b8206000", 13151 => x"48010007",
    13152 => x"29620000", 13153 => x"2b810010", 13154 => x"3443ff38",
    13155 => x"54610003", 13156 => x"344200c8", 13157 => x"50410012",
    13158 => x"34020001", 13159 => x"b9600800", 13160 => x"f80001c1",
    13161 => x"78030001", 13162 => x"b8206000", 13163 => x"29620000",
    13164 => x"386337ac", 13165 => x"4c200003", 13166 => x"78030001",
    13167 => x"386337a4", 13168 => x"78010001", 13169 => x"382137b4",
    13170 => x"fbfff802", 13171 => x"e0000004", 13172 => x"b9600800",
    13173 => x"fbfffee4", 13174 => x"b8206000", 13175 => x"29610000",
    13176 => x"fbfff396", 13177 => x"b9800800", 13178 => x"2b9d0004",
    13179 => x"2b8b000c", 13180 => x"2b8c0008", 13181 => x"379c0010",
    13182 => x"c3a00000", 13183 => x"379cfffc", 13184 => x"5b9d0004",
    13185 => x"34010800", 13186 => x"34020001", 13187 => x"fbfffa60",
    13188 => x"34010400", 13189 => x"34020000", 13190 => x"fbfffa5d",
    13191 => x"34011000", 13192 => x"34020000", 13193 => x"fbfffa5a",
    13194 => x"2b9d0004", 13195 => x"379c0004", 13196 => x"c3a00000",
    13197 => x"40440000", 13198 => x"78030001", 13199 => x"40450001",
    13200 => x"38636dc0", 13201 => x"28630000", 13202 => x"3c840008",
    13203 => x"b8a42000", 13204 => x"58640010", 13205 => x"40450002",
    13206 => x"40440003", 13207 => x"3ca50018", 13208 => x"3c840010",
    13209 => x"b8a42800", 13210 => x"40440005", 13211 => x"b8a42800",
    13212 => x"40440004", 13213 => x"3c840008", 13214 => x"b8a41000",
    13215 => x"58620014", 13216 => x"40240000", 13217 => x"40220003",
    13218 => x"3c840018", 13219 => x"b8442000", 13220 => x"40220001",
    13221 => x"3c420010", 13222 => x"b8822000", 13223 => x"40220002",
    13224 => x"3c420008", 13225 => x"b8820800", 13226 => x"58610018",
    13227 => x"3801ea60", 13228 => x"5861001c", 13229 => x"78020001",
    13230 => x"34210001", 13231 => x"38423d2c", 13232 => x"58610020",
    13233 => x"34210001", 13234 => x"58610024", 13235 => x"28410000",
    13236 => x"78020001", 13237 => x"38423d30", 13238 => x"58610028",
    13239 => x"38019890", 13240 => x"5861002c", 13241 => x"28410000",
    13242 => x"58610030", 13243 => x"34011f40", 13244 => x"58610034",
    13245 => x"c3a00000", 13246 => x"379cffe0", 13247 => x"5b8b001c",
    13248 => x"5b8c0018", 13249 => x"5b8d0014", 13250 => x"5b8e0010",
    13251 => x"5b8f000c", 13252 => x"5b900008", 13253 => x"5b9d0004",
    13254 => x"b8205800", 13255 => x"78010001", 13256 => x"38216a58",
    13257 => x"b8406000", 13258 => x"40220000", 13259 => x"b8607000",
    13260 => x"b8807800", 13261 => x"b8a06800", 13262 => x"3401ffff",
    13263 => x"4440002b", 13264 => x"3d8c0001", 13265 => x"b9600800",
    13266 => x"fbfffa1f", 13267 => x"218200fe", 13268 => x"b9600800",
    13269 => x"fbfffa64", 13270 => x"01c20008", 13271 => x"b9600800",
    13272 => x"204200ff", 13273 => x"fbfffa60", 13274 => x"21c200ff",
    13275 => x"b9600800", 13276 => x"fbfffa5d", 13277 => x"b9600800",
    13278 => x"fbfffa27", 13279 => x"39820001", 13280 => x"b9600800",
    13281 => x"204200ff", 13282 => x"fbfffa57", 13283 => x"340c0000",
    13284 => x"35aeffff", 13285 => x"37900023", 13286 => x"e0000009",
    13287 => x"b9600800", 13288 => x"ba001000", 13289 => x"34030000",
    13290 => x"fbfffa8c", 13291 => x"43820023", 13292 => x"b5ec0800",
    13293 => x"358c0001", 13294 => x"30220000", 13295 => x"55ccfff8",
    13296 => x"b9600800", 13297 => x"ba001000", 13298 => x"34030001",
    13299 => x"fbfffa83", 13300 => x"43810023", 13301 => x"b5ee7000",
    13302 => x"31c10000", 13303 => x"b9600800", 13304 => x"fbfffa29",
    13305 => x"b9a00800", 13306 => x"2b9d0004", 13307 => x"2b8b001c",
    13308 => x"2b8c0018", 13309 => x"2b8d0014", 13310 => x"2b8e0010",
    13311 => x"2b8f000c", 13312 => x"2b900008", 13313 => x"379c0020",
    13314 => x"c3a00000", 13315 => x"379cffe0", 13316 => x"5b8b0020",
    13317 => x"5b8c001c", 13318 => x"5b8d0018", 13319 => x"5b8e0014",
    13320 => x"5b8f0010", 13321 => x"5b90000c", 13322 => x"5b910008",
    13323 => x"5b9d0004", 13324 => x"b8205800", 13325 => x"78010001",
    13326 => x"38216a58", 13327 => x"b8606800", 13328 => x"40230000",
    13329 => x"3c4f0001", 13330 => x"b8808000", 13331 => x"b8a07000",
    13332 => x"3401ffff", 13333 => x"21ef00ff", 13334 => x"340c0000",
    13335 => x"5c60001f", 13336 => x"e0000020", 13337 => x"b9600800",
    13338 => x"fbfff9d7", 13339 => x"b9e01000", 13340 => x"b9600800",
    13341 => x"fbfffa1c", 13342 => x"01a20008", 13343 => x"b9600800",
    13344 => x"204200ff", 13345 => x"fbfffa18", 13346 => x"21a200ff",
    13347 => x"b9600800", 13348 => x"fbfffa15", 13349 => x"b60c1000",
    13350 => x"40420000", 13351 => x"b9600800", 13352 => x"35ad0001",
    13353 => x"fbfffa10", 13354 => x"b9600800", 13355 => x"fbfff9f6",
    13356 => x"b9600800", 13357 => x"fbfff9c4", 13358 => x"b9600800",
    13359 => x"b9e01000", 13360 => x"fbfffa09", 13361 => x"b8208800",
    13362 => x"b9600800", 13363 => x"fbfff9ee", 13364 => x"5e20fff8",
    13365 => x"358c0001", 13366 => x"55ccffe3", 13367 => x"b9c00800",
    13368 => x"2b9d0004", 13369 => x"2b8b0020", 13370 => x"2b8c001c",
    13371 => x"2b8d0018", 13372 => x"2b8e0014", 13373 => x"2b8f0010",
    13374 => x"2b90000c", 13375 => x"2b910008", 13376 => x"379c0020",
    13377 => x"c3a00000", 13378 => x"379cffec", 13379 => x"5b8b0014",
    13380 => x"5b8c0010", 13381 => x"5b8d000c", 13382 => x"5b8e0008",
    13383 => x"5b9d0004", 13384 => x"780d0001", 13385 => x"780c0001",
    13386 => x"39ad6a5c", 13387 => x"398c6a60", 13388 => x"780b0001",
    13389 => x"59a10000", 13390 => x"59820000", 13391 => x"34030001",
    13392 => x"396b6a58", 13393 => x"202100ff", 13394 => x"204200ff",
    13395 => x"31630000", 13396 => x"fbfffa80", 13397 => x"b8207000",
    13398 => x"5c200006", 13399 => x"41a10003", 13400 => x"41820003",
    13401 => x"fbfffa7b", 13402 => x"5c2e0002", 13403 => x"31600000",
    13404 => x"2b9d0004", 13405 => x"2b8b0014", 13406 => x"2b8c0010",
    13407 => x"2b8d000c", 13408 => x"2b8e0008", 13409 => x"379c0014",
    13410 => x"c3a00000", 13411 => x"379cfff8", 13412 => x"5b9d0004",
    13413 => x"78010001", 13414 => x"78020001", 13415 => x"38216a5c",
    13416 => x"38426a60", 13417 => x"40420003", 13418 => x"40210003",
    13419 => x"34031004", 13420 => x"3784000b", 13421 => x"34050001",
    13422 => x"3380000b", 13423 => x"fbffff94", 13424 => x"34030001",
    13425 => x"3402ffff", 13426 => x"5c230002", 13427 => x"4382000b",
    13428 => x"b8400800", 13429 => x"2b9d0004", 13430 => x"379c0008",
    13431 => x"c3a00000", 13432 => x"379cffec", 13433 => x"5b8b0014",
    13434 => x"5b8c0010", 13435 => x"5b8d000c", 13436 => x"5b8e0008",
    13437 => x"5b9d0004", 13438 => x"b8205800", 13439 => x"206d00ff",
    13440 => x"34010003", 13441 => x"204c00ff", 13442 => x"3405fffc",
    13443 => x"55a1005d", 13444 => x"5da0000f", 13445 => x"78010001",
    13446 => x"78020001", 13447 => x"38216a5c", 13448 => x"38426a60",
    13449 => x"40420003", 13450 => x"40210003", 13451 => x"78040001",
    13452 => x"34050001", 13453 => x"34031004", 13454 => x"38846a68",
    13455 => x"fbffff2f", 13456 => x"34020001", 13457 => x"3405ffff",
    13458 => x"5c22004e", 13459 => x"45800007", 13460 => x"78010001",
    13461 => x"38216a68", 13462 => x"40220000", 13463 => x"34010004",
    13464 => x"3405fffe", 13465 => x"44410047", 13466 => x"b9ac0800",
    13467 => x"5c200007", 13468 => x"78010001", 13469 => x"38216a68",
    13470 => x"40210000", 13471 => x"34050000", 13472 => x"5c250006",
    13473 => x"e000003f", 13474 => x"3562001c", 13475 => x"b9600800",
    13476 => x"34030000", 13477 => x"5d80001b", 13478 => x"78010001",
    13479 => x"78020001", 13480 => x"38216a5c", 13481 => x"38426a60",
    13482 => x"09a3001d", 13483 => x"40420003", 13484 => x"40210003",
    13485 => x"3405001d", 13486 => x"34631005", 13487 => x"b9602000",
    13488 => x"fbffff0e", 13489 => x"3402001d", 13490 => x"b9606000",
    13491 => x"3405ffff", 13492 => x"5c22002c", 13493 => x"3562001c",
    13494 => x"34010000", 13495 => x"41830000", 13496 => x"358c0001",
    13497 => x"b4230800", 13498 => x"202100ff", 13499 => x"5d82fffc",
    13500 => x"4162001c", 13501 => x"3405fffd", 13502 => x"5c410022",
    13503 => x"e000001e", 13504 => x"40240000", 13505 => x"34210001",
    13506 => x"b4641800", 13507 => x"206300ff", 13508 => x"5c22fffc",
    13509 => x"780c0001", 13510 => x"3163001c", 13511 => x"398c6a68",
    13512 => x"41830000", 13513 => x"780e0001", 13514 => x"780d0001",
    13515 => x"39ce6a5c", 13516 => x"39ad6a60", 13517 => x"0863001d",
    13518 => x"41a20003", 13519 => x"41c10003", 13520 => x"34631005",
    13521 => x"b9602000", 13522 => x"3405001d", 13523 => x"fbffff30",
    13524 => x"41810000", 13525 => x"41a20003", 13526 => x"34031004",
    13527 => x"34210001", 13528 => x"31810000", 13529 => x"41c10003",
    13530 => x"b9802000", 13531 => x"34050001", 13532 => x"fbffff27",
    13533 => x"78010001", 13534 => x"38216a68", 13535 => x"40250000",
    13536 => x"b8a00800", 13537 => x"2b9d0004", 13538 => x"2b8b0014",
    13539 => x"2b8c0010", 13540 => x"2b8d000c", 13541 => x"2b8e0008",
    13542 => x"379c0014", 13543 => x"c3a00000", 13544 => x"379cffc8",
    13545 => x"5b8b0018", 13546 => x"5b8c0014", 13547 => x"5b8d0010",
    13548 => x"5b8e000c", 13549 => x"5b8f0008", 13550 => x"5b9d0004",
    13551 => x"340c0000", 13552 => x"b8205800", 13553 => x"340d0001",
    13554 => x"378e001c", 13555 => x"340f00fd", 13556 => x"e000002b",
    13557 => x"34020000", 13558 => x"b9c00800", 13559 => x"b9801800",
    13560 => x"fbffff80", 13561 => x"b1801000", 13562 => x"5c400005",
    13563 => x"202d00ff", 13564 => x"35a1ffff", 13565 => x"202100ff",
    13566 => x"542f0022", 13567 => x"b9c00800", 13568 => x"b9601000",
    13569 => x"34030010", 13570 => x"f800107d", 13571 => x"358c0001",
    13572 => x"5c20001b", 13573 => x"2b810030", 13574 => x"00220018",
    13575 => x"31610017", 13576 => x"31620014", 13577 => x"00220010",
    13578 => x"31620015", 13579 => x"00220008", 13580 => x"2b810034",
    13581 => x"31620016", 13582 => x"00220018", 13583 => x"3161001b",
    13584 => x"31620018", 13585 => x"00220010", 13586 => x"31620019",
    13587 => x"00220008", 13588 => x"2b81002c", 13589 => x"3162001a",
    13590 => x"00220018", 13591 => x"31610013", 13592 => x"31620010",
    13593 => x"00220010", 13594 => x"31620011", 13595 => x"00220008",
    13596 => x"34010001", 13597 => x"31620012", 13598 => x"e0000003",
    13599 => x"49acffd6", 13600 => x"34010000", 13601 => x"2b9d0004",
    13602 => x"2b8b0018", 13603 => x"2b8c0014", 13604 => x"2b8d0010",
    13605 => x"2b8e000c", 13606 => x"2b8f0008", 13607 => x"379c0038",
    13608 => x"c3a00000", 13609 => x"379cfff8", 13610 => x"5b8b0008",
    13611 => x"5b9d0004", 13612 => x"78030001", 13613 => x"b8205800",
    13614 => x"204200ff", 13615 => x"78010001", 13616 => x"38216a5c",
    13617 => x"38636a60", 13618 => x"44400015", 13619 => x"29640000",
    13620 => x"78028000", 13621 => x"34050004", 13622 => x"b8821000",
    13623 => x"59620000", 13624 => x"40620003", 13625 => x"40210003",
    13626 => x"34031000", 13627 => x"b9602000", 13628 => x"fbfffec7",
    13629 => x"7c210004", 13630 => x"78040001", 13631 => x"38843d20",
    13632 => x"c8011000", 13633 => x"29630000", 13634 => x"28810000",
    13635 => x"38420001", 13636 => x"a0610800", 13637 => x"59610000",
    13638 => x"e0000013", 13639 => x"40620003", 13640 => x"40210003",
    13641 => x"34031000", 13642 => x"b9602000", 13643 => x"34050004",
    13644 => x"fbfffe72", 13645 => x"34030004", 13646 => x"3402ffff",
    13647 => x"5c23000a", 13648 => x"29610000", 13649 => x"34020000",
    13650 => x"4c200007", 13651 => x"78030001", 13652 => x"38633d20",
    13653 => x"28620000", 13654 => x"a0220800", 13655 => x"59610000",
    13656 => x"34020001", 13657 => x"b8400800", 13658 => x"2b9d0004",
    13659 => x"2b8b0008", 13660 => x"379c0008", 13661 => x"c3a00000",
    13662 => x"379cfff8", 13663 => x"5b9d0004", 13664 => x"78010001",
    13665 => x"78020001", 13666 => x"38216a5c", 13667 => x"38426a60",
    13668 => x"40420003", 13669 => x"40210003", 13670 => x"34031074",
    13671 => x"3784000a", 13672 => x"34050002", 13673 => x"0f80000a",
    13674 => x"fbfffe99", 13675 => x"34030002", 13676 => x"3402ffff",
    13677 => x"5c230002", 13678 => x"2f82000a", 13679 => x"b8400800",
    13680 => x"2b9d0004", 13681 => x"379c0008", 13682 => x"c3a00000",
    13683 => x"379cffcc", 13684 => x"5b8b002c", 13685 => x"5b8c0028",
    13686 => x"5b8d0024", 13687 => x"5b8e0020", 13688 => x"5b8f001c",
    13689 => x"5b900018", 13690 => x"5b910014", 13691 => x"5b920010",
    13692 => x"5b93000c", 13693 => x"5b940008", 13694 => x"5b9d0004",
    13695 => x"78030001", 13696 => x"78020001", 13697 => x"38636a5c",
    13698 => x"b8208800", 13699 => x"38426a60", 13700 => x"34010020",
    13701 => x"33810037", 13702 => x"40420003", 13703 => x"40610003",
    13704 => x"37840034", 13705 => x"34031074", 13706 => x"34050002",
    13707 => x"fbfffe33", 13708 => x"34020002", 13709 => x"340bffff",
    13710 => x"5c220051", 13711 => x"2f820034", 13712 => x"3801ffff",
    13713 => x"5c410002", 13714 => x"0f800034", 13715 => x"780d0001",
    13716 => x"780c0001", 13717 => x"340b0001", 13718 => x"39ad6a5c",
    13719 => x"398c6a60", 13720 => x"37900037", 13721 => x"e0000023",
    13722 => x"41b40003", 13723 => x"41930003", 13724 => x"b9c00800",
    13725 => x"34721076", 13726 => x"f8000fb2", 13727 => x"b8202800",
    13728 => x"b9c02000", 13729 => x"ba800800", 13730 => x"ba601000",
    13731 => x"ba401800", 13732 => x"fbfffe5f", 13733 => x"b8207000",
    13734 => x"29e10000", 13735 => x"f8000fa9", 13736 => x"5dc10036",
    13737 => x"29e10000", 13738 => x"2f8e0034", 13739 => x"f8000fa5",
    13740 => x"b5c11800", 13741 => x"41820003", 13742 => x"41a10003",
    13743 => x"2063ffff", 13744 => x"0f830034", 13745 => x"ba002000",
    13746 => x"34631076", 13747 => x"34050001", 13748 => x"fbfffe4f",
    13749 => x"34020001", 13750 => x"5c220028", 13751 => x"2f810034",
    13752 => x"356b0001", 13753 => x"216b00ff", 13754 => x"34210001",
    13755 => x"0f810034", 13756 => x"3d6f0002", 13757 => x"2f830034",
    13758 => x"b62f7800", 13759 => x"29ee0000", 13760 => x"5dc0ffda",
    13761 => x"3401000a", 13762 => x"33810037", 13763 => x"41820003",
    13764 => x"41a10003", 13765 => x"34631075", 13766 => x"37840037",
    13767 => x"34050001", 13768 => x"fbfffe3b", 13769 => x"34020001",
    13770 => x"340bffff", 13771 => x"5c220014", 13772 => x"41a10003",
    13773 => x"41820003", 13774 => x"34031074", 13775 => x"37840034",
    13776 => x"34050002", 13777 => x"fbfffe32", 13778 => x"b8207000",
    13779 => x"34010002", 13780 => x"5dc1000b", 13781 => x"41a10003",
    13782 => x"41820003", 13783 => x"34031074", 13784 => x"37840032",
    13785 => x"34050002", 13786 => x"fbfffde4", 13787 => x"e42e5800",
    13788 => x"356bffff", 13789 => x"e0000002", 13790 => x"340bffff",
    13791 => x"b9600800", 13792 => x"2b9d0004", 13793 => x"2b8b002c",
    13794 => x"2b8c0028", 13795 => x"2b8d0024", 13796 => x"2b8e0020",
    13797 => x"2b8f001c", 13798 => x"2b900018", 13799 => x"2b910014",
    13800 => x"2b920010", 13801 => x"2b93000c", 13802 => x"2b940008",
    13803 => x"379c0034", 13804 => x"c3a00000", 13805 => x"379cffe4",
    13806 => x"5b8b0018", 13807 => x"5b8c0014", 13808 => x"5b8d0010",
    13809 => x"5b8e000c", 13810 => x"5b8f0008", 13811 => x"5b9d0004",
    13812 => x"78010001", 13813 => x"78020001", 13814 => x"38216a5c",
    13815 => x"38426a60", 13816 => x"40420003", 13817 => x"40210003",
    13818 => x"34031074", 13819 => x"3784001c", 13820 => x"34050002",
    13821 => x"fbfffdc1", 13822 => x"34030002", 13823 => x"3402ffff",
    13824 => x"5c230025", 13825 => x"2f81001c", 13826 => x"3802fffd",
    13827 => x"3421ffff", 13828 => x"2021ffff", 13829 => x"50410005",
    13830 => x"78010001", 13831 => x"38212fdc", 13832 => x"0f80001c",
    13833 => x"fbfff56b", 13834 => x"780e0001", 13835 => x"780d0001",
    13836 => x"780c0001", 13837 => x"340b0000", 13838 => x"39ce6a5c",
    13839 => x"39ad6a60", 13840 => x"378f001f", 13841 => x"398c2fd8",
    13842 => x"e000000e", 13843 => x"41a20003", 13844 => x"41c10003",
    13845 => x"35631076", 13846 => x"b9e02000", 13847 => x"34050001",
    13848 => x"fbfffda6", 13849 => x"34020001", 13850 => x"5c22000a",
    13851 => x"4382001f", 13852 => x"b9800800", 13853 => x"356b0001",
    13854 => x"fbfff556", 13855 => x"216bffff", 13856 => x"2f81001c",
    13857 => x"542bfff2", 13858 => x"34020000", 13859 => x"e0000002",
    13860 => x"3402ffff", 13861 => x"b8400800", 13862 => x"2b9d0004",
    13863 => x"2b8b0018", 13864 => x"2b8c0014", 13865 => x"2b8d0010",
    13866 => x"2b8e000c", 13867 => x"2b8f0008", 13868 => x"379c001c",
    13869 => x"c3a00000", 13870 => x"379cffdc", 13871 => x"5b8b0024",
    13872 => x"5b8c0020", 13873 => x"5b8d001c", 13874 => x"5b8e0018",
    13875 => x"5b8f0014", 13876 => x"5b900010", 13877 => x"5b91000c",
    13878 => x"5b920008", 13879 => x"5b9d0004", 13880 => x"206300ff",
    13881 => x"b8208800", 13882 => x"205200ff", 13883 => x"5c600012",
    13884 => x"78040001", 13885 => x"78030001", 13886 => x"38846a5c",
    13887 => x"38636a60", 13888 => x"40620003", 13889 => x"40810003",
    13890 => x"78040001", 13891 => x"34031074", 13892 => x"38846a64",
    13893 => x"34050002", 13894 => x"fbfffd78", 13895 => x"34020002",
    13896 => x"3403ffff", 13897 => x"5c22002b", 13898 => x"78030001",
    13899 => x"38636a66", 13900 => x"0c610000", 13901 => x"78040001",
    13902 => x"38846a66", 13903 => x"78030001", 13904 => x"38636a64",
    13905 => x"2c820000", 13906 => x"2c610000", 13907 => x"34030000",
    13908 => x"3442fffe", 13909 => x"5041001f", 13910 => x"780d0001",
    13911 => x"780c0001", 13912 => x"340b0000", 13913 => x"b8807000",
    13914 => x"39ad6a5c", 13915 => x"398c6a60", 13916 => x"3410000a",
    13917 => x"2dc30000", 13918 => x"3461fffe", 13919 => x"54320012",
    13920 => x"41820003", 13921 => x"41a10003", 13922 => x"34640001",
    13923 => x"b62b7800", 13924 => x"0dc40000", 13925 => x"34631074",
    13926 => x"b9e02000", 13927 => x"34050001", 13928 => x"fbfffd56",
    13929 => x"34020001", 13930 => x"5c220009", 13931 => x"41e10000",
    13932 => x"356b0001", 13933 => x"216b00ff", 13934 => x"5c30ffef",
    13935 => x"b9601800", 13936 => x"e0000004", 13937 => x"3403fffd",
    13938 => x"e0000002", 13939 => x"3403ffff", 13940 => x"b8600800",
    13941 => x"2b9d0004", 13942 => x"2b8b0024", 13943 => x"2b8c0020",
    13944 => x"2b8d001c", 13945 => x"2b8e0018", 13946 => x"2b8f0014",
    13947 => x"2b900010", 13948 => x"2b91000c", 13949 => x"2b920008",
    13950 => x"379c0024", 13951 => x"c3a00000", 13952 => x"379cfffc",
    13953 => x"5b9d0004", 13954 => x"78010001", 13955 => x"382137d8",
    13956 => x"fbfff4f0", 13957 => x"3401ffff", 13958 => x"2b9d0004",
    13959 => x"379c0004", 13960 => x"c3a00000", 13961 => x"379cfff8",
    13962 => x"5b8b0008", 13963 => x"5b9d0004", 13964 => x"78010001",
    13965 => x"b8405800", 13966 => x"78020001", 13967 => x"3842408c",
    13968 => x"382137fc", 13969 => x"fbfff4e3", 13970 => x"78020001",
    13971 => x"78010001", 13972 => x"38426d18", 13973 => x"38216d28",
    13974 => x"34460090", 13975 => x"34050022", 13976 => x"34040033",
    13977 => x"28220004", 13978 => x"204300ff", 13979 => x"7c670042",
    13980 => x"7c630028", 13981 => x"a0e31800", 13982 => x"5c60000b",
    13983 => x"28230000", 13984 => x"31650000", 13985 => x"31640001",
    13986 => x"31630002", 13987 => x"00430018", 13988 => x"31630003",
    13989 => x"00430010", 13990 => x"00420008", 13991 => x"31630004",
    13992 => x"31620005", 13993 => x"34210010", 13994 => x"5c26ffef",
    13995 => x"34010000", 13996 => x"2b9d0004", 13997 => x"2b8b0008",
    13998 => x"379c0008", 13999 => x"c3a00000", 14000 => x"379cffe8",
    14001 => x"5b8b0018", 14002 => x"5b8c0014", 14003 => x"5b8d0010",
    14004 => x"5b8e000c", 14005 => x"5b8f0008", 14006 => x"5b9d0004",
    14007 => x"780b0001", 14008 => x"b8207800", 14009 => x"b8407000",
    14010 => x"340d0008", 14011 => x"340c0001", 14012 => x"396b4d40",
    14013 => x"a18e1800", 14014 => x"29640008", 14015 => x"7c620000",
    14016 => x"b9e00800", 14017 => x"35adffff", 14018 => x"d8800000",
    14019 => x"3d8c0001", 14020 => x"5da0fff9", 14021 => x"2b9d0004",
    14022 => x"2b8b0018", 14023 => x"2b8c0014", 14024 => x"2b8d0010",
    14025 => x"2b8e000c", 14026 => x"2b8f0008", 14027 => x"379c0018",
    14028 => x"c3a00000", 14029 => x"379cffe8", 14030 => x"5b8b0018",
    14031 => x"5b8c0014", 14032 => x"5b8d0010", 14033 => x"5b8e000c",
    14034 => x"5b8f0008", 14035 => x"5b9d0004", 14036 => x"780b0001",
    14037 => x"b8207800", 14038 => x"340e0008", 14039 => x"340c0000",
    14040 => x"340d0001", 14041 => x"396b4d40", 14042 => x"29620004",
    14043 => x"b9e00800", 14044 => x"35ceffff", 14045 => x"d8400000",
    14046 => x"7c220000", 14047 => x"c8021000", 14048 => x"a1a21000",
    14049 => x"b9826000", 14050 => x"3dad0001", 14051 => x"5dc0fff7",
    14052 => x"34010064", 14053 => x"fbfff009", 14054 => x"b9800800",
    14055 => x"2b9d0004", 14056 => x"2b8b0018", 14057 => x"2b8c0014",
    14058 => x"2b8d0010", 14059 => x"2b8e000c", 14060 => x"2b8f0008",
    14061 => x"379c0018", 14062 => x"c3a00000", 14063 => x"379cffc0",
    14064 => x"5b8b0040", 14065 => x"5b8c003c", 14066 => x"5b8d0038",
    14067 => x"5b8e0034", 14068 => x"5b8f0030", 14069 => x"5b90002c",
    14070 => x"5b910028", 14071 => x"5b920024", 14072 => x"5b930020",
    14073 => x"5b94001c", 14074 => x"5b950018", 14075 => x"5b960014",
    14076 => x"5b970010", 14077 => x"5b98000c", 14078 => x"5b990008",
    14079 => x"5b9d0004", 14080 => x"34020000", 14081 => x"b8206000",
    14082 => x"34030080", 14083 => x"34210008", 14084 => x"780d0001",
    14085 => x"f8000dc5", 14086 => x"39ad4d40", 14087 => x"29a10000",
    14088 => x"340f0000", 14089 => x"44200061", 14090 => x"b9805800",
    14091 => x"34120000", 14092 => x"34110000", 14093 => x"78194000",
    14094 => x"34160001", 14095 => x"34180008", 14096 => x"596c0008",
    14097 => x"45e00022", 14098 => x"29610000", 14099 => x"78028000",
    14100 => x"34030000", 14101 => x"59610010", 14102 => x"29610004",
    14103 => x"59610014", 14104 => x"a0590800", 14105 => x"44200003",
    14106 => x"78024000", 14107 => x"34030000", 14108 => x"a0710800",
    14109 => x"a0522800", 14110 => x"b8a12800", 14111 => x"29640010",
    14112 => x"29610014", 14113 => x"5ca0000e", 14114 => x"a4603000",
    14115 => x"a0260800", 14116 => x"59610014", 14117 => x"00630001",
    14118 => x"3c41001f", 14119 => x"a4403800", 14120 => x"00420001",
    14121 => x"a0872000", 14122 => x"b8231800", 14123 => x"59640010",
    14124 => x"b8430800", 14125 => x"5c25ffeb", 14126 => x"e000003c",
    14127 => x"b8821000", 14128 => x"b8231800", 14129 => x"59620010",
    14130 => x"59630014", 14131 => x"35ee0001", 14132 => x"29a20000",
    14133 => x"3dce0004", 14134 => x"b9800800", 14135 => x"b58e7000",
    14136 => x"d8400000", 14137 => x"5c360031", 14138 => x"b9800800",
    14139 => x"340200f0", 14140 => x"fbffff74", 14141 => x"34140040",
    14142 => x"34130000", 14143 => x"34100001", 14144 => x"34120000",
    14145 => x"34110000", 14146 => x"29a20004", 14147 => x"b9800800",
    14148 => x"29d70004", 14149 => x"d8400000", 14150 => x"29a20004",
    14151 => x"b820a800", 14152 => x"b9800800", 14153 => x"a2f0b800",
    14154 => x"d8400000", 14155 => x"46a10008", 14156 => x"29a30008",
    14157 => x"baa01000", 14158 => x"7eb50000", 14159 => x"b9800800",
    14160 => x"d8600000", 14161 => x"5eb60011", 14162 => x"e0000007",
    14163 => x"29a30008", 14164 => x"b9800800", 14165 => x"bae01000",
    14166 => x"d8600000", 14167 => x"46e00009", 14168 => x"e000000a",
    14169 => x"29c10000", 14170 => x"b8330800", 14171 => x"59c10000",
    14172 => x"29c10004", 14173 => x"b8300800", 14174 => x"59c10004",
    14175 => x"e0000003", 14176 => x"ba539000", 14177 => x"ba308800",
    14178 => x"3e010001", 14179 => x"3e730001", 14180 => x"f6018000",
    14181 => x"3694ffff", 14182 => x"b6139800", 14183 => x"b8208000",
    14184 => x"5e80ffda", 14185 => x"e0000014", 14186 => x"b9e00800",
    14187 => x"2b9d0004", 14188 => x"2b8b0040", 14189 => x"2b8c003c",
    14190 => x"2b8d0038", 14191 => x"2b8e0034", 14192 => x"2b8f0030",
    14193 => x"2b90002c", 14194 => x"2b910028", 14195 => x"2b920024",
    14196 => x"2b930020", 14197 => x"2b94001c", 14198 => x"2b950018",
    14199 => x"2b960014", 14200 => x"2b970010", 14201 => x"2b98000c",
    14202 => x"2b990008", 14203 => x"379c0040", 14204 => x"c3a00000",
    14205 => x"35ef0001", 14206 => x"356b0010", 14207 => x"5df8ff91",
    14208 => x"e3ffffea", 14209 => x"379cfff0", 14210 => x"5b8b0010",
    14211 => x"5b8c000c", 14212 => x"5b8d0008", 14213 => x"5b9d0004",
    14214 => x"b8205800", 14215 => x"78010001", 14216 => x"38214d40",
    14217 => x"28220000", 14218 => x"29610000", 14219 => x"340c0000",
    14220 => x"340d0040", 14221 => x"d8400000", 14222 => x"29610000",
    14223 => x"34020055", 14224 => x"fbffff20", 14225 => x"29610008",
    14226 => x"2962000c", 14227 => x"b9801800", 14228 => x"358c0008",
    14229 => x"f8000bfa", 14230 => x"29610000", 14231 => x"fbffff19",
    14232 => x"5d8dfff9", 14233 => x"2b9d0004", 14234 => x"2b8b0010",
    14235 => x"2b8c000c", 14236 => x"2b8d0008", 14237 => x"379c0010",
    14238 => x"c3a00000", 14239 => x"28210000", 14240 => x"78020001",
    14241 => x"38426da0", 14242 => x"28420000", 14243 => x"3c210008",
    14244 => x"3821000a", 14245 => x"58410000", 14246 => x"28410000",
    14247 => x"20230008", 14248 => x"5c60fffe", 14249 => x"20210001",
    14250 => x"18210001", 14251 => x"c3a00000", 14252 => x"28210000",
    14253 => x"78020001", 14254 => x"38426da0", 14255 => x"28420000",
    14256 => x"3c210008", 14257 => x"38210009", 14258 => x"58410000",
    14259 => x"28410000", 14260 => x"20230008", 14261 => x"5c60fffe",
    14262 => x"20210001", 14263 => x"c3a00000", 14264 => x"28210000",
    14265 => x"78030001", 14266 => x"38636da0", 14267 => x"3c210008",
    14268 => x"28630000", 14269 => x"7c420000", 14270 => x"38210008",
    14271 => x"b8221000", 14272 => x"58620000", 14273 => x"28610000",
    14274 => x"20210008", 14275 => x"5c20fffe", 14276 => x"c3a00000",
    14277 => x"78010001", 14278 => x"78030001", 14279 => x"38216da0",
    14280 => x"38633d34", 14281 => x"28210000", 14282 => x"28620000",
    14283 => x"58220004", 14284 => x"c3a00000", 14285 => x"379cffc4",
    14286 => x"5b8b001c", 14287 => x"5b8c0018", 14288 => x"5b8d0014",
    14289 => x"5b8e0010", 14290 => x"5b8f000c", 14291 => x"5b900008",
    14292 => x"5b9d0004", 14293 => x"b8206000", 14294 => x"28210000",
    14295 => x"340bffff", 14296 => x"4420002a", 14297 => x"29820004",
    14298 => x"44400028", 14299 => x"fbffeec7", 14300 => x"780e0001",
    14301 => x"b8206800", 14302 => x"340b0000", 14303 => x"3410001f",
    14304 => x"378f0020", 14305 => x"39ce3818", 14306 => x"e000000b",
    14307 => x"fbffeebf", 14308 => x"202400ff", 14309 => x"b56d1000",
    14310 => x"b5eb0800", 14311 => x"30240000", 14312 => x"b8401800",
    14313 => x"b9c00800", 14314 => x"b8802800", 14315 => x"fbfff389",
    14316 => x"356b0001", 14317 => x"29810004", 14318 => x"ee0b1800",
    14319 => x"358c0004", 14320 => x"7c220000", 14321 => x"a0621000",
    14322 => x"5c40fff1", 14323 => x"78010001", 14324 => x"b9602000",
    14325 => x"b9a01000", 14326 => x"b9e01800", 14327 => x"38216d18",
    14328 => x"f80001cc", 14329 => x"b8206000", 14330 => x"b9601800",
    14331 => x"78010001", 14332 => x"fd8b5800", 14333 => x"3821383c",
    14334 => x"b9a01000", 14335 => x"b9802000", 14336 => x"fbfff374",
    14337 => x"c80b5800", 14338 => x"b9600800", 14339 => x"2b9d0004",
    14340 => x"2b8b001c", 14341 => x"2b8c0018", 14342 => x"2b8d0014",
    14343 => x"2b8e0010", 14344 => x"2b8f000c", 14345 => x"2b900008",
    14346 => x"379c003c", 14347 => x"c3a00000", 14348 => x"379cffc8",
    14349 => x"5b8b0018", 14350 => x"5b8c0014", 14351 => x"5b8d0010",
    14352 => x"5b8e000c", 14353 => x"5b8f0008", 14354 => x"5b9d0004",
    14355 => x"b8205800", 14356 => x"28210000", 14357 => x"3405ffff",
    14358 => x"4420002c", 14359 => x"29620004", 14360 => x"4440002a",
    14361 => x"fbffee89", 14362 => x"b8207000", 14363 => x"29610004",
    14364 => x"fbffee86", 14365 => x"b8205800", 14366 => x"34010020",
    14367 => x"4c2b0002", 14368 => x"340b0020", 14369 => x"378d001c",
    14370 => x"78010001", 14371 => x"b9602000", 14372 => x"b9c01000",
    14373 => x"b9a01800", 14374 => x"38216d18", 14375 => x"f8000189",
    14376 => x"b8206000", 14377 => x"78010001", 14378 => x"b9601800",
    14379 => x"3821385c", 14380 => x"b9c01000", 14381 => x"b9802000",
    14382 => x"fbfff346", 14383 => x"e98b5800", 14384 => x"ec0c0800",
    14385 => x"3405ffff", 14386 => x"b9615800", 14387 => x"5d60000f",
    14388 => x"b9a07800", 14389 => x"780d0001", 14390 => x"39ad3818",
    14391 => x"b5eb0800", 14392 => x"40240000", 14393 => x"b56e1000",
    14394 => x"b9a00800", 14395 => x"b8401800", 14396 => x"b8802800",
    14397 => x"356b0001", 14398 => x"fbfff336", 14399 => x"498bfff8",
    14400 => x"fd8b2800", 14401 => x"c8052800", 14402 => x"b8a00800",
    14403 => x"2b9d0004", 14404 => x"2b8b0018", 14405 => x"2b8c0014",
    14406 => x"2b8d0010", 14407 => x"2b8e000c", 14408 => x"2b8f0008",
    14409 => x"379c0038", 14410 => x"c3a00000", 14411 => x"379cffe4",
    14412 => x"5b8b001c", 14413 => x"5b8c0018", 14414 => x"5b8d0014",
    14415 => x"5b8e0010", 14416 => x"5b8f000c", 14417 => x"5b900008",
    14418 => x"5b9d0004", 14419 => x"780d0001", 14420 => x"39ad6d18",
    14421 => x"b9a00800", 14422 => x"780b0001", 14423 => x"780f0001",
    14424 => x"780e0001", 14425 => x"fbfffe96", 14426 => x"396b6d28",
    14427 => x"340c0000", 14428 => x"39ef387c", 14429 => x"39ce3894",
    14430 => x"34100008", 14431 => x"29630000", 14432 => x"29640004",
    14433 => x"b8640800", 14434 => x"44200010", 14435 => x"b9801000",
    14436 => x"b9e00800", 14437 => x"fbfff30f", 14438 => x"3d810004",
    14439 => x"34020000", 14440 => x"34210008", 14441 => x"b5a10800",
    14442 => x"f8000015", 14443 => x"2023ffff", 14444 => x"08632710",
    14445 => x"b8201000", 14446 => x"14420010", 14447 => x"14630010",
    14448 => x"b9c00800", 14449 => x"fbfff303", 14450 => x"358c0001",
    14451 => x"356b0010", 14452 => x"5d90ffeb", 14453 => x"34010000",
    14454 => x"2b9d0004", 14455 => x"2b8b001c", 14456 => x"2b8c0018",
    14457 => x"2b8d0014", 14458 => x"2b8e0010", 14459 => x"2b8f000c",
    14460 => x"2b900008", 14461 => x"379c001c", 14462 => x"c3a00000",
    14463 => x"379cffec", 14464 => x"5b8b0014", 14465 => x"5b8c0010",
    14466 => x"5b8d000c", 14467 => x"5b8e0008", 14468 => x"5b9d0004",
    14469 => x"402d000f", 14470 => x"b8206000", 14471 => x"34010028",
    14472 => x"b8407000", 14473 => x"45a10005", 14474 => x"34010042",
    14475 => x"45a10003", 14476 => x"34010010", 14477 => x"5da10034",
    14478 => x"21cb0002", 14479 => x"5d60000f", 14480 => x"b9800800",
    14481 => x"fbfffef0", 14482 => x"29810000", 14483 => x"34020044",
    14484 => x"21ce0001", 14485 => x"fbfffe1b", 14486 => x"34010000",
    14487 => x"5dcb002d", 14488 => x"780b0001", 14489 => x"396b4d40",
    14490 => x"29620004", 14491 => x"29810000", 14492 => x"d8400000",
    14493 => x"4420fffd", 14494 => x"b9800800", 14495 => x"fbfffee2",
    14496 => x"29810000", 14497 => x"780b0001", 14498 => x"340200be",
    14499 => x"396b6a6c", 14500 => x"fbfffe0c", 14501 => x"356e0008",
    14502 => x"e0000005", 14503 => x"29810000", 14504 => x"fbfffe25",
    14505 => x"31610000", 14506 => x"356b0001", 14507 => x"5d6efffc",
    14508 => x"78020001", 14509 => x"38426a6c", 14510 => x"40410001",
    14511 => x"40430000", 14512 => x"3c210008", 14513 => x"b8230800",
    14514 => x"34030028", 14515 => x"dc200800", 14516 => x"45a3000b",
    14517 => x"34030042", 14518 => x"45a30009", 14519 => x"34030010",
    14520 => x"5da3000b", 14521 => x"40420006", 14522 => x"3c21000f",
    14523 => x"3c42000c", 14524 => x"3421c000", 14525 => x"b8220800",
    14526 => x"e0000006", 14527 => x"3c21000c", 14528 => x"e0000004",
    14529 => x"78018000", 14530 => x"e0000002", 14531 => x"34010000",
    14532 => x"2b9d0004", 14533 => x"2b8b0014", 14534 => x"2b8c0010",
    14535 => x"2b8d000c", 14536 => x"2b8e0008", 14537 => x"379c0014",
    14538 => x"c3a00000", 14539 => x"379cfffc", 14540 => x"5b9d0004",
    14541 => x"34030000", 14542 => x"b8202000", 14543 => x"34090028",
    14544 => x"34080042", 14545 => x"34070010", 14546 => x"34060008",
    14547 => x"40850017", 14548 => x"44a90003", 14549 => x"44a80002",
    14550 => x"5ca70006", 14551 => x"3c630004", 14552 => x"34630008",
    14553 => x"b4230800", 14554 => x"fbffffa5", 14555 => x"e0000005",
    14556 => x"34630001", 14557 => x"34840010", 14558 => x"5c66fff5",
    14559 => x"78018000", 14560 => x"2b9d0004", 14561 => x"379c0004",
    14562 => x"c3a00000", 14563 => x"379cffe0", 14564 => x"5b8b0020",
    14565 => x"5b8c001c", 14566 => x"5b8d0018", 14567 => x"5b8e0014",
    14568 => x"5b8f0010", 14569 => x"5b90000c", 14570 => x"5b910008",
    14571 => x"5b9d0004", 14572 => x"b8205800", 14573 => x"b8408800",
    14574 => x"b8608000", 14575 => x"b8806000", 14576 => x"fbfffe91",
    14577 => x"29610000", 14578 => x"3402000f", 14579 => x"222e00ff",
    14580 => x"fbfffdbc", 14581 => x"29610000", 14582 => x"b9c01000",
    14583 => x"2231ff00", 14584 => x"fbfffdb8", 14585 => x"16310008",
    14586 => x"29610000", 14587 => x"ba201000", 14588 => x"340d0000",
    14589 => x"fbfffdb3", 14590 => x"e0000006", 14591 => x"b60d1000",
    14592 => x"29610000", 14593 => x"40420000", 14594 => x"35ad0001",
    14595 => x"fbfffdad", 14596 => x"498dfffb", 14597 => x"b9600800",
    14598 => x"fbfffe7b", 14599 => x"29610000", 14600 => x"340200aa",
    14601 => x"fbfffda7", 14602 => x"29610000", 14603 => x"fbfffdc2",
    14604 => x"b8207800", 14605 => x"5c2e0022", 14606 => x"29610000",
    14607 => x"fbfffdbe", 14608 => x"b8207000", 14609 => x"5c310020",
    14610 => x"29610000", 14611 => x"340d0000", 14612 => x"fbfffdb9",
    14613 => x"b8208800", 14614 => x"e0000007", 14615 => x"29610000",
    14616 => x"fbfffdb5", 14617 => x"b60d1000", 14618 => x"40420000",
    14619 => x"5c220018", 14620 => x"35ad0001", 14621 => x"498dfffa",
    14622 => x"b9600800", 14623 => x"fbfffe62", 14624 => x"29610000",
    14625 => x"34020055", 14626 => x"fbfffd8e", 14627 => x"29610000",
    14628 => x"b9e01000", 14629 => x"fbfffd8b", 14630 => x"29610000",
    14631 => x"b9c01000", 14632 => x"fbfffd88", 14633 => x"29610000",
    14634 => x"ba201000", 14635 => x"fbfffd85", 14636 => x"34012710",
    14637 => x"fbffedc1", 14638 => x"e0000006", 14639 => x"340cffff",
    14640 => x"e0000004", 14641 => x"340cfffe", 14642 => x"e0000002",
    14643 => x"340cfffd", 14644 => x"b9800800", 14645 => x"2b9d0004",
    14646 => x"2b8b0020", 14647 => x"2b8c001c", 14648 => x"2b8d0018",
    14649 => x"2b8e0014", 14650 => x"2b8f0010", 14651 => x"2b90000c",
    14652 => x"2b910008", 14653 => x"379c0020", 14654 => x"c3a00000",
    14655 => x"379cffe4", 14656 => x"5b8b001c", 14657 => x"5b8c0018",
    14658 => x"5b8d0014", 14659 => x"5b8e0010", 14660 => x"5b8f000c",
    14661 => x"5b900008", 14662 => x"5b9d0004", 14663 => x"b8208000",
    14664 => x"2041001f", 14665 => x"b8405800", 14666 => x"b8607000",
    14667 => x"b8806000", 14668 => x"340d0000", 14669 => x"44200030",
    14670 => x"3441ffff", 14671 => x"b4240800", 14672 => x"1422001f",
    14673 => x"b8807800", 14674 => x"0042001b", 14675 => x"b4410800",
    14676 => x"1562001f", 14677 => x"14210005", 14678 => x"0042001b",
    14679 => x"b44b1000", 14680 => x"14420005", 14681 => x"4422000c",
    14682 => x"78010001", 14683 => x"38213d38", 14684 => x"28220000",
    14685 => x"a1621000", 14686 => x"4c400005", 14687 => x"3442ffff",
    14688 => x"3401ffe0", 14689 => x"b8411000", 14690 => x"34420001",
    14691 => x"340f0020", 14692 => x"c9e27800", 14693 => x"ba000800",
    14694 => x"b9601000", 14695 => x"b9c01800", 14696 => x"b9e02000",
    14697 => x"fbffff7a", 14698 => x"b8206800", 14699 => x"48010016",
    14700 => x"b5cf7000", 14701 => x"b56f5800", 14702 => x"c98f6000",
    14703 => x"e000000e", 14704 => x"b9802000", 14705 => x"4dec0002",
    14706 => x"34040020", 14707 => x"ba000800", 14708 => x"b9601000",
    14709 => x"b9c01800", 14710 => x"fbffff6d", 14711 => x"48010009",
    14712 => x"b5a16800", 14713 => x"35ce0020", 14714 => x"356b0020",
    14715 => x"358cffe0", 14716 => x"e0000002", 14717 => x"340f0020",
    14718 => x"4980fff2", 14719 => x"e0000002", 14720 => x"b8206800",
    14721 => x"b9a00800", 14722 => x"2b9d0004", 14723 => x"2b8b001c",
    14724 => x"2b8c0018", 14725 => x"2b8d0014", 14726 => x"2b8e0010",
    14727 => x"2b8f000c", 14728 => x"2b900008", 14729 => x"379c001c",
    14730 => x"c3a00000", 14731 => x"379cffec", 14732 => x"5b8b0014",
    14733 => x"5b8c0010", 14734 => x"5b8d000c", 14735 => x"5b8e0008",
    14736 => x"5b9d0004", 14737 => x"b8405800", 14738 => x"b8206000",
    14739 => x"b8607000", 14740 => x"b8806800", 14741 => x"fbfffdec",
    14742 => x"29810000", 14743 => x"340200f0", 14744 => x"fbfffd18",
    14745 => x"29810000", 14746 => x"216200ff", 14747 => x"fbfffd15",
    14748 => x"2162ff00", 14749 => x"29810000", 14750 => x"00420008",
    14751 => x"340b0000", 14752 => x"fbfffd10", 14753 => x"e0000006",
    14754 => x"29810000", 14755 => x"fbfffd2a", 14756 => x"b5cb1000",
    14757 => x"30410000", 14758 => x"356b0001", 14759 => x"49abfffb",
    14760 => x"b9a00800", 14761 => x"2b9d0004", 14762 => x"2b8b0014",
    14763 => x"2b8c0010", 14764 => x"2b8d000c", 14765 => x"2b8e0008",
    14766 => x"379c0014", 14767 => x"c3a00000", 14768 => x"379cfffc",
    14769 => x"5b9d0004", 14770 => x"34050000", 14771 => x"b8203000",
    14772 => x"34080043", 14773 => x"34070008", 14774 => x"40c90017",
    14775 => x"5d280006", 14776 => x"3ca50004", 14777 => x"34a50008",
    14778 => x"b4250800", 14779 => x"fbffffd0", 14780 => x"e0000005",
    14781 => x"34a50001", 14782 => x"34c60010", 14783 => x"5ca7fff7",
    14784 => x"3401ffff", 14785 => x"2b9d0004", 14786 => x"379c0004",
    14787 => x"c3a00000", 14788 => x"379cfffc", 14789 => x"5b9d0004",
    14790 => x"34050000", 14791 => x"b8203000", 14792 => x"34080043",
    14793 => x"34070008", 14794 => x"40c90017", 14795 => x"5d280006",
    14796 => x"3ca50004", 14797 => x"34a50008", 14798 => x"b4250800",
    14799 => x"fbffff70", 14800 => x"e0000005", 14801 => x"34a50001",
    14802 => x"34c60010", 14803 => x"5ca7fff7", 14804 => x"3401ffff",
    14805 => x"2b9d0004", 14806 => x"379c0004", 14807 => x"c3a00000",
    14808 => x"78010001", 14809 => x"38216da4", 14810 => x"28220000",
    14811 => x"78010001", 14812 => x"38216dc4", 14813 => x"58220000",
    14814 => x"340103c6", 14815 => x"58410004", 14816 => x"c3a00000",
    14817 => x"c3a00000", 14818 => x"379cfff8", 14819 => x"5b8b0008",
    14820 => x"5b9d0004", 14821 => x"b8205800", 14822 => x"3401000a",
    14823 => x"5d610003", 14824 => x"3401000d", 14825 => x"fbfffff9",
    14826 => x"78020001", 14827 => x"38426dc4", 14828 => x"28420000",
    14829 => x"28410000", 14830 => x"20210001", 14831 => x"5c20fffe",
    14832 => x"584b0008", 14833 => x"2b9d0004", 14834 => x"2b8b0008",
    14835 => x"379c0008", 14836 => x"c3a00000", 14837 => x"379cfff4",
    14838 => x"5b8b000c", 14839 => x"5b8c0008", 14840 => x"5b9d0004",
    14841 => x"b8206000", 14842 => x"b8205800", 14843 => x"e0000004",
    14844 => x"b8400800", 14845 => x"356b0001", 14846 => x"fbffffe4",
    14847 => x"41620000", 14848 => x"5c40fffc", 14849 => x"c96c0800",
    14850 => x"2b9d0004", 14851 => x"2b8b000c", 14852 => x"2b8c0008",
    14853 => x"379c000c", 14854 => x"c3a00000", 14855 => x"78010001",
    14856 => x"38216dc4", 14857 => x"28220000", 14858 => x"3401ffff",
    14859 => x"28430000", 14860 => x"20630002", 14861 => x"44600003",
    14862 => x"2841000c", 14863 => x"202100ff", 14864 => x"c3a00000",
    14865 => x"28250008", 14866 => x"28240000", 14867 => x"28260004",
    14868 => x"b4451800", 14869 => x"88642000", 14870 => x"5822001c",
    14871 => x"88461000", 14872 => x"b4821000", 14873 => x"2824000c",
    14874 => x"1442000c", 14875 => x"b4442000", 14876 => x"28220014",
    14877 => x"4c820005", 14878 => x"28240010", 14879 => x"44800008",
    14880 => x"4ca3000b", 14881 => x"e0000006", 14882 => x"28220018",
    14883 => x"4c440006", 14884 => x"28240010", 14885 => x"44800002",
    14886 => x"4c650005", 14887 => x"58230008", 14888 => x"e0000003",
    14889 => x"58230008", 14890 => x"b8801000", 14891 => x"58220020",
    14892 => x"b8400800", 14893 => x"c3a00000", 14894 => x"2822000c",
    14895 => x"58200008", 14896 => x"58220020", 14897 => x"c3a00000",
    14898 => x"379cfff8", 14899 => x"5b8b0008", 14900 => x"5b9d0004",
    14901 => x"b8205800", 14902 => x"58200014", 14903 => x"b8400800",
    14904 => x"f80009ef", 14905 => x"2963000c", 14906 => x"29620000",
    14907 => x"4823000b", 14908 => x"29610004", 14909 => x"4c410003",
    14910 => x"34420001", 14911 => x"59620000", 14912 => x"29620000",
    14913 => x"5c410011", 14914 => x"34010001", 14915 => x"59610014",
    14916 => x"59610010", 14917 => x"e000000e", 14918 => x"29610008",
    14919 => x"4c220003", 14920 => x"3442ffff", 14921 => x"59620000",
    14922 => x"29620000", 14923 => x"5c410007", 14924 => x"34010001",
    14925 => x"59610014", 14926 => x"59600000", 14927 => x"59600010",
    14928 => x"3401ffff", 14929 => x"e0000002", 14930 => x"29610010",
    14931 => x"2b9d0004", 14932 => x"2b8b0008", 14933 => x"379c0008",
    14934 => x"c3a00000", 14935 => x"58200010", 14936 => x"58200000",
    14937 => x"58200014", 14938 => x"c3a00000", 14939 => x"379cfff4",
    14940 => x"5b8b000c", 14941 => x"5b8c0008", 14942 => x"5b9d0004",
    14943 => x"b8205800", 14944 => x"b8406000", 14945 => x"78020001",
    14946 => x"34010000", 14947 => x"384238b0", 14948 => x"b9601800",
    14949 => x"b9802000", 14950 => x"fbffc61f", 14951 => x"78010001",
    14952 => x"38216db0", 14953 => x"28220000", 14954 => x"484b0013",
    14955 => x"78050001", 14956 => x"38a56d08", 14957 => x"c9621000",
    14958 => x"45800007", 14959 => x"28a10000", 14960 => x"34040001",
    14961 => x"bc821000", 14962 => x"28230028", 14963 => x"b8431000",
    14964 => x"e0000007", 14965 => x"28a10000", 14966 => x"34040001",
    14967 => x"bc821000", 14968 => x"28230028", 14969 => x"a4401000",
    14970 => x"a0431000", 14971 => x"58220028", 14972 => x"e0000011",
    14973 => x"78050001", 14974 => x"38a56d08", 14975 => x"45800007",
    14976 => x"28a10000", 14977 => x"34020001", 14978 => x"bc4b1000",
    14979 => x"28230024", 14980 => x"b8431000", 14981 => x"e0000007",
    14982 => x"28a10000", 14983 => x"34020001", 14984 => x"bc4b1000",
    14985 => x"28230024", 14986 => x"a4401000", 14987 => x"a0431000",
    14988 => x"58220024", 14989 => x"78010001", 14990 => x"38216d08",
    14991 => x"28210000", 14992 => x"78020001", 14993 => x"78030001",
    14994 => x"28250028", 14995 => x"28260024", 14996 => x"384238c4",
    14997 => x"34010000", 14998 => x"386340a0", 14999 => x"b9602000",
    15000 => x"fbffc5ed", 15001 => x"2b9d0004", 15002 => x"2b8b000c",
    15003 => x"2b8c0008", 15004 => x"379c000c", 15005 => x"c3a00000",
    15006 => x"379cfff0", 15007 => x"5b8b0010", 15008 => x"5b8c000c",
    15009 => x"5b8d0008", 15010 => x"5b9d0004", 15011 => x"b8406800",
    15012 => x"b8606000", 15013 => x"34020000", 15014 => x"34030028",
    15015 => x"b8205800", 15016 => x"f8000a22", 15017 => x"b9600800",
    15018 => x"b9a01000", 15019 => x"34030014", 15020 => x"f80009a0",
    15021 => x"596c0014", 15022 => x"2b9d0004", 15023 => x"2b8b0010",
    15024 => x"2b8c000c", 15025 => x"2b8d0008", 15026 => x"379c0010",
    15027 => x"c3a00000", 15028 => x"b8201800", 15029 => x"e0000004",
    15030 => x"28840000", 15031 => x"34630008", 15032 => x"44820006",
    15033 => x"28610004", 15034 => x"b8602000", 15035 => x"5c20fffb",
    15036 => x"78010001", 15037 => x"382138e8", 15038 => x"c3a00000",
    15039 => x"78020001", 15040 => x"38426d08", 15041 => x"28420000",
    15042 => x"b8201800", 15043 => x"34010000", 15044 => x"28440008",
    15045 => x"20840002", 15046 => x"4480000c", 15047 => x"34040002",
    15048 => x"58440008", 15049 => x"78060001", 15050 => x"28420010",
    15051 => x"38c63d3c", 15052 => x"28c40000", 15053 => x"3445ff9b",
    15054 => x"54a40004", 15055 => x"08420064", 15056 => x"34010001",
    15057 => x"58620000", 15058 => x"c3a00000", 15059 => x"379cfff0",
    15060 => x"5b8b0010", 15061 => x"5b8c000c", 15062 => x"5b8d0008",
    15063 => x"5b9d0004", 15064 => x"780b0001", 15065 => x"b8206000",
    15066 => x"78010001", 15067 => x"396b6db0", 15068 => x"38216da8",
    15069 => x"28210000", 15070 => x"296d0000", 15071 => x"b42d6800",
    15072 => x"29810000", 15073 => x"b9a01000", 15074 => x"f8000116",
    15075 => x"29810004", 15076 => x"29630000", 15077 => x"b9a01000",
    15078 => x"f800019b", 15079 => x"5980000c", 15080 => x"59800008",
    15081 => x"2b9d0004", 15082 => x"2b8b0010", 15083 => x"2b8c000c",
    15084 => x"2b8d0008", 15085 => x"379c0010", 15086 => x"c3a00000",
    15087 => x"379cfff8", 15088 => x"5b8b0008", 15089 => x"5b9d0004",
    15090 => x"b8205800", 15091 => x"28210000", 15092 => x"f800016e",
    15093 => x"78010001", 15094 => x"38216d08", 15095 => x"28210000",
    15096 => x"34020001", 15097 => x"34030009", 15098 => x"58220004",
    15099 => x"5963000c", 15100 => x"78030001", 15101 => x"38633d40",
    15102 => x"59620008", 15103 => x"28620000", 15104 => x"5822004c",
    15105 => x"2b9d0004", 15106 => x"2b8b0008", 15107 => x"379c0008",
    15108 => x"c3a00000", 15109 => x"b8201000", 15110 => x"28210000",
    15111 => x"2823004c", 15112 => x"34010000", 15113 => x"44600016",
    15114 => x"28430004", 15115 => x"28630038", 15116 => x"44600013",
    15117 => x"78030001", 15118 => x"38636d08", 15119 => x"28630000",
    15120 => x"28640004", 15121 => x"20840004", 15122 => x"4480000d",
    15123 => x"28630004", 15124 => x"20630008", 15125 => x"5c60000a",
    15126 => x"2842000c", 15127 => x"3403000a", 15128 => x"34010001",
    15129 => x"54430006", 15130 => x"78010001", 15131 => x"3c420002",
    15132 => x"382140dc", 15133 => x"b4220800", 15134 => x"28210000",
    15135 => x"c3a00000", 15136 => x"379cfff0", 15137 => x"5b8b000c",
    15138 => x"5b8c0008", 15139 => x"5b9d0004", 15140 => x"2822000c",
    15141 => x"b8205800", 15142 => x"34010009", 15143 => x"3442ffff",
    15144 => x"544100a9", 15145 => x"78010001", 15146 => x"3c420002",
    15147 => x"382140b4", 15148 => x"b4220800", 15149 => x"28210000",
    15150 => x"c0200000", 15151 => x"78010001", 15152 => x"38216d08",
    15153 => x"28210000", 15154 => x"28220004", 15155 => x"20420008",
    15156 => x"5c40009d", 15157 => x"28230004", 15158 => x"78028000",
    15159 => x"b8621000", 15160 => x"58220004", 15161 => x"3401000a",
    15162 => x"e0000096", 15163 => x"78010001", 15164 => x"38216d08",
    15165 => x"28210000", 15166 => x"78040001", 15167 => x"38843d20",
    15168 => x"28230004", 15169 => x"28820000", 15170 => x"a0621000",
    15171 => x"58220004", 15172 => x"28220004", 15173 => x"20420008",
    15174 => x"5c400089", 15175 => x"28210004", 15176 => x"20210004",
    15177 => x"44220088", 15178 => x"34010001", 15179 => x"e0000085",
    15180 => x"29610000", 15181 => x"2821004c", 15182 => x"44200083",
    15183 => x"fbffc523", 15184 => x"29610004", 15185 => x"f800015e",
    15186 => x"fbffc529", 15187 => x"34010008", 15188 => x"e000007c",
    15189 => x"78010001", 15190 => x"38216d08", 15191 => x"28210000",
    15192 => x"34020002", 15193 => x"58220008", 15194 => x"29610000",
    15195 => x"2821004c", 15196 => x"44200075", 15197 => x"29610004",
    15198 => x"28210038", 15199 => x"44200072", 15200 => x"78010001",
    15201 => x"38216d0c", 15202 => x"28210000", 15203 => x"340300a2",
    15204 => x"58230000", 15205 => x"34030003", 15206 => x"58230010",
    15207 => x"34030001", 15208 => x"5823001c", 15209 => x"5962000c",
    15210 => x"78020001", 15211 => x"34010000", 15212 => x"384238f4",
    15213 => x"e0000017", 15214 => x"78010001", 15215 => x"38216d0c",
    15216 => x"28210000", 15217 => x"2822001c", 15218 => x"20420001",
    15219 => x"4440005e", 15220 => x"34020002", 15221 => x"5822001c",
    15222 => x"fbfff630", 15223 => x"342107d0", 15224 => x"59610010",
    15225 => x"34010003", 15226 => x"e0000056", 15227 => x"fbfff62b",
    15228 => x"29620010", 15229 => x"54410054", 15230 => x"34010007",
    15231 => x"5961000c", 15232 => x"78020001", 15233 => x"5960001c",
    15234 => x"34010000", 15235 => x"38423908", 15236 => x"fbffc501",
    15237 => x"e000004c", 15238 => x"37810010", 15239 => x"fbffff38",
    15240 => x"44200049", 15241 => x"78030001", 15242 => x"38633cfc",
    15243 => x"2b810010", 15244 => x"28620000", 15245 => x"f800083e",
    15246 => x"3802c34f", 15247 => x"e8221000", 15248 => x"5b810010",
    15249 => x"64210000", 15250 => x"b8410800", 15251 => x"44200005",
    15252 => x"34010064", 15253 => x"59610014", 15254 => x"3401ff9c",
    15255 => x"e0000003", 15256 => x"59600014", 15257 => x"34010064",
    15258 => x"59610018", 15259 => x"29630014", 15260 => x"29640018",
    15261 => x"78020001", 15262 => x"34010000", 15263 => x"38423920",
    15264 => x"fbffc4e5", 15265 => x"34010004", 15266 => x"e000002e",
    15267 => x"29610004", 15268 => x"f80001e9", 15269 => x"b8206000",
    15270 => x"5c20002b", 15271 => x"37810010", 15272 => x"fbffff17",
    15273 => x"442c0028", 15274 => x"78040001", 15275 => x"38843cfc",
    15276 => x"2b810010", 15277 => x"28820000", 15278 => x"f800081d",
    15279 => x"29620014", 15280 => x"5b810010", 15281 => x"44220009",
    15282 => x"2961001c", 15283 => x"29620018", 15284 => x"b4410800",
    15285 => x"5961001c", 15286 => x"29610004", 15287 => x"2962001c",
    15288 => x"f80001b3", 15289 => x"e0000018", 15290 => x"29620014",
    15291 => x"5c220016", 15292 => x"2961001c", 15293 => x"34217530",
    15294 => x"5961001c", 15295 => x"29610004", 15296 => x"2962001c",
    15297 => x"f80001aa", 15298 => x"34010005", 15299 => x"e000000d",
    15300 => x"29610004", 15301 => x"f80001c8", 15302 => x"5c20000b",
    15303 => x"78020001", 15304 => x"38423940", 15305 => x"fbffc4bc",
    15306 => x"34010006", 15307 => x"e0000005", 15308 => x"b9600800",
    15309 => x"fbffff38", 15310 => x"5c200003", 15311 => x"34010009",
    15312 => x"5961000c", 15313 => x"2b9d0004", 15314 => x"2b8b000c",
    15315 => x"2b8c0008", 15316 => x"379c0010", 15317 => x"c3a00000",
    15318 => x"78040001", 15319 => x"64630000", 15320 => x"38846d08",
    15321 => x"28850000", 15322 => x"c8031800", 15323 => x"78048000",
    15324 => x"78060001", 15325 => x"a0641800", 15326 => x"38c63d44",
    15327 => x"b4641800", 15328 => x"28c40000", 15329 => x"3c210018",
    15330 => x"a0441000", 15331 => x"b8410800", 15332 => x"b8231800",
    15333 => x"58a3004c", 15334 => x"c3a00000", 15335 => x"78040001",
    15336 => x"64630000", 15337 => x"38846d08", 15338 => x"28850000",
    15339 => x"c8031800", 15340 => x"78048000", 15341 => x"78060001",
    15342 => x"a0641800", 15343 => x"38c63d44", 15344 => x"b4641800",
    15345 => x"28c40000", 15346 => x"3c210018", 15347 => x"a0441000",
    15348 => x"b8410800", 15349 => x"b8231800", 15350 => x"58a3004c",
    15351 => x"c3a00000", 15352 => x"34030005", 15353 => x"5823002c",
    15354 => x"3803fffb", 15355 => x"58230030", 15356 => x"3403ff6a",
    15357 => x"5823001c", 15358 => x"3403fffe", 15359 => x"58230018",
    15360 => x"34030001", 15361 => x"58230028", 15362 => x"340300c8",
    15363 => x"58230048", 15364 => x"34032710", 15365 => x"58230040",
    15366 => x"34030064", 15367 => x"58230044", 15368 => x"5822000c",
    15369 => x"58200014", 15370 => x"c3a00000", 15371 => x"379cfff0",
    15372 => x"5b8b0010", 15373 => x"5b8c000c", 15374 => x"5b8d0008",
    15375 => x"5b9d0004", 15376 => x"b8205800", 15377 => x"2821000c",
    15378 => x"b8406800", 15379 => x"340c0000", 15380 => x"5c610047",
    15381 => x"34010022", 15382 => x"34030000", 15383 => x"fbffffbf",
    15384 => x"29620004", 15385 => x"34010025", 15386 => x"34030000",
    15387 => x"fbffffbb", 15388 => x"29610008", 15389 => x"4c200004",
    15390 => x"596d0004", 15391 => x"596d0008", 15392 => x"e000003b",
    15393 => x"4da10005", 15394 => x"29620000", 15395 => x"78010040",
    15396 => x"b4410800", 15397 => x"59610000", 15398 => x"29630000",
    15399 => x"78050001", 15400 => x"29620004", 15401 => x"38a53d48",
    15402 => x"28a10000", 15403 => x"b5a32000", 15404 => x"c8826000",
    15405 => x"482c0006", 15406 => x"78050001", 15407 => x"38a53d4c",
    15408 => x"28a10000", 15409 => x"49810002", 15410 => x"e0000002",
    15411 => x"b8206000", 15412 => x"78050001", 15413 => x"38a53d50",
    15414 => x"28a10000", 15415 => x"4c240006", 15416 => x"4c220005",
    15417 => x"c8611800", 15418 => x"c8410800", 15419 => x"59630000",
    15420 => x"59610004", 15421 => x"29610004", 15422 => x"b9801000",
    15423 => x"596d0008", 15424 => x"34214000", 15425 => x"59610004",
    15426 => x"35610018", 15427 => x"fbfffdce", 15428 => x"78030001",
    15429 => x"38636d08", 15430 => x"29620010", 15431 => x"b8206800",
    15432 => x"28610000", 15433 => x"34030000", 15434 => x"582d0040",
    15435 => x"34410001", 15436 => x"59610010", 15437 => x"34010026",
    15438 => x"fbffff88", 15439 => x"34010020", 15440 => x"b9a01000",
    15441 => x"34030000", 15442 => x"fbffff84", 15443 => x"b9801000",
    15444 => x"34010021", 15445 => x"34030001", 15446 => x"fbffff80",
    15447 => x"b9801000", 15448 => x"3561003c", 15449 => x"fbfffdd9",
    15450 => x"7c2c0000", 15451 => x"b9800800", 15452 => x"2b9d0004",
    15453 => x"2b8b0010", 15454 => x"2b8c000c", 15455 => x"2b8d0008",
    15456 => x"379c0010", 15457 => x"c3a00000", 15458 => x"379cfff8",
    15459 => x"5b8b0008", 15460 => x"5b9d0004", 15461 => x"b8205800",
    15462 => x"2821002c", 15463 => x"59600004", 15464 => x"59600000",
    15465 => x"59610024", 15466 => x"3401ffff", 15467 => x"59610008",
    15468 => x"59600010", 15469 => x"35610018", 15470 => x"fbfffdc0",
    15471 => x"3561003c", 15472 => x"fbfffde7", 15473 => x"78020001",
    15474 => x"35610054", 15475 => x"34030010", 15476 => x"38424108",
    15477 => x"fbfffe29", 15478 => x"2961000c", 15479 => x"34020001",
    15480 => x"fbfffde3", 15481 => x"34010024", 15482 => x"34020001",
    15483 => x"34030001", 15484 => x"fbffff5a", 15485 => x"2b9d0004",
    15486 => x"2b8b0008", 15487 => x"379c0008", 15488 => x"c3a00000",
    15489 => x"379cfff8", 15490 => x"5b8b0008", 15491 => x"5b9d0004",
    15492 => x"b8205800", 15493 => x"34010005", 15494 => x"59610018",
    15495 => x"3801fffa", 15496 => x"5961001c", 15497 => x"34010001",
    15498 => x"59610014", 15499 => x"34017530", 15500 => x"59610010",
    15501 => x"3401fbb4", 15502 => x"59610008", 15503 => x"3401ffe2",
    15504 => x"59610004", 15505 => x"340104b0", 15506 => x"59610034",
    15507 => x"340103e8", 15508 => x"5961002c", 15509 => x"34010064",
    15510 => x"59610030", 15511 => x"78010001", 15512 => x"38216db0",
    15513 => x"28250000", 15514 => x"b8403000", 15515 => x"59620070",
    15516 => x"c8652800", 15517 => x"78020001", 15518 => x"b8602000",
    15519 => x"59650080", 15520 => x"38423954", 15521 => x"59630074",
    15522 => x"5960007c", 15523 => x"b8c01800", 15524 => x"59600084",
    15525 => x"34010000", 15526 => x"fbffc3df", 15527 => x"35610004",
    15528 => x"fbfffd86", 15529 => x"35610028", 15530 => x"fbfffdad",
    15531 => x"2b9d0004", 15532 => x"2b8b0008", 15533 => x"379c0008",
    15534 => x"c3a00000", 15535 => x"379cfff8", 15536 => x"5b8b0008",
    15537 => x"5b9d0004", 15538 => x"b8205800", 15539 => x"29630080",
    15540 => x"78020001", 15541 => x"3842396c", 15542 => x"34010000",
    15543 => x"fbffc3ce", 15544 => x"3401ffff", 15545 => x"59610048",
    15546 => x"5961004c", 15547 => x"59610050", 15548 => x"59610054",
    15549 => x"34010001", 15550 => x"59610084", 15551 => x"59600044",
    15552 => x"35610004", 15553 => x"59600040", 15554 => x"59600058",
    15555 => x"5960005c", 15556 => x"59600060", 15557 => x"59600068",
    15558 => x"5960006c", 15559 => x"59600078", 15560 => x"fbfffd66",
    15561 => x"35610028", 15562 => x"fbfffd8d", 15563 => x"29610070",
    15564 => x"34020001", 15565 => x"fbfffd8e", 15566 => x"29610074",
    15567 => x"34020001", 15568 => x"fbfffd8b", 15569 => x"34010004",
    15570 => x"34020001", 15571 => x"34030001", 15572 => x"fbffff13",
    15573 => x"2b9d0004", 15574 => x"2b8b0008", 15575 => x"379c0008",
    15576 => x"c3a00000", 15577 => x"379cfff8", 15578 => x"5b8b0008",
    15579 => x"5b9d0004", 15580 => x"b8205800", 15581 => x"28210074",
    15582 => x"34020000", 15583 => x"fbfffd7c", 15584 => x"59600084",
    15585 => x"2b9d0004", 15586 => x"2b8b0008", 15587 => x"379c0008",
    15588 => x"c3a00000", 15589 => x"379cfff0", 15590 => x"5b8b0010",
    15591 => x"5b8c000c", 15592 => x"5b8d0008", 15593 => x"5b9d0004",
    15594 => x"28240084", 15595 => x"b8205800", 15596 => x"34010001",
    15597 => x"44800078", 15598 => x"29610070", 15599 => x"5c610002",
    15600 => x"59620048", 15601 => x"29610074", 15602 => x"5c610002",
    15603 => x"5962004c", 15604 => x"29610048", 15605 => x"48010009",
    15606 => x"29620050", 15607 => x"48020006", 15608 => x"4c220005",
    15609 => x"29630040", 15610 => x"78020040", 15611 => x"b4621000",
    15612 => x"59620040", 15613 => x"59610050", 15614 => x"2961004c",
    15615 => x"48010009", 15616 => x"29620054", 15617 => x"48020006",
    15618 => x"4c220005", 15619 => x"29630044", 15620 => x"78020040",
    15621 => x"b4621000", 15622 => x"59620044", 15623 => x"59610054",
    15624 => x"29630048", 15625 => x"34010000", 15626 => x"4803005b",
    15627 => x"2962004c", 15628 => x"48020059", 15629 => x"296c0040",
    15630 => x"29610038", 15631 => x"b46c1800", 15632 => x"296c0044",
    15633 => x"c8621000", 15634 => x"c84c6000", 15635 => x"44200006",
    15636 => x"218c3fff", 15637 => x"21812000", 15638 => x"44200003",
    15639 => x"3401c000", 15640 => x"b9816000", 15641 => x"b9801000",
    15642 => x"35610004", 15643 => x"fbfffcf6", 15644 => x"29620080",
    15645 => x"78030001", 15646 => x"38636d08", 15647 => x"2042000f",
    15648 => x"b8206800", 15649 => x"3c420010", 15650 => x"28610000",
    15651 => x"21a3ffff", 15652 => x"b8621000", 15653 => x"58220044",
    15654 => x"29630040", 15655 => x"29620048", 15656 => x"34010005",
    15657 => x"b4621000", 15658 => x"34030000", 15659 => x"fbfffebc",
    15660 => x"29630044", 15661 => x"2962004c", 15662 => x"34010002",
    15663 => x"b4621000", 15664 => x"34030000", 15665 => x"fbfffeb6",
    15666 => x"34010001", 15667 => x"b9801000", 15668 => x"34030000",
    15669 => x"fbfffeb2", 15670 => x"29620078", 15671 => x"34030000",
    15672 => x"34410001", 15673 => x"59610078", 15674 => x"34010006",
    15675 => x"fbfffeac", 15676 => x"34010000", 15677 => x"b9a01000",
    15678 => x"34030001", 15679 => x"fbfffea8", 15680 => x"78020001",
    15681 => x"3401ffff", 15682 => x"38423d54", 15683 => x"5961004c",
    15684 => x"59610048", 15685 => x"29630040", 15686 => x"28410000",
    15687 => x"4c23000a", 15688 => x"29620044", 15689 => x"4c220008",
    15690 => x"78040001", 15691 => x"38843d58", 15692 => x"28810000",
    15693 => x"b4611800", 15694 => x"b4410800", 15695 => x"59630040",
    15696 => x"59610044", 15697 => x"29610038", 15698 => x"4420000f",
    15699 => x"2961006c", 15700 => x"29620068", 15701 => x"4c220006",
    15702 => x"34210001", 15703 => x"5961006c", 15704 => x"29610040",
    15705 => x"3421ffff", 15706 => x"e0000006", 15707 => x"4c410006",
    15708 => x"3421ffff", 15709 => x"5961006c", 15710 => x"29610040",
    15711 => x"34210001", 15712 => x"59610040", 15713 => x"35610028",
    15714 => x"b9801000", 15715 => x"fbfffccf", 15716 => x"7c210000",
    15717 => x"2b9d0004", 15718 => x"2b8b0010", 15719 => x"2b8c000c",
    15720 => x"2b8d0008", 15721 => x"379c0010", 15722 => x"c3a00000",
    15723 => x"379cfff0", 15724 => x"5b8b0008", 15725 => x"5b9d0004",
    15726 => x"b8205800", 15727 => x"1443001f", 15728 => x"3781000c",
    15729 => x"4802000b", 15730 => x"00440012", 15731 => x"3c63000e",
    15732 => x"3c42000e", 15733 => x"b8641800", 15734 => x"5b820010",
    15735 => x"34021f40", 15736 => x"5b83000c", 15737 => x"fbffcbec",
    15738 => x"2b820010", 15739 => x"e0000009", 15740 => x"0842c000",
    15741 => x"5b820010", 15742 => x"1442001f", 15743 => x"5b82000c",
    15744 => x"34021f40", 15745 => x"fbffcbe4", 15746 => x"2b820010",
    15747 => x"c8021000", 15748 => x"0041001f", 15749 => x"b4221000",
    15750 => x"14420001", 15751 => x"34010000", 15752 => x"59620068",
    15753 => x"2b9d0004", 15754 => x"2b8b0008", 15755 => x"379c0010",
    15756 => x"c3a00000", 15757 => x"28220068", 15758 => x"2821006c",
    15759 => x"fc410800", 15760 => x"c3a00000", 15761 => x"58220004",
    15762 => x"5820001c", 15763 => x"58230008", 15764 => x"5820000c",
    15765 => x"58200010", 15766 => x"58200000", 15767 => x"c3a00000",
    15768 => x"379cfffc", 15769 => x"5b9d0004", 15770 => x"34020001",
    15771 => x"58220000", 15772 => x"58200014", 15773 => x"5820001c",
    15774 => x"5820000c", 15775 => x"58200010", 15776 => x"28210004",
    15777 => x"fbfffcba", 15778 => x"78010001", 15779 => x"38216db0",
    15780 => x"28210000", 15781 => x"34020001", 15782 => x"fbfffcb5",
    15783 => x"2b9d0004", 15784 => x"379c0004", 15785 => x"c3a00000",
    15786 => x"379cffb0", 15787 => x"5b8b0010", 15788 => x"5b8c000c",
    15789 => x"5b8d0008", 15790 => x"5b9d0004", 15791 => x"b8205800",
    15792 => x"b8406000", 15793 => x"b8606800", 15794 => x"37810014",
    15795 => x"34020000", 15796 => x"34030040", 15797 => x"f8000715",
    15798 => x"3401c000", 15799 => x"78040001", 15800 => x"5b810020",
    15801 => x"38846db0", 15802 => x"34014000", 15803 => x"5b810044",
    15804 => x"28810000", 15805 => x"5da10005", 15806 => x"78030001",
    15807 => x"38634d4c", 15808 => x"586c0000", 15809 => x"e0000027",
    15810 => x"3dad0005", 15811 => x"b56d5800", 15812 => x"29610000",
    15813 => x"44200023", 15814 => x"78030001", 15815 => x"38634d4c",
    15816 => x"28610000", 15817 => x"29620010", 15818 => x"c9810800",
    15819 => x"20213fff", 15820 => x"1423000c", 15821 => x"5c400007",
    15822 => x"3c630002", 15823 => x"5961000c", 15824 => x"34010001",
    15825 => x"59630014", 15826 => x"59610010", 15827 => x"e0000015",
    15828 => x"2964000c", 15829 => x"34420001", 15830 => x"b4240800",
    15831 => x"29640014", 15832 => x"b4641800", 15833 => x"3c630002",
    15834 => x"37840050", 15835 => x"b4831800", 15836 => x"2863ffc4",
    15837 => x"59620010", 15838 => x"b4230800", 15839 => x"29630008",
    15840 => x"5961000c", 15841 => x"5c430007", 15842 => x"f80005bc",
    15843 => x"59610018", 15844 => x"34010001", 15845 => x"5961001c",
    15846 => x"5960000c", 15847 => x"59600010", 15848 => x"34010000",
    15849 => x"2b9d0004", 15850 => x"2b8b0010", 15851 => x"2b8c000c",
    15852 => x"2b8d0008", 15853 => x"379c0050", 15854 => x"c3a00000",
    15855 => x"78030001", 15856 => x"38636d08", 15857 => x"5c40000a",
    15858 => x"34040001", 15859 => x"28620000", 15860 => x"bc810800",
    15861 => x"202100ff", 15862 => x"28430020", 15863 => x"3c210010",
    15864 => x"a4200800", 15865 => x"a0230800", 15866 => x"e0000008",
    15867 => x"28620000", 15868 => x"34040001", 15869 => x"bc810800",
    15870 => x"28430020", 15871 => x"202100ff", 15872 => x"3c210010",
    15873 => x"b8230800", 15874 => x"58410020", 15875 => x"c3a00000",
    15876 => x"379cffe0", 15877 => x"5b8b0010", 15878 => x"5b8c000c",
    15879 => x"5b8d0008", 15880 => x"5b9d0004", 15881 => x"b8406000",
    15882 => x"c8231000", 15883 => x"1441001f", 15884 => x"b8605800",
    15885 => x"48010002", 15886 => x"e0000020", 15887 => x"c9836000",
    15888 => x"1583001f", 15889 => x"5c60001d", 15890 => x"4583001c",
    15891 => x"78050001", 15892 => x"38a53d5c", 15893 => x"28a40000",
    15894 => x"3403ffff", 15895 => x"f8000560", 15896 => x"5b81001c",
    15897 => x"5b820020", 15898 => x"3781001c", 15899 => x"b9601000",
    15900 => x"fbffcb49", 15901 => x"78050001", 15902 => x"38a53ccc",
    15903 => x"28a40000", 15904 => x"34030000", 15905 => x"34010000",
    15906 => x"b9801000", 15907 => x"f8000554", 15908 => x"5b810014",
    15909 => x"5b820018", 15910 => x"37810014", 15911 => x"b9601000",
    15912 => x"2b8d0020", 15913 => x"fbffcb3c", 15914 => x"2b810018",
    15915 => x"4da10004", 15916 => x"b9a00800", 15917 => x"e0000002",
    15918 => x"3401ffff", 15919 => x"2b9d0004", 15920 => x"2b8b0010",
    15921 => x"2b8c000c", 15922 => x"2b8d0008", 15923 => x"379c0020",
    15924 => x"c3a00000", 15925 => x"379cfff8", 15926 => x"5b8b0008",
    15927 => x"5b9d0004", 15928 => x"34020001", 15929 => x"44220009",
    15930 => x"34020002", 15931 => x"4422000c", 15932 => x"5c200017",
    15933 => x"78010001", 15934 => x"38216d08", 15935 => x"282b0000",
    15936 => x"356b0018", 15937 => x"e000000a", 15938 => x"78010001",
    15939 => x"38216d08", 15940 => x"282b0000", 15941 => x"356b0014",
    15942 => x"e0000005", 15943 => x"78010001", 15944 => x"38216d08",
    15945 => x"282b0000", 15946 => x"356b001c", 15947 => x"340107d0",
    15948 => x"fbfff35f", 15949 => x"78030001", 15950 => x"38633d14",
    15951 => x"29620000", 15952 => x"28610000", 15953 => x"a0410800",
    15954 => x"e0000002", 15955 => x"34010000", 15956 => x"2b9d0004",
    15957 => x"2b8b0008", 15958 => x"379c0008", 15959 => x"c3a00000",
    15960 => x"379cfff8", 15961 => x"5b8b0008", 15962 => x"5b9d0004",
    15963 => x"78030001", 15964 => x"b8405800", 15965 => x"38636b2c",
    15966 => x"44200007", 15967 => x"3421ffff", 15968 => x"08230090",
    15969 => x"78010001", 15970 => x"38216a78", 15971 => x"b4610800",
    15972 => x"34230144", 15973 => x"b8600800", 15974 => x"b9601000",
    15975 => x"fbffff04", 15976 => x"78010001", 15977 => x"38216a78",
    15978 => x"582b0014", 15979 => x"2b9d0004", 15980 => x"2b8b0008",
    15981 => x"379c0008", 15982 => x"c3a00000", 15983 => x"379cffec",
    15984 => x"5b8b0014", 15985 => x"5b8c0010", 15986 => x"5b8d000c",
    15987 => x"5b8e0008", 15988 => x"5b9d0004", 15989 => x"780c0001",
    15990 => x"780d0001", 15991 => x"b8207000", 15992 => x"340b0000",
    15993 => x"398c6db0", 15994 => x"39ad6cf4", 15995 => x"e000000a",
    15996 => x"29a10000", 15997 => x"942b0800", 15998 => x"20210001",
    15999 => x"44200005", 16000 => x"3d620005", 16001 => x"b5c21000",
    16002 => x"3441025c", 16003 => x"fbffff15", 16004 => x"356b0001",
    16005 => x"29810000", 16006 => x"482bfff6", 16007 => x"2b9d0004",
    16008 => x"2b8b0014", 16009 => x"2b8c0010", 16010 => x"2b8d000c",
    16011 => x"2b8e0008", 16012 => x"379c0014", 16013 => x"c3a00000",
    16014 => x"379cffb8", 16015 => x"5b8b0044", 16016 => x"5b8c0040",
    16017 => x"5b8d003c", 16018 => x"5b8e0038", 16019 => x"5b8f0034",
    16020 => x"5b900030", 16021 => x"5b91002c", 16022 => x"5b920028",
    16023 => x"5b930024", 16024 => x"5b940020", 16025 => x"5b95001c",
    16026 => x"5b960018", 16027 => x"5b970014", 16028 => x"5b980010",
    16029 => x"5b99000c", 16030 => x"5b9b0008", 16031 => x"5b9d0004",
    16032 => x"78010001", 16033 => x"78190001", 16034 => x"38213d44",
    16035 => x"780b0001", 16036 => x"78180001", 16037 => x"780d0001",
    16038 => x"78110001", 16039 => x"78100001", 16040 => x"780c0001",
    16041 => x"78160001", 16042 => x"780f0001", 16043 => x"3b396d08",
    16044 => x"283b0000", 16045 => x"396b6a78", 16046 => x"34130009",
    16047 => x"3b18411c", 16048 => x"34170001", 16049 => x"34120003",
    16050 => x"39ad6b0c", 16051 => x"3a316b2c", 16052 => x"3a106a90",
    16053 => x"398c6db0", 16054 => x"3ad66cd4", 16055 => x"39ef6da8",
    16056 => x"e000007b", 16057 => x"2861007c", 16058 => x"5b810048",
    16059 => x"2b8e0048", 16060 => x"2b940048", 16061 => x"29610004",
    16062 => x"01ce0018", 16063 => x"a29ba000", 16064 => x"3421ffff",
    16065 => x"21ce007f", 16066 => x"54330050", 16067 => x"3c210002",
    16068 => x"b7010800", 16069 => x"28210000", 16070 => x"c0200000",
    16071 => x"29610048", 16072 => x"58610040", 16073 => x"296100d0",
    16074 => x"296200cc", 16075 => x"b4410800", 16076 => x"0022001f",
    16077 => x"b4410800", 16078 => x"14210001", 16079 => x"34020001",
    16080 => x"58610044", 16081 => x"29810000", 16082 => x"fbfffb89",
    16083 => x"fbfff2d3", 16084 => x"34210032", 16085 => x"59610008",
    16086 => x"3401000a", 16087 => x"e0000011", 16088 => x"29750008",
    16089 => x"fbfff2cd", 16090 => x"caa10800", 16091 => x"4c200037",
    16092 => x"29610000", 16093 => x"5c370003", 16094 => x"59770004",
    16095 => x"e0000033", 16096 => x"59720004", 16097 => x"e0000031",
    16098 => x"29810000", 16099 => x"34020000", 16100 => x"fbfffb77",
    16101 => x"b9a00800", 16102 => x"fbfffc09", 16103 => x"34010002",
    16104 => x"59610004", 16105 => x"e0000029", 16106 => x"b9a00800",
    16107 => x"fbfffc1a", 16108 => x"e0000012", 16109 => x"ba000800",
    16110 => x"fbfffd74", 16111 => x"34010004", 16112 => x"e3fffff8",
    16113 => x"29610064", 16114 => x"44200020", 16115 => x"29610068",
    16116 => x"4420001e", 16117 => x"29610000", 16118 => x"5c320009",
    16119 => x"34010005", 16120 => x"e3fffff0", 16121 => x"ba200800",
    16122 => x"fbfffdb5", 16123 => x"34010006", 16124 => x"e3ffffec",
    16125 => x"296100ec", 16126 => x"44200014", 16127 => x"b9600800",
    16128 => x"fbffff6f", 16129 => x"34010008", 16130 => x"e3ffffe6",
    16131 => x"29610000", 16132 => x"5c370004", 16133 => x"b9a00800",
    16134 => x"fbfffbff", 16135 => x"44200007", 16136 => x"29610064",
    16137 => x"44200005", 16138 => x"29610000", 16139 => x"5c320007",
    16140 => x"296100ec", 16141 => x"5c200005", 16142 => x"29610010",
    16143 => x"34210001", 16144 => x"59610010", 16145 => x"59730004",
    16146 => x"ba000800", 16147 => x"ba801000", 16148 => x"b9c01800",
    16149 => x"fbfffcf6", 16150 => x"29610064", 16151 => x"4420001c",
    16152 => x"ba801000", 16153 => x"ba200800", 16154 => x"b9c01800",
    16155 => x"fbfffdca", 16156 => x"29620004", 16157 => x"34010008",
    16158 => x"5c410015", 16159 => x"29610000", 16160 => x"34150000",
    16161 => x"5c32000c", 16162 => x"e0000008", 16163 => x"0aa10090",
    16164 => x"ba801000", 16165 => x"b9c01800", 16166 => x"b5610800",
    16167 => x"34210144", 16168 => x"fbfffdbd", 16169 => x"36b50001",
    16170 => x"29e10000", 16171 => x"3421ffff", 16172 => x"4835fff7",
    16173 => x"29810000", 16174 => x"49c10005", 16175 => x"bac00800",
    16176 => x"ba801000", 16177 => x"b9c01800", 16178 => x"fbfffe78",
    16179 => x"2b230000", 16180 => x"78020002", 16181 => x"28610080",
    16182 => x"a0220800", 16183 => x"4420ff82", 16184 => x"78010001",
    16185 => x"38216a74", 16186 => x"28220000", 16187 => x"34420001",
    16188 => x"58220000", 16189 => x"34010001", 16190 => x"d0410000",
    16191 => x"2b9d0004", 16192 => x"2b8b0044", 16193 => x"2b8c0040",
    16194 => x"2b8d003c", 16195 => x"2b8e0038", 16196 => x"2b8f0034",
    16197 => x"2b900030", 16198 => x"2b91002c", 16199 => x"2b920028",
    16200 => x"2b930024", 16201 => x"2b940020", 16202 => x"2b95001c",
    16203 => x"2b960018", 16204 => x"2b970014", 16205 => x"2b980010",
    16206 => x"2b99000c", 16207 => x"2b9b0008", 16208 => x"379c0048",
    16209 => x"c3a00000", 16210 => x"78010001", 16211 => x"38216d10",
    16212 => x"28220000", 16213 => x"78030001", 16214 => x"78010001",
    16215 => x"38216d0c", 16216 => x"38633d60", 16217 => x"58220000",
    16218 => x"28610000", 16219 => x"58410000", 16220 => x"c3a00000",
    16221 => x"379cffd4", 16222 => x"5b8b0028", 16223 => x"5b8c0024",
    16224 => x"5b8d0020", 16225 => x"5b8e001c", 16226 => x"5b8f0018",
    16227 => x"5b900014", 16228 => x"5b910010", 16229 => x"5b92000c",
    16230 => x"5b930008", 16231 => x"5b9d0004", 16232 => x"b8205800",
    16233 => x"b8408000", 16234 => x"b8609000", 16235 => x"fbffc107",
    16236 => x"78010001", 16237 => x"38216dd4", 16238 => x"28240000",
    16239 => x"78010001", 16240 => x"38216d08", 16241 => x"58240000",
    16242 => x"78010001", 16243 => x"28860000", 16244 => x"38216d10",
    16245 => x"28220000", 16246 => x"78010001", 16247 => x"38216d0c",
    16248 => x"00c50010", 16249 => x"58220000", 16250 => x"78010001",
    16251 => x"38216db0", 16252 => x"20a5003f", 16253 => x"00c60018",
    16254 => x"58250000", 16255 => x"78010001", 16256 => x"38216da8",
    16257 => x"20c60007", 16258 => x"58260000", 16259 => x"78010001",
    16260 => x"38216a78", 16261 => x"582b0000", 16262 => x"58200010",
    16263 => x"58800040", 16264 => x"58800044", 16265 => x"58800000",
    16266 => x"58800028", 16267 => x"58800024", 16268 => x"58800004",
    16269 => x"58800020", 16270 => x"340303e8", 16271 => x"58830048",
    16272 => x"78040001", 16273 => x"38843d24", 16274 => x"28830000",
    16275 => x"5840001c", 16276 => x"58430000", 16277 => x"34020004",
    16278 => x"5d620004", 16279 => x"34020007", 16280 => x"58220004",
    16281 => x"e0000006", 16282 => x"34020009", 16283 => x"58220004",
    16284 => x"34010003", 16285 => x"5d610002", 16286 => x"ba002800",
    16287 => x"78010001", 16288 => x"b8a01000", 16289 => x"38216a90",
    16290 => x"780d0001", 16291 => x"fbfffc55", 16292 => x"39ad6db0",
    16293 => x"29a30000", 16294 => x"78010001", 16295 => x"38216b2c",
    16296 => x"ba001000", 16297 => x"780f0001", 16298 => x"780e0001",
    16299 => x"fbfffcd6", 16300 => x"340c0000", 16301 => x"39ef6da8",
    16302 => x"39ce6a78", 16303 => x"34130001", 16304 => x"e000000c",
    16305 => x"09910090", 16306 => x"29a40000", 16307 => x"ba001000",
    16308 => x"b5d10800", 16309 => x"34840001", 16310 => x"b48c1800",
    16311 => x"34210144", 16312 => x"b5d18800", 16313 => x"fbfffcc8",
    16314 => x"358c0001", 16315 => x"5a33013c", 16316 => x"29e10000",
    16317 => x"3421ffff", 16318 => x"482cfff3", 16319 => x"34010002",
    16320 => x"5d610006", 16321 => x"78010001", 16322 => x"38216d0c",
    16323 => x"28210000", 16324 => x"34020006", 16325 => x"5822001c",
    16326 => x"780e0001", 16327 => x"780d0001", 16328 => x"340c0000",
    16329 => x"39ce6db0", 16330 => x"39ad6a78", 16331 => x"e0000008",
    16332 => x"3d810005", 16333 => x"b9801000", 16334 => x"b5a10800",
    16335 => x"3421025c", 16336 => x"34030200", 16337 => x"fbfffdc0",
    16338 => x"358c0001", 16339 => x"29c20000", 16340 => x"484cfff8",
    16341 => x"34010001", 16342 => x"5d61001d", 16343 => x"78010001",
    16344 => x"38216d08", 16345 => x"28210000", 16346 => x"28210004",
    16347 => x"20210002", 16348 => x"44200012", 16349 => x"78010001",
    16350 => x"78040001", 16351 => x"38216a78", 16352 => x"38846a90",
    16353 => x"58240094", 16354 => x"78040001", 16355 => x"38846b2c",
    16356 => x"58240098", 16357 => x"78010001", 16358 => x"38216da8",
    16359 => x"28240000", 16360 => x"78010001", 16361 => x"38216b0c",
    16362 => x"b4441000", 16363 => x"ba401800", 16364 => x"fbfffae7",
    16365 => x"e0000006", 16366 => x"78020001", 16367 => x"34010000",
    16368 => x"38423984", 16369 => x"fbffc094", 16370 => x"e0000020",
    16371 => x"78010001", 16372 => x"3d6b0002", 16373 => x"3821419c",
    16374 => x"78040001", 16375 => x"78050001", 16376 => x"b42b5800",
    16377 => x"38846db0", 16378 => x"38a56da8", 16379 => x"29630000",
    16380 => x"28840000", 16381 => x"28a50000", 16382 => x"78020001",
    16383 => x"34010000", 16384 => x"384239c0", 16385 => x"fbffc084",
    16386 => x"78010001", 16387 => x"38216d08", 16388 => x"28210000",
    16389 => x"78020002", 16390 => x"e0000003", 16391 => x"2823007c",
    16392 => x"5b83002c", 16393 => x"28230080", 16394 => x"a0621800",
    16395 => x"4460fffc", 16396 => x"34020001", 16397 => x"58220064",
    16398 => x"28220028", 16399 => x"38420001", 16400 => x"58220028",
    16401 => x"fbffc06a", 16402 => x"2b9d0004", 16403 => x"2b8b0028",
    16404 => x"2b8c0024", 16405 => x"2b8d0020", 16406 => x"2b8e001c",
    16407 => x"2b8f0018", 16408 => x"2b900014", 16409 => x"2b910010",
    16410 => x"2b92000c", 16411 => x"2b930008", 16412 => x"379c002c",
    16413 => x"c3a00000", 16414 => x"379cfffc", 16415 => x"5b9d0004",
    16416 => x"78020001", 16417 => x"38426a78", 16418 => x"b8201800",
    16419 => x"28410004", 16420 => x"64640000", 16421 => x"7c210008",
    16422 => x"b8810800", 16423 => x"44200006", 16424 => x"78020001",
    16425 => x"34010000", 16426 => x"384239f4", 16427 => x"fbffc05a",
    16428 => x"e0000006", 16429 => x"3463ffff", 16430 => x"08630090",
    16431 => x"b4431000", 16432 => x"34410144", 16433 => x"fbfffc7e",
    16434 => x"2b9d0004", 16435 => x"379c0004", 16436 => x"c3a00000",
    16437 => x"379cfffc", 16438 => x"5b9d0004", 16439 => x"44200008",
    16440 => x"3421ffff", 16441 => x"08210090", 16442 => x"78020001",
    16443 => x"38426a78", 16444 => x"b4220800", 16445 => x"34210144",
    16446 => x"fbfffc9b", 16447 => x"2b9d0004", 16448 => x"379c0004",
    16449 => x"c3a00000", 16450 => x"78020001", 16451 => x"b8201800",
    16452 => x"38426a78", 16453 => x"5c200004", 16454 => x"28410004",
    16455 => x"64210008", 16456 => x"c3a00000", 16457 => x"28450004",
    16458 => x"34040008", 16459 => x"34010000", 16460 => x"5ca40006",
    16461 => x"3463ffff", 16462 => x"08630090", 16463 => x"b4431000",
    16464 => x"2841017c", 16465 => x"7c210000", 16466 => x"c3a00000",
    16467 => x"379cffe8", 16468 => x"5b8b0018", 16469 => x"5b8c0014",
    16470 => x"5b8d0010", 16471 => x"5b8e000c", 16472 => x"5b8f0008",
    16473 => x"5b9d0004", 16474 => x"3403ffff", 16475 => x"b8407800",
    16476 => x"5c230016", 16477 => x"34010000", 16478 => x"780c0001",
    16479 => x"780d0001", 16480 => x"fbfffff3", 16481 => x"340b0000",
    16482 => x"398c6da8", 16483 => x"39ad6a78", 16484 => x"340e0004",
    16485 => x"e0000009", 16486 => x"09610090", 16487 => x"b5a10800",
    16488 => x"2821013c", 16489 => x"5c2e0004", 16490 => x"35610001",
    16491 => x"b9e01000", 16492 => x"fbfffdec", 16493 => x"356b0001",
    16494 => x"29810000", 16495 => x"3421ffff", 16496 => x"482bfff6",
    16497 => x"e0000002", 16498 => x"fbfffde6", 16499 => x"2b9d0004",
    16500 => x"2b8b0018", 16501 => x"2b8c0014", 16502 => x"2b8d0010",
    16503 => x"2b8e000c", 16504 => x"2b8f0008", 16505 => x"379c0018",
    16506 => x"c3a00000", 16507 => x"379cfff0", 16508 => x"5b8b0010",
    16509 => x"5b8c000c", 16510 => x"5b8d0008", 16511 => x"5b9d0004",
    16512 => x"780b0001", 16513 => x"b8406800", 16514 => x"b8606000",
    16515 => x"396b6b2c", 16516 => x"44200007", 16517 => x"3421ffff",
    16518 => x"082b0090", 16519 => x"78010001", 16520 => x"38216a78",
    16521 => x"b5610800", 16522 => x"342b0144", 16523 => x"45a0000b",
    16524 => x"2962006c", 16525 => x"34041f40", 16526 => x"34030000",
    16527 => x"3c420001", 16528 => x"1441001f", 16529 => x"f80002e6",
    16530 => x"3c210012", 16531 => x"0044000e", 16532 => x"b8242000",
    16533 => x"59a40000", 16534 => x"4580000b", 16535 => x"29620068",
    16536 => x"34030000", 16537 => x"34041f40", 16538 => x"3c420001",
    16539 => x"1441001f", 16540 => x"f80002db", 16541 => x"3c210012",
    16542 => x"0042000e", 16543 => x"b8221000", 16544 => x"59820000",
    16545 => x"2b9d0004", 16546 => x"2b8b0010", 16547 => x"2b8c000c",
    16548 => x"2b8d0008", 16549 => x"379c0010", 16550 => x"c3a00000",
    16551 => x"379cfff0", 16552 => x"5b8b0010", 16553 => x"5b8c000c",
    16554 => x"5b8d0008", 16555 => x"5b9d0004", 16556 => x"b8205800",
    16557 => x"b8406800", 16558 => x"78010001", 16559 => x"3d620005",
    16560 => x"38216a78", 16561 => x"b4220800", 16562 => x"28240274",
    16563 => x"b8606000", 16564 => x"4c800003", 16565 => x"34844000",
    16566 => x"e0000004", 16567 => x"34013fff", 16568 => x"4c240002",
    16569 => x"3484c000", 16570 => x"3c840001", 16571 => x"34010000",
    16572 => x"20823ffe", 16573 => x"34030000", 16574 => x"34041f40",
    16575 => x"f80002b8", 16576 => x"3c210012", 16577 => x"0044000e",
    16578 => x"b8242000", 16579 => x"59a40000", 16580 => x"4580000c",
    16581 => x"78010001", 16582 => x"38216cf4", 16583 => x"28220000",
    16584 => x"3d630005", 16585 => x"78010001", 16586 => x"38216a78",
    16587 => x"b4230800", 16588 => x"28210260", 16589 => x"94410800",
    16590 => x"20210001", 16591 => x"59810000", 16592 => x"3d6b0005",
    16593 => x"78020001", 16594 => x"38426a78", 16595 => x"b44b1000",
    16596 => x"28410278", 16597 => x"2b9d0004", 16598 => x"2b8b0010",
    16599 => x"2b8c000c", 16600 => x"2b8d0008", 16601 => x"379c0010",
    16602 => x"c3a00000", 16603 => x"379cffec", 16604 => x"5b8b0014",
    16605 => x"5b8c0010", 16606 => x"5b9d000c", 16607 => x"780b0001",
    16608 => x"396b6a78", 16609 => x"29610000", 16610 => x"4c010016",
    16611 => x"78010001", 16612 => x"38216a74", 16613 => x"282c0000",
    16614 => x"29620004", 16615 => x"78010001", 16616 => x"38214144",
    16617 => x"fbfff9cb", 16618 => x"29640000", 16619 => x"b8201800",
    16620 => x"296500a0", 16621 => x"29660064", 16622 => x"296700ec",
    16623 => x"29680050", 16624 => x"296200d8", 16625 => x"29610010",
    16626 => x"5b820004", 16627 => x"5b810008", 16628 => x"78010001",
    16629 => x"38213a24", 16630 => x"b9801000", 16631 => x"fbffea7d",
    16632 => x"2b9d000c", 16633 => x"2b8b0014", 16634 => x"2b8c0010",
    16635 => x"379c0014", 16636 => x"c3a00000", 16637 => x"379cfffc",
    16638 => x"5b9d0004", 16639 => x"5c200004", 16640 => x"78010001",
    16641 => x"38216b2c", 16642 => x"e0000007", 16643 => x"3421ffff",
    16644 => x"08210090", 16645 => x"78020001", 16646 => x"38426a78",
    16647 => x"b4220800", 16648 => x"34210144", 16649 => x"fbfffc84",
    16650 => x"2b9d0004", 16651 => x"379c0004", 16652 => x"c3a00000",
    16653 => x"379cfff0", 16654 => x"5b8b0010", 16655 => x"5b8c000c",
    16656 => x"5b8d0008", 16657 => x"5b9d0004", 16658 => x"780d0001",
    16659 => x"780c0001", 16660 => x"b8205800", 16661 => x"39ad6a78",
    16662 => x"398c6cf4", 16663 => x"44400010", 16664 => x"34020001",
    16665 => x"fbfff942", 16666 => x"3d610005", 16667 => x"b5a16800",
    16668 => x"35a1025c", 16669 => x"fbfffc7b", 16670 => x"29820000",
    16671 => x"34010001", 16672 => x"bc2b0800", 16673 => x"b8220800",
    16674 => x"78020001", 16675 => x"59810000", 16676 => x"38423a78",
    16677 => x"34010000", 16678 => x"e000000d", 16679 => x"34030001",
    16680 => x"29840000", 16681 => x"bc611800", 16682 => x"a4601800",
    16683 => x"a0641800", 16684 => x"59830000", 16685 => x"29a30124",
    16686 => x"44230002", 16687 => x"fbfff92c", 16688 => x"78020001",
    16689 => x"34010000", 16690 => x"38423a98", 16691 => x"b9601800",
    16692 => x"fbffbf51", 16693 => x"2b9d0004", 16694 => x"2b8b0010",
    16695 => x"2b8c000c", 16696 => x"2b8d0008", 16697 => x"379c0010",
    16698 => x"c3a00000", 16699 => x"08210090", 16700 => x"78020001",
    16701 => x"38426a78", 16702 => x"b4411000", 16703 => x"2841013c",
    16704 => x"2843013c", 16705 => x"34020004", 16706 => x"7c210001",
    16707 => x"5c620002", 16708 => x"38210002", 16709 => x"c3a00000",
    16710 => x"4c200005", 16711 => x"78010001", 16712 => x"38216a78",
    16713 => x"28210050", 16714 => x"c3a00000", 16715 => x"78020001",
    16716 => x"38426a78", 16717 => x"5c200003", 16718 => x"284100d8",
    16719 => x"c3a00000", 16720 => x"3421ffff", 16721 => x"08210090",
    16722 => x"b4411000", 16723 => x"28410168", 16724 => x"c3a00000",
    16725 => x"78030001", 16726 => x"38636d08", 16727 => x"4c200007",
    16728 => x"78010001", 16729 => x"38216a78", 16730 => x"58220050",
    16731 => x"28610000", 16732 => x"58220040", 16733 => x"c3a00000",
    16734 => x"2024000f", 16735 => x"28630000", 16736 => x"3c840010",
    16737 => x"2045ffff", 16738 => x"b8a42000", 16739 => x"58640044",
    16740 => x"78030001", 16741 => x"38636a78", 16742 => x"5c200003",
    16743 => x"586200d8", 16744 => x"c3a00000", 16745 => x"3421ffff",
    16746 => x"08210090", 16747 => x"b4611800", 16748 => x"58620168",
    16749 => x"c3a00000", 16750 => x"379cffc0", 16751 => x"5b8b0040",
    16752 => x"5b8c003c", 16753 => x"5b8d0038", 16754 => x"5b8e0034",
    16755 => x"5b8f0030", 16756 => x"5b90002c", 16757 => x"5b910028",
    16758 => x"5b920024", 16759 => x"5b930020", 16760 => x"5b94001c",
    16761 => x"5b950018", 16762 => x"5b960014", 16763 => x"5b970010",
    16764 => x"5b98000c", 16765 => x"5b990008", 16766 => x"5b9d0004",
    16767 => x"78010001", 16768 => x"38216a78", 16769 => x"28220000",
    16770 => x"34010001", 16771 => x"5c410004", 16772 => x"78010001",
    16773 => x"38216b0c", 16774 => x"fbfff99a", 16775 => x"78100001",
    16776 => x"780c0001", 16777 => x"780d0001", 16778 => x"78160001",
    16779 => x"78140001", 16780 => x"78130001", 16781 => x"78120001",
    16782 => x"78110001", 16783 => x"340b0001", 16784 => x"3a106da8",
    16785 => x"398c6a78", 16786 => x"340e0001", 16787 => x"39ad6d08",
    16788 => x"3ad63acc", 16789 => x"34150002", 16790 => x"3a943b14",
    16791 => x"34190003", 16792 => x"3a733b44", 16793 => x"34180004",
    16794 => x"3a523b68", 16795 => x"3a313af0", 16796 => x"e0000058",
    16797 => x"3577ffff", 16798 => x"0aef0090", 16799 => x"b58f7800",
    16800 => x"29e1013c", 16801 => x"442e0011", 16802 => x"29a10000",
    16803 => x"bdcb1000", 16804 => x"28210020", 16805 => x"00210008",
    16806 => x"202100ff", 16807 => x"a0220800", 16808 => x"5c20000a",
    16809 => x"bac01000", 16810 => x"b9601800", 16811 => x"fbffbeda",
    16812 => x"b9600800", 16813 => x"fbfffe88", 16814 => x"b9600800",
    16815 => x"34020000", 16816 => x"fbfffc3f", 16817 => x"59ee013c",
    16818 => x"0ae10090", 16819 => x"b5817800", 16820 => x"29e3013c",
    16821 => x"44750018", 16822 => x"48750003", 16823 => x"5c6e003c",
    16824 => x"e0000004", 16825 => x"44790020", 16826 => x"5c780039",
    16827 => x"e000002a", 16828 => x"298100ec", 16829 => x"44200036",
    16830 => x"29a10000", 16831 => x"bdcb1000", 16832 => x"28210020",
    16833 => x"00210008", 16834 => x"202100ff", 16835 => x"a0220800",
    16836 => x"4420002f", 16837 => x"34010000", 16838 => x"ba201000",
    16839 => x"b9601800", 16840 => x"fbffbebd", 16841 => x"b9600800",
    16842 => x"fbfffe54", 16843 => x"59f5013c", 16844 => x"e0000027",
    16845 => x"29e1017c", 16846 => x"44200025", 16847 => x"29840014",
    16848 => x"34010000", 16849 => x"ba801000", 16850 => x"b9601800",
    16851 => x"fbffbeb2", 16852 => x"29820014", 16853 => x"b9600800",
    16854 => x"fbfffc82", 16855 => x"59f9013c", 16856 => x"e000001b",
    16857 => x"b5810800", 16858 => x"34210144", 16859 => x"fbfffbb2",
    16860 => x"5c200017", 16861 => x"ba601000", 16862 => x"b9601800",
    16863 => x"fbffbea6", 16864 => x"b9600800", 16865 => x"34020001",
    16866 => x"fbfffc0d", 16867 => x"59f8013c", 16868 => x"e000000f",
    16869 => x"298100ec", 16870 => x"44200003", 16871 => x"29e1017c",
    16872 => x"5c20000b", 16873 => x"0af70090", 16874 => x"34010000",
    16875 => x"ba401000", 16876 => x"b9601800", 16877 => x"fbffbe98",
    16878 => x"b9600800", 16879 => x"34020000", 16880 => x"b597b800",
    16881 => x"fbfffbfe", 16882 => x"5aee013c", 16883 => x"356b0001",
    16884 => x"2a010000", 16885 => x"482bffa8", 16886 => x"2b9d0004",
    16887 => x"2b8b0040", 16888 => x"2b8c003c", 16889 => x"2b8d0038",
    16890 => x"2b8e0034", 16891 => x"2b8f0030", 16892 => x"2b90002c",
    16893 => x"2b910028", 16894 => x"2b920024", 16895 => x"2b930020",
    16896 => x"2b94001c", 16897 => x"2b950018", 16898 => x"2b960014",
    16899 => x"2b970010", 16900 => x"2b98000c", 16901 => x"2b990008",
    16902 => x"379c0040", 16903 => x"c3a00000", 16904 => x"379cfff0",
    16905 => x"5b8b0010", 16906 => x"5b8c000c", 16907 => x"5b8d0008",
    16908 => x"5b9d0004", 16909 => x"fbffbe65", 16910 => x"78020001",
    16911 => x"34010000", 16912 => x"38423b94", 16913 => x"fbffbe74",
    16914 => x"34020000", 16915 => x"3401ffff", 16916 => x"fbffff41",
    16917 => x"34010001", 16918 => x"fbfffc1f", 16919 => x"380bffff",
    16920 => x"b8206800", 16921 => x"b9601000", 16922 => x"3401ffff",
    16923 => x"fbffff3a", 16924 => x"34010001", 16925 => x"fbfffc18",
    16926 => x"78040001", 16927 => x"38843d64", 16928 => x"28830000",
    16929 => x"b8206000", 16930 => x"b9801000", 16931 => x"b9a00800",
    16932 => x"fbfffbe0", 16933 => x"78020001", 16934 => x"b8202800",
    16935 => x"b9a01800", 16936 => x"b9802000", 16937 => x"34010000",
    16938 => x"38423bb8", 16939 => x"fbffbe5a", 16940 => x"34020000",
    16941 => x"34010000", 16942 => x"fbffff27", 16943 => x"34010000",
    16944 => x"fbfffc05", 16945 => x"b8206000", 16946 => x"b9601000",
    16947 => x"34010000", 16948 => x"fbffff21", 16949 => x"34010000",
    16950 => x"fbfffbff", 16951 => x"78040001", 16952 => x"38843d68",
    16953 => x"28830000", 16954 => x"b8205800", 16955 => x"b9601000",
    16956 => x"b9800800", 16957 => x"fbfffbc7", 16958 => x"78020001",
    16959 => x"b8202800", 16960 => x"b9801800", 16961 => x"b9602000",
    16962 => x"38423be8", 16963 => x"34010000", 16964 => x"fbffbe41",
    16965 => x"34010002", 16966 => x"fbfffbef", 16967 => x"78020001",
    16968 => x"b8201800", 16969 => x"38423c18", 16970 => x"34010000",
    16971 => x"fbffbe3a", 16972 => x"2b9d0004", 16973 => x"2b8b0010",
    16974 => x"2b8c000c", 16975 => x"2b8d0008", 16976 => x"379c0010",
    16977 => x"c3a00000", 16978 => x"379cfff0", 16979 => x"5b8b0010",
    16980 => x"5b8c000c", 16981 => x"5b8d0008", 16982 => x"5b9d0004",
    16983 => x"78010001", 16984 => x"780b0001", 16985 => x"38213cc0",
    16986 => x"780c0001", 16987 => x"396bf800", 16988 => x"282d0000",
    16989 => x"398c3cac", 16990 => x"e0000005", 16991 => x"b9800800",
    16992 => x"fbffe914", 16993 => x"340103e8", 16994 => x"fbffef49",
    16995 => x"29610000", 16996 => x"5c2dfffb", 16997 => x"2b9d0004",
    16998 => x"2b8b0010", 16999 => x"2b8c000c", 17000 => x"2b8d0008",
    17001 => x"379c0010", 17002 => x"c3a00000", 17003 => x"c3a00000",
    17004 => x"379cfff8", 17005 => x"5b8b0008", 17006 => x"5b9d0004",
    17007 => x"28240014", 17008 => x"b8201800", 17009 => x"b8403000",
    17010 => x"44800015", 17011 => x"28250010", 17012 => x"20a50002",
    17013 => x"5ca00007", 17014 => x"b4862000", 17015 => x"b8800800",
    17016 => x"2b9d0004", 17017 => x"2b8b0008", 17018 => x"379c0008",
    17019 => x"c3a00000", 17020 => x"346b0030", 17021 => x"b4861000",
    17022 => x"b9600800", 17023 => x"34030040", 17024 => x"f80001cc",
    17025 => x"b9602000", 17026 => x"b8800800", 17027 => x"2b9d0004",
    17028 => x"2b8b0008", 17029 => x"379c0008", 17030 => x"c3a00000",
    17031 => x"28250010", 17032 => x"20a70004", 17033 => x"5ce4ffeb",
    17034 => x"2825001c", 17035 => x"34040000", 17036 => x"44a7ffeb",
    17037 => x"342b0030", 17038 => x"34040040", 17039 => x"b9601800",
    17040 => x"d8a00000", 17041 => x"b9602000", 17042 => x"e3fffff0",
    17043 => x"379cfff4", 17044 => x"5b8b0008", 17045 => x"5b9d0004",
    17046 => x"28220014", 17047 => x"b8205800", 17048 => x"44400013",
    17049 => x"2961000c", 17050 => x"b4411000", 17051 => x"28430000",
    17052 => x"78040001", 17053 => x"38843d6c", 17054 => x"28820000",
    17055 => x"3401ffec", 17056 => x"5c620007", 17057 => x"78020001",
    17058 => x"38426cf8", 17059 => x"28430000", 17060 => x"34010000",
    17061 => x"584b0000", 17062 => x"5963007c", 17063 => x"2b9d0004",
    17064 => x"2b8b0008", 17065 => x"379c000c", 17066 => x"c3a00000",
    17067 => x"28230010", 17068 => x"20630004", 17069 => x"5c62ffec",
    17070 => x"2825001c", 17071 => x"2822000c", 17072 => x"3783000c",
    17073 => x"34040004", 17074 => x"d8a00000", 17075 => x"2b83000c",
    17076 => x"e3ffffe8", 17077 => x"379cfff0", 17078 => x"5b8b0010",
    17079 => x"5b8c000c", 17080 => x"5b8d0008", 17081 => x"5b9d0004",
    17082 => x"b8205800", 17083 => x"44400047", 17084 => x"2822000c",
    17085 => x"58200080", 17086 => x"582000b0", 17087 => x"58220090",
    17088 => x"340c0000", 17089 => x"b9600800", 17090 => x"fbffffaa",
    17091 => x"59610028", 17092 => x"4022003f", 17093 => x"5c400006",
    17094 => x"78040001", 17095 => x"38843d6c", 17096 => x"28230000",
    17097 => x"28820000", 17098 => x"4462005d", 17099 => x"34010000",
    17100 => x"45800030", 17101 => x"3583ffff", 17102 => x"346c0028",
    17103 => x"b58c0800", 17104 => x"b4210800", 17105 => x"b5610800",
    17106 => x"28220000", 17107 => x"5c40000f", 17108 => x"34010000",
    17109 => x"44620027", 17110 => x"34620027", 17111 => x"b4421000",
    17112 => x"b4421000", 17113 => x"b5621000", 17114 => x"e0000002",
    17115 => x"44610044", 17116 => x"28410000", 17117 => x"3463ffff",
    17118 => x"3442fffc", 17119 => x"4420fffc", 17120 => x"596300b0",
    17121 => x"346c0028", 17122 => x"346d0024", 17123 => x"b5ad6800",
    17124 => x"b5ad6800", 17125 => x"b56d6800", 17126 => x"29a20000",
    17127 => x"b9600800", 17128 => x"b58c6000", 17129 => x"fbffff83",
    17130 => x"b58c6000", 17131 => x"b56c1000", 17132 => x"29a40000",
    17133 => x"28430000", 17134 => x"296c00b0", 17135 => x"34840040",
    17136 => x"3463ffff", 17137 => x"59610028", 17138 => x"59a40000",
    17139 => x"58430000", 17140 => x"35830020", 17141 => x"b4631800",
    17142 => x"b4631800", 17143 => x"b5631800", 17144 => x"2824000c",
    17145 => x"28620000", 17146 => x"b4441000", 17147 => x"59620074",
    17148 => x"2b9d0004", 17149 => x"2b8b0010", 17150 => x"2b8c000c",
    17151 => x"2b8d0008", 17152 => x"379c0010", 17153 => x"c3a00000",
    17154 => x"28210028", 17155 => x"296300b0", 17156 => x"34050002",
    17157 => x"4024003f", 17158 => x"eca32800", 17159 => x"64840002",
    17160 => x"a0852000", 17161 => x"4482ffc5", 17162 => x"34620020",
    17163 => x"b4421000", 17164 => x"b4421000", 17165 => x"b5621000",
    17166 => x"28450000", 17167 => x"34640025", 17168 => x"28220004",
    17169 => x"b4842000", 17170 => x"b4842000", 17171 => x"b4a21000",
    17172 => x"b5642000", 17173 => x"58820000", 17174 => x"2824000c",
    17175 => x"34610021", 17176 => x"b4210800", 17177 => x"b4210800",
    17178 => x"b5610800", 17179 => x"b4852800", 17180 => x"346c0001",
    17181 => x"58250000", 17182 => x"e3ffffa3", 17183 => x"34010000",
    17184 => x"596000b0", 17185 => x"2b9d0004", 17186 => x"2b8b0010",
    17187 => x"2b8c000c", 17188 => x"2b8d0008", 17189 => x"379c0010",
    17190 => x"c3a00000", 17191 => x"35820024", 17192 => x"b4421000",
    17193 => x"b4421000", 17194 => x"b5621800", 17195 => x"2c250004",
    17196 => x"28640000", 17197 => x"35820028", 17198 => x"b4421000",
    17199 => x"b4421000", 17200 => x"b5621000", 17201 => x"34a5ffff",
    17202 => x"34840040", 17203 => x"58450000", 17204 => x"58640000",
    17205 => x"596c00b0", 17206 => x"e3ffffbe", 17207 => x"379cffec",
    17208 => x"5b8b0014", 17209 => x"5b8c0010", 17210 => x"5b8d000c",
    17211 => x"5b8e0008", 17212 => x"5b9d0004", 17213 => x"b8406000",
    17214 => x"34020001", 17215 => x"b8205800", 17216 => x"b8607000",
    17217 => x"b8806800", 17218 => x"fbffff73", 17219 => x"b9600800",
    17220 => x"34020000", 17221 => x"fbffff70", 17222 => x"b8202800",
    17223 => x"4420001e", 17224 => x"28a10018", 17225 => x"5c2cfffa",
    17226 => x"28a1001c", 17227 => x"5c2efff8", 17228 => x"28a10020",
    17229 => x"5c2dfff6", 17230 => x"296100b0", 17231 => x"59650028",
    17232 => x"28a2000c", 17233 => x"34210020", 17234 => x"b4210800",
    17235 => x"b4210800", 17236 => x"b5610800", 17237 => x"28230000",
    17238 => x"34010000", 17239 => x"b4431800", 17240 => x"59630074",
    17241 => x"28a30014", 17242 => x"59600078", 17243 => x"34630001",
    17244 => x"c8621000", 17245 => x"59620070", 17246 => x"2b9d0004",
    17247 => x"2b8b0014", 17248 => x"2b8c0010", 17249 => x"2b8d000c",
    17250 => x"2b8e0008", 17251 => x"379c0014", 17252 => x"c3a00000",
    17253 => x"3401fffe", 17254 => x"e3fffff8", 17255 => x"379cfff8",
    17256 => x"5b8b0008", 17257 => x"5b9d0004", 17258 => x"b8205800",
    17259 => x"fbffffcc", 17260 => x"4c200005", 17261 => x"2b9d0004",
    17262 => x"2b8b0008", 17263 => x"379c0008", 17264 => x"c3a00000",
    17265 => x"29610074", 17266 => x"59600028", 17267 => x"2b9d0004",
    17268 => x"2b8b0008", 17269 => x"379c0008", 17270 => x"c3a00000",
    17271 => x"2045ffff", 17272 => x"00460010", 17273 => x"2088ffff",
    17274 => x"00890010", 17275 => x"89053800", 17276 => x"89064000",
    17277 => x"89252800", 17278 => x"00ea0010", 17279 => x"89263000",
    17280 => x"b5052800", 17281 => x"b4aa2800", 17282 => x"50a80003",
    17283 => x"78080001", 17284 => x"b4c83000", 17285 => x"88431000",
    17286 => x"88812000", 17287 => x"00a10010", 17288 => x"3ca50010",
    17289 => x"b4c13000", 17290 => x"20e7ffff", 17291 => x"b4440800",
    17292 => x"b4260800", 17293 => x"b4a71000", 17294 => x"c3a00000",
    17295 => x"44600008", 17296 => x"34040020", 17297 => x"c8832000",
    17298 => x"48800006", 17299 => x"c8041000", 17300 => x"34030000",
    17301 => x"80221000", 17302 => x"b8600800", 17303 => x"c3a00000",
    17304 => x"bc242000", 17305 => x"80431000", 17306 => x"80231800",
    17307 => x"b8821000", 17308 => x"b8600800", 17309 => x"e3fffffa",
    17310 => x"379cfff8", 17311 => x"5b8b0008", 17312 => x"5b9d0004",
    17313 => x"44400022", 17314 => x"b8412000", 17315 => x"3403000f",
    17316 => x"5483000b", 17317 => x"78030001", 17318 => x"386341b0",
    17319 => x"3c210004", 17320 => x"b4621000", 17321 => x"b4410800",
    17322 => x"40210000", 17323 => x"2b9d0004", 17324 => x"2b8b0008",
    17325 => x"379c0008", 17326 => x"c3a00000", 17327 => x"340b0000",
    17328 => x"4c200003", 17329 => x"c8010800", 17330 => x"340b0001",
    17331 => x"4c400003", 17332 => x"c8021000", 17333 => x"196b0001",
    17334 => x"90c01800", 17335 => x"20630002", 17336 => x"44600008",
    17337 => x"8c220800", 17338 => x"45600002", 17339 => x"c8010800",
    17340 => x"2b9d0004", 17341 => x"2b8b0008", 17342 => x"379c0008",
    17343 => x"c3a00000", 17344 => x"34030000", 17345 => x"f800004a",
    17346 => x"e3fffff8", 17347 => x"90000800", 17348 => x"20210001",
    17349 => x"3c210001", 17350 => x"d0010000", 17351 => x"90e00800",
    17352 => x"bba0f000", 17353 => x"342100a0", 17354 => x"c0200000",
    17355 => x"379cfff8", 17356 => x"5b8b0008", 17357 => x"5b9d0004",
    17358 => x"44400015", 17359 => x"340b0000", 17360 => x"4c200003",
    17361 => x"c8010800", 17362 => x"340b0001", 17363 => x"1443001f",
    17364 => x"90c02000", 17365 => x"98621000", 17366 => x"20840002",
    17367 => x"c8431000", 17368 => x"44800008", 17369 => x"c4220800",
    17370 => x"45600002", 17371 => x"c8010800", 17372 => x"2b9d0004",
    17373 => x"2b8b0008", 17374 => x"379c0008", 17375 => x"c3a00000",
    17376 => x"34030001", 17377 => x"f800002a", 17378 => x"e3fffff8",
    17379 => x"90000800", 17380 => x"20210001", 17381 => x"3c210001",
    17382 => x"d0010000", 17383 => x"90e00800", 17384 => x"bba0f000",
    17385 => x"342100a0", 17386 => x"c0200000", 17387 => x"379cfffc",
    17388 => x"5b9d0004", 17389 => x"44400006", 17390 => x"34030000",
    17391 => x"f800001c", 17392 => x"2b9d0004", 17393 => x"379c0004",
    17394 => x"c3a00000", 17395 => x"90000800", 17396 => x"20210001",
    17397 => x"3c210001", 17398 => x"d0010000", 17399 => x"90e00800",
    17400 => x"bba0f000", 17401 => x"342100a0", 17402 => x"c0200000",
    17403 => x"379cfffc", 17404 => x"5b9d0004", 17405 => x"44400006",
    17406 => x"34030001", 17407 => x"f800000c", 17408 => x"2b9d0004",
    17409 => x"379c0004", 17410 => x"c3a00000", 17411 => x"90000800",
    17412 => x"20210001", 17413 => x"3c210001", 17414 => x"d0010000",
    17415 => x"90e00800", 17416 => x"bba0f000", 17417 => x"342100a0",
    17418 => x"c0200000", 17419 => x"f4222000", 17420 => x"44800018",
    17421 => x"34040001", 17422 => x"4c40000b", 17423 => x"34050000",
    17424 => x"54410003", 17425 => x"c8220800", 17426 => x"b8a42800",
    17427 => x"00840001", 17428 => x"00420001", 17429 => x"5c80fffb",
    17430 => x"5c600002", 17431 => x"b8a00800", 17432 => x"c3a00000",
    17433 => x"3c420001", 17434 => x"3c840001", 17435 => x"f4222800",
    17436 => x"7c860000", 17437 => x"a0c52800", 17438 => x"44a00002",
    17439 => x"4c40fffa", 17440 => x"34050000", 17441 => x"4480fff5",
    17442 => x"34050000", 17443 => x"e3ffffed", 17444 => x"34040001",
    17445 => x"34050000", 17446 => x"e3ffffea", 17447 => x"1422001f",
    17448 => x"98410800", 17449 => x"c8220800", 17450 => x"c3a00000",
    17451 => x"34060003", 17452 => x"b8202000", 17453 => x"b8402800",
    17454 => x"50c3000c", 17455 => x"b8413000", 17456 => x"20c60003",
    17457 => x"5cc0000b", 17458 => x"34010003", 17459 => x"28860000",
    17460 => x"28a20000", 17461 => x"5cc20005", 17462 => x"3463fffc",
    17463 => x"34840004", 17464 => x"34a50004", 17465 => x"5461fffa",
    17466 => x"34010000", 17467 => x"4460000e", 17468 => x"40860000",
    17469 => x"40a10000", 17470 => x"3462ffff", 17471 => x"44c10006",
    17472 => x"e000000a", 17473 => x"40860000", 17474 => x"40a10000",
    17475 => x"3442ffff", 17476 => x"5cc10006", 17477 => x"34840001",
    17478 => x"34a50001", 17479 => x"5c40fffa", 17480 => x"34010000",
    17481 => x"c3a00000", 17482 => x"c8c10800", 17483 => x"c3a00000",
    17484 => x"3404000f", 17485 => x"b8203800", 17486 => x"b8403000",
    17487 => x"5083002d", 17488 => x"b8412000", 17489 => x"20840003",
    17490 => x"5c80002b", 17491 => x"b8402000", 17492 => x"b8202800",
    17493 => x"b8603000", 17494 => x"3407000f", 17495 => x"28880000",
    17496 => x"34c6fff0", 17497 => x"58a80000", 17498 => x"28880004",
    17499 => x"58a80004", 17500 => x"28880008", 17501 => x"58a80008",
    17502 => x"2888000c", 17503 => x"34840010", 17504 => x"58a8000c",
    17505 => x"34a50010", 17506 => x"54c7fff5", 17507 => x"3463fff0",
    17508 => x"00660004", 17509 => x"2063000f", 17510 => x"34c60001",
    17511 => x"3cc60004", 17512 => x"b4263800", 17513 => x"b4463000",
    17514 => x"34020003", 17515 => x"50430011", 17516 => x"34020000",
    17517 => x"34080003", 17518 => x"b4c22000", 17519 => x"28850000",
    17520 => x"b4e22000", 17521 => x"34420004", 17522 => x"58850000",
    17523 => x"c8622000", 17524 => x"5488fffa", 17525 => x"3463fffc",
    17526 => x"00620002", 17527 => x"20630003", 17528 => x"34420001",
    17529 => x"3c420002", 17530 => x"b4e23800", 17531 => x"b4c23000",
    17532 => x"44600008", 17533 => x"34020000", 17534 => x"b4c22000",
    17535 => x"40850000", 17536 => x"b4e22000", 17537 => x"34420001",
    17538 => x"30850000", 17539 => x"5c43fffb", 17540 => x"c3a00000",
    17541 => x"b8203800", 17542 => x"b8403000", 17543 => x"5041000c",
    17544 => x"b4432000", 17545 => x"5024000a", 17546 => x"4460003f",
    17547 => x"b4231000", 17548 => x"3484ffff", 17549 => x"40850000",
    17550 => x"3442ffff", 17551 => x"3463ffff", 17552 => x"30450000",
    17553 => x"5c60fffb", 17554 => x"c3a00000", 17555 => x"3404000f",
    17556 => x"5083002d", 17557 => x"b8412000", 17558 => x"20840003",
    17559 => x"5c80002b", 17560 => x"b8402000", 17561 => x"b8202800",
    17562 => x"b8603000", 17563 => x"3407000f", 17564 => x"28880000",
    17565 => x"34c6fff0", 17566 => x"58a80000", 17567 => x"28880004",
    17568 => x"58a80004", 17569 => x"28880008", 17570 => x"58a80008",
    17571 => x"2888000c", 17572 => x"34840010", 17573 => x"58a8000c",
    17574 => x"34a50010", 17575 => x"54c7fff5", 17576 => x"3463fff0",
    17577 => x"00660004", 17578 => x"2063000f", 17579 => x"34c60001",
    17580 => x"3cc60004", 17581 => x"b4263800", 17582 => x"b4463000",
    17583 => x"34020003", 17584 => x"50430011", 17585 => x"34020000",
    17586 => x"34080003", 17587 => x"b4c22000", 17588 => x"28850000",
    17589 => x"b4e22000", 17590 => x"34420004", 17591 => x"58850000",
    17592 => x"c8622000", 17593 => x"5488fffa", 17594 => x"3463fffc",
    17595 => x"00620002", 17596 => x"20630003", 17597 => x"34420001",
    17598 => x"3c420002", 17599 => x"b4e23800", 17600 => x"b4c23000",
    17601 => x"44600008", 17602 => x"34020000", 17603 => x"b4c22000",
    17604 => x"40850000", 17605 => x"b4e22000", 17606 => x"34420001",
    17607 => x"30850000", 17608 => x"5c43fffb", 17609 => x"c3a00000",
    17610 => x"20250003", 17611 => x"b8202000", 17612 => x"44a0000b",
    17613 => x"4460002c", 17614 => x"3463ffff", 17615 => x"204600ff",
    17616 => x"e0000003", 17617 => x"44600028", 17618 => x"3463ffff",
    17619 => x"30860000", 17620 => x"34840001", 17621 => x"20850003",
    17622 => x"5ca0fffb", 17623 => x"34050003", 17624 => x"50a3001a",
    17625 => x"204500ff", 17626 => x"3ca60008", 17627 => x"340a000f",
    17628 => x"b8c52800", 17629 => x"3ca60010", 17630 => x"b8804000",
    17631 => x"b8c53000", 17632 => x"b8603800", 17633 => x"b8802800",
    17634 => x"3409000f", 17635 => x"546a0017", 17636 => x"34040000",
    17637 => x"34070003", 17638 => x"b5042800", 17639 => x"34840004",
    17640 => x"58a60000", 17641 => x"c8642800", 17642 => x"54a7fffc",
    17643 => x"3463fffc", 17644 => x"00640002", 17645 => x"20630003",
    17646 => x"34840001", 17647 => x"3c840002", 17648 => x"b5044000",
    17649 => x"b9002000", 17650 => x"44600007", 17651 => x"204200ff",
    17652 => x"34050000", 17653 => x"b4853000", 17654 => x"30c20000",
    17655 => x"34a50001", 17656 => x"5c65fffd", 17657 => x"c3a00000",
    17658 => x"58a60000", 17659 => x"58a60004", 17660 => x"58a60008",
    17661 => x"58a6000c", 17662 => x"34e7fff0", 17663 => x"34a50010",
    17664 => x"54e9fffa", 17665 => x"3463fff0", 17666 => x"00680004",
    17667 => x"2063000f", 17668 => x"35080001", 17669 => x"3d080004",
    17670 => x"b4884000", 17671 => x"34040003", 17672 => x"5464ffdc",
    17673 => x"b9002000", 17674 => x"e3ffffe8", 17675 => x"78030001",
    17676 => x"38634d50", 17677 => x"28670000", 17678 => x"b8204800",
    17679 => x"34030000", 17680 => x"34060001", 17681 => x"e0000009",
    17682 => x"40840000", 17683 => x"b4e44000", 17684 => x"41080001",
    17685 => x"21080003", 17686 => x"45060012", 17687 => x"c8a40800",
    17688 => x"5c200013", 17689 => x"44810012", 17690 => x"b5232800",
    17691 => x"40a50000", 17692 => x"b4432000", 17693 => x"34630001",
    17694 => x"b4e54000", 17695 => x"41080001", 17696 => x"21080003",
    17697 => x"5d06fff1", 17698 => x"40840000", 17699 => x"34a50020",
    17700 => x"b4e44000", 17701 => x"41080001", 17702 => x"21080003",
    17703 => x"5d06fff0", 17704 => x"34840020", 17705 => x"c8a40800",
    17706 => x"4420ffef", 17707 => x"c3a00000", 17708 => x"b8412800",
    17709 => x"20a50003", 17710 => x"b8403800", 17711 => x"b8202000",
    17712 => x"5ca00018", 17713 => x"78040001", 17714 => x"388442b0",
    17715 => x"28430000", 17716 => x"28880000", 17717 => x"78040001",
    17718 => x"388442b4", 17719 => x"28870000", 17720 => x"a4603000",
    17721 => x"b4682000", 17722 => x"a0c43000", 17723 => x"a0c73000",
    17724 => x"b8202000", 17725 => x"5cc5000a", 17726 => x"58830000",
    17727 => x"34420004", 17728 => x"28430000", 17729 => x"34840004",
    17730 => x"a4603000", 17731 => x"b4682800", 17732 => x"a0c52800",
    17733 => x"a0a72800", 17734 => x"44a0fff8", 17735 => x"b8403800",
    17736 => x"34030000", 17737 => x"b4e32800", 17738 => x"40a50000",
    17739 => x"b4833000", 17740 => x"34630001", 17741 => x"30c50000",
    17742 => x"5ca0fffb", 17743 => x"c3a00000", 17744 => x"20220003",
    17745 => x"4440002c", 17746 => x"40230000", 17747 => x"34020000",
    17748 => x"44600027", 17749 => x"b8201000", 17750 => x"e0000003",
    17751 => x"40430000", 17752 => x"44600022", 17753 => x"34420001",
    17754 => x"20430003", 17755 => x"5c60fffc", 17756 => x"78040001",
    17757 => x"388442b0", 17758 => x"28430000", 17759 => x"28860000",
    17760 => x"78040001", 17761 => x"388442b4", 17762 => x"28850000",
    17763 => x"a4602000", 17764 => x"b4661800", 17765 => x"a0641800",
    17766 => x"a0651800", 17767 => x"5c600011", 17768 => x"34420004",
    17769 => x"28430000", 17770 => x"b4662000", 17771 => x"a4601800",
    17772 => x"a0831800", 17773 => x"a0651800", 17774 => x"5c60000a",
    17775 => x"34420004", 17776 => x"28430000", 17777 => x"b4662000",
    17778 => x"a4601800", 17779 => x"a0831800", 17780 => x"a0651800",
    17781 => x"4460fff3", 17782 => x"e0000002", 17783 => x"34420001",
    17784 => x"40430000", 17785 => x"5c60fffe", 17786 => x"c8411000",
    17787 => x"b8400800", 17788 => x"c3a00000", 17789 => x"b8201000",
    17790 => x"e3ffffde", 17791 => x"34060000", 17792 => x"44600017",
    17793 => x"b8413800", 17794 => x"20e70003", 17795 => x"3464ffff",
    17796 => x"44e00015", 17797 => x"40230000", 17798 => x"40450000",
    17799 => x"5c65000f", 17800 => x"34060000", 17801 => x"4480000e",
    17802 => x"34210001", 17803 => x"34420001", 17804 => x"5c600004",
    17805 => x"e000000a", 17806 => x"44800033", 17807 => x"44600032",
    17808 => x"40230000", 17809 => x"40450000", 17810 => x"3484ffff",
    17811 => x"34210001", 17812 => x"34420001", 17813 => x"4465fff9",
    17814 => x"c8653000", 17815 => x"b8c00800", 17816 => x"c3a00000",
    17817 => x"b8202800", 17818 => x"34010003", 17819 => x"b8402000",
    17820 => x"50230028", 17821 => x"28a10000", 17822 => x"28420000",
    17823 => x"5c220025", 17824 => x"3463fffc", 17825 => x"b8e03000",
    17826 => x"4460fff5", 17827 => x"78020001", 17828 => x"384242b0",
    17829 => x"28490000", 17830 => x"78020001", 17831 => x"384242b4",
    17832 => x"28480000", 17833 => x"a4201000", 17834 => x"b4290800",
    17835 => x"a0220800", 17836 => x"a0280800", 17837 => x"34070003",
    17838 => x"5c20ffe9", 17839 => x"34a50004", 17840 => x"34840004",
    17841 => x"54670006", 17842 => x"b8a00800", 17843 => x"b8801000",
    17844 => x"44600014", 17845 => x"3464ffff", 17846 => x"e3ffffcf",
    17847 => x"28a10000", 17848 => x"288a0000", 17849 => x"b4293000",
    17850 => x"a4201000", 17851 => x"a0c21000", 17852 => x"a0481000",
    17853 => x"5c2a0007", 17854 => x"3463fffc", 17855 => x"44600002",
    17856 => x"4440ffef", 17857 => x"34060000", 17858 => x"b8c00800",
    17859 => x"c3a00000", 17860 => x"b8801000", 17861 => x"b8a00800",
    17862 => x"3464ffff", 17863 => x"e3ffffbe", 17864 => x"40a30000",
    17865 => x"40850000", 17866 => x"c8653000", 17867 => x"e3ffffcc",
    17868 => x"b8412000", 17869 => x"20840003", 17870 => x"74650003",
    17871 => x"64840000", 17872 => x"b8403000", 17873 => x"a0852000",
    17874 => x"b8202800", 17875 => x"44800015", 17876 => x"78040001",
    17877 => x"388442b0", 17878 => x"28890000", 17879 => x"78040001",
    17880 => x"388442b4", 17881 => x"28880000", 17882 => x"340a0003",
    17883 => x"e0000006", 17884 => x"58a40000", 17885 => x"3463fffc",
    17886 => x"34a50004", 17887 => x"34420004", 17888 => x"51430007",
    17889 => x"28440000", 17890 => x"a4803800", 17891 => x"b4893000",
    17892 => x"a0e63000", 17893 => x"a0c83000", 17894 => x"44c0fff6",
    17895 => x"b8403000", 17896 => x"44600014", 17897 => x"40c20000",
    17898 => x"3463ffff", 17899 => x"34a40001", 17900 => x"30a20000",
    17901 => x"44400009", 17902 => x"34c20001", 17903 => x"4460000e",
    17904 => x"40450000", 17905 => x"3463ffff", 17906 => x"34420001",
    17907 => x"30850000", 17908 => x"34840001", 17909 => x"5ca0fffa",
    17910 => x"34020000", 17911 => x"44600007", 17912 => x"b4822800",
    17913 => x"30a00000", 17914 => x"34420001", 17915 => x"5c62fffd",
    17916 => x"c3a00000", 17917 => x"c3a00000", 17918 => x"c3a00000",
    17919 => x"57522043", 17920 => x"6f72653a", 17921 => x"20737461",
    17922 => x"7274696e", 17923 => x"67207570", 17924 => x"2e2e2e0a",
    17925 => x"00000000", 17926 => x"556e6162", 17927 => x"6c652074",
    17928 => x"6f206465", 17929 => x"7465726d", 17930 => x"696e6520",
    17931 => x"4d414320", 17932 => x"61646472", 17933 => x"6573730a",
    17934 => x"00000000", 17935 => x"4c6f6361", 17936 => x"6c204d41",
    17937 => x"43206164", 17938 => x"64726573", 17939 => x"733a2025",
    17940 => x"3032783a", 17941 => x"25303278", 17942 => x"3a253032",
    17943 => x"783a2530", 17944 => x"32783a25", 17945 => x"3032783a",
    17946 => x"25303278", 17947 => x"0a000000", 17948 => x"4c696e6b",
    17949 => x"2075702e", 17950 => x"0a000000", 17951 => x"4c696e6b",
    17952 => x"20646f77", 17953 => x"6e2e0a00", 17954 => x"25750000",
    17955 => x"25752575", 17956 => x"00000000", 17957 => x"0a0a5054",
    17958 => x"50207374", 17959 => x"61747573", 17960 => x"3a200000",
    17961 => x"25730000", 17962 => x"0a0a5379", 17963 => x"6e632069",
    17964 => x"6e666f20", 17965 => x"6e6f7420", 17966 => x"76616c69",
    17967 => x"640a0a00", 17968 => x"0a0a5379", 17969 => x"6e636872",
    17970 => x"6f6e697a", 17971 => x"6174696f", 17972 => x"6e207374",
    17973 => x"61747573", 17974 => x"3a0a0a00", 17975 => x"57522050",
    17976 => x"54502043", 17977 => x"6f726520", 17978 => x"53796e63",
    17979 => x"204d6f6e", 17980 => x"69746f72", 17981 => x"20762031",
    17982 => x"2e300000", 17983 => x"45736320", 17984 => x"3d206578",
    17985 => x"69740000", 17986 => x"0a0a5441", 17987 => x"49205469",
    17988 => x"6d653a20", 17989 => x"20202020", 17990 => x"20202020",
    17991 => x"20202020", 17992 => x"20202020", 17993 => x"20000000",
    17994 => x"0a0a4c69", 17995 => x"6e6b2073", 17996 => x"74617475",
    17997 => x"733a0000", 17998 => x"25733a20", 17999 => x"00000000",
    18000 => x"77727531", 18001 => x"00000000", 18002 => x"4c696e6b",
    18003 => x"20757020", 18004 => x"20200000", 18005 => x"4c696e6b",
    18006 => x"20646f77", 18007 => x"6e200000", 18008 => x"2852583a",
    18009 => x"2025642c", 18010 => x"2054583a", 18011 => x"20256429",
    18012 => x"2c206d6f", 18013 => x"64653a20", 18014 => x"00000000",
    18015 => x"5752204f", 18016 => x"66660000", 18017 => x"436c6f63",
    18018 => x"6b206f66", 18019 => x"66736574", 18020 => x"3a202020",
    18021 => x"20202020", 18022 => x"20202020", 18023 => x"20202020",
    18024 => x"20200000", 18025 => x"2532692e", 18026 => x"25303969",
    18027 => x"20730000", 18028 => x"25396920", 18029 => x"6e730000",
    18030 => x"0a4f6e65", 18031 => x"2d776179", 18032 => x"2064656c",
    18033 => x"61792061", 18034 => x"76657261", 18035 => x"6765643a",
    18036 => x"20202020", 18037 => x"20202000", 18038 => x"0a4f6273",
    18039 => x"65727665", 18040 => x"64206472", 18041 => x"6966743a",
    18042 => x"20202020", 18043 => x"20202020", 18044 => x"20202020",
    18045 => x"20202000", 18046 => x"5752204d", 18047 => x"61737465",
    18048 => x"72202000", 18049 => x"57522053", 18050 => x"6c617665",
    18051 => x"20202000", 18052 => x"57522055", 18053 => x"6e6b6e6f",
    18054 => x"776e2020", 18055 => x"20000000", 18056 => x"4c6f636b",
    18057 => x"65642020", 18058 => x"00000000", 18059 => x"4e6f4c6f",
    18060 => x"636b2020", 18061 => x"00000000", 18062 => x"43616c69",
    18063 => x"62726174", 18064 => x"65642020", 18065 => x"00000000",
    18066 => x"556e6361", 18067 => x"6c696272", 18068 => x"61746564",
    18069 => x"20200000", 18070 => x"0a495076", 18071 => x"343a2000",
    18072 => x"424f4f54", 18073 => x"50207275", 18074 => x"6e6e696e",
    18075 => x"67000000", 18076 => x"25642e25", 18077 => x"642e2564",
    18078 => x"2e256400", 18079 => x"53657276", 18080 => x"6f207374",
    18081 => x"6174653a", 18082 => x"20202020", 18083 => x"20202020",
    18084 => x"20202020", 18085 => x"20202000", 18086 => x"50686173",
    18087 => x"65207472", 18088 => x"61636b69", 18089 => x"6e673a20",
    18090 => x"20202020", 18091 => x"20202020", 18092 => x"20202000",
    18093 => x"4f4e0a00", 18094 => x"4f46460a", 18095 => x"00000000",
    18096 => x"41757820", 18097 => x"636c6f63", 18098 => x"6b207374",
    18099 => x"61747573", 18100 => x"3a202020", 18101 => x"20202020",
    18102 => x"20202000", 18103 => x"656e6162", 18104 => x"6c656400",
    18105 => x"2c206c6f", 18106 => x"636b6564", 18107 => x"00000000",
    18108 => x"0a54696d", 18109 => x"696e6720", 18110 => x"70617261",
    18111 => x"6d657465", 18112 => x"72733a0a", 18113 => x"0a000000",
    18114 => x"526f756e", 18115 => x"642d7472", 18116 => x"69702074",
    18117 => x"696d6520", 18118 => x"286d7529", 18119 => x"3a202020",
    18120 => x"20000000", 18121 => x"25732070", 18122 => x"730a0000",
    18123 => x"4d617374", 18124 => x"65722d73", 18125 => x"6c617665",
    18126 => x"2064656c", 18127 => x"61793a20", 18128 => x"20202020",
    18129 => x"20000000", 18130 => x"4d617374", 18131 => x"65722050",
    18132 => x"48592064", 18133 => x"656c6179", 18134 => x"733a2020",
    18135 => x"20202020", 18136 => x"20000000", 18137 => x"54583a20",
    18138 => x"25642070", 18139 => x"732c2052", 18140 => x"583a2025",
    18141 => x"64207073", 18142 => x"0a000000", 18143 => x"536c6176",
    18144 => x"65205048", 18145 => x"59206465", 18146 => x"6c617973",
    18147 => x"3a202020", 18148 => x"20202020", 18149 => x"20000000",
    18150 => x"546f7461", 18151 => x"6c206c69", 18152 => x"6e6b2061",
    18153 => x"73796d6d", 18154 => x"65747279", 18155 => x"3a202020",
    18156 => x"20000000", 18157 => x"25396420", 18158 => x"70730a00",
    18159 => x"4361626c", 18160 => x"65207274", 18161 => x"74206465",
    18162 => x"6c61793a", 18163 => x"20202020", 18164 => x"20202020",
    18165 => x"20000000", 18166 => x"436c6f63", 18167 => x"6b206f66",
    18168 => x"66736574", 18169 => x"3a202020", 18170 => x"20202020",
    18171 => x"20202020", 18172 => x"20000000", 18173 => x"50686173",
    18174 => x"65207365", 18175 => x"74706f69", 18176 => x"6e743a20",
    18177 => x"20202020", 18178 => x"20202020", 18179 => x"20000000",
    18180 => x"536b6577", 18181 => x"3a202020", 18182 => x"20202020",
    18183 => x"20202020", 18184 => x"20202020", 18185 => x"20202020",
    18186 => x"20000000", 18187 => x"4d616e75", 18188 => x"616c2070",
    18189 => x"68617365", 18190 => x"2061646a", 18191 => x"7573746d",
    18192 => x"656e743a", 18193 => x"20000000", 18194 => x"55706461",
    18195 => x"74652063", 18196 => x"6f756e74", 18197 => x"65723a20",
    18198 => x"20202020", 18199 => x"20202020", 18200 => x"20000000",
    18201 => x"2539640a", 18202 => x"00000000", 18203 => x"2d2d0000",
    18204 => x"6c6e6b3a", 18205 => x"25642072", 18206 => x"783a2564",
    18207 => x"2074783a", 18208 => x"25642000", 18209 => x"6c6f636b",
    18210 => x"3a256420", 18211 => x"00000000", 18212 => x"7074703a",
    18213 => x"25732000", 18214 => x"73763a25", 18215 => x"64200000",
    18216 => x"73733a27", 18217 => x"25732720", 18218 => x"00000000",
    18219 => x"6175783a", 18220 => x"25782000", 18221 => x"7365633a",
    18222 => x"2564206e", 18223 => x"7365633a", 18224 => x"25642000",
    18225 => x"6d753a25", 18226 => x"73200000", 18227 => x"646d733a",
    18228 => x"25732000", 18229 => x"6474786d", 18230 => x"3a256420",
    18231 => x"6472786d", 18232 => x"3a256420", 18233 => x"00000000",
    18234 => x"64747873", 18235 => x"3a256420", 18236 => x"64727873",
    18237 => x"3a256420", 18238 => x"00000000", 18239 => x"6173796d",
    18240 => x"3a256420", 18241 => x"00000000", 18242 => x"63727474",
    18243 => x"3a257320", 18244 => x"00000000", 18245 => x"636b6f3a",
    18246 => x"25642000", 18247 => x"73657470", 18248 => x"3a256420",
    18249 => x"00000000", 18250 => x"75636e74", 18251 => x"3a256420",
    18252 => x"00000000", 18253 => x"68643a25", 18254 => x"64206d64",
    18255 => x"3a256420", 18256 => x"61643a25", 18257 => x"64200000",
    18258 => x"74656d70", 18259 => x"3a202564", 18260 => x"2e253034",
    18261 => x"64204300", 18262 => x"756e6b6e", 18263 => x"6f776e00",
    18264 => x"64696167", 18265 => x"2d66736d", 18266 => x"2d312d25",
    18267 => x"733a2025", 18268 => x"3039642e", 18269 => x"25303364",
    18270 => x"3a200000", 18271 => x"454e5445", 18272 => x"52202573",
    18273 => x"2c207061", 18274 => x"636b6574", 18275 => x"206c656e",
    18276 => x"2025690a", 18277 => x"00000000", 18278 => x"25733a20",
    18279 => x"7265656e", 18280 => x"74657220", 18281 => x"696e2025",
    18282 => x"69206d73", 18283 => x"0a000000", 18284 => x"4c454156",
    18285 => x"45202573", 18286 => x"20286e65", 18287 => x"78743a20",
    18288 => x"25336929", 18289 => x"0a0a0000", 18290 => x"52454356",
    18291 => x"20253032", 18292 => x"64206279", 18293 => x"74657320",
    18294 => x"61742025", 18295 => x"642e2530", 18296 => x"39642028",
    18297 => x"74797065", 18298 => x"2025782c", 18299 => x"20257329",
    18300 => x"0a000000", 18301 => x"66736d20", 18302 => x"666f7220",
    18303 => x"25733a20", 18304 => x"4572726f", 18305 => x"72202569",
    18306 => x"20696e20", 18307 => x"25730a00", 18308 => x"66736d3a",
    18309 => x"20556e6b", 18310 => x"6e6f776e", 18311 => x"20737461",
    18312 => x"74652066", 18313 => x"6f722070", 18314 => x"6f727420",
    18315 => x"25730a00", 18316 => x"70707369", 18317 => x"00000000",
    18318 => x"25732d25", 18319 => x"692d2573", 18320 => x"3a200000",
    18321 => x"25733a20", 18322 => x"6572726f", 18323 => x"72207061",
    18324 => x"7273696e", 18325 => x"67202225", 18326 => x"73220a00",
    18327 => x"64696167", 18328 => x"2d636f6e", 18329 => x"66696700",
    18330 => x"64696167", 18331 => x"2d657874", 18332 => x"656e7369",
    18333 => x"6f6e0000", 18334 => x"64696167", 18335 => x"2d626d63",
    18336 => x"00000000", 18337 => x"64696167", 18338 => x"2d736572",
    18339 => x"766f0000", 18340 => x"64696167", 18341 => x"2d667261",
    18342 => x"6d657300", 18343 => x"64696167", 18344 => x"2d74696d",
    18345 => x"65000000", 18346 => x"64696167", 18347 => x"2d66736d",
    18348 => x"00000000", 18349 => x"50505369", 18350 => x"20666f72",
    18351 => x"20575250", 18352 => x"432e2043", 18353 => x"6f6d6d69",
    18354 => x"74202573", 18355 => x"2c206275", 18356 => x"696c7420",
    18357 => x"6f6e204a", 18358 => x"756e2031", 18359 => x"34203230",
    18360 => x"31360a00", 18361 => x"70707369", 18362 => x"2d763230",
    18363 => x"31342e30", 18364 => x"372d3137", 18365 => x"332d6762",
    18366 => x"32303363", 18367 => x"63390000", 18368 => x"4c6f636b",
    18369 => x"696e6720", 18370 => x"504c4c00", 18371 => x"0a4c6f63",
    18372 => x"6b207469", 18373 => x"6d656f75", 18374 => x"742e0000",
    18375 => x"2e000000", 18376 => x"4c696e6b", 18377 => x"20646f77",
    18378 => x"6e3a2050", 18379 => x"54502073", 18380 => x"746f700a",
    18381 => x"00000000", 18382 => x"4c696e6b", 18383 => x"2075703a",
    18384 => x"20505450", 18385 => x"20737461", 18386 => x"72740a00",
    18387 => x"77723100", 18388 => x"25732573", 18389 => x"25303278",
    18390 => x"2d253032", 18391 => x"782d2530", 18392 => x"32782d25",
    18393 => x"3032782d", 18394 => x"25303278", 18395 => x"2d253032",
    18396 => x"782d2530", 18397 => x"32782d25", 18398 => x"3032782d",
    18399 => x"25303278", 18400 => x"2d253032", 18401 => x"780a0000",
    18402 => x"25732573", 18403 => x"25732028", 18404 => x"73697a65",
    18405 => x"20256929", 18406 => x"0a000000", 18407 => x"25732573",
    18408 => x"00000000", 18409 => x"25303278", 18410 => x"00000000",
    18411 => x"25735645", 18412 => x"5253494f", 18413 => x"4e3a2075",
    18414 => x"6e737570", 18415 => x"706f7274", 18416 => x"65642028",
    18417 => x"2569290a", 18418 => x"00000000", 18419 => x"25735645",
    18420 => x"5253494f", 18421 => x"4e3a2025", 18422 => x"69202874",
    18423 => x"79706520", 18424 => x"25692c20", 18425 => x"6c656e20",
    18426 => x"25692c20", 18427 => x"646f6d61", 18428 => x"696e2025",
    18429 => x"69290a00", 18430 => x"2573464c", 18431 => x"4147533a",
    18432 => x"20307825", 18433 => x"30347820", 18434 => x"28636f72",
    18435 => x"72656374", 18436 => x"696f6e20", 18437 => x"2530386c",
    18438 => x"75290a00", 18439 => x"504f5254", 18440 => x"3a200000",
    18441 => x"25735245", 18442 => x"53543a20", 18443 => x"73657120",
    18444 => x"25692c20", 18445 => x"6374726c", 18446 => x"2025692c",
    18447 => x"206c6f67", 18448 => x"2d696e74", 18449 => x"65727661",
    18450 => x"6c202569", 18451 => x"0a000000", 18452 => x"25734d45",
    18453 => x"53534147", 18454 => x"453a2028", 18455 => x"45292053",
    18456 => x"594e430a", 18457 => x"00000000", 18458 => x"25732573",
    18459 => x"256c752e", 18460 => x"25303969", 18461 => x"0a000000",
    18462 => x"4d53472d", 18463 => x"53594e43", 18464 => x"3a200000",
    18465 => x"25734d45", 18466 => x"53534147", 18467 => x"453a2028",
    18468 => x"45292044", 18469 => x"454c4159", 18470 => x"5f524551",
    18471 => x"0a000000", 18472 => x"4d53472d", 18473 => x"44454c41",
    18474 => x"595f5245", 18475 => x"513a2000", 18476 => x"25734d45",
    18477 => x"53534147", 18478 => x"453a2028", 18479 => x"47292046",
    18480 => x"4f4c4c4f", 18481 => x"575f5550", 18482 => x"0a000000",
    18483 => x"4d53472d", 18484 => x"464f4c4c", 18485 => x"4f575f55",
    18486 => x"503a2000", 18487 => x"25734d45", 18488 => x"53534147",
    18489 => x"453a2028", 18490 => x"47292044", 18491 => x"454c4159",
    18492 => x"5f524553", 18493 => x"500a0000", 18494 => x"4d53472d",
    18495 => x"44454c41", 18496 => x"595f5245", 18497 => x"53503a20",
    18498 => x"00000000", 18499 => x"25734d45", 18500 => x"53534147",
    18501 => x"453a2028", 18502 => x"47292041", 18503 => x"4e4e4f55",
    18504 => x"4e43450a", 18505 => x"00000000", 18506 => x"4d53472d",
    18507 => x"414e4e4f", 18508 => x"554e4345", 18509 => x"3a207374",
    18510 => x"616d7020", 18511 => x"00000000", 18512 => x"25732573",
    18513 => x"25303278", 18514 => x"2d253032", 18515 => x"782d2530",
    18516 => x"34780a00", 18517 => x"4d53472d", 18518 => x"414e4e4f",
    18519 => x"554e4345", 18520 => x"3a206772", 18521 => x"616e646d",
    18522 => x"61737465", 18523 => x"722d7175", 18524 => x"616c6974",
    18525 => x"79200000", 18526 => x"25734d53", 18527 => x"472d414e",
    18528 => x"4e4f554e", 18529 => x"43453a20", 18530 => x"6772616e",
    18531 => x"646d6173", 18532 => x"7465722d", 18533 => x"7072696f",
    18534 => x"20256920", 18535 => x"25690a00", 18536 => x"25732573",
    18537 => x"25303278", 18538 => x"2d253032", 18539 => x"782d2530",
    18540 => x"32782d25", 18541 => x"3032782d", 18542 => x"25303278",
    18543 => x"2d253032", 18544 => x"782d2530", 18545 => x"32782d25",
    18546 => x"3032780a", 18547 => x"00000000", 18548 => x"4d53472d",
    18549 => x"414e4e4f", 18550 => x"554e4345", 18551 => x"3a206772",
    18552 => x"616e646d", 18553 => x"61737465", 18554 => x"722d6964",
    18555 => x"20000000", 18556 => x"25734d45", 18557 => x"53534147",
    18558 => x"453a2028", 18559 => x"47292053", 18560 => x"49474e41",
    18561 => x"4c494e47", 18562 => x"0a000000", 18563 => x"4d53472d",
    18564 => x"5349474e", 18565 => x"414c494e", 18566 => x"473a2074",
    18567 => x"61726765", 18568 => x"742d706f", 18569 => x"72742000",
    18570 => x"2573544c", 18571 => x"563a2074", 18572 => x"6f6f2073",
    18573 => x"686f7274", 18574 => x"20282569", 18575 => x"202d2025",
    18576 => x"69203d20", 18577 => x"2569290a", 18578 => x"00000000",
    18579 => x"2573544c", 18580 => x"563a2074", 18581 => x"79706520",
    18582 => x"25303478", 18583 => x"206c656e", 18584 => x"20256920",
    18585 => x"6f756920", 18586 => x"25303278", 18587 => x"3a253032",
    18588 => x"783a2530", 18589 => x"32782073", 18590 => x"75622025",
    18591 => x"3032783a", 18592 => x"25303278", 18593 => x"3a253032",
    18594 => x"780a0000", 18595 => x"2573544c", 18596 => x"563a2074",
    18597 => x"6f6f2073", 18598 => x"686f7274", 18599 => x"20286578",
    18600 => x"70656374", 18601 => x"65642025", 18602 => x"692c2074",
    18603 => x"6f74616c", 18604 => x"20256929", 18605 => x"0a000000",
    18606 => x"544c563a", 18607 => x"20000000", 18608 => x"746c762d",
    18609 => x"636f6e74", 18610 => x"656e7400", 18611 => x"44554d50",
    18612 => x"3a200000", 18613 => x"7061796c", 18614 => x"6f616400",
    18615 => x"20696e76", 18616 => x"616c6964", 18617 => x"00000000",
    18618 => x"25735449", 18619 => x"4d453a20", 18620 => x"28256c69",
    18621 => x"202d2030", 18622 => x"78256c78", 18623 => x"2920256c",
    18624 => x"692e2530", 18625 => x"366c6925", 18626 => x"730a0000",
    18627 => x"2573564c", 18628 => x"414e2025", 18629 => x"690a0000",
    18630 => x"25734554", 18631 => x"483a2025", 18632 => x"30347820",
    18633 => x"28253032", 18634 => x"783a2530", 18635 => x"32783a25",
    18636 => x"3032783a", 18637 => x"25303278", 18638 => x"3a253032",
    18639 => x"783a2530", 18640 => x"3278202d", 18641 => x"3e202530",
    18642 => x"32783a25", 18643 => x"3032783a", 18644 => x"25303278",
    18645 => x"3a253032", 18646 => x"783a2530", 18647 => x"32783a25",
    18648 => x"30327829", 18649 => x"0a000000", 18650 => x"25734950",
    18651 => x"3a202569", 18652 => x"20282569", 18653 => x"2e25692e",
    18654 => x"25692e25", 18655 => x"69202d3e", 18656 => x"2025692e",
    18657 => x"25692e25", 18658 => x"692e2569", 18659 => x"29206c65",
    18660 => x"6e202569", 18661 => x"0a000000", 18662 => x"25735544",
    18663 => x"503a2028", 18664 => x"2569202d", 18665 => x"3e202569",
    18666 => x"29206c65", 18667 => x"6e202569", 18668 => x"0a000000",
    18669 => x"25733a20", 18670 => x"256c690a", 18671 => x"00000000",
    18672 => x"5761726e", 18673 => x"696e673a", 18674 => x"2025733a",
    18675 => x"2063616e", 18676 => x"206e6f74", 18677 => x"2061646a",
    18678 => x"75737420", 18679 => x"66726571", 18680 => x"5f707062",
    18681 => x"20256c69", 18682 => x"0a000000", 18683 => x"25733a20",
    18684 => x"25396c75", 18685 => x"2e253039", 18686 => x"6c690a00",
    18687 => x"25733a20", 18688 => x"736e743d", 18689 => x"25642c20",
    18690 => x"7365633d", 18691 => x"25642c20", 18692 => x"6e736563",
    18693 => x"3d25640a", 18694 => x"00000000", 18695 => x"73656e64",
    18696 => x"3a200000", 18697 => x"72656376", 18698 => x"3a200000",
    18699 => x"696e6974", 18700 => x"69616c69", 18701 => x"7a696e67",
    18702 => x"00000000", 18703 => x"6661756c", 18704 => x"74790000",
    18705 => x"64697361", 18706 => x"626c6564", 18707 => x"00000000",
    18708 => x"6c697374", 18709 => x"656e696e", 18710 => x"67000000",
    18711 => x"756e6361", 18712 => x"6c696272", 18713 => x"61746564",
    18714 => x"00000000", 18715 => x"736c6176", 18716 => x"65000000",
    18717 => x"756e6361", 18718 => x"6c696272", 18719 => x"61746564",
    18720 => x"2f77722d", 18721 => x"70726573", 18722 => x"656e7400",
    18723 => x"6d617374", 18724 => x"65722f77", 18725 => x"722d6d2d",
    18726 => x"6c6f636b", 18727 => x"00000000", 18728 => x"756e6361",
    18729 => x"6c696272", 18730 => x"61746564", 18731 => x"2f77722d",
    18732 => x"732d6c6f", 18733 => x"636b0000", 18734 => x"756e6361",
    18735 => x"6c696272", 18736 => x"61746564", 18737 => x"2f77722d",
    18738 => x"6c6f636b", 18739 => x"65640000", 18740 => x"77722d63",
    18741 => x"616c6962", 18742 => x"72617469", 18743 => x"6f6e0000",
    18744 => x"77722d63", 18745 => x"616c6962", 18746 => x"72617465",
    18747 => x"64000000", 18748 => x"77722d72", 18749 => x"6573702d",
    18750 => x"63616c69", 18751 => x"622d7265", 18752 => x"71000000",
    18753 => x"77722d6c", 18754 => x"696e6b2d", 18755 => x"6f6e0000",
    18756 => x"686f6f6b", 18757 => x"3a202573", 18758 => x"0a000000",
    18759 => x"5432206f", 18760 => x"72205433", 18761 => x"20696e63",
    18762 => x"6f727265", 18763 => x"63742c20", 18764 => x"64697363",
    18765 => x"61726469", 18766 => x"6e672074", 18767 => x"75706c65",
    18768 => x"0a000000", 18769 => x"48616e64", 18770 => x"7368616b",
    18771 => x"65206661", 18772 => x"696c7572", 18773 => x"653a206e",
    18774 => x"6f77206e", 18775 => x"6f6e2d77", 18776 => x"72202573",
    18777 => x"0a000000", 18778 => x"52657472", 18779 => x"79206f6e",
    18780 => x"2074696d", 18781 => x"656f7574", 18782 => x"0a000000",
    18783 => x"25733a20", 18784 => x"73756273", 18785 => x"74617465",
    18786 => x"2025690a", 18787 => x"00000000", 18788 => x"54783d3e",
    18789 => x"3e736361", 18790 => x"6c656450", 18791 => x"69636f73",
    18792 => x"65636f6e", 18793 => x"64732e6d", 18794 => x"7362203d",
    18795 => x"20307825", 18796 => x"780a0000", 18797 => x"54783d3e",
    18798 => x"3e736361", 18799 => x"6c656450", 18800 => x"69636f73",
    18801 => x"65636f6e", 18802 => x"64732e6c", 18803 => x"7362203d",
    18804 => x"20307825", 18805 => x"780a0000", 18806 => x"52782066",
    18807 => x"69786564", 18808 => x"2064656c", 18809 => x"6179203d",
    18810 => x"2025640a", 18811 => x"00000000", 18812 => x"52783d3e",
    18813 => x"3e736361", 18814 => x"6c656450", 18815 => x"69636f73",
    18816 => x"65636f6e", 18817 => x"64732e6d", 18818 => x"7362203d",
    18819 => x"20307825", 18820 => x"780a0000", 18821 => x"52783d3e",
    18822 => x"3e736361", 18823 => x"6c656450", 18824 => x"69636f73",
    18825 => x"65636f6e", 18826 => x"64732e6c", 18827 => x"7362203d",
    18828 => x"20307825", 18829 => x"780a0000", 18830 => x"4552524f",
    18831 => x"523a204e", 18832 => x"65772063", 18833 => x"6c617373",
    18834 => x"2025690a", 18835 => x"00000000", 18836 => x"4255473a",
    18837 => x"20547279", 18838 => x"696e6720", 18839 => x"746f2073",
    18840 => x"656e6420", 18841 => x"696e7661", 18842 => x"6c696420",
    18843 => x"77725f6d", 18844 => x"7367206d", 18845 => x"6f64653d",
    18846 => x"25782069", 18847 => x"643d2578", 18848 => x"00000000",
    18849 => x"68616e64", 18850 => x"6c652053", 18851 => x"69676e61",
    18852 => x"6c696e67", 18853 => x"206d7367", 18854 => x"2c206661",
    18855 => x"696c6564", 18856 => x"2c205468", 18857 => x"69732069",
    18858 => x"73206e6f", 18859 => x"74206f72", 18860 => x"67616e69",
    18861 => x"7a617469", 18862 => x"6f6e2065", 18863 => x"7874656e",
    18864 => x"73696f6e", 18865 => x"20544c56", 18866 => x"203d2030",
    18867 => x"7825780a", 18868 => x"00000000", 18869 => x"68616e64",
    18870 => x"6c652053", 18871 => x"69676e61", 18872 => x"6c696e67",
    18873 => x"206d7367", 18874 => x"2c206661", 18875 => x"696c6564",
    18876 => x"2c206e6f", 18877 => x"74204345", 18878 => x"524e2773",
    18879 => x"204f5549", 18880 => x"203d2030", 18881 => x"7825780a",
    18882 => x"00000000", 18883 => x"68616e64", 18884 => x"6c652053",
    18885 => x"69676e61", 18886 => x"6c696e67", 18887 => x"206d7367",
    18888 => x"2c206661", 18889 => x"696c6564", 18890 => x"2c206e6f",
    18891 => x"74205768", 18892 => x"69746520", 18893 => x"52616262",
    18894 => x"6974206d", 18895 => x"61676963", 18896 => x"206e756d",
    18897 => x"62657220", 18898 => x"3d203078", 18899 => x"25780a00",
    18900 => x"68616e64", 18901 => x"6c652053", 18902 => x"69676e61",
    18903 => x"6c696e67", 18904 => x"206d7367", 18905 => x"2c206661",
    18906 => x"696c6564", 18907 => x"2c206e6f", 18908 => x"74207375",
    18909 => x"70706f72", 18910 => x"74656420", 18911 => x"76657273",
    18912 => x"696f6e20", 18913 => x"6e756d62", 18914 => x"6572203d",
    18915 => x"20307825", 18916 => x"780a0000", 18917 => x"25732825",
    18918 => x"6429204d", 18919 => x"65737361", 18920 => x"67652063",
    18921 => x"616e2774", 18922 => x"20626520", 18923 => x"73656e74",
    18924 => x"0a000000", 18925 => x"53454e54", 18926 => x"20253032",
    18927 => x"64206279", 18928 => x"74657320", 18929 => x"61742025",
    18930 => x"642e2530", 18931 => x"39642028", 18932 => x"2573290a",
    18933 => x"00000000", 18934 => x"556e696e", 18935 => x"69746961",
    18936 => x"6c697a65", 18937 => x"64000000", 18938 => x"20287761",
    18939 => x"69742066", 18940 => x"6f722068", 18941 => x"77290000",
    18942 => x"4552524f", 18943 => x"523a2025", 18944 => x"733a2054",
    18945 => x"696d6573", 18946 => x"74616d70", 18947 => x"73496e63",
    18948 => x"6f727265", 18949 => x"63743a20", 18950 => x"25642025",
    18951 => x"64202564", 18952 => x"2025640a", 18953 => x"00000000",
    18954 => x"2573203d", 18955 => x"2025643a", 18956 => x"25643a25",
    18957 => x"640a0000", 18958 => x"73657276", 18959 => x"6f3a7431",
    18960 => x"00000000", 18961 => x"73657276", 18962 => x"6f3a7432",
    18963 => x"00000000", 18964 => x"73657276", 18965 => x"6f3a7433",
    18966 => x"00000000", 18967 => x"73657276", 18968 => x"6f3a7434",
    18969 => x"00000000", 18970 => x"2d3e6d64", 18971 => x"656c6179",
    18972 => x"00000000", 18973 => x"504c4c20", 18974 => x"4f75744f",
    18975 => x"664c6f63", 18976 => x"6b2c2073", 18977 => x"686f756c",
    18978 => x"64207265", 18979 => x"73746172", 18980 => x"74207379",
    18981 => x"6e630a00", 18982 => x"73657276", 18983 => x"6f3a6275",
    18984 => x"73790a00", 18985 => x"6f666673", 18986 => x"65745f68",
    18987 => x"773a2025", 18988 => x"6c692e25", 18989 => x"30396c69",
    18990 => x"20282b25", 18991 => x"6c69290a", 18992 => x"00000000",
    18993 => x"77725f73", 18994 => x"6572766f", 18995 => x"20737461",
    18996 => x"74653a20", 18997 => x"25732573", 18998 => x"0a000000",
    18999 => x"6f6c6473", 19000 => x"65747020", 19001 => x"25692c20",
    19002 => x"6f666673", 19003 => x"65742025", 19004 => x"693a2530",
    19005 => x"34690a00", 19006 => x"61646a75", 19007 => x"73742070",
    19008 => x"68617365", 19009 => x"2025690a", 19010 => x"00000000",
    19011 => x"53594e43", 19012 => x"5f4e5345", 19013 => x"43000000",
    19014 => x"53594e43", 19015 => x"5f534543", 19016 => x"00000000",
    19017 => x"53594e43", 19018 => x"5f504841", 19019 => x"53450000",
    19020 => x"54524143", 19021 => x"4b5f5048", 19022 => x"41534500",
    19023 => x"57414954", 19024 => x"5f4f4646", 19025 => x"5345545f",
    19026 => x"53544142", 19027 => x"4c450000", 19028 => x"7072652d",
    19029 => x"6d617374", 19030 => x"65720000", 19031 => x"70617373",
    19032 => x"69766500", 19033 => x"25733a20", 19034 => x"63616e27",
    19035 => x"7420696e", 19036 => x"69742065", 19037 => x"7874656e",
    19038 => x"73696f6e", 19039 => x"0a000000", 19040 => x"636c6f63",
    19041 => x"6b20636c", 19042 => x"61737320", 19043 => x"3d202564",
    19044 => x"0a000000", 19045 => x"636c6f63", 19046 => x"6b206163",
    19047 => x"63757261", 19048 => x"6379203d", 19049 => x"2025640a",
    19050 => x"00000000", 19051 => x"70705f73", 19052 => x"6c617665",
    19053 => x"203a2044", 19054 => x"656c6179", 19055 => x"20526573",
    19056 => x"7020646f", 19057 => x"65736e27", 19058 => x"74206d61",
    19059 => x"74636820", 19060 => x"44656c61", 19061 => x"79205265",
    19062 => x"710a0000", 19063 => x"4e657720", 19064 => x"666f7265",
    19065 => x"69676e20", 19066 => x"4d617374", 19067 => x"65722025",
    19068 => x"69206164", 19069 => x"6465640a", 19070 => x"00000000",
    19071 => x"4552524f", 19072 => x"523a2025", 19073 => x"733a2046",
    19074 => x"6f6c6c6f", 19075 => x"77207570", 19076 => x"206d6573",
    19077 => x"73616765", 19078 => x"20697320", 19079 => x"6e6f7420",
    19080 => x"66726f6d", 19081 => x"20637572", 19082 => x"72656e74",
    19083 => x"20706172", 19084 => x"656e740a", 19085 => x"00000000",
    19086 => x"4552524f", 19087 => x"523a2025", 19088 => x"733a2053",
    19089 => x"6c617665", 19090 => x"20776173", 19091 => x"206e6f74",
    19092 => x"20776169", 19093 => x"74696e67", 19094 => x"20612066",
    19095 => x"6f6c6c6f", 19096 => x"77207570", 19097 => x"206d6573",
    19098 => x"73616765", 19099 => x"0a000000", 19100 => x"4552524f",
    19101 => x"523a2025", 19102 => x"733a2053", 19103 => x"65717565",
    19104 => x"6e636549", 19105 => x"44202564", 19106 => x"20646f65",
    19107 => x"736e2774", 19108 => x"206d6174", 19109 => x"6368206c",
    19110 => x"61737420", 19111 => x"53796e63", 19112 => x"206d6573",
    19113 => x"73616765", 19114 => x"2025640a", 19115 => x"00000000",
    19116 => x"416e6e6f", 19117 => x"756e6365", 19118 => x"206d6573",
    19119 => x"73616765", 19120 => x"2066726f", 19121 => x"6d20616e",
    19122 => x"6f746865", 19123 => x"7220666f", 19124 => x"72656967",
    19125 => x"6e206d61", 19126 => x"73746572", 19127 => x"0a000000",
    19128 => x"25733a25", 19129 => x"693a2045", 19130 => x"72726f72",
    19131 => x"20310a00", 19132 => x"25733a25", 19133 => x"693a2045",
    19134 => x"72726f72", 19135 => x"20320a00", 19136 => x"42657374",
    19137 => x"20666f72", 19138 => x"6569676e", 19139 => x"206d6173",
    19140 => x"74657220", 19141 => x"69732025", 19142 => x"692f2569",
    19143 => x"0a000000", 19144 => x"25733a20", 19145 => x"6572726f",
    19146 => x"720a0000", 19147 => x"25733a20", 19148 => x"70617373",
    19149 => x"6976650a", 19150 => x"00000000", 19151 => x"25733a20",
    19152 => x"6d617374", 19153 => x"65720a00", 19154 => x"4e657720",
    19155 => x"55544320", 19156 => x"6f666673", 19157 => x"65743a20",
    19158 => x"25690a00", 19159 => x"25733a20", 19160 => x"736c6176",
    19161 => x"650a0000", 19162 => x"73796e63", 19163 => x"00000000",
    19164 => x"64656c61", 19165 => x"795f7265", 19166 => x"71000000",
    19167 => x"7064656c", 19168 => x"61795f72", 19169 => x"65710000",
    19170 => x"7064656c", 19171 => x"61795f72", 19172 => x"65737000",
    19173 => x"64656c61", 19174 => x"795f7265", 19175 => x"73700000",
    19176 => x"7064656c", 19177 => x"61795f72", 19178 => x"6573705f",
    19179 => x"666f6c6c", 19180 => x"6f775f75", 19181 => x"70000000",
    19182 => x"616e6e6f", 19183 => x"756e6365", 19184 => x"00000000",
    19185 => x"7369676e", 19186 => x"616c696e", 19187 => x"67000000",
    19188 => x"6d616e61", 19189 => x"67656d65", 19190 => x"6e740000",
    19191 => x"4552524f", 19192 => x"523a2042", 19193 => x"55473a20",
    19194 => x"25732064", 19195 => x"6f65736e", 19196 => x"27742073",
    19197 => x"7570706f", 19198 => x"7274206e", 19199 => x"65676174",
    19200 => x"69766573", 19201 => x"0a000000", 19202 => x"4552524f",
    19203 => x"523a204e", 19204 => x"65676174", 19205 => x"69766520",
    19206 => x"76616c75", 19207 => x"65206361", 19208 => x"6e6e6f74",
    19209 => x"20626520", 19210 => x"636f6e76", 19211 => x"65727465",
    19212 => x"6420696e", 19213 => x"746f2074", 19214 => x"696d6573",
    19215 => x"74616d70", 19216 => x"0a000000", 19217 => x"4552524f",
    19218 => x"523a2074", 19219 => x"6f5f5469", 19220 => x"6d65496e",
    19221 => x"7465726e", 19222 => x"616c3a20", 19223 => x"7365636f",
    19224 => x"6e647320", 19225 => x"6669656c", 19226 => x"64206973",
    19227 => x"20686967", 19228 => x"68657220", 19229 => x"7468616e",
    19230 => x"20736967", 19231 => x"6e656420", 19232 => x"696e7465",
    19233 => x"67657220", 19234 => x"28333262", 19235 => x"69747329",
    19236 => x"0a000000", 19237 => x"2d000000", 19238 => x"25732564",
    19239 => x"2e253039", 19240 => x"64000000", 19241 => x"6572726f",
    19242 => x"7220696e", 19243 => x"20745f6f", 19244 => x"70732d3e",
    19245 => x"73657276", 19246 => x"6f5f696e", 19247 => x"69740000",
    19248 => x"496e6974", 19249 => x"69616c69", 19250 => x"7a65643a",
    19251 => x"206f6273", 19252 => x"5f647269", 19253 => x"66742025",
    19254 => x"6c6c690a", 19255 => x"00000000", 19256 => x"636f7272",
    19257 => x"65637469", 19258 => x"6f6e2066", 19259 => x"69656c64",
    19260 => x"20313a20", 19261 => x"25730a00", 19262 => x"64697363",
    19263 => x"61726420", 19264 => x"54332f54", 19265 => x"343a2077",
    19266 => x"65206d69", 19267 => x"73732054", 19268 => x"312f5432",
    19269 => x"0a000000", 19270 => x"636f7272", 19271 => x"65637469",
    19272 => x"6f6e2066", 19273 => x"69656c64", 19274 => x"20323a20",
    19275 => x"25730a00", 19276 => x"54313a20", 19277 => x"25730a00",
    19278 => x"54323a20", 19279 => x"25730a00", 19280 => x"54333a20",
    19281 => x"25730a00", 19282 => x"54343a20", 19283 => x"25730a00",
    19284 => x"4d617374", 19285 => x"65722074", 19286 => x"6f20736c",
    19287 => x"6176653a", 19288 => x"2025730a", 19289 => x"00000000",
    19290 => x"536c6176", 19291 => x"6520746f", 19292 => x"206d6173",
    19293 => x"7465723a", 19294 => x"2025730a", 19295 => x"00000000",
    19296 => x"6d65616e", 19297 => x"50617468", 19298 => x"44656c61",
    19299 => x"793a2025", 19300 => x"730a0000", 19301 => x"73657276",
    19302 => x"6f206162", 19303 => x"6f727465", 19304 => x"642c2064",
    19305 => x"656c6179", 19306 => x"20677265", 19307 => x"61746572",
    19308 => x"20746861", 19309 => x"6e203120", 19310 => x"7365636f",
    19311 => x"6e640a00", 19312 => x"73657276", 19313 => x"6f206162",
    19314 => x"6f727465", 19315 => x"642c2064", 19316 => x"656c6179",
    19317 => x"20256420", 19318 => x"6f722025", 19319 => x"64206772",
    19320 => x"65617465", 19321 => x"72207468", 19322 => x"616e2063",
    19323 => x"6f6e6669", 19324 => x"67757265", 19325 => x"64206d61",
    19326 => x"78696d75", 19327 => x"6d202564", 19328 => x"0a000000",
    19329 => x"5472696d", 19330 => x"20746f6f", 19331 => x"2d6c6f6e",
    19332 => x"67206d70", 19333 => x"643a2025", 19334 => x"690a0000",
    19335 => x"41667465", 19336 => x"72206176", 19337 => x"67282569",
    19338 => x"292c206d", 19339 => x"65616e50", 19340 => x"61746844",
    19341 => x"656c6179", 19342 => x"3a202569", 19343 => x"0a000000",
    19344 => x"4f666673", 19345 => x"65742066", 19346 => x"726f6d20",
    19347 => x"6d617374", 19348 => x"65723a20", 19349 => x"20202020",
    19350 => x"25730a00", 19351 => x"73657276", 19352 => x"6f206162",
    19353 => x"6f727465", 19354 => x"642c206f", 19355 => x"66667365",
    19356 => x"74206772", 19357 => x"65617465", 19358 => x"72207468",
    19359 => x"616e2031", 19360 => x"20736563", 19361 => x"6f6e640a",
    19362 => x"00000000", 19363 => x"73657276", 19364 => x"6f206162",
    19365 => x"6f727465", 19366 => x"642c206f", 19367 => x"66667365",
    19368 => x"74206772", 19369 => x"65617465", 19370 => x"72207468",
    19371 => x"616e2063", 19372 => x"6f6e6669", 19373 => x"67757265",
    19374 => x"64206d61", 19375 => x"78696d75", 19376 => x"6d202564",
    19377 => x"0a000000", 19378 => x"4f627365", 19379 => x"72766564",
    19380 => x"20647269", 19381 => x"66743a20", 19382 => x"2539690a",
    19383 => x"00000000", 19384 => x"74696d65", 19385 => x"6f757420",
    19386 => x"65787069", 19387 => x"7265643a", 19388 => x"2025730a",
    19389 => x"00000000", 19390 => x"50505f54", 19391 => x"4f5f4445",
    19392 => x"4c415952", 19393 => x"45510000", 19394 => x"50505f54",
    19395 => x"4f5f5359", 19396 => x"4e430000", 19397 => x"50505f54",
    19398 => x"4f5f414e", 19399 => x"4e5f5245", 19400 => x"43454950",
    19401 => x"54000000", 19402 => x"50505f54", 19403 => x"4f5f414e",
    19404 => x"4e5f494e", 19405 => x"54455256", 19406 => x"414c0000",
    19407 => x"50505f54", 19408 => x"4f5f4641", 19409 => x"554c5459",
    19410 => x"00000000", 19411 => x"50505f54", 19412 => x"4f5f4558",
    19413 => x"545f3000", 19414 => x"50505f54", 19415 => x"4f5f4558",
    19416 => x"545f3100", 19417 => x"50505f54", 19418 => x"4f5f4558",
    19419 => x"545f3200", 19420 => x"536c6176", 19421 => x"65204f6e",
    19422 => x"6c792c20", 19423 => x"636c6f63", 19424 => x"6b20636c",
    19425 => x"61737320", 19426 => x"73657420", 19427 => x"746f2032",
    19428 => x"35350a00", 19429 => x"1b5b3125", 19430 => x"63000000",
    19431 => x"436f6d6d", 19432 => x"616e6420", 19433 => x"22257322",
    19434 => x"3a206572", 19435 => x"726f7220", 19436 => x"25640a00",
    19437 => x"556e7265", 19438 => x"636f676e", 19439 => x"697a6564",
    19440 => x"20636f6d", 19441 => x"6d616e64", 19442 => x"20222573",
    19443 => x"222e0a00", 19444 => x"77726323", 19445 => x"20000000",
    19446 => x"25630000", 19447 => x"456d7074", 19448 => x"7920696e",
    19449 => x"69742073", 19450 => x"63726970", 19451 => x"742e2e2e",
    19452 => x"0a000000", 19453 => x"65786563", 19454 => x"7574696e",
    19455 => x"673a2025", 19456 => x"730a0000", 19457 => x"57522043",
    19458 => x"6f726520", 19459 => x"6275696c", 19460 => x"643a2025",
    19461 => x"7325730a", 19462 => x"00000000", 19463 => x"2028756e",
    19464 => x"73757070", 19465 => x"6f727465", 19466 => x"64206465",
    19467 => x"76656c6f", 19468 => x"70657220", 19469 => x"6275696c",
    19470 => x"64290000", 19471 => x"4275696c", 19472 => x"743a2025",
    19473 => x"73202573", 19474 => x"0a000000", 19475 => x"4275696c",
    19476 => x"7420666f", 19477 => x"72202564", 19478 => x"206b4220",
    19479 => x"52414d2c", 19480 => x"20737461", 19481 => x"636b2069",
    19482 => x"73202564", 19483 => x"20627974", 19484 => x"65730a00",
    19485 => x"5741524e", 19486 => x"494e473a", 19487 => x"20686172",
    19488 => x"64776172", 19489 => x"65207361", 19490 => x"79732025",
    19491 => x"696b4220", 19492 => x"3c3d2052", 19493 => x"414d203c",
    19494 => x"2025696b", 19495 => x"420a0000", 19496 => x"76657200",
    19497 => x"696e6974", 19498 => x"00000000", 19499 => x"636c0000",
    19500 => x"73746174", 19501 => x"00000000", 19502 => x"73707300",
    19503 => x"67707300", 19504 => x"25642025", 19505 => x"640a0000",
    19506 => x"73746172", 19507 => x"74000000", 19508 => x"73746f70",
    19509 => x"00000000", 19510 => x"73646163", 19511 => x"00000000",
    19512 => x"67646163", 19513 => x"00000000", 19514 => x"63686563",
    19515 => x"6b76636f", 19516 => x"00000000", 19517 => x"706c6c00",
    19518 => x"64657465", 19519 => x"63740000", 19520 => x"4e6f2053",
    19521 => x"46502e0a", 19522 => x"00000000", 19523 => x"65726173",
    19524 => x"65000000", 19525 => x"436f756c", 19526 => x"64206e6f",
    19527 => x"74206572", 19528 => x"61736520", 19529 => x"44420a00",
    19530 => x"61646400", 19531 => x"53465020", 19532 => x"44422069",
    19533 => x"73206675", 19534 => x"6c6c0a00", 19535 => x"49324320",
    19536 => x"6572726f", 19537 => x"720a0000", 19538 => x"25642053",
    19539 => x"46507320", 19540 => x"696e2044", 19541 => x"420a0000",
    19542 => x"73686f77", 19543 => x"00000000", 19544 => x"53465020",
    19545 => x"64617461", 19546 => x"62617365", 19547 => x"20656d70",
    19548 => x"74792e2e", 19549 => x"2e0a0000", 19550 => x"53465020",
    19551 => x"64617461", 19552 => x"62617365", 19553 => x"20636f72",
    19554 => x"72757074", 19555 => x"65642e2e", 19556 => x"2e0a0000",
    19557 => x"25643a20", 19558 => x"504e3a00", 19559 => x"20645478",
    19560 => x"3a202564", 19561 => x"2c206452", 19562 => x"783a2025",
    19563 => x"642c2061", 19564 => x"6c706861", 19565 => x"3a202564",
    19566 => x"0a000000", 19567 => x"6d617463", 19568 => x"68000000",
    19569 => x"52756e20", 19570 => x"73667020", 19571 => x"64657465",
    19572 => x"63742066", 19573 => x"69727374", 19574 => x"0a000000",
    19575 => x"53465020", 19576 => x"6d617463", 19577 => x"6865642c",
    19578 => x"20645478", 19579 => x"3d25642c", 19580 => x"20645278",
    19581 => x"3d25642c", 19582 => x"20616c70", 19583 => x"68613d25",
    19584 => x"640a0000", 19585 => x"436f756c", 19586 => x"64206e6f",
    19587 => x"74206d61", 19588 => x"74636820", 19589 => x"746f2044",
    19590 => x"420a0000", 19591 => x"656e6100", 19592 => x"73667000",
    19593 => x"73746174", 19594 => x"69737469", 19595 => x"6373206e",
    19596 => x"6f77206f", 19597 => x"66660a00", 19598 => x"62747300",
    19599 => x"6f666600", 19600 => x"70747000", 19601 => x"676d0000",
    19602 => x"6d6f6465", 19603 => x"00000000", 19604 => x"6772616e",
    19605 => x"646d6173", 19606 => x"74657200", 19607 => x"666f7263",
    19608 => x"65000000", 19609 => x"466f756e", 19610 => x"64207068",
    19611 => x"61736520", 19612 => x"7472616e", 19613 => x"73697469",
    19614 => x"6f6e2069", 19615 => x"6e204545", 19616 => x"50524f4d",
    19617 => x"3a202564", 19618 => x"70730a00", 19619 => x"4d656173",
    19620 => x"7572696e", 19621 => x"67207432", 19622 => x"2f743420",
    19623 => x"70686173", 19624 => x"65207472", 19625 => x"616e7369",
    19626 => x"74696f6e", 19627 => x"2e2e2e0a", 19628 => x"00000000",
    19629 => x"63616c69", 19630 => x"62726174", 19631 => x"696f6e00",
    19632 => x"73657400", 19633 => x"73657473", 19634 => x"65630000",
    19635 => x"7365746e", 19636 => x"73656300", 19637 => x"72617700",
    19638 => x"2573202b", 19639 => x"2564206e", 19640 => x"616e6f73",
    19641 => x"65636f6e", 19642 => x"64732e0a", 19643 => x"00000000",
    19644 => x"74696d65", 19645 => x"00000000", 19646 => x"67756900",
    19647 => x"73646200", 19648 => x"67657400", 19649 => x"67657470",
    19650 => x"00000000", 19651 => x"73657470", 19652 => x"00000000",
    19653 => x"4d41432d", 19654 => x"61646472", 19655 => x"6573733a",
    19656 => x"20253032", 19657 => x"783a2530", 19658 => x"32783a25",
    19659 => x"3032783a", 19660 => x"25303278", 19661 => x"3a253032",
    19662 => x"783a2530", 19663 => x"32780a00", 19664 => x"6d616300",
    19665 => x"45455052", 19666 => x"4f4d206e", 19667 => x"6f742066",
    19668 => x"6f756e64", 19669 => x"2e2e0a00", 19670 => x"436f756c",
    19671 => x"64206e6f", 19672 => x"74206572", 19673 => x"61736520",
    19674 => x"696e6974", 19675 => x"20736372", 19676 => x"6970740a",
    19677 => x"00000000", 19678 => x"436f756c", 19679 => x"64206e6f",
    19680 => x"74206164", 19681 => x"64207468", 19682 => x"6520636f",
    19683 => x"6d6d616e", 19684 => x"640a0000", 19685 => x"4f4b2e0a",
    19686 => x"00000000", 19687 => x"626f6f74", 19688 => x"00000000",
    19689 => x"4f4e0000", 19690 => x"4f464600", 19691 => x"656e6162",
    19692 => x"6c650000", 19693 => x"64697361", 19694 => x"626c6500",
    19695 => x"70686173", 19696 => x"65207472", 19697 => x"61636b69",
    19698 => x"6e672025", 19699 => x"730a0000", 19700 => x"70747261",
    19701 => x"636b0000", 19702 => x"41766169", 19703 => x"6c61626c",
    19704 => x"6520636f", 19705 => x"6d6d616e", 19706 => x"64733a0a",
    19707 => x"00000000", 19708 => x"20202573", 19709 => x"0a000000",
    19710 => x"68656c70", 19711 => x"00000000", 19712 => x"55736167",
    19713 => x"653a2072", 19714 => x"65667265", 19715 => x"7368203c",
    19716 => x"7365636f", 19717 => x"6e64733e", 19718 => x"0a000000",
    19719 => x"72656672", 19720 => x"65736800", 19721 => x"49502d61",
    19722 => x"64647265", 19723 => x"73733a20", 19724 => x"696e2074",
    19725 => x"7261696e", 19726 => x"696e670a", 19727 => x"00000000",
    19728 => x"49502d61", 19729 => x"64647265", 19730 => x"73733a20",
    19731 => x"25642e25", 19732 => x"642e2564", 19733 => x"2e25640a",
    19734 => x"00000000", 19735 => x"69700000", 19736 => x"50505349",
    19737 => x"20766572", 19738 => x"626f7369", 19739 => x"74793a20",
    19740 => x"2530386c", 19741 => x"780a0000", 19742 => x"76657262",
    19743 => x"6f736500", 19744 => x"25732c20", 19745 => x"25732025",
    19746 => x"642c2025", 19747 => x"642c2025", 19748 => x"3032643a",
    19749 => x"25303264", 19750 => x"3a253032", 19751 => x"64000000",
    19752 => x"1b5b3025", 19753 => x"643b3325", 19754 => x"646d0000",
    19755 => x"1b5b6d00", 19756 => x"1b5b2564", 19757 => x"3b256466",
    19758 => x"00000000", 19759 => x"1b5b324a", 19760 => x"1b5b313b",
    19761 => x"31480000", 19762 => x"53756e00", 19763 => x"4d6f6e00",
    19764 => x"54756500", 19765 => x"57656400", 19766 => x"54687500",
    19767 => x"46726900", 19768 => x"53617400", 19769 => x"4a616e00",
    19770 => x"46656200", 19771 => x"4d617200", 19772 => x"41707200",
    19773 => x"4d617900", 19774 => x"4a756e00", 19775 => x"4a756c00",
    19776 => x"41756700", 19777 => x"53657000", 19778 => x"4f637400",
    19779 => x"4e6f7600", 19780 => x"44656300", 19781 => x"4c6f6f70",
    19782 => x"73207065", 19783 => x"72206a69", 19784 => x"6666793a",
    19785 => x"2025690a", 19786 => x"00000000", 19787 => x"77723000",
    19788 => x"44697363", 19789 => x"6f766572", 19790 => x"65642049",
    19791 => x"50206164", 19792 => x"64726573", 19793 => x"73202825",
    19794 => x"642e2564", 19795 => x"2e25642e", 19796 => x"25642921",
    19797 => x"0a000000", 19798 => x"30313233", 19799 => x"34353637",
    19800 => x"38396162", 19801 => x"63646566", 19802 => x"00000000",
    19803 => x"49443a20", 19804 => x"25780a00", 19805 => x"7066696c",
    19806 => x"7465723a", 19807 => x"2077726f", 19808 => x"6e67206d",
    19809 => x"61676963", 19810 => x"206e756d", 19811 => x"62657220",
    19812 => x"28676f74", 19813 => x"20307825", 19814 => x"78290a00",
    19815 => x"7066696c", 19816 => x"7465723a", 19817 => x"2077726f",
    19818 => x"6e672072", 19819 => x"756c652d", 19820 => x"7365742c",
    19821 => x"2063616e", 19822 => x"27742061", 19823 => x"70706c79",
    19824 => x"0a000000", 19825 => x"696e7661", 19826 => x"6c696420",
    19827 => x"64657363", 19828 => x"72697074", 19829 => x"6f722040",
    19830 => x"2578203d", 19831 => x"2025780a", 19832 => x"00000000",
    19833 => x"5761726e", 19834 => x"696e673a", 19835 => x"20747820",
    19836 => x"6e6f7420", 19837 => x"7465726d", 19838 => x"696e6174",
    19839 => x"65642069", 19840 => x"6e66696e", 19841 => x"69746520",
    19842 => x"6d63723d", 19843 => x"30782578", 19844 => x"0a000000",
    19845 => x"5761726e", 19846 => x"696e673a", 19847 => x"20747820",
    19848 => x"74696d65", 19849 => x"7374616d", 19850 => x"70206e65",
    19851 => x"76657220", 19852 => x"62656361", 19853 => x"6d652061",
    19854 => x"7661696c", 19855 => x"61626c65", 19856 => x"0a000000",
    19857 => x"6d696e69", 19858 => x"635f7478", 19859 => x"5f667261",
    19860 => x"6d653a20", 19861 => x"756e6d61", 19862 => x"74636865",
    19863 => x"64206669", 19864 => x"64202564", 19865 => x"20767320",
    19866 => x"25640a00", 19867 => x"6e616e6f", 19868 => x"7365636f",
    19869 => x"6e647300", 19870 => x"41646a75", 19871 => x"73743a20",
    19872 => x"636f756e", 19873 => x"74657220", 19874 => x"3d202573",
    19875 => x"205b2563", 19876 => x"25645d0a", 19877 => x"00000000",
    19878 => x"64657620", 19879 => x"20307825", 19880 => x"30386c78",
    19881 => x"20402025", 19882 => x"30366c78", 19883 => x"2c202573",
    19884 => x"0a000000", 19885 => x"66706761", 19886 => x"2d617265",
    19887 => x"61000000", 19888 => x"4572726f", 19889 => x"72202564",
    19890 => x"20776869", 19891 => x"6c652072", 19892 => x"65616469",
    19893 => x"6e672074", 19894 => x"32347020", 19895 => x"66726f6d",
    19896 => x"2073746f", 19897 => x"72616765", 19898 => x"0a000000",
    19899 => x"74323470", 19900 => x"20726561", 19901 => x"64206672",
    19902 => x"6f6d2073", 19903 => x"746f7261", 19904 => x"67653a20",
    19905 => x"25642070", 19906 => x"730a0000", 19907 => x"52585453",
    19908 => x"2063616c", 19909 => x"69627261", 19910 => x"74696f6e",
    19911 => x"20657272", 19912 => x"6f722e0a", 19913 => x"00000000",
    19914 => x"52585453", 19915 => x"2063616c", 19916 => x"69627261",
    19917 => x"74696f6e", 19918 => x"3a205240", 19919 => x"25647073",
    19920 => x"2c204640", 19921 => x"25647073", 19922 => x"2c207472",
    19923 => x"616e7369", 19924 => x"74696f6e", 19925 => x"40256470",
    19926 => x"730a0000", 19927 => x"57616974", 19928 => x"696e6720",
    19929 => x"666f7220", 19930 => x"6c696e6b", 19931 => x"2e2e2e0a",
    19932 => x"00000000", 19933 => x"4c6f636b", 19934 => x"696e6720",
    19935 => x"504c4c2e", 19936 => x"2e2e0a00", 19937 => x"43616c69",
    19938 => x"62726174", 19939 => x"696e6720", 19940 => x"52582074",
    19941 => x"696d6573", 19942 => x"74616d70", 19943 => x"65722e2e",
    19944 => x"2e0a0000", 19945 => x"4661696c", 19946 => x"65640000",
    19947 => x"53756363", 19948 => x"65737300", 19949 => x"57726f74",
    19950 => x"65206e65", 19951 => x"77207432", 19952 => x"34702076",
    19953 => x"616c7565", 19954 => x"3a202564", 19955 => x"20707320",
    19956 => x"28257329", 19957 => x"0a000000", 19958 => x"43616e27",
    19959 => x"74207361", 19960 => x"76652070", 19961 => x"65727369",
    19962 => x"7374656e", 19963 => x"74204d41", 19964 => x"43206164",
    19965 => x"64726573", 19966 => x"730a0000", 19967 => x"25733a20",
    19968 => x"5573696e", 19969 => x"67205731", 19970 => x"20736572",
    19971 => x"69616c20", 19972 => x"6e756d62", 19973 => x"65720a00",
    19974 => x"6f666673", 19975 => x"65742025", 19976 => x"34692028",
    19977 => x"30782530", 19978 => x"3378293a", 19979 => x"20253369",
    19980 => x"20283078", 19981 => x"25303278", 19982 => x"290a0000",
    19983 => x"77726974", 19984 => x"65283078", 19985 => x"25782c20",
    19986 => x"2569293a", 19987 => x"20726573", 19988 => x"756c7420",
    19989 => x"3d202569", 19990 => x"0a000000", 19991 => x"72656164",
    19992 => x"28307825", 19993 => x"782c2025", 19994 => x"69293a20",
    19995 => x"72657375", 19996 => x"6c74203d", 19997 => x"2025690a",
    19998 => x"00000000", 19999 => x"64657669", 20000 => x"63652025",
    20001 => x"693a2025", 20002 => x"30387825", 20003 => x"3038780a",
    20004 => x"00000000", 20005 => x"74656d70", 20006 => x"3a202564",
    20007 => x"2e253034", 20008 => x"640a0000", 20009 => x"77310000",
    20010 => x"77317200", 20011 => x"77317700", 20012 => x"456e6162",
    20013 => x"6c655461", 20014 => x"67676572", 20015 => x"20256420",
    20016 => x"25640a00", 20017 => x"25733a20", 20018 => x"63682025",
    20019 => x"642c204f", 20020 => x"43455220", 20021 => x"30782578",
    20022 => x"2c205243", 20023 => x"45522030", 20024 => x"7825780a",
    20025 => x"00000000", 20026 => x"3c756e6b", 20027 => x"6e6f776e",
    20028 => x"3e000000", 20029 => x"4558543a", 20030 => x"20444d54",
    20031 => x"44206c6f", 20032 => x"636b6564", 20033 => x"2e0a0000",
    20034 => x"4558543a", 20035 => x"20435379", 20036 => x"6e632063",
    20037 => x"6f6d706c", 20038 => x"6574652e", 20039 => x"0a000000",
    20040 => x"4558543a", 20041 => x"20416c69", 20042 => x"676e2074",
    20043 => x"61726765", 20044 => x"74202564", 20045 => x"2c207374",
    20046 => x"65702025", 20047 => x"642e0a00", 20048 => x"4558543a",
    20049 => x"20416c69", 20050 => x"676e2064", 20051 => x"6f6e652e",
    20052 => x"0a000000", 20053 => x"72656620", 20054 => x"2564206f",
    20055 => x"75742025", 20056 => x"64206964", 20057 => x"78202578",
    20058 => x"200a0000", 20059 => x"4d504c4c", 20060 => x"5f537461",
    20061 => x"7274205b", 20062 => x"64616320", 20063 => x"25645d0a",
    20064 => x"00000000", 20065 => x"736f6674", 20066 => x"706c6c3a",
    20067 => x"20617474", 20068 => x"656d7074", 20069 => x"696e6720",
    20070 => x"746f2065", 20071 => x"6e61626c", 20072 => x"6520474d",
    20073 => x"206d6f64", 20074 => x"65206f6e", 20075 => x"206e6f6e",
    20076 => x"2d474d20", 20077 => x"68617264", 20078 => x"77617265",
    20079 => x"2e0a0000", 20080 => x"736f6674", 20081 => x"706c6c3a",
    20082 => x"206d6f64", 20083 => x"65202573", 20084 => x"2c202564",
    20085 => x"20726566", 20086 => x"20636861", 20087 => x"6e6e656c",
    20088 => x"732c2025", 20089 => x"64206f75", 20090 => x"74206368",
    20091 => x"616e6e65", 20092 => x"6c730a00", 20093 => x"43616e27",
    20094 => x"74207374", 20095 => x"61727420", 20096 => x"6368616e",
    20097 => x"6e656c20", 20098 => x"25642c20", 20099 => x"74686520",
    20100 => x"504c4c20", 20101 => x"6973206e", 20102 => x"6f742072",
    20103 => x"65616479", 20104 => x"0a000000", 20105 => x"736f6674",
    20106 => x"706c6c3a", 20107 => x"20697271", 20108 => x"73202564",
    20109 => x"20736571", 20110 => x"20257320", 20111 => x"6d6f6465",
    20112 => x"20256420", 20113 => x"616c6967", 20114 => x"6e6d656e",
    20115 => x"745f7374", 20116 => x"61746520", 20117 => x"25642048",
    20118 => x"4c256420", 20119 => x"4d4c2564", 20120 => x"2048593d",
    20121 => x"2564204d", 20122 => x"593d2564", 20123 => x"2044656c",
    20124 => x"436e743d", 20125 => x"25640a00", 20126 => x"456e6162",
    20127 => x"6c696e67", 20128 => x"20707472", 20129 => x"61636b65",
    20130 => x"72206368", 20131 => x"616e6e65", 20132 => x"6c3a2025",
    20133 => x"640a0000", 20134 => x"44697361", 20135 => x"626c696e",
    20136 => x"67207074", 20137 => x"7261636b", 20138 => x"65722074",
    20139 => x"61676765", 20140 => x"723a2025", 20141 => x"640a0000",
    20142 => x"6c6f636b", 20143 => x"696e6700", 20144 => x"616c6967",
    20145 => x"6e696e67", 20146 => x"00000000", 20147 => x"736f6674",
    20148 => x"706c6c3a", 20149 => x"20646973", 20150 => x"61626c65",
    20151 => x"64206175", 20152 => x"78206368", 20153 => x"616e6e65",
    20154 => x"6c202564", 20155 => x"0a000000", 20156 => x"736f6674",
    20157 => x"706c6c3a", 20158 => x"20656e61", 20159 => x"626c6564",
    20160 => x"20617578", 20161 => x"20636861", 20162 => x"6e6e656c",
    20163 => x"2025640a", 20164 => x"00000000", 20165 => x"736f6674",
    20166 => x"706c6c3a", 20167 => x"20636861", 20168 => x"6e6e656c",
    20169 => x"20256420", 20170 => x"6c6f636b", 20171 => x"6564205b",
    20172 => x"616c6967", 20173 => x"6e696e67", 20174 => x"20402025",
    20175 => x"64207073", 20176 => x"5d0a0000", 20177 => x"736f6674",
    20178 => x"706c6c3a", 20179 => x"20636861", 20180 => x"6e6e656c",
    20181 => x"20256420", 20182 => x"70686173", 20183 => x"6520616c",
    20184 => x"69676e65", 20185 => x"640a0000", 20186 => x"736f6674",
    20187 => x"706c6c3a", 20188 => x"20617578", 20189 => x"20636861",
    20190 => x"6e6e656c", 20191 => x"20256420", 20192 => x"6f72206d",
    20193 => x"706c6c20", 20194 => x"6c6f7374", 20195 => x"206c6f63",
    20196 => x"6b0a0000", 20197 => x"536f6674", 20198 => x"504c4c20",
    20199 => x"56434f20", 20200 => x"46726571", 20201 => x"75656e63",
    20202 => x"792f4150", 20203 => x"52207465", 20204 => x"73743a0a",
    20205 => x"00000000", 20206 => x"444d5444", 20207 => x"2056434f",
    20208 => x"3a20204c", 20209 => x"6f773d25", 20210 => x"6420487a",
    20211 => x"2048693d", 20212 => x"25642048", 20213 => x"7a2c2041",
    20214 => x"5052203d", 20215 => x"20256420", 20216 => x"70706d2e",
    20217 => x"0a000000", 20218 => x"52454620", 20219 => x"56434f3a",
    20220 => x"2020204c", 20221 => x"6f773d25", 20222 => x"6420487a",
    20223 => x"2048693d", 20224 => x"25642048", 20225 => x"7a2c2041",
    20226 => x"5052203d", 20227 => x"20256420", 20228 => x"70706d2e",
    20229 => x"0a000000", 20230 => x"45585420", 20231 => x"636c6f63",
    20232 => x"6b3a2046", 20233 => x"7265713d", 20234 => x"25642048",
    20235 => x"7a0a0000", 20236 => x"73746172", 20237 => x"742d6578",
    20238 => x"74000000", 20239 => x"77616974", 20240 => x"2d657874",
    20241 => x"00000000", 20242 => x"73746172", 20243 => x"742d6865",
    20244 => x"6c706572", 20245 => x"00000000", 20246 => x"77616974",
    20247 => x"2d68656c", 20248 => x"70657200", 20249 => x"73746172",
    20250 => x"742d6d61", 20251 => x"696e0000", 20252 => x"77616974",
    20253 => x"2d6d6169", 20254 => x"6e000000", 20255 => x"72656164",
    20256 => x"79000000", 20257 => x"636c6561", 20258 => x"722d6461",
    20259 => x"63730000", 20260 => x"77616974", 20261 => x"2d636c65",
    20262 => x"61722d64", 20263 => x"61637300", 20264 => x"66726565",
    20265 => x"6d617374", 20266 => x"65720000", 20267 => x"53746163",
    20268 => x"6b206f76", 20269 => x"6572666c", 20270 => x"6f77210a",
    20271 => x"00000000", 20272 => x"badc0ffe", 20273 => x"3b9ac9ff",
    20274 => x"3b9aca00", 20275 => x"000f4240", 20276 => x"00080030",
    20277 => x"d4a51000", 20278 => x"c4653600", 20279 => x"7ffffffe",
    20280 => x"80000001", 20281 => x"fff06000", 20282 => x"0007d000",
    20283 => x"41c64e6d", 20284 => x"00010043", 20285 => x"00010044",
    20286 => x"00015180", 20287 => x"000186a0", 20288 => x"00062000",
    20289 => x"005ee000", 20290 => x"01000001", 20291 => x"11223344",
    20292 => x"e0001fff", 20293 => x"0fffffff", 20294 => x"059682f0",
    20295 => x"0ee6b27f", 20296 => x"7fffffff", 20297 => x"01312d02",
    20298 => x"01312d0a", 20299 => x"c0a80001", 20300 => x"96aa9e04",
    20301 => x"003d0137", 20302 => x"8000001f", 20303 => x"009895b6",
    20304 => x"c4000001", 20305 => x"00ffffff", 20306 => x"fffdb610",
    20307 => x"000249f0", 20308 => x"05f5e100", 20309 => x"0bebc200",
    20310 => x"fa0a1f00", 20311 => x"fff0bdc0", 20312 => x"01312d03",
    20313 => x"03b9aca0", 20314 => x"07735940", 20315 => x"5344422d",
    20316 => x"011b1900", 20317 => x"00000000", 20318 => x"70705f64",
    20319 => x"6961675f", 20320 => x"70617273", 20321 => x"65000000",
    20322 => x"00000000", 20323 => x"00011e5c", 20324 => x"00011e68",
    20325 => x"00011e78", 20326 => x"00011e84", 20327 => x"00011e90",
    20328 => x"00011e9c", 20329 => x"00011ea8", 20330 => x"00002088",
    20331 => x"000020f8", 20332 => x"000023b0", 20333 => x"000023b0",
    20334 => x"000023b0", 20335 => x"000023b0", 20336 => x"000023b0",
    20337 => x"000023b0", 20338 => x"00002174", 20339 => x"000021e4",
    20340 => x"000023b0", 20341 => x"00002278", 20342 => x"00002384",
    20343 => x"77727063", 20344 => x"5f74696d", 20345 => x"655f6164",
    20346 => x"6a757374", 20347 => x"5f6f6666", 20348 => x"73657400",
    20349 => x"77727063", 20350 => x"5f74696d", 20351 => x"655f6164",
    20352 => x"6a757374", 20353 => x"00000000", 20354 => x"77727063",
    20355 => x"5f74696d", 20356 => x"655f7365", 20357 => x"74000000",
    20358 => x"77727063", 20359 => x"5f74696d", 20360 => x"655f6765",
    20361 => x"74000000", 20362 => x"77727063", 20363 => x"5f6e6574",
    20364 => x"5f73656e", 20365 => x"64000000", 20366 => x"77725f75",
    20367 => x"6e706163", 20368 => x"6b5f616e", 20369 => x"6e6f756e",
    20370 => x"63650000", 20371 => x"77725f70", 20372 => x"61636b5f",
    20373 => x"616e6e6f", 20374 => x"756e6365", 20375 => x"00000000",
    20376 => x"77725f68", 20377 => x"616e646c", 20378 => x"655f666f",
    20379 => x"6c6c6f77", 20380 => x"75700000", 20381 => x"77725f68",
    20382 => x"616e646c", 20383 => x"655f616e", 20384 => x"6e6f756e",
    20385 => x"63650000", 20386 => x"77725f65", 20387 => x"78656375",
    20388 => x"74655f73", 20389 => x"6c617665", 20390 => x"00000000",
    20391 => x"77725f73", 20392 => x"31000000", 20393 => x"77725f68",
    20394 => x"616e646c", 20395 => x"655f7265", 20396 => x"73700000",
    20397 => x"77725f6e", 20398 => x"65775f73", 20399 => x"6c617665",
    20400 => x"00000000", 20401 => x"77725f6d", 20402 => x"61737465",
    20403 => x"725f6d73", 20404 => x"67000000", 20405 => x"77725f6c",
    20406 => x"69737465", 20407 => x"6e696e67", 20408 => x"00000000",
    20409 => x"77725f6f", 20410 => x"70656e00", 20411 => x"77725f69",
    20412 => x"6e697400", 20413 => x"00003980", 20414 => x"000039a8",
    20415 => x"000039c8", 20416 => x"00003a38", 20417 => x"00003a58",
    20418 => x"00003a74", 20419 => x"00003a94", 20420 => x"00003b20",
    20421 => x"00003b40", 20422 => x"77725f63", 20423 => x"616c6962",
    20424 => x"72617469", 20425 => x"6f6e0000", 20426 => x"00004f24",
    20427 => x"00004f0c", 20428 => x"00004f4c", 20429 => x"0000505c",
    20430 => x"00004fa0", 20431 => x"000127d8", 20432 => x"0001290c",
    20433 => x"00012918", 20434 => x"00012924", 20435 => x"00012930",
    20436 => x"0001293c", 20437 => x"77725f73", 20438 => x"6572766f",
    20439 => x"5f757064", 20440 => x"61746500", 20441 => x"70705f69",
    20442 => x"6e697469", 20443 => x"616c697a", 20444 => x"696e6700",
    20445 => x"73745f63", 20446 => x"6f6d5f73", 20447 => x"6c617665",
    20448 => x"5f68616e", 20449 => x"646c655f", 20450 => x"666f6c6c",
    20451 => x"6f777570", 20452 => x"00000000", 20453 => x"626d635f",
    20454 => x"64617461", 20455 => x"7365745f", 20456 => x"636d7000",
    20457 => x"626d635f", 20458 => x"73746174", 20459 => x"655f6465",
    20460 => x"63697369", 20461 => x"6f6e0000", 20462 => x"63466965",
    20463 => x"6c645f74", 20464 => x"6f5f5469", 20465 => x"6d65496e",
    20466 => x"7465726e", 20467 => x"616c0000", 20468 => x"00011d58",
    20469 => x"00013250", 20470 => x"00012954", 20471 => x"0001246c",
    20472 => x"0000001f", 20473 => x"0000001c", 20474 => x"0000001f",
    20475 => x"0000001e", 20476 => x"0000001f", 20477 => x"0000001e",
    20478 => x"0000001f", 20479 => x"0000001f", 20480 => x"0000001e",
    20481 => x"0000001f", 20482 => x"0000001e", 20483 => x"0000001f",
    20484 => x"0000001f", 20485 => x"0000001d", 20486 => x"0000001f",
    20487 => x"0000001e", 20488 => x"0000001f", 20489 => x"0000001e",
    20490 => x"0000001f", 20491 => x"0000001f", 20492 => x"0000001e",
    20493 => x"0000001f", 20494 => x"0000001e", 20495 => x"0000001f",
    20496 => x"000134c8", 20497 => x"000134cc", 20498 => x"000134d0",
    20499 => x"000134d4", 20500 => x"000134d8", 20501 => x"000134dc",
    20502 => x"000134e0", 20503 => x"000134e4", 20504 => x"000134e8",
    20505 => x"000134ec", 20506 => x"000134f0", 20507 => x"000134f4",
    20508 => x"000134f8", 20509 => x"000134fc", 20510 => x"00013500",
    20511 => x"00013504", 20512 => x"00013508", 20513 => x"0001350c",
    20514 => x"00013510", 20515 => x"6765745f", 20516 => x"70657273",
    20517 => x"69737465", 20518 => x"6e745f6d", 20519 => x"61630000",
    20520 => x"73706c6c", 20521 => x"5f656e61", 20522 => x"626c655f",
    20523 => x"74616767", 20524 => x"65720000", 20525 => x"0000ed30",
    20526 => x"0000edb8", 20527 => x"0000edec", 20528 => x"0000ee8c",
    20529 => x"0000ef10", 20530 => x"0000ef30", 20531 => x"0000ee18",
    20532 => x"0000ed54", 20533 => x"0000ecbc", 20534 => x"0000ecec",
    20535 => x"00000000", 20536 => x"00000000", 20537 => x"00000000",
    20538 => x"00000000", 20539 => x"00000001", 20540 => x"00000001",
    20541 => x"00000001", 20542 => x"00000001", 20543 => x"00000000",
    20544 => x"00000000", 20545 => x"00000000", 20546 => x"0000ece8",
    20547 => x"0000ece8", 20548 => x"00000000", 20549 => x"0000d9d0",
    20550 => x"00000000", 20551 => x"0000fb88", 20552 => x"0000fba8",
    20553 => x"0000fbb4", 20554 => x"0000fbc4", 20555 => x"0000fbe4",
    20556 => x"0000fbf4", 20557 => x"0000fc48", 20558 => x"0000fc0c",
    20559 => x"0000fb1c", 20560 => x"0000fb60", 20561 => x"00000001",
    20562 => x"00013c30", 20563 => x"00000002", 20564 => x"00013c3c",
    20565 => x"00000003", 20566 => x"00013c48", 20567 => x"00000004",
    20568 => x"00013c58", 20569 => x"00000005", 20570 => x"00013c64",
    20571 => x"00000006", 20572 => x"00013c70", 20573 => x"00000007",
    20574 => x"00012444", 20575 => x"00000008", 20576 => x"00013c7c",
    20577 => x"00000009", 20578 => x"00013c84", 20579 => x"0000000a",
    20580 => x"00013c90", 20581 => x"00000000", 20582 => x"00000000",
    20583 => x"00013cbc", 20584 => x"00013250", 20585 => x"00013ca0",
    20586 => x"0001246c", 20587 => x"00012444", 20588 => x"00000000",
    20589 => x"00000000", 20590 => x"00000000", 20591 => x"00000000",
    20592 => x"00010000", 20593 => x"00000000", 20594 => x"00000000",
    20595 => x"00000000", 20596 => x"00020100", 20597 => x"00000000",
    20598 => x"00000000", 20599 => x"00000000", 20600 => x"00030101",
    20601 => x"00000000", 20602 => x"00000000", 20603 => x"00000000",
    20604 => x"00040201", 20605 => x"01000000", 20606 => x"00000000",
    20607 => x"00000000", 20608 => x"00050201", 20609 => x"01010000",
    20610 => x"00000000", 20611 => x"00000000", 20612 => x"00060302",
    20613 => x"01010100", 20614 => x"00000000", 20615 => x"00000000",
    20616 => x"00070302", 20617 => x"01010101", 20618 => x"00000000",
    20619 => x"00000000", 20620 => x"00080402", 20621 => x"02010101",
    20622 => x"01000000", 20623 => x"00000000", 20624 => x"00090403",
    20625 => x"02010101", 20626 => x"01010000", 20627 => x"00000000",
    20628 => x"000a0503", 20629 => x"02020101", 20630 => x"01010100",
    20631 => x"00000000", 20632 => x"000b0503", 20633 => x"02020101",
    20634 => x"01010101", 20635 => x"00000000", 20636 => x"000c0604",
    20637 => x"03020201", 20638 => x"01010101", 20639 => x"01000000",
    20640 => x"000d0604", 20641 => x"03020201", 20642 => x"01010101",
    20643 => x"01010000", 20644 => x"000e0704", 20645 => x"03020202",
    20646 => x"01010101", 20647 => x"01010100", 20648 => x"000f0705",
    20649 => x"03030202", 20650 => x"01010101", 20651 => x"01010101",
    20652 => x"fefefeff", 20653 => x"80808080", 20654 => x"00202020",
    20655 => x"20202020", 20656 => x"20202828", 20657 => x"28282820",
    20658 => x"20202020", 20659 => x"20202020", 20660 => x"20202020",
    20661 => x"20202020", 20662 => x"20881010", 20663 => x"10101010",
    20664 => x"10101010", 20665 => x"10101010", 20666 => x"10040404",
    20667 => x"04040404", 20668 => x"04040410", 20669 => x"10101010",
    20670 => x"10104141", 20671 => x"41414141", 20672 => x"01010101",
    20673 => x"01010101", 20674 => x"01010101", 20675 => x"01010101",
    20676 => x"01010101", 20677 => x"10101010", 20678 => x"10104242",
    20679 => x"42424242", 20680 => x"02020202", 20681 => x"02020202",
    20682 => x"02020202", 20683 => x"02020202", 20684 => x"02020202",
    20685 => x"10101010", 20686 => x"20000000", 20687 => x"00000000",
    20688 => x"00000000", 20689 => x"00000000", 20690 => x"00000000",
    20691 => x"00000000", 20692 => x"00000000", 20693 => x"00000000",
    20694 => x"00000000", 20695 => x"00000000", 20696 => x"00000000",
    20697 => x"00000000", 20698 => x"00000000", 20699 => x"00000000",
    20700 => x"00000000", 20701 => x"00000000", 20702 => x"00000000",
    20703 => x"00000000", 20704 => x"00000000", 20705 => x"00000000",
    20706 => x"00000000", 20707 => x"00000000", 20708 => x"00000000",
    20709 => x"00000000", 20710 => x"00000000", 20711 => x"00000000",
    20712 => x"00000000", 20713 => x"00000000", 20714 => x"00000000",
    20715 => x"00000000", 20716 => x"00000000", 20717 => x"00000000",
    20718 => x"00000000", 20719 => x"00000000", 20720 => x"00014d88",
    20721 => x"00014da8", 20722 => x"00014db8", 20723 => x"000003e8",
    20724 => x"00000001", 20725 => x"046362a0", 20726 => x"00000955",
    20727 => x"ffffffff", 20728 => x"000143e4", 20729 => x"00000000",
    20730 => x"00000000", 20731 => x"00000000", 20732 => x"00000000",
    20733 => x"00000000", 20734 => x"00000000", 20735 => x"00000000",
    20736 => x"00000000", 20737 => x"00014758", 20738 => x"00014878",
    20739 => x"0001485c", 20740 => x"00014f34", 20741 => x"00014fb4",
    20742 => x"00000000", 20743 => x"00000000", 20744 => x"00000000",
    20745 => x"00000000", 20746 => x"00000000", 20747 => x"00000000",
    20748 => x"00000000", 20749 => x"00000000", 20750 => x"00000000",
    20751 => x"00000000", 20752 => x"00000000", 20753 => x"00000000",
    20754 => x"00000000", 20755 => x"00000000", 20756 => x"00000000",
    20757 => x"00000000", 20758 => x"00000000", 20759 => x"00000000",
    20760 => x"00000000", 20761 => x"00000000", 20762 => x"00000000",
    20763 => x"00000000", 20764 => x"00000000", 20765 => x"00000000",
    20766 => x"00000000", 20767 => x"00000000", 20768 => x"00000000",
    20769 => x"00000000", 20770 => x"00000000", 20771 => x"00000000",
    20772 => x"00000000", 20773 => x"00000000", 20774 => x"00000000",
    20775 => x"00000000", 20776 => x"00000000", 20777 => x"00000000",
    20778 => x"00000000", 20779 => x"00000000", 20780 => x"00000000",
    20781 => x"00000000", 20782 => x"00000000", 20783 => x"00000000",
    20784 => x"00000000", 20785 => x"00000000", 20786 => x"00000000",
    20787 => x"00000000", 20788 => x"00000000", 20789 => x"00000000",
    20790 => x"00000000", 20791 => x"00000000", 20792 => x"00000000",
    20793 => x"00000000", 20794 => x"00000000", 20795 => x"00000000",
    20796 => x"00000000", 20797 => x"00000000", 20798 => x"00000000",
    20799 => x"00000000", 20800 => x"00000000", 20801 => x"00000000",
    20802 => x"00000000", 20803 => x"00000000", 20804 => x"00000000",
    20805 => x"00000000", 20806 => x"00000000", 20807 => x"00000000",
    20808 => x"00000000", 20809 => x"00000000", 20810 => x"00000000",
    20811 => x"00000000", 20812 => x"00000000", 20813 => x"00000000",
    20814 => x"00000000", 20815 => x"00000000", 20816 => x"00000000",
    20817 => x"00000000", 20818 => x"00000000", 20819 => x"00000000",
    20820 => x"00000000", 20821 => x"00000000", 20822 => x"00000000",
    20823 => x"00000000", 20824 => x"00000000", 20825 => x"00000000",
    20826 => x"00000000", 20827 => x"00000000", 20828 => x"00000000",
    20829 => x"00000000", 20830 => x"00000000", 20831 => x"00000000",
    20832 => x"00000000", 20833 => x"00000000", 20834 => x"00000000",
    20835 => x"00000000", 20836 => x"00000000", 20837 => x"00000000",
    20838 => x"00000000", 20839 => x"00000000", 20840 => x"00000000",
    20841 => x"00000000", 20842 => x"00000000", 20843 => x"00000000",
    20844 => x"00000000", 20845 => x"00000000", 20846 => x"00000000",
    20847 => x"00000000", 20848 => x"00000000", 20849 => x"00000000",
    20850 => x"00000000", 20851 => x"00000000", 20852 => x"00000000",
    20853 => x"00000000", 20854 => x"00000000", 20855 => x"00000000",
    20856 => x"00000000", 20857 => x"00000000", 20858 => x"00000000",
    20859 => x"00000000", 20860 => x"00000000", 20861 => x"00000000",
    20862 => x"00000000", 20863 => x"00000000", 20864 => x"00000000",
    20865 => x"00000000", 20866 => x"00000000", 20867 => x"00000000",
    20868 => x"00000000", 20869 => x"00000000", 20870 => x"00000000",
    20871 => x"00000000", 20872 => x"00000000", 20873 => x"00000000",
    20874 => x"00000000", 20875 => x"00000000", 20876 => x"00000000",
    20877 => x"00000000", 20878 => x"00000000", 20879 => x"00000000",
    20880 => x"00000000", 20881 => x"00000000", 20882 => x"00000000",
    20883 => x"00000000", 20884 => x"00000000", 20885 => x"00000000",
    20886 => x"00000000", 20887 => x"00000000", 20888 => x"00000000",
    20889 => x"00000000", 20890 => x"00000000", 20891 => x"00000000",
    20892 => x"00000000", 20893 => x"00000000", 20894 => x"00000000",
    20895 => x"00000000", 20896 => x"00000000", 20897 => x"00000000",
    20898 => x"00000000", 20899 => x"00000000", 20900 => x"00000000",
    20901 => x"00000000", 20902 => x"00000000", 20903 => x"00000000",
    20904 => x"00000000", 20905 => x"00000000", 20906 => x"00000000",
    20907 => x"000147a0", 20908 => x"00000000", 20909 => x"00000000",
    20910 => x"00000000", 20911 => x"00000000", 20912 => x"00000000",
    20913 => x"00000000", 20914 => x"00000000", 20915 => x"00000000",
    20916 => x"00000000", 20917 => x"00000000", 20918 => x"00000000",
    20919 => x"00000000", 20920 => x"00000000", 20921 => x"00000000",
    20922 => x"00000000", 20923 => x"00000000", 20924 => x"00000000",
    20925 => x"00000000", 20926 => x"00000000", 20927 => x"00000000",
    20928 => x"00000000", 20929 => x"00000000", 20930 => x"00000000",
    20931 => x"00000000", 20932 => x"00000000", 20933 => x"00011f4c",
    20934 => x"00011f4c", 20935 => x"00000000", 20936 => x"00000001",
    20937 => x"00000000", 20938 => x"00000000", 20939 => x"00000000",
    20940 => x"00000000", 20941 => x"00000000", 20942 => x"00000000",
    20943 => x"00000000", 20944 => x"00000000", 20945 => x"00000000",
    20946 => x"00000000", 20947 => x"00000000", 20948 => x"00000000",
    20949 => x"00000000", 20950 => x"000143e4", 20951 => x"00015038",
    20952 => x"00000000", 20953 => x"00015078", 20954 => x"00015094",
    20955 => x"000150c4", 20956 => x"000150e4", 20957 => x"00000000",
    20958 => x"00000000", 20959 => x"00000000", 20960 => x"00000000",
    20961 => x"00000000", 20962 => x"00000000", 20963 => x"00000000",
    20964 => x"00000000", 20965 => x"00000000", 20966 => x"00015108",
    20967 => x"000003e8", 20968 => x"00000000", 20969 => x"00000000",
    20970 => x"00000000", 20971 => x"00000000", 20972 => x"000147b4",
    20973 => x"00014820", 20974 => x"00000000", 20975 => x"00000000",
    20976 => x"00000000", 20977 => x"00000000", 20978 => x"00000000",
    20979 => x"00000000", 20980 => x"00000000", 20981 => x"00000000",
    20982 => x"00000000", 20983 => x"00000000", 20984 => x"00000000",
    20985 => x"00000000", 20986 => x"00000000", 20987 => x"00000000",
    20988 => x"00000000", 20989 => x"00000000", 20990 => x"00000000",
    20991 => x"00000000", 20992 => x"00000000", 20993 => x"00000000",
    20994 => x"00000000", 20995 => x"00000000", 20996 => x"00000000",
    20997 => x"00000000", 20998 => x"00000000", 20999 => x"00000000",
    21000 => x"000015c0", 21001 => x"000015f4", 21002 => x"00001674",
    21003 => x"0000167c", 21004 => x"000016d4", 21005 => x"00001700",
    21006 => x"00001758", 21007 => x"0000177c", 21008 => x"00001840",
    21009 => x"00001848", 21010 => x"00001850", 21011 => x"000018b4",
    21012 => x"000018d0", 21013 => x"000016a0", 21014 => x"00000000",
    21015 => x"00002838", 21016 => x"000027bc", 21017 => x"00002760",
    21018 => x"00002708", 21019 => x"00000000", 21020 => x"00000000",
    21021 => x"000026d8", 21022 => x"00002ac4", 21023 => x"00002aa4",
    21024 => x"000029d4", 21025 => x"000028b8", 21026 => x"00000000",
    21027 => x"00000001", 21028 => x"0001242c", 21029 => x"00005238",
    21030 => x"00000002", 21031 => x"0001243c", 21032 => x"00005404",
    21033 => x"00000003", 21034 => x"00012444", 21035 => x"000054c0",
    21036 => x"00000004", 21037 => x"00012450", 21038 => x"000054d0",
    21039 => x"00000006", 21040 => x"00012954", 21041 => x"0000567c",
    21042 => x"00000008", 21043 => x"0001245c", 21044 => x"000059bc",
    21045 => x"00000009", 21046 => x"0001246c", 21047 => x"00005a30",
    21048 => x"00000064", 21049 => x"00012474", 21050 => x"000033b8",
    21051 => x"00000066", 21052 => x"0001248c", 21053 => x"00003530",
    21054 => x"00000065", 21055 => x"000124a0", 21056 => x"0000365c",
    21057 => x"00000067", 21058 => x"000124b8", 21059 => x"00003760",
    21060 => x"00000068", 21061 => x"000124d0", 21062 => x"0000388c",
    21063 => x"00000069", 21064 => x"000124e0", 21065 => x"00003ba8",
    21066 => x"0000006a", 21067 => x"000124f0", 21068 => x"00003cbc",
    21069 => x"0000006b", 21070 => x"00012504", 21071 => x"00003e40",
    21072 => x"00000000", 21073 => x"00000000", 21074 => x"00000000",
    21075 => x"00000001", 21076 => x"0001242c", 21077 => x"00005238",
    21078 => x"00000002", 21079 => x"0001243c", 21080 => x"00005404",
    21081 => x"00000003", 21082 => x"00012444", 21083 => x"000054c0",
    21084 => x"00000004", 21085 => x"00012450", 21086 => x"000054d0",
    21087 => x"00000005", 21088 => x"00012950", 21089 => x"000055e8",
    21090 => x"00000006", 21091 => x"00012954", 21092 => x"0000567c",
    21093 => x"00000007", 21094 => x"0001295c", 21095 => x"000058f8",
    21096 => x"00000008", 21097 => x"0001245c", 21098 => x"000059bc",
    21099 => x"00000009", 21100 => x"0001246c", 21101 => x"00005a30",
    21102 => x"00000000", 21103 => x"00000000", 21104 => x"00000000",
    21105 => x"00002dbc", 21106 => x"00002cdc", 21107 => x"00000000",
    21108 => x"00002c94", 21109 => x"00003154", 21110 => x"0000310c",
    21111 => x"00003020", 21112 => x"00002c04", 21113 => x"00002b78",
    21114 => x"00002fa8", 21115 => x"00002f30", 21116 => x"00002ec8",
    21117 => x"00002e5c", 21118 => x"00000001", 21119 => x"00012b68",
    21120 => x"00012b70", 21121 => x"00012b7c", 21122 => x"00012b88",
    21123 => x"00000000", 21124 => x"00000000", 21125 => x"00000000",
    21126 => x"00000000", 21127 => x"00012bac", 21128 => x"00012b94",
    21129 => x"00012ba0", 21130 => x"00012bb8", 21131 => x"00012bc4",
    21132 => x"00012bd0", 21133 => x"00000000", 21134 => x"00000000",
    21135 => x"00012ef8", 21136 => x"00012f08", 21137 => x"00012f14",
    21138 => x"00012f28", 21139 => x"00012f3c", 21140 => x"00012f4c",
    21141 => x"00012f58", 21142 => x"00012f64", 21143 => x"bbfef060",
    21144 => x"00000000", 21145 => x"00000000", 21146 => x"00000000",
    21147 => x"00000000", 21148 => x"00000000", 21149 => x"00000000",
    21150 => x"00000000", 21151 => x"00000000", 21152 => x"00000000",
    21153 => x"00000000", 21154 => x"00000000", 21155 => x"00000000",
    21156 => x"00000001", 21157 => x"00000000", 21158 => x"000a03e8",
    21159 => x"00060100", 21160 => x"80800000", 21161 => x"00000000",
    21162 => x"00000000", 21163 => x"00000000", 21164 => x"00000000",
    21165 => x"00000000", 21166 => x"00000000", 21167 => x"44332211",
    21168 => x"00000000", 21169 => x"04000000", 21170 => x"1b8046e2",
    21171 => x"01000000", 21172 => x"9800cfea", 21173 => x"01000000",
    21174 => x"188157f3", 21175 => x"01000000", 21176 => x"0be0ffff",
    21177 => x"01000000", 21178 => x"88e0ffff", 21179 => x"01000000",
    21180 => x"08e1ffff", 21181 => x"01000000", 21182 => x"136023e0",
    21183 => x"01000000", 21184 => x"900020e3", 21185 => x"01000000",
    21186 => x"100100e0", 21187 => x"01000000", 21188 => x"230300e1",
    21189 => x"01000000", 21190 => x"2be31ef1", 21191 => x"01000000",
    21192 => x"33c300e1", 21193 => x"01000000", 21194 => x"4be37ffb",
    21195 => x"01000000", 21196 => x"bb250060", 21197 => x"00000000",
    21198 => x"c3250260", 21199 => x"00000000", 21200 => x"59031000",
    21201 => x"04000000", 21202 => x"61611000", 21203 => x"04000000",
    21204 => x"78c19400", 21205 => x"04000000", 21206 => x"80ebbc00",
    21207 => x"04000000", 21208 => x"7b8908e0", 21209 => x"01000000",
    21210 => x"780f3100", 21211 => x"04000000", 21212 => x"810f8201",
    21213 => x"04000000", 21214 => x"53097afd", 21215 => x"01000000",
    21216 => x"c3108001", 21217 => x"04000000", 21218 => x"e90a8001",
    21219 => x"04000000", 21220 => x"f9508103", 21221 => x"04000000",
    21222 => x"00000000", 21223 => x"08000000", 21224 => x"00000004",
    21225 => x"00000008", 21226 => x"00000100", 21227 => x"00000200",
    21228 => x"00016dcc", 21229 => x"00000000", 21230 => x"00000000",
    21231 => x"0000ce42", 21232 => x"ab28633a", 21233 => x"00000000",
    21234 => x"00016d00", 21235 => x"00000000", 21236 => x"00000000",
    21237 => x"0000ce42", 21238 => x"650c2d4f", 21239 => x"00000000",
    21240 => x"00016dd4", 21241 => x"00000000", 21242 => x"00000000",
    21243 => x"0000ce42", 21244 => x"65158dc0", 21245 => x"00000000",
    21246 => x"00016d10", 21247 => x"00000000", 21248 => x"00000000",
    21249 => x"0000ce42", 21250 => x"de0d8ced", 21251 => x"00000000",
    21252 => x"00016dd0", 21253 => x"00000000", 21254 => x"00000000",
    21255 => x"0000ce42", 21256 => x"ff07fc47", 21257 => x"00000000",
    21258 => x"00016da4", 21259 => x"00000000", 21260 => x"00000000",
    21261 => x"0000ce42", 21262 => x"e2d13d04", 21263 => x"00000000",
    21264 => x"00016da0", 21265 => x"00000000", 21266 => x"00000000",
    21267 => x"0000ce42", 21268 => x"779c5443", 21269 => x"00000000",
    21270 => x"00016dc8", 21271 => x"00000000", 21272 => x"00000000",
    21273 => x"00000651", 21274 => x"68202b22", 21275 => x"00000000",
    21276 => x"00016dc0", 21277 => x"00000000", 21278 => x"00000000",
    21279 => x"00001103", 21280 => x"c0413599", 21281 => x"00000000",
    21282 => x"000136b4", 21283 => x"00000000", 21284 => x"00000001",
    21285 => x"00030000", 21286 => x"00000004", 21287 => x"00000000",
    21288 => x"00000000", 21289 => x"00000000", 21290 => x"00000000",
    21291 => x"00000000", 21292 => x"00000000", 21293 => x"00000000",
    21294 => x"00000000", 21295 => x"00000000", 21296 => x"00000000",
    21297 => x"00000000", 21298 => x"00000000", 21299 => x"00000000",
    21300 => x"00000000", 21301 => x"00000000", 21302 => x"00000000",
    21303 => x"00000000", 21304 => x"00000000", 21305 => x"00000000",
    21306 => x"00000000", 21307 => x"00000000", 21308 => x"00000000",
    21309 => x"00000000", 21310 => x"00000000", 21311 => x"00000000",
    21312 => x"00000000", 21313 => x"00000000", 21314 => x"00000000",
    21315 => x"00000000", 21316 => x"00000000", 21317 => x"00000000",
    21318 => x"00000000", 21319 => x"00000000", 21320 => x"00000000",
    21321 => x"00000000", 21322 => x"00000000", 21323 => x"00000000",
    21324 => x"00000000", 21325 => x"00000000", 21326 => x"00000000",
    21327 => x"00000000", 21328 => x"0000de7c", 21329 => x"0000deb0",
    21330 => x"0000dee0", 21331 => x"ffffffff", 21332 => x"000142b8",
    21333 => x"5b1157a7", 21334 => x"00000002", 21335 => x"00000000",
    21336 => x"00000000", 21337 => x"00000000", 21338 => x"00000000",
    21339 => x"00000000", 21340 => x"00000000", 21341 => x"00000000",
    21342 => x"00000000", 21343 => x"00000000", 21344 => x"00000000",
    21345 => x"00000000", 21346 => x"77727063", 21347 => x"2d76332e",
    21348 => x"302d342d", 21349 => x"67313934", 21350 => x"64626231",
    21351 => x"2d646972", 21352 => x"74790000", 21353 => x"00000000",
    21354 => x"4a756e20", 21355 => x"31342032", 21356 => x"30313600",
    21357 => x"00000000", 21358 => x"31313a34", 21359 => x"313a3336",
    21360 => x"00000000", 21361 => x"00000000", 21362 => x"000130a0",
    21363 => x"000086b4", 21364 => x"000130f4", 21365 => x"00008768",
    21366 => x"00013220", 21367 => x"000089d0", 21368 => x"000130b0",
    21369 => x"00008d80", 21370 => x"00013240", 21371 => x"00008e84",
    21372 => x"00013248", 21373 => x"00008ee4", 21374 => x"000132b4",
    21375 => x"00008f80", 21376 => x"000132f0", 21377 => x"00009058",
    21378 => x"000132f8", 21379 => x"000091b4", 21380 => x"000132fc",
    21381 => x"000091cc", 21382 => x"00013340", 21383 => x"00009248",
    21384 => x"000130a4", 21385 => x"00009360", 21386 => x"000133d0",
    21387 => x"00009470", 21388 => x"000133f8", 21389 => x"0000951c",
    21390 => x"0001341c", 21391 => x"00009588", 21392 => x"0001345c",
    21393 => x"000095e8", 21394 => x"00013478", 21395 => x"000096dc",
    21396 => x"000138a4", 21397 => x"0000e12c", 21398 => x"000138a8",
    21399 => x"0000e030", 21400 => x"000138ac", 21401 => x"0000df34",
    21402 => x"00000000", 21403 => x"00000000", 21404 => x"00000000",
    21405 => x"00000000", 21406 => x"00000000", 21407 => x"00000000",
    21408 => x"00000000", 21409 => x"00000000", 21410 => x"00000000",
    21411 => x"00000000", 21412 => x"00000000", 21413 => x"00000000",
    21414 => x"00000000", 21415 => x"00000000", 21416 => x"00000000",
    21417 => x"00000000", 21418 => x"00000000", 21419 => x"00000000",
    21420 => x"00000000", 21421 => x"00000000", 21422 => x"00000000",
    21423 => x"00000000", 21424 => x"00000000", 21425 => x"00000000",
    21426 => x"00000000", 21427 => x"00000000", 21428 => x"00000000",
    21429 => x"00000000", 21430 => x"00000000", 21431 => x"00000000",
    21432 => x"00000000", 21433 => x"00000000", 21434 => x"00000000",
    21435 => x"00000000", 21436 => x"00000000", 21437 => x"00000000",
    21438 => x"00000000", 21439 => x"00000000", 21440 => x"00000000",
    21441 => x"00000000", 21442 => x"00000000", 21443 => x"00000000",
    21444 => x"00000000", 21445 => x"00000000", 21446 => x"00000000",
    21447 => x"00000000", 21448 => x"00000000", 21449 => x"00000000",
    21450 => x"00000000", 21451 => x"00000000", 21452 => x"00000000",
    21453 => x"00000000", 21454 => x"00000000", 21455 => x"00000000",
    21456 => x"00000000", 21457 => x"00000000", 21458 => x"00000000",
    21459 => x"00000000", 21460 => x"00000000", 21461 => x"00000000",
    21462 => x"00000000", 21463 => x"00000000", 21464 => x"00000000",
    21465 => x"00000000", 21466 => x"00000000", 21467 => x"00000000",
    21468 => x"00000000", 21469 => x"00000000", 21470 => x"00000000",
    21471 => x"00000000", 21472 => x"00000000", 21473 => x"00000000",
    21474 => x"00000000", 21475 => x"00000000", 21476 => x"00000000",
    21477 => x"00000000", 21478 => x"00000000", 21479 => x"00000000",
    21480 => x"00000000", 21481 => x"00000000", 21482 => x"00000000",
    21483 => x"00000000", 21484 => x"00000000", 21485 => x"00000000",
    21486 => x"00000000", 21487 => x"00000000", 21488 => x"00000000",
    21489 => x"00000000", 21490 => x"00000000", 21491 => x"00000000",
    21492 => x"00000000", 21493 => x"00000000", 21494 => x"00000000",
    21495 => x"00000000", 21496 => x"00000000", 21497 => x"00000000",
    21498 => x"00000000", 21499 => x"00000000", 21500 => x"00000000",
    21501 => x"00000000", 21502 => x"00000000", 21503 => x"00000000",
    21504 => x"00000000", 21505 => x"00000000", 21506 => x"00000000",
    21507 => x"00000000", 21508 => x"00000000", 21509 => x"00000000",
    21510 => x"00000000", 21511 => x"00000000", 21512 => x"00000000",
    21513 => x"00000000", 21514 => x"00000000", 21515 => x"00000000",
    21516 => x"00000000", 21517 => x"00000000", 21518 => x"00000000",
    21519 => x"00000000", 21520 => x"00000000", 21521 => x"00000000",
    21522 => x"00000000", 21523 => x"00000000", 21524 => x"00000000",
    21525 => x"00000000", 21526 => x"00000000", 21527 => x"00000000",
    21528 => x"00000000", 21529 => x"00000000", 21530 => x"00000000",
    21531 => x"00000000", 21532 => x"00000000", 21533 => x"00000000",
    21534 => x"00000000", 21535 => x"00000000", 21536 => x"00000000",
    21537 => x"00000000", 21538 => x"00000000", 21539 => x"00000000",
    21540 => x"00000000", 21541 => x"00000000", 21542 => x"00000000",
    21543 => x"00000000", 21544 => x"00000000", 21545 => x"00000000",
    21546 => x"00000000", 21547 => x"00000000", 21548 => x"00000000",
    21549 => x"00000000", 21550 => x"00000000", 21551 => x"00000000",
    21552 => x"00000000", 21553 => x"00000000", 21554 => x"00000000",
    21555 => x"00000000", 21556 => x"00000000", 21557 => x"00000000",
    21558 => x"00000000", 21559 => x"00000000", 21560 => x"00000000",
    21561 => x"00000000", 21562 => x"00000000", 21563 => x"00000000",
    21564 => x"00000000", 21565 => x"00000000", 21566 => x"00000000",
    21567 => x"00000000", 21568 => x"00000000", 21569 => x"00000000",
    21570 => x"00000000", 21571 => x"00000000", 21572 => x"00000000",
    21573 => x"00000000", 21574 => x"00000000", 21575 => x"00000000",
    21576 => x"00000000", 21577 => x"00000000", 21578 => x"00000000",
    21579 => x"00000000", 21580 => x"00000000", 21581 => x"00000000",
    21582 => x"00000000", 21583 => x"00000000", 21584 => x"00000000",
    21585 => x"00000000", 21586 => x"00000000", 21587 => x"00000000",
    21588 => x"00000000", 21589 => x"00000000", 21590 => x"00000000",
    21591 => x"00000000", 21592 => x"00000000", 21593 => x"00000000",
    21594 => x"00000000", 21595 => x"00000000", 21596 => x"00000000",
    21597 => x"00000000", 21598 => x"00000000", 21599 => x"00000000",
    21600 => x"00000000", 21601 => x"00000000", 21602 => x"00000000",
    21603 => x"00000000", 21604 => x"00000000", 21605 => x"00000000",
    21606 => x"00000000", 21607 => x"00000000", 21608 => x"00000000",
    21609 => x"00000000", 21610 => x"00000000", 21611 => x"00000000",
    21612 => x"00000000", 21613 => x"00000000", 21614 => x"00000000",
    21615 => x"00000000", 21616 => x"00000000", 21617 => x"00000000",
    21618 => x"00000000", 21619 => x"00000000", 21620 => x"00000000",
    21621 => x"00000000", 21622 => x"00000000", 21623 => x"00000000",
    21624 => x"00000000", 21625 => x"00000000", 21626 => x"00000000",
    21627 => x"00000000", 21628 => x"00000000", 21629 => x"00000000",
    21630 => x"00000000", 21631 => x"00000000", 21632 => x"00000000",
    21633 => x"00000000", 21634 => x"00000000", 21635 => x"00000000",
    21636 => x"00000000", 21637 => x"00000000", 21638 => x"00000000",
    21639 => x"00000000", 21640 => x"00000000", 21641 => x"00000000",
    21642 => x"00000000", 21643 => x"00000000", 21644 => x"00000000",
    21645 => x"00000000", 21646 => x"00000000", 21647 => x"00000000",
    21648 => x"00000000", 21649 => x"00000000", 21650 => x"00000000",
    21651 => x"00000000", 21652 => x"00000000", 21653 => x"00000000",
    21654 => x"00000000", 21655 => x"00000000", 21656 => x"00000000",
    21657 => x"00000000", 21658 => x"00000000", 21659 => x"00000000",
    21660 => x"00000000", 21661 => x"00000000", 21662 => x"00000000",
    21663 => x"00000000", 21664 => x"00000000", 21665 => x"00000000",
    21666 => x"00000000", 21667 => x"00000000", 21668 => x"00000000",
    21669 => x"00000000", 21670 => x"00000000", 21671 => x"00000000",
    21672 => x"00000000", 21673 => x"00000000", 21674 => x"00000000",
    21675 => x"00000000", 21676 => x"00000000", 21677 => x"00000000",
    21678 => x"00000000", 21679 => x"00000000", 21680 => x"00000000",
    21681 => x"00000000", 21682 => x"00000000", 21683 => x"00000000",
    21684 => x"00000000", 21685 => x"00000000", 21686 => x"00000000",
    21687 => x"00000000", 21688 => x"00000000", 21689 => x"00000000",
    21690 => x"00000000", 21691 => x"00000000", 21692 => x"00000000",
    21693 => x"00000000", 21694 => x"00000000", 21695 => x"00000000",
    21696 => x"00000000", 21697 => x"00000000", 21698 => x"00000000",
    21699 => x"00000000", 21700 => x"00000000", 21701 => x"00000000",
    21702 => x"00000000", 21703 => x"00000000", 21704 => x"00000000",
    21705 => x"00000000", 21706 => x"00000000", 21707 => x"00000000",
    21708 => x"00000000", 21709 => x"00000000", 21710 => x"00000000",
    21711 => x"00000000", 21712 => x"00000000", 21713 => x"00000000",
    21714 => x"00000000", 21715 => x"00000000", 21716 => x"00000000",
    21717 => x"00000000", 21718 => x"00000000", 21719 => x"00000000",
    21720 => x"00000000", 21721 => x"00000000", 21722 => x"00000000",
    21723 => x"00000000", 21724 => x"00000000", 21725 => x"00000000",
    21726 => x"00000000", 21727 => x"00000000", 21728 => x"00000000",
    21729 => x"00000000", 21730 => x"00000000", 21731 => x"00000000",
    21732 => x"00000000", 21733 => x"00000000", 21734 => x"00000000",
    21735 => x"00000000", 21736 => x"00000000", 21737 => x"00000000",
    21738 => x"00000000", 21739 => x"00000000", 21740 => x"00000000",
    21741 => x"00000000", 21742 => x"00000000", 21743 => x"00000000",
    21744 => x"00000000", 21745 => x"00000000", 21746 => x"00000000",
    21747 => x"00000000", 21748 => x"00000000", 21749 => x"00000000",
    21750 => x"00000000", 21751 => x"00000000", 21752 => x"00000000",
    21753 => x"00000000", 21754 => x"00000000", 21755 => x"00000000",
    21756 => x"00000000", 21757 => x"00000000", 21758 => x"00000000",
    21759 => x"00000000", 21760 => x"00000000", 21761 => x"00000000",
    21762 => x"00000000", 21763 => x"00000000", 21764 => x"00000000",
    21765 => x"00000000", 21766 => x"00000000", 21767 => x"00000000",
    21768 => x"00000000", 21769 => x"00000000", 21770 => x"00000000",
    21771 => x"00000000", 21772 => x"00000000", 21773 => x"00000000",
    21774 => x"00000000", 21775 => x"00000000", 21776 => x"00000000",
    21777 => x"00000000", 21778 => x"00000000", 21779 => x"00000000",
    21780 => x"00000000", 21781 => x"00000000", 21782 => x"00000000",
    21783 => x"00000000", 21784 => x"00000000", 21785 => x"00000000",
    21786 => x"00000000", 21787 => x"00000000", 21788 => x"00000000",
    21789 => x"00000000", 21790 => x"00000000", 21791 => x"00000000",
    21792 => x"00000000", 21793 => x"00000000", 21794 => x"00000000",
    21795 => x"00000000", 21796 => x"00000000", 21797 => x"00000000",
    21798 => x"00000000", 21799 => x"00000000", 21800 => x"00000000",
    21801 => x"00000000", 21802 => x"00000000", 21803 => x"00000000",
    21804 => x"00000000", 21805 => x"00000000", 21806 => x"00000000",
    21807 => x"00000000", 21808 => x"00000000", 21809 => x"00000000",
    21810 => x"00000000", 21811 => x"00000000", 21812 => x"00000000",
    21813 => x"00000000", 21814 => x"00000000", 21815 => x"00000000",
    21816 => x"00000000", 21817 => x"00000000", 21818 => x"00000000",
    21819 => x"00000000", 21820 => x"00000000", 21821 => x"00000000",
    21822 => x"00000000", 21823 => x"00000000", 21824 => x"00000000",
    21825 => x"00000000", 21826 => x"00000000", 21827 => x"00000000",
    21828 => x"00000000", 21829 => x"00000000", 21830 => x"00000000",
    21831 => x"00000000", 21832 => x"00000000", 21833 => x"00000000",
    21834 => x"00000000", 21835 => x"00000000", 21836 => x"00000000",
    21837 => x"00000000", 21838 => x"00000000", 21839 => x"00000000",
    21840 => x"00000000", 21841 => x"00000000", 21842 => x"00000000",
    21843 => x"00000000", 21844 => x"00000000", 21845 => x"00000000",
    21846 => x"00000000", 21847 => x"00000000", 21848 => x"00000000",
    21849 => x"00000000", 21850 => x"00000000", 21851 => x"00000000",
    21852 => x"00000000", 21853 => x"00000000", 21854 => x"00000000",
    21855 => x"00000000", 21856 => x"00000000", 21857 => x"00000000",
    21858 => x"00000000", 21859 => x"00000000", 21860 => x"00000000",
    21861 => x"00000000", 21862 => x"00000000", 21863 => x"00000000",
    21864 => x"00000000", 21865 => x"00000000", 21866 => x"00000000",
    21867 => x"00000000", 21868 => x"00000000", 21869 => x"00000000",
    21870 => x"00000000", 21871 => x"00000000", 21872 => x"00000000",
    21873 => x"00000000", 21874 => x"00000000", 21875 => x"00000000",
    21876 => x"00000000", 21877 => x"00000000", 21878 => x"00000000",
    21879 => x"00000000", 21880 => x"00000000", 21881 => x"00000000",
    21882 => x"00000000", 21883 => x"00000000", 21884 => x"00000000",
    21885 => x"00000000", 21886 => x"00000000", 21887 => x"00000000",
    21888 => x"00000000", 21889 => x"00000000", 21890 => x"00000000",
    21891 => x"00000000", 21892 => x"00000000", 21893 => x"00000000",
    21894 => x"00000000", 21895 => x"00000000", 21896 => x"00000000",
    21897 => x"00000000", 21898 => x"00000000", 21899 => x"00000000",
    21900 => x"00000000", 21901 => x"00000000", 21902 => x"00000000",
    21903 => x"00000000", 21904 => x"00000000", 21905 => x"00000000",
    21906 => x"00000000", 21907 => x"00000000", 21908 => x"00000000",
    21909 => x"00000000", 21910 => x"00000000", 21911 => x"00000000",
    21912 => x"00000000", 21913 => x"00000000", 21914 => x"00000000",
    21915 => x"00000000", 21916 => x"00000000", 21917 => x"00000000",
    21918 => x"00000000", 21919 => x"00000000", 21920 => x"00000000",
    21921 => x"00000000", 21922 => x"00000000", 21923 => x"00000000",
    21924 => x"00000000", 21925 => x"00000000", 21926 => x"00000000",
    21927 => x"00000000", 21928 => x"00000000", 21929 => x"00000000",
    21930 => x"00000000", 21931 => x"00000000", 21932 => x"00000000",
    21933 => x"00000000", 21934 => x"00000000", 21935 => x"00000000",
    21936 => x"00000000", 21937 => x"00000000", 21938 => x"00000000",
    21939 => x"00000000", 21940 => x"00000000", 21941 => x"00000000",
    21942 => x"00000000", 21943 => x"00000000", 21944 => x"00000000",
    21945 => x"00000000", 21946 => x"00000000", 21947 => x"00000000",
    21948 => x"00000000", 21949 => x"00000000", 21950 => x"00000000",
    21951 => x"00000000", 21952 => x"00000000", 21953 => x"00000000",
    21954 => x"00000000", 21955 => x"00000000", 21956 => x"00000000",
    21957 => x"00000000", 21958 => x"00000000", 21959 => x"00000000",
    21960 => x"00000000", 21961 => x"00000000", 21962 => x"00000000",
    21963 => x"00000000", 21964 => x"00000000", 21965 => x"00000000",
    21966 => x"00000000", 21967 => x"00000000", 21968 => x"00000000",
    21969 => x"00000000", 21970 => x"00000000", 21971 => x"00000000",
    21972 => x"00000000", 21973 => x"00000000", 21974 => x"00000000",
    21975 => x"00000000", 21976 => x"00000000", 21977 => x"00000000",
    21978 => x"00000000", 21979 => x"00000000", 21980 => x"00000000",
    21981 => x"00000000", 21982 => x"00000000", 21983 => x"00000000",
    21984 => x"00000000", 21985 => x"00000000", 21986 => x"00000000",
    21987 => x"00000000", 21988 => x"00000000", 21989 => x"00000000",
    21990 => x"00000000", 21991 => x"00000000", 21992 => x"00000000",
    21993 => x"00000000", 21994 => x"00000000", 21995 => x"00000000",
    21996 => x"00000000", 21997 => x"00000000", 21998 => x"00000000",
    21999 => x"00000000", 22000 => x"00000000", 22001 => x"00000000",
    22002 => x"00000000", 22003 => x"00000000", 22004 => x"00000000",
    22005 => x"00000000", 22006 => x"00000000", 22007 => x"00000000",
    22008 => x"00000000", 22009 => x"00000000", 22010 => x"00000000",
    22011 => x"00000000", 22012 => x"00000000", 22013 => x"00000000",
    22014 => x"00000000", 22015 => x"00000000", 22016 => x"00000000",
    22017 => x"00000000", 22018 => x"00000000", 22019 => x"00000000",
    22020 => x"00000000", 22021 => x"00000000", 22022 => x"00000000",
    22023 => x"00000000", 22024 => x"00000000", 22025 => x"00000000",
    22026 => x"00000000", 22027 => x"00000000", 22028 => x"00000000",
    22029 => x"00000000", 22030 => x"00000000", 22031 => x"00000000",
    22032 => x"00000000", 22033 => x"00000000", 22034 => x"00000000",
    22035 => x"00000000", 22036 => x"00000000", 22037 => x"00000000",
    22038 => x"00000000", 22039 => x"00000000", 22040 => x"00000000",
    22041 => x"00000000", 22042 => x"00000000", 22043 => x"00000000",
    22044 => x"00000000", 22045 => x"00000000", 22046 => x"00000000",
    22047 => x"00000000", 22048 => x"00000000", 22049 => x"00000000",
    22050 => x"00000000", 22051 => x"00000000", 22052 => x"00000000",
    22053 => x"00000000", 22054 => x"00000000", 22055 => x"00000000",
    22056 => x"00000000", 22057 => x"00000000", 22058 => x"00000000",
    22059 => x"00000000", 22060 => x"00000000", 22061 => x"00000000",
    22062 => x"00000000", 22063 => x"00000000", 22064 => x"00000000",
    22065 => x"00000000", 22066 => x"00000000", 22067 => x"00000000",
    22068 => x"00000000", 22069 => x"00000000", 22070 => x"00000000",
    22071 => x"00000000", 22072 => x"00000000", 22073 => x"00000000",
    22074 => x"00000000", 22075 => x"00000000", 22076 => x"00000000",
    22077 => x"00000000", 22078 => x"00000000", 22079 => x"00000000",
    22080 => x"00000000", 22081 => x"00000000", 22082 => x"00000000",
    22083 => x"00000000", 22084 => x"00000000", 22085 => x"00000000",
    22086 => x"00000000", 22087 => x"00000000", 22088 => x"00000000",
    22089 => x"00000000", 22090 => x"00000000", 22091 => x"00000000",
    22092 => x"00000000", 22093 => x"00000000", 22094 => x"00000000",
    22095 => x"00000000", 22096 => x"00000000", 22097 => x"00000000",
    22098 => x"00000000", 22099 => x"00000000", 22100 => x"00000000",
    22101 => x"00000000", 22102 => x"00000000", 22103 => x"00000000",
    22104 => x"00000000", 22105 => x"00000000", 22106 => x"00000000",
    22107 => x"00000000", 22108 => x"00000000", 22109 => x"00000000",
    22110 => x"00000000", 22111 => x"00000000", 22112 => x"00000000",
    22113 => x"00000000", 22114 => x"00000000", 22115 => x"00000000",
    22116 => x"00000000", 22117 => x"00000000", 22118 => x"00000000",
    22119 => x"00000000", 22120 => x"00000000", 22121 => x"00000000",
    22122 => x"00000000", 22123 => x"00000000", 22124 => x"00000000",
    22125 => x"00000000", 22126 => x"00000000", 22127 => x"00000000",
    22128 => x"00000000", 22129 => x"00000000", 22130 => x"00000000",
    22131 => x"00000000", 22132 => x"00000000", 22133 => x"00000000",
    22134 => x"00000000", 22135 => x"00000000", 22136 => x"00000000",
    22137 => x"00000000", 22138 => x"00000000", 22139 => x"00000000",
    22140 => x"00000000", 22141 => x"00000000", 22142 => x"00000000",
    22143 => x"00000000", 22144 => x"00000000", 22145 => x"00000000",
    22146 => x"00000000", 22147 => x"00000000", 22148 => x"00000000",
    22149 => x"00000000", 22150 => x"00000000", 22151 => x"00000000",
    22152 => x"00000000", 22153 => x"00000000", 22154 => x"00000000",
    22155 => x"00000000", 22156 => x"00000000", 22157 => x"00000000",
    22158 => x"00000000", 22159 => x"00000000", 22160 => x"00000000",
    22161 => x"00000000", 22162 => x"00000000", 22163 => x"00000000",
    22164 => x"00000000", 22165 => x"00000000", 22166 => x"00000000",
    22167 => x"00000000", 22168 => x"00000000", 22169 => x"00000000",
    22170 => x"00000000", 22171 => x"00000000", 22172 => x"00000000",
    22173 => x"00000000", 22174 => x"00000000", 22175 => x"00000000",
    22176 => x"00000000", 22177 => x"00000000", 22178 => x"00000000",
    22179 => x"00000000", 22180 => x"00000000", 22181 => x"00000000",
    22182 => x"00000000", 22183 => x"00000000", 22184 => x"00000000",
    22185 => x"00000000", 22186 => x"00000000", 22187 => x"00000000",
    22188 => x"00000000", 22189 => x"00000000", 22190 => x"00000000",
    22191 => x"00000000", 22192 => x"00000000", 22193 => x"00000000",
    22194 => x"00000000", 22195 => x"00000000", 22196 => x"00000000",
    22197 => x"00000000", 22198 => x"00000000", 22199 => x"00000000",
    22200 => x"00000000", 22201 => x"00000000", 22202 => x"00000000",
    22203 => x"00000000", 22204 => x"00000000", 22205 => x"00000000",
    22206 => x"00000000", 22207 => x"00000000", 22208 => x"00000000",
    22209 => x"00000000", 22210 => x"00000000", 22211 => x"00000000",
    22212 => x"00000000", 22213 => x"00000000", 22214 => x"00000000",
    22215 => x"00000000", 22216 => x"00000000", 22217 => x"00000000",
    22218 => x"00000000", 22219 => x"00000000", 22220 => x"00000000",
    22221 => x"00000000", 22222 => x"00000000", 22223 => x"00000000",
    22224 => x"00000000", 22225 => x"00000000", 22226 => x"00000000",
    22227 => x"00000000", 22228 => x"00000000", 22229 => x"00000000",
    22230 => x"00000000", 22231 => x"00000000", 22232 => x"00000000",
    22233 => x"00000000", 22234 => x"00000000", 22235 => x"00000000",
    22236 => x"00000000", 22237 => x"00000000", 22238 => x"00000000",
    22239 => x"00000000", 22240 => x"00000000", 22241 => x"00000000",
    22242 => x"00000000", 22243 => x"00000000", 22244 => x"00000000",
    22245 => x"00000000", 22246 => x"00000000", 22247 => x"00000000",
    22248 => x"00000000", 22249 => x"00000000", 22250 => x"00000000",
    22251 => x"00000000", 22252 => x"00000000", 22253 => x"00000000",
    22254 => x"00000000", 22255 => x"00000000", 22256 => x"00000000",
    22257 => x"00000000", 22258 => x"00000000", 22259 => x"00000000",
    22260 => x"00000000", 22261 => x"00000000", 22262 => x"00000000",
    22263 => x"00000000", 22264 => x"00000000", 22265 => x"00000000",
    22266 => x"00000000", 22267 => x"00000000", 22268 => x"00000000",
    22269 => x"00000000", 22270 => x"00000000", 22271 => x"00000000",
    22272 => x"00000000", 22273 => x"00000000", 22274 => x"00000000",
    22275 => x"00000000", 22276 => x"00000000", 22277 => x"00000000",
    22278 => x"00000000", 22279 => x"00000000", 22280 => x"00000000",
    22281 => x"00000000", 22282 => x"00000000", 22283 => x"00000000",
    22284 => x"00000000", 22285 => x"00000000", 22286 => x"00000000",
    22287 => x"00000000", 22288 => x"00000000", 22289 => x"00000000",
    22290 => x"00000000", 22291 => x"00000000", 22292 => x"00000000",
    22293 => x"00000000", 22294 => x"00000000", 22295 => x"00000000",
    22296 => x"00000000", 22297 => x"00000000", 22298 => x"00000000",
    22299 => x"00000000", 22300 => x"00000000", 22301 => x"00000000",
    22302 => x"00000000", 22303 => x"00000000", 22304 => x"00000000",
    22305 => x"00000000", 22306 => x"00000000", 22307 => x"00000000",
    22308 => x"00000000", 22309 => x"00000000", 22310 => x"00000000",
    22311 => x"00000000", 22312 => x"00000000", 22313 => x"00000000",
    22314 => x"00000000", 22315 => x"00000000", 22316 => x"00000000",
    22317 => x"00000000", 22318 => x"00000000", 22319 => x"00000000",
    22320 => x"00000000", 22321 => x"00000000", 22322 => x"00000000",
    22323 => x"00000000", 22324 => x"00000000", 22325 => x"00000000",
    22326 => x"00000000", 22327 => x"00000000", 22328 => x"00000000",
    22329 => x"00000000", 22330 => x"00000000", 22331 => x"00000000",
    22332 => x"00000000", 22333 => x"00000000", 22334 => x"00000000",
    22335 => x"00000000", 22336 => x"00000000", 22337 => x"00000000",
    22338 => x"00000000", 22339 => x"00000000", 22340 => x"00000000",
    22341 => x"00000000", 22342 => x"00000000", 22343 => x"00000000",
    22344 => x"00000000", 22345 => x"00000000", 22346 => x"00000000",
    22347 => x"00000000", 22348 => x"00000000", 22349 => x"00000000",
    22350 => x"00000000", 22351 => x"00000000", 22352 => x"00000000",
    22353 => x"00000000", 22354 => x"00000000", 22355 => x"00000000",
    22356 => x"00000000", 22357 => x"00000000", 22358 => x"00000000",
    22359 => x"00000000", 22360 => x"00000000", 22361 => x"00000000",
    22362 => x"00000000", 22363 => x"00000000", 22364 => x"00000000",
    22365 => x"00000000", 22366 => x"00000000", 22367 => x"00000000",
    22368 => x"00000000", 22369 => x"00000000", 22370 => x"00000000",
    22371 => x"00000000", 22372 => x"00000000", 22373 => x"00000000",
    22374 => x"00000000", 22375 => x"00000000", 22376 => x"00000000",
    22377 => x"00000000", 22378 => x"00000000", 22379 => x"00000000",
    22380 => x"00000000", 22381 => x"00000000", 22382 => x"00000000",
    22383 => x"00000000", 22384 => x"00000000", 22385 => x"00000000",
    22386 => x"00000000", 22387 => x"00000000", 22388 => x"00000000",
    22389 => x"00000000", 22390 => x"00000000", 22391 => x"00000000",
    22392 => x"00000000", 22393 => x"00000000", 22394 => x"00000000",
    22395 => x"00000000", 22396 => x"00000000", 22397 => x"00000000",
    22398 => x"00000000", 22399 => x"00000000", 22400 => x"00000000",
    22401 => x"00000000", 22402 => x"00000000", 22403 => x"00000000",
    22404 => x"00000000", 22405 => x"00000000", 22406 => x"00000000",
    22407 => x"00000000", 22408 => x"00000000", 22409 => x"00000000",
    22410 => x"00000000", 22411 => x"00000000", 22412 => x"00000000",
    22413 => x"00000000", 22414 => x"00000000", 22415 => x"00000000",
    22416 => x"00000000", 22417 => x"00000000", 22418 => x"00000000",
    22419 => x"00000000", 22420 => x"00000000", 22421 => x"00000000",
    22422 => x"00000000", 22423 => x"00000000", 22424 => x"00000000",
    22425 => x"00000000", 22426 => x"00000000", 22427 => x"00000000",
    22428 => x"00000000", 22429 => x"00000000", 22430 => x"00000000",
    22431 => x"00000000", 22432 => x"00000000", 22433 => x"00000000",
    22434 => x"00000000", 22435 => x"00000000", 22436 => x"00000000",
    22437 => x"00000000", 22438 => x"00000000", 22439 => x"00000000",
    22440 => x"00000000", 22441 => x"00000000", 22442 => x"00000000",
    22443 => x"00000000", 22444 => x"00000000", 22445 => x"00000000",
    22446 => x"00000000", 22447 => x"00000000", 22448 => x"00000000",
    22449 => x"00000000", 22450 => x"00000000", 22451 => x"00000000",
    22452 => x"00000000", 22453 => x"00000000", 22454 => x"00000000",
    22455 => x"00000000", 22456 => x"00000000", 22457 => x"00000000",
    22458 => x"00000000", 22459 => x"00000000", 22460 => x"00000000",
    22461 => x"00000000", 22462 => x"00000000", 22463 => x"00000000",
    22464 => x"00000000", 22465 => x"00000000", 22466 => x"00000000",
    22467 => x"00000000", 22468 => x"00000000", 22469 => x"00000000",
    22470 => x"00000000", 22471 => x"00000000", 22472 => x"00000000",
    22473 => x"00000000", 22474 => x"00000000", 22475 => x"00000000",
    22476 => x"00000000", 22477 => x"00000000", 22478 => x"00000000",
    22479 => x"00000000", 22480 => x"00000000", 22481 => x"00000000",
    22482 => x"00000000", 22483 => x"00000000", 22484 => x"00000000",
    22485 => x"00000000", 22486 => x"00000000", 22487 => x"00000000",
    22488 => x"00000000", 22489 => x"00000000", 22490 => x"00000000",
    22491 => x"00000000", 22492 => x"00000000", 22493 => x"00000000",
    22494 => x"00000000", 22495 => x"00000000", 22496 => x"00000000",
    22497 => x"00000000", 22498 => x"00000000", 22499 => x"00000000",
    22500 => x"00000000", 22501 => x"00000000", 22502 => x"00000000",
    22503 => x"00000000", 22504 => x"00000000", 22505 => x"00000000",
    22506 => x"00000000", 22507 => x"00000000", 22508 => x"00000000",
    22509 => x"00000000", 22510 => x"00000000", 22511 => x"00000000",
    22512 => x"00000000", 22513 => x"00000000", 22514 => x"00000000",
    22515 => x"00000000", 22516 => x"00000000", 22517 => x"00000000",
    22518 => x"00000000", 22519 => x"00000000", 22520 => x"00000000",
    22521 => x"00000000", 22522 => x"00000000", 22523 => x"00000000",
    22524 => x"00000000", 22525 => x"00000000", 22526 => x"00000000",
    22527 => x"00000000", 22528 => x"00000000", 22529 => x"00000000",
    22530 => x"00000000", 22531 => x"00000000", 22532 => x"00000000",
    22533 => x"00000000", 22534 => x"00000000", 22535 => x"00000000",
    22536 => x"00000000", 22537 => x"00000000", 22538 => x"00000000",
    22539 => x"00000000", 22540 => x"00000000", 22541 => x"00000000",
    22542 => x"00000000", 22543 => x"00000000", 22544 => x"00000000",
    22545 => x"00000000", 22546 => x"00000000", 22547 => x"00000000",
    22548 => x"00000000", 22549 => x"00000000", 22550 => x"00000000",
    22551 => x"00000000", 22552 => x"00000000", 22553 => x"00000000",
    22554 => x"00000000", 22555 => x"00000000", 22556 => x"00000000",
    22557 => x"00000000", 22558 => x"00000000", 22559 => x"00000000",
    22560 => x"00000000", 22561 => x"00000000", 22562 => x"00000000",
    22563 => x"00000000", 22564 => x"00000000", 22565 => x"00000000",
    22566 => x"00000000", 22567 => x"00000000", 22568 => x"00000000",
    22569 => x"00000000", 22570 => x"00000000", 22571 => x"00000000",
    22572 => x"00000000", 22573 => x"00000000", 22574 => x"00000000",
    22575 => x"00000000", 22576 => x"00000000", 22577 => x"00000000",
    22578 => x"00000000", 22579 => x"00000000", 22580 => x"00000000",
    22581 => x"00000000", 22582 => x"00000000", 22583 => x"00000000",
    22584 => x"00000000", 22585 => x"00000000", 22586 => x"00000000",
    22587 => x"00000000", 22588 => x"00000000", 22589 => x"00000000",
    22590 => x"00000000", 22591 => x"00000000", 22592 => x"00000000",
    22593 => x"00000000", 22594 => x"00000000", 22595 => x"00000000",
    22596 => x"00000000", 22597 => x"00000000", 22598 => x"00000000",
    22599 => x"00000000", 22600 => x"00000000", 22601 => x"00000000",
    22602 => x"00000000", 22603 => x"00000000", 22604 => x"00000000",
    22605 => x"00000000", 22606 => x"00000000", 22607 => x"00000000",
    22608 => x"00000000", 22609 => x"00000000", 22610 => x"00000000",
    22611 => x"00000000", 22612 => x"00000000", 22613 => x"00000000",
    22614 => x"00000000", 22615 => x"00000000", 22616 => x"00000000",
    22617 => x"00000000", 22618 => x"00000000", 22619 => x"00000000",
    22620 => x"00000000", 22621 => x"00000000", 22622 => x"00000000",
    22623 => x"00000000", 22624 => x"00000000", 22625 => x"00000000",
    22626 => x"00000000", 22627 => x"00000000", 22628 => x"00000000",
    22629 => x"00000000", 22630 => x"00000000", 22631 => x"00000000",
    22632 => x"00000000", 22633 => x"00000000", 22634 => x"00000000",
    22635 => x"00000000", 22636 => x"00000000", 22637 => x"00000000",
    22638 => x"00000000", 22639 => x"00000000", 22640 => x"00000000",
    22641 => x"00000000", 22642 => x"00000000", 22643 => x"00000000",
    22644 => x"00000000", 22645 => x"00000000", 22646 => x"00000000",
    22647 => x"00000000", 22648 => x"00000000", 22649 => x"00000000",
    22650 => x"00000000", 22651 => x"00000000", 22652 => x"00000000",
    22653 => x"00000000", 22654 => x"00000000", 22655 => x"00000000",
    22656 => x"00000000", 22657 => x"00000000", 22658 => x"00000000",
    22659 => x"00000000", 22660 => x"00000000", 22661 => x"00000000",
    22662 => x"00000000", 22663 => x"00000000", 22664 => x"00000000",
    22665 => x"00000000", 22666 => x"00000000", 22667 => x"00000000",
    22668 => x"00000000", 22669 => x"00000000", 22670 => x"00000000",
    22671 => x"00000000", 22672 => x"00000000", 22673 => x"00000000",
    22674 => x"00000000", 22675 => x"00000000", 22676 => x"00000000",
    22677 => x"00000000", 22678 => x"00000000", 22679 => x"00000000",
    22680 => x"00000000", 22681 => x"00000000", 22682 => x"00000000",
    22683 => x"00000000", 22684 => x"00000000", 22685 => x"00000000",
    22686 => x"00000000", 22687 => x"00000000", 22688 => x"00000000",
    22689 => x"00000000", 22690 => x"00000000", 22691 => x"00000000",
    22692 => x"00000000", 22693 => x"00000000", 22694 => x"00000000",
    22695 => x"00000000", 22696 => x"00000000", 22697 => x"00000000",
    22698 => x"00000000", 22699 => x"00000000", 22700 => x"00000000",
    22701 => x"00000000", 22702 => x"00000000", 22703 => x"00000000",
    22704 => x"00000000", 22705 => x"00000000", 22706 => x"00000000",
    22707 => x"00000000", 22708 => x"00000000", 22709 => x"00000000",
    22710 => x"00000000", 22711 => x"00000000", 22712 => x"00000000",
    22713 => x"00000000", 22714 => x"00000000", 22715 => x"00000000",
    22716 => x"00000000", 22717 => x"00000000", 22718 => x"00000000",
    22719 => x"00000000", 22720 => x"00000000", 22721 => x"00000000",
    22722 => x"00000000", 22723 => x"00000000", 22724 => x"00000000",
    22725 => x"00000000", 22726 => x"00000000", 22727 => x"00000000",
    22728 => x"00000000", 22729 => x"00000000", 22730 => x"00000000",
    22731 => x"00000000", 22732 => x"00000000", 22733 => x"00000000",
    22734 => x"00000000", 22735 => x"00000000", 22736 => x"00000000",
    22737 => x"00000000", 22738 => x"00000000", 22739 => x"00000000",
    22740 => x"00000000", 22741 => x"00000000", 22742 => x"00000000",
    22743 => x"00000000", 22744 => x"00000000", 22745 => x"00000000",
    22746 => x"00000000", 22747 => x"00000000", 22748 => x"00000000",
    22749 => x"00000000", 22750 => x"00000000", 22751 => x"00000000",
    22752 => x"00000000", 22753 => x"00000000", 22754 => x"00000000",
    22755 => x"00000000", 22756 => x"00000000", 22757 => x"00000000",
    22758 => x"00000000", 22759 => x"00000000", 22760 => x"00000000",
    22761 => x"00000000", 22762 => x"00000000", 22763 => x"00000000",
    22764 => x"00000000", 22765 => x"00000000", 22766 => x"00000000",
    22767 => x"00000000", 22768 => x"00000000", 22769 => x"00000000",
    22770 => x"00000000", 22771 => x"00000000", 22772 => x"00000000",
    22773 => x"00000000", 22774 => x"00000000", 22775 => x"00000000",
    22776 => x"00000000", 22777 => x"00000000", 22778 => x"00000000",
    22779 => x"00000000", 22780 => x"00000000", 22781 => x"00000000",
    22782 => x"00000000", 22783 => x"00000000", 22784 => x"00000000",
    22785 => x"00000000", 22786 => x"00000000", 22787 => x"00000000",
    22788 => x"00000000", 22789 => x"00000000", 22790 => x"00000000",
    22791 => x"00000000", 22792 => x"00000000", 22793 => x"00000000",
    22794 => x"00000000", 22795 => x"00000000", 22796 => x"00000000",
    22797 => x"00000000", 22798 => x"00000000", 22799 => x"00000000",
    22800 => x"00000000", 22801 => x"00000000", 22802 => x"00000000",
    22803 => x"00000000", 22804 => x"00000000", 22805 => x"00000000",
    22806 => x"00000000", 22807 => x"00000000", 22808 => x"00000000",
    22809 => x"00000000", 22810 => x"00000000", 22811 => x"00000000",
    22812 => x"00000000", 22813 => x"00000000", 22814 => x"00000000",
    22815 => x"00000000", 22816 => x"00000000", 22817 => x"00000000",
    22818 => x"00000000", 22819 => x"00000000", 22820 => x"00000000",
    22821 => x"00000000", 22822 => x"00000000", 22823 => x"00000000",
    22824 => x"00000000", 22825 => x"00000000", 22826 => x"00000000",
    22827 => x"00000000", 22828 => x"00000000", 22829 => x"00000000",
    22830 => x"00000000", 22831 => x"00000000", 22832 => x"00000000",
    22833 => x"00000000", 22834 => x"00000000", 22835 => x"00000000",
    22836 => x"00000000", 22837 => x"00000000", 22838 => x"00000000",
    22839 => x"00000000", 22840 => x"00000000", 22841 => x"00000000",
    22842 => x"00000000", 22843 => x"00000000", 22844 => x"00000000",
    22845 => x"00000000", 22846 => x"00000000", 22847 => x"00000000",
    22848 => x"00000000", 22849 => x"00000000", 22850 => x"00000000",
    22851 => x"00000000", 22852 => x"00000000", 22853 => x"00000000",
    22854 => x"00000000", 22855 => x"00000000", 22856 => x"00000000",
    22857 => x"00000000", 22858 => x"00000000", 22859 => x"00000000",
    22860 => x"00000000", 22861 => x"00000000", 22862 => x"00000000",
    22863 => x"00000000", 22864 => x"00000000", 22865 => x"00000000",
    22866 => x"00000000", 22867 => x"00000000", 22868 => x"00000000",
    22869 => x"00000000", 22870 => x"00000000", 22871 => x"00000000",
    22872 => x"00000000", 22873 => x"00000000", 22874 => x"00000000",
    22875 => x"00000000", 22876 => x"00000000", 22877 => x"00000000",
    22878 => x"00000000", 22879 => x"00000000", 22880 => x"00000000",
    22881 => x"00000000", 22882 => x"00000000", 22883 => x"00000000",
    22884 => x"00000000", 22885 => x"00000000", 22886 => x"00000000",
    22887 => x"00000000", 22888 => x"00000000", 22889 => x"00000000",
    22890 => x"00000000", 22891 => x"00000000", 22892 => x"00000000",
    22893 => x"00000000", 22894 => x"00000000", 22895 => x"00000000",
    22896 => x"00000000", 22897 => x"00000000", 22898 => x"00000000",
    22899 => x"00000000", 22900 => x"00000000", 22901 => x"00000000",
    22902 => x"00000000", 22903 => x"00000000", 22904 => x"00000000",
    22905 => x"00000000", 22906 => x"00000000", 22907 => x"00000000",
    22908 => x"00000000", 22909 => x"00000000", 22910 => x"00000000",
    22911 => x"00000000", 22912 => x"00000000", 22913 => x"00000000",
    22914 => x"00000000", 22915 => x"00000000", 22916 => x"00000000",
    22917 => x"00000000", 22918 => x"00000000", 22919 => x"00000000",
    22920 => x"00000000", 22921 => x"00000000", 22922 => x"00000000",
    22923 => x"00000000", 22924 => x"00000000", 22925 => x"00000000",
    22926 => x"00000000", 22927 => x"00000000", 22928 => x"00000000",
    22929 => x"00000000", 22930 => x"00000000", 22931 => x"00000000",
    22932 => x"00000000", 22933 => x"00000000", 22934 => x"00000000",
    22935 => x"00000000", 22936 => x"00000000", 22937 => x"00000000",
    22938 => x"00000000", 22939 => x"00000000", 22940 => x"00000000",
    22941 => x"00000000", 22942 => x"00000000", 22943 => x"00000000",
    22944 => x"00000000", 22945 => x"00000000", 22946 => x"00000000",
    22947 => x"00000000", 22948 => x"00000000", 22949 => x"00000000",
    22950 => x"00000000", 22951 => x"00000000", 22952 => x"00000000",
    22953 => x"00000000", 22954 => x"00000000", 22955 => x"00000000",
    22956 => x"00000000", 22957 => x"00000000", 22958 => x"00000000",
    22959 => x"00000000", 22960 => x"00000000", 22961 => x"00000000",
    22962 => x"00000000", 22963 => x"00000000", 22964 => x"00000000",
    22965 => x"00000000", 22966 => x"00000000", 22967 => x"00000000",
    22968 => x"00000000", 22969 => x"00000000", 22970 => x"00000000",
    22971 => x"00000000", 22972 => x"00000000", 22973 => x"00000000",
    22974 => x"00000000", 22975 => x"00000000", 22976 => x"00000000",
    22977 => x"00000000", 22978 => x"00000000", 22979 => x"00000000",
    22980 => x"00000000", 22981 => x"00000000", 22982 => x"00000000",
    22983 => x"00000000", 22984 => x"00000000", 22985 => x"00000000",
    22986 => x"00000000", 22987 => x"00000000", 22988 => x"00000000",
    22989 => x"00000000", 22990 => x"00000000", 22991 => x"00000000",
    22992 => x"00000000", 22993 => x"00000000", 22994 => x"00000000",
    22995 => x"00000000", 22996 => x"00000000", 22997 => x"00000000",
    22998 => x"00000000", 22999 => x"00000000", 23000 => x"00000000",
    23001 => x"00000000", 23002 => x"00000000", 23003 => x"00000000",
    23004 => x"00000000", 23005 => x"00000000", 23006 => x"00000000",
    23007 => x"00000000", 23008 => x"00000000", 23009 => x"00000000",
    23010 => x"00000000", 23011 => x"00000000", 23012 => x"00000000",
    23013 => x"00000000", 23014 => x"00000000", 23015 => x"00000000",
    23016 => x"00000000", 23017 => x"00000000", 23018 => x"00000000",
    23019 => x"00000000", 23020 => x"00000000", 23021 => x"00000000",
    23022 => x"00000000", 23023 => x"00000000", 23024 => x"00000000",
    23025 => x"00000000", 23026 => x"00000000", 23027 => x"00000000",
    23028 => x"00000000", 23029 => x"00000000", 23030 => x"00000000",
    23031 => x"00000000", 23032 => x"00000000", 23033 => x"00000000",
    23034 => x"00000000", 23035 => x"00000000", 23036 => x"00000000",
    23037 => x"00000000", 23038 => x"00000000", 23039 => x"00000000",
    23040 => x"00000000", 23041 => x"00000000", 23042 => x"00000000",
    23043 => x"00000000", 23044 => x"00000000", 23045 => x"00000000",
    23046 => x"00000000", 23047 => x"00000000", 23048 => x"00000000",
    23049 => x"00000000", 23050 => x"00000000", 23051 => x"00000000",
    23052 => x"00000000", 23053 => x"00000000", 23054 => x"00000000",
    23055 => x"00000000", 23056 => x"00000000", 23057 => x"00000000",
    23058 => x"00000000", 23059 => x"00000000", 23060 => x"00000000",
    23061 => x"00000000", 23062 => x"00000000", 23063 => x"00000000",
    23064 => x"00000000", 23065 => x"00000000", 23066 => x"00000000",
    23067 => x"00000000", 23068 => x"00000000", 23069 => x"00000000",
    23070 => x"00000000", 23071 => x"00000000", 23072 => x"00000000",
    23073 => x"00000000", 23074 => x"00000000", 23075 => x"00000000",
    23076 => x"00000000", 23077 => x"00000000", 23078 => x"00000000",
    23079 => x"00000000", 23080 => x"00000000", 23081 => x"00000000",
    23082 => x"00000000", 23083 => x"00000000", 23084 => x"00000000",
    23085 => x"00000000", 23086 => x"00000000", 23087 => x"00000000",
    23088 => x"00000000", 23089 => x"00000000", 23090 => x"00000000",
    23091 => x"00000000", 23092 => x"00000000", 23093 => x"00000000",
    23094 => x"00000000", 23095 => x"00000000", 23096 => x"00000000",
    23097 => x"00000000", 23098 => x"00000000", 23099 => x"00000000",
    23100 => x"00000000", 23101 => x"00000000", 23102 => x"00000000",
    23103 => x"00000000", 23104 => x"00000000", 23105 => x"00000000",
    23106 => x"00000000", 23107 => x"00000000", 23108 => x"00000000",
    23109 => x"00000000", 23110 => x"00000000", 23111 => x"00000000",
    23112 => x"00000000", 23113 => x"00000000", 23114 => x"00000000",
    23115 => x"00000000", 23116 => x"00000000", 23117 => x"00000000",
    23118 => x"00000000", 23119 => x"00000000", 23120 => x"00000000",
    23121 => x"00000000", 23122 => x"00000000", 23123 => x"00000000",
    23124 => x"00000000", 23125 => x"00000000", 23126 => x"00000000",
    23127 => x"00000000", 23128 => x"00000000", 23129 => x"00000000",
    23130 => x"00000000", 23131 => x"00000000", 23132 => x"00000000",
    23133 => x"00000000", 23134 => x"00000000", 23135 => x"00000000",
    23136 => x"00000000", 23137 => x"00000000", 23138 => x"00000000",
    23139 => x"00000000", 23140 => x"00000000", 23141 => x"00000000",
    23142 => x"00000000", 23143 => x"00000000", 23144 => x"00000000",
    23145 => x"00000000", 23146 => x"00000000", 23147 => x"00000000",
    23148 => x"00000000", 23149 => x"00000000", 23150 => x"00000000",
    23151 => x"00000000", 23152 => x"00000000", 23153 => x"00000000",
    23154 => x"00000000", 23155 => x"00000000", 23156 => x"00000000",
    23157 => x"00000000", 23158 => x"00000000", 23159 => x"00000000",
    23160 => x"00000000", 23161 => x"00000000", 23162 => x"00000000",
    23163 => x"00000000", 23164 => x"00000000", 23165 => x"00000000",
    23166 => x"00000000", 23167 => x"00000000", 23168 => x"00000000",
    23169 => x"00000000", 23170 => x"00000000", 23171 => x"00000000",
    23172 => x"00000000", 23173 => x"00000000", 23174 => x"00000000",
    23175 => x"00000000", 23176 => x"00000000", 23177 => x"00000000",
    23178 => x"00000000", 23179 => x"00000000", 23180 => x"00000000",
    23181 => x"00000000", 23182 => x"00000000", 23183 => x"00000000",
    23184 => x"00000000", 23185 => x"00000000", 23186 => x"00000000",
    23187 => x"00000000", 23188 => x"00000000", 23189 => x"00000000",
    23190 => x"00000000", 23191 => x"00000000", 23192 => x"00000000",
    23193 => x"00000000", 23194 => x"00000000", 23195 => x"00000000",
    23196 => x"00000000", 23197 => x"00000000", 23198 => x"00000000",
    23199 => x"00000000", 23200 => x"00000000", 23201 => x"00000000",
    23202 => x"00000000", 23203 => x"00000000", 23204 => x"00000000",
    23205 => x"00000000", 23206 => x"00000000", 23207 => x"00000000",
    23208 => x"00000000", 23209 => x"00000000", 23210 => x"00000000",
    23211 => x"00000000", 23212 => x"00000000", 23213 => x"00000000",
    23214 => x"00000000", 23215 => x"00000000", 23216 => x"00000000",
    23217 => x"00000000", 23218 => x"00000000", 23219 => x"00000000",
    23220 => x"00000000", 23221 => x"00000000", 23222 => x"00000000",
    23223 => x"00000000", 23224 => x"00000000", 23225 => x"00000000",
    23226 => x"00000000", 23227 => x"00000000", 23228 => x"00000000",
    23229 => x"00000000", 23230 => x"00000000", 23231 => x"00000000",
    23232 => x"00000000", 23233 => x"00000000", 23234 => x"00000000",
    23235 => x"00000000", 23236 => x"00000000", 23237 => x"00000000",
    23238 => x"00000000", 23239 => x"00000000", 23240 => x"00000000",
    23241 => x"00000000", 23242 => x"00000000", 23243 => x"00000000",
    23244 => x"00000000", 23245 => x"00000000", 23246 => x"00000000",
    23247 => x"00000000", 23248 => x"00000000", 23249 => x"00000000",
    23250 => x"00000000", 23251 => x"00000000", 23252 => x"00000000",
    23253 => x"00000000", 23254 => x"00000000", 23255 => x"00000000",
    23256 => x"00000000", 23257 => x"00000000", 23258 => x"00000000",
    23259 => x"00000000", 23260 => x"00000000", 23261 => x"00000000",
    23262 => x"00000000", 23263 => x"00000000", 23264 => x"00000000",
    23265 => x"00000000", 23266 => x"00000000", 23267 => x"00000000",
    23268 => x"00000000", 23269 => x"00000000", 23270 => x"00000000",
    23271 => x"00000000", 23272 => x"00000000", 23273 => x"00000000",
    23274 => x"00000000", 23275 => x"00000000", 23276 => x"00000000",
    23277 => x"00000000", 23278 => x"00000000", 23279 => x"00000000",
    23280 => x"00000000", 23281 => x"00000000", 23282 => x"00000000",
    23283 => x"00000000", 23284 => x"00000000", 23285 => x"00000000",
    23286 => x"00000000", 23287 => x"00000000", 23288 => x"00000000",
    23289 => x"00000000", 23290 => x"00000000", 23291 => x"00000000",
    23292 => x"00000000", 23293 => x"00000000", 23294 => x"00000000",
    23295 => x"00000000", 23296 => x"00000000", 23297 => x"00000000",
    23298 => x"00000000", 23299 => x"00000000", 23300 => x"00000000",
    23301 => x"00000000", 23302 => x"00000000", 23303 => x"00000000",
    23304 => x"00000000", 23305 => x"00000000", 23306 => x"00000000",
    23307 => x"00000000", 23308 => x"00000000", 23309 => x"00000000",
    23310 => x"00000000", 23311 => x"00000000", 23312 => x"00000000",
    23313 => x"00000000", 23314 => x"00000000", 23315 => x"00000000",
    23316 => x"00000000", 23317 => x"00000000", 23318 => x"00000000",
    23319 => x"00000000", 23320 => x"00000000", 23321 => x"00000000",
    23322 => x"00000000", 23323 => x"00000000", 23324 => x"00000000",
    23325 => x"00000000", 23326 => x"00000000", 23327 => x"00000000",
    23328 => x"00000000", 23329 => x"00000000", 23330 => x"00000000",
    23331 => x"00000000", 23332 => x"00000000", 23333 => x"00000000",
    23334 => x"00000000", 23335 => x"00000000", 23336 => x"00000000",
    23337 => x"00000000", 23338 => x"00000000", 23339 => x"00000000",
    23340 => x"00000000", 23341 => x"00000000", 23342 => x"00000000",
    23343 => x"00000000", 23344 => x"00000000", 23345 => x"00000000",
    23346 => x"00000000", 23347 => x"00000000", 23348 => x"00000000",
    23349 => x"00000000", 23350 => x"00000000", 23351 => x"00000000",
    23352 => x"00000000", 23353 => x"00000000", 23354 => x"00000000",
    23355 => x"00000000", 23356 => x"00000000", 23357 => x"00000000",
    23358 => x"00000000", 23359 => x"00000000", 23360 => x"00000000",
    23361 => x"00000000", 23362 => x"00000000", 23363 => x"00000000",
    23364 => x"00000000", 23365 => x"00000000", 23366 => x"00000000",
    23367 => x"00000000", 23368 => x"00000000", 23369 => x"00000000",
    23370 => x"00000000", 23371 => x"00000000", 23372 => x"00000000",
    23373 => x"00000000", 23374 => x"00000000", 23375 => x"00000000",
    23376 => x"00000000", 23377 => x"00000000", 23378 => x"00000000",
    23379 => x"00000000", 23380 => x"00000000", 23381 => x"00000000",
    23382 => x"00000000", 23383 => x"00000000", 23384 => x"00000000",
    23385 => x"00000000", 23386 => x"00000000", 23387 => x"00000000",
    23388 => x"00000000", 23389 => x"00000000", 23390 => x"00000000",
    23391 => x"00000000", 23392 => x"00000000", 23393 => x"00000000",
    23394 => x"00000000", 23395 => x"00000000", 23396 => x"00000000",
    23397 => x"00000000", 23398 => x"00000000", 23399 => x"00000000",
    23400 => x"00000000", 23401 => x"00000000", 23402 => x"00000000",
    23403 => x"00000000", 23404 => x"00000000", 23405 => x"00000000",
    23406 => x"00000000", 23407 => x"00000000", 23408 => x"00000000",
    23409 => x"00000000", 23410 => x"00000000", 23411 => x"00000000",
    23412 => x"00000000", 23413 => x"00000000", 23414 => x"00000000",
    23415 => x"00000000", 23416 => x"00000000", 23417 => x"00000000",
    23418 => x"00000000", 23419 => x"00000000", 23420 => x"00000000",
    23421 => x"00000000", 23422 => x"00000000", 23423 => x"00000000",
    23424 => x"00000000", 23425 => x"00000000", 23426 => x"00000000",
    23427 => x"00000000", 23428 => x"00000000", 23429 => x"00000000",
    23430 => x"00000000", 23431 => x"00000000", 23432 => x"00000000",
    23433 => x"00000000", 23434 => x"00000000", 23435 => x"00000000",
    23436 => x"00000000", 23437 => x"00000000", 23438 => x"00000000",
    23439 => x"00000000", 23440 => x"00000000", 23441 => x"00000000",
    23442 => x"00000000", 23443 => x"00000000", 23444 => x"00000000",
    23445 => x"00000000", 23446 => x"00000000", 23447 => x"00000000",
    23448 => x"00000000", 23449 => x"00000000", 23450 => x"00000000",
    23451 => x"00000000", 23452 => x"00000000", 23453 => x"00000000",
    23454 => x"00000000", 23455 => x"00000000", 23456 => x"00000000",
    23457 => x"00000000", 23458 => x"00000000", 23459 => x"00000000",
    23460 => x"00000000", 23461 => x"00000000", 23462 => x"00000000",
    23463 => x"00000000", 23464 => x"00000000", 23465 => x"00000000",
    23466 => x"00000000", 23467 => x"00000000", 23468 => x"00000000",
    23469 => x"00000000", 23470 => x"00000000", 23471 => x"00000000",
    23472 => x"00000000", 23473 => x"00000000", 23474 => x"00000000",
    23475 => x"00000000", 23476 => x"00000000", 23477 => x"00000000",
    23478 => x"00000000", 23479 => x"00000000", 23480 => x"00000000",
    23481 => x"00000000", 23482 => x"00000000", 23483 => x"00000000",
    23484 => x"00000000", 23485 => x"00000000", 23486 => x"00000000",
    23487 => x"00000000", 23488 => x"00000000", 23489 => x"00000000",
    23490 => x"00000000", 23491 => x"00000000", 23492 => x"00000000",
    23493 => x"00000000", 23494 => x"00000000", 23495 => x"00000000",
    23496 => x"00000000", 23497 => x"00000000", 23498 => x"00000000",
    23499 => x"00000000", 23500 => x"00000000", 23501 => x"00000000",
    23502 => x"00000000", 23503 => x"00000000", 23504 => x"00000000",
    23505 => x"00000000", 23506 => x"00000000", 23507 => x"00000000",
    23508 => x"00000000", 23509 => x"00000000", 23510 => x"00000000",
    23511 => x"00000000", 23512 => x"00000000", 23513 => x"00000000",
    23514 => x"00000000", 23515 => x"00000000", 23516 => x"00000000",
    23517 => x"00000000", 23518 => x"00000000", 23519 => x"00000000",
    23520 => x"00000000", 23521 => x"00000000", 23522 => x"00000000",
    23523 => x"00000000", 23524 => x"00000000", 23525 => x"00000000",
    23526 => x"00000000", 23527 => x"00000000", 23528 => x"00000000",
    23529 => x"00000000", 23530 => x"00000000", 23531 => x"00000000",
    23532 => x"00000000", 23533 => x"00000000", 23534 => x"00000000",
    23535 => x"00000000", 23536 => x"00000000", 23537 => x"00000000",
    23538 => x"00000000", 23539 => x"00000000", 23540 => x"00000000",
    23541 => x"00000000", 23542 => x"00000000", 23543 => x"00000000",
    23544 => x"00000000", 23545 => x"00000000", 23546 => x"00000000",
    23547 => x"00000000", 23548 => x"00000000", 23549 => x"00000000",
    23550 => x"00000000", 23551 => x"00000000", 23552 => x"00000000",
    23553 => x"00000000", 23554 => x"00000000", 23555 => x"00000000",
    23556 => x"00000000", 23557 => x"00000000", 23558 => x"00000000",
    23559 => x"00000000", 23560 => x"00000000", 23561 => x"00000000",
    23562 => x"00000000", 23563 => x"00000000", 23564 => x"00000000",
    23565 => x"00000000", 23566 => x"00000000", 23567 => x"00000000",
    23568 => x"00000000", 23569 => x"00000000", 23570 => x"00000000",
    23571 => x"00000000", 23572 => x"00000000", 23573 => x"00000000",
    23574 => x"00000000", 23575 => x"00000000", 23576 => x"00000000",
    23577 => x"00000000", 23578 => x"00000000", 23579 => x"00000000",
    23580 => x"00000000", 23581 => x"00000000", 23582 => x"00000000",
    23583 => x"00000000", 23584 => x"00000000", 23585 => x"00000000",
    23586 => x"00000000", 23587 => x"00000000", 23588 => x"00000000",
    23589 => x"00000000", 23590 => x"00000000", 23591 => x"00000000",
    23592 => x"00000000", 23593 => x"00000000", 23594 => x"00000000",
    23595 => x"00000000", 23596 => x"00000000", 23597 => x"00000000",
    23598 => x"00000000", 23599 => x"00000000", 23600 => x"00000000",
    23601 => x"00000000", 23602 => x"00000000", 23603 => x"00000000",
    23604 => x"00000000", 23605 => x"00000000", 23606 => x"00000000",
    23607 => x"00000000", 23608 => x"00000000", 23609 => x"00000000",
    23610 => x"00000000", 23611 => x"00000000", 23612 => x"00000000",
    23613 => x"00000000", 23614 => x"00000000", 23615 => x"00000000",
    23616 => x"00000000", 23617 => x"00000000", 23618 => x"00000000",
    23619 => x"00000000", 23620 => x"00000000", 23621 => x"00000000",
    23622 => x"00000000", 23623 => x"00000000", 23624 => x"00000000",
    23625 => x"00000000", 23626 => x"00000000", 23627 => x"00000000",
    23628 => x"00000000", 23629 => x"00000000", 23630 => x"00000000",
    23631 => x"00000000", 23632 => x"00000000", 23633 => x"00000000",
    23634 => x"00000000", 23635 => x"00000000", 23636 => x"00000000",
    23637 => x"00000000", 23638 => x"00000000", 23639 => x"00000000",
    23640 => x"00000000", 23641 => x"00000000", 23642 => x"00000000",
    23643 => x"00000000", 23644 => x"00000000", 23645 => x"00000000",
    23646 => x"00000000", 23647 => x"00000000", 23648 => x"00000000",
    23649 => x"00000000", 23650 => x"00000000", 23651 => x"00000000",
    23652 => x"00000000", 23653 => x"00000000", 23654 => x"00000000",
    23655 => x"00000000", 23656 => x"00000000", 23657 => x"00000000",
    23658 => x"00000000", 23659 => x"00000000", 23660 => x"00000000",
    23661 => x"00000000", 23662 => x"00000000", 23663 => x"00000000",
    23664 => x"00000000", 23665 => x"00000000", 23666 => x"00000000",
    23667 => x"00000000", 23668 => x"00000000", 23669 => x"00000000",
    23670 => x"00000000", 23671 => x"00000000", 23672 => x"00000000",
    23673 => x"00000000", 23674 => x"00000000", 23675 => x"00000000",
    23676 => x"00000000", 23677 => x"00000000", 23678 => x"00000000",
    23679 => x"00000000", 23680 => x"00000000", 23681 => x"00000000",
    23682 => x"00000000", 23683 => x"00000000", 23684 => x"00000000",
    23685 => x"00000000", 23686 => x"00000000", 23687 => x"00000000",
    23688 => x"00000000", 23689 => x"00000000", 23690 => x"00000000",
    23691 => x"00000000", 23692 => x"00000000", 23693 => x"00000000",
    23694 => x"00000000", 23695 => x"00000000", 23696 => x"00000000",
    23697 => x"00000000", 23698 => x"00000000", 23699 => x"00000000",
    23700 => x"00000000", 23701 => x"00000000", 23702 => x"00000000",
    23703 => x"00000000", 23704 => x"00000000", 23705 => x"00000000",
    23706 => x"00000000", 23707 => x"00000000", 23708 => x"00000000",
    23709 => x"00000000", 23710 => x"00000000", 23711 => x"00000000",
    23712 => x"00000000", 23713 => x"00000000", 23714 => x"00000000",
    23715 => x"00000000", 23716 => x"00000000", 23717 => x"00000000",
    23718 => x"00000000", 23719 => x"00000000", 23720 => x"00000000",
    23721 => x"00000000", 23722 => x"00000000", 23723 => x"00000000",
    23724 => x"00000000", 23725 => x"00000000", 23726 => x"00000000",
    23727 => x"00000000", 23728 => x"00000000", 23729 => x"00000000",
    23730 => x"00000000", 23731 => x"00000000", 23732 => x"00000000",
    23733 => x"00000000", 23734 => x"00000000", 23735 => x"00000000",
    23736 => x"00000000", 23737 => x"00000000", 23738 => x"00000000",
    23739 => x"00000000", 23740 => x"00000000", 23741 => x"00000000",
    23742 => x"00000000", 23743 => x"00000000", 23744 => x"00000000",
    23745 => x"00000000", 23746 => x"00000000", 23747 => x"00000000",
    23748 => x"00000000", 23749 => x"00000000", 23750 => x"00000000",
    23751 => x"00000000", 23752 => x"00000000", 23753 => x"00000000",
    23754 => x"00000000", 23755 => x"00000000", 23756 => x"00000000",
    23757 => x"00000000", 23758 => x"00000000", 23759 => x"00000000",
    23760 => x"00000000", 23761 => x"00000000", 23762 => x"00000000",
    23763 => x"00000000", 23764 => x"00000000", 23765 => x"00000000",
    23766 => x"00000000", 23767 => x"00000000", 23768 => x"00000000",
    23769 => x"00000000", 23770 => x"00000000", 23771 => x"00000000",
    23772 => x"00000000", 23773 => x"00000000", 23774 => x"00000000",
    23775 => x"00000000", 23776 => x"00000000", 23777 => x"00000000",
    23778 => x"00000000", 23779 => x"00000000", 23780 => x"00000000",
    23781 => x"00000000", 23782 => x"00000000", 23783 => x"00000000",
    23784 => x"00000000", 23785 => x"00000000", 23786 => x"00000000",
    23787 => x"00000000", 23788 => x"00000000", 23789 => x"00000000",
    23790 => x"00000000", 23791 => x"00000000", 23792 => x"00000000",
    23793 => x"00000000", 23794 => x"00000000", 23795 => x"00000000",
    23796 => x"00000000", 23797 => x"00000000", 23798 => x"00000000",
    23799 => x"00000000", 23800 => x"00000000", 23801 => x"00000000",
    23802 => x"00000000", 23803 => x"00000000", 23804 => x"00000000",
    23805 => x"00000000", 23806 => x"00000000", 23807 => x"00000000",
    23808 => x"00000000", 23809 => x"00000000", 23810 => x"00000000",
    23811 => x"00000000", 23812 => x"00000000", 23813 => x"00000000",
    23814 => x"00000000", 23815 => x"00000000", 23816 => x"00000000",
    23817 => x"00000000", 23818 => x"00000000", 23819 => x"00000000",
    23820 => x"00000000", 23821 => x"00000000", 23822 => x"00000000",
    23823 => x"00000000", 23824 => x"00000000", 23825 => x"00000000",
    23826 => x"00000000", 23827 => x"00000000", 23828 => x"00000000",
    23829 => x"00000000", 23830 => x"00000000", 23831 => x"00000000",
    23832 => x"00000000", 23833 => x"00000000", 23834 => x"00000000",
    23835 => x"00000000", 23836 => x"00000000", 23837 => x"00000000",
    23838 => x"00000000", 23839 => x"00000000", 23840 => x"00000000",
    23841 => x"00000000", 23842 => x"00000000", 23843 => x"00000000",
    23844 => x"00000000", 23845 => x"00000000", 23846 => x"00000000",
    23847 => x"00000000", 23848 => x"00000000", 23849 => x"00000000",
    23850 => x"00000000", 23851 => x"00000000", 23852 => x"00000000",
    23853 => x"00000000", 23854 => x"00000000", 23855 => x"00000000",
    23856 => x"00000000", 23857 => x"00000000", 23858 => x"00000000",
    23859 => x"00000000", 23860 => x"00000000", 23861 => x"00000000",
    23862 => x"00000000", 23863 => x"00000000", 23864 => x"00000000",
    23865 => x"00000000", 23866 => x"00000000", 23867 => x"00000000",
    23868 => x"00000000", 23869 => x"00000000", 23870 => x"00000000",
    23871 => x"00000000", 23872 => x"00000000", 23873 => x"00000000",
    23874 => x"00000000", 23875 => x"00000000", 23876 => x"00000000",
    23877 => x"00000000", 23878 => x"00000000", 23879 => x"00000000",
    23880 => x"00000000", 23881 => x"00000000", 23882 => x"00000000",
    23883 => x"00000000", 23884 => x"00000000", 23885 => x"00000000",
    23886 => x"00000000", 23887 => x"00000000", 23888 => x"00000000",
    23889 => x"00000000", 23890 => x"00000000", 23891 => x"00000000",
    23892 => x"00000000", 23893 => x"00000000", 23894 => x"00000000",
    23895 => x"00000000", 23896 => x"00000000", 23897 => x"00000000",
    23898 => x"00000000", 23899 => x"00000000", 23900 => x"00000000",
    23901 => x"00000000", 23902 => x"00000000", 23903 => x"00000000",
    23904 => x"00000000", 23905 => x"00000000", 23906 => x"00000000",
    23907 => x"00000000", 23908 => x"00000000", 23909 => x"00000000",
    23910 => x"00000000", 23911 => x"00000000", 23912 => x"00000000",
    23913 => x"00000000", 23914 => x"00000000", 23915 => x"00000000",
    23916 => x"00000000", 23917 => x"00000000", 23918 => x"00000000",
    23919 => x"00000000", 23920 => x"00000000", 23921 => x"00000000",
    23922 => x"00000000", 23923 => x"00000000", 23924 => x"00000000",
    23925 => x"00000000", 23926 => x"00000000", 23927 => x"00000000",
    23928 => x"00000000", 23929 => x"00000000", 23930 => x"00000000",
    23931 => x"00000000", 23932 => x"00000000", 23933 => x"00000000",
    23934 => x"00000000", 23935 => x"00000000", 23936 => x"00000000",
    23937 => x"00000000", 23938 => x"00000000", 23939 => x"00000000",
    23940 => x"00000000", 23941 => x"00000000", 23942 => x"00000000",
    23943 => x"00000000", 23944 => x"00000000", 23945 => x"00000000",
    23946 => x"00000000", 23947 => x"00000000", 23948 => x"00000000",
    23949 => x"00000000", 23950 => x"00000000", 23951 => x"00000000",
    23952 => x"00000000", 23953 => x"00000000", 23954 => x"00000000",
    23955 => x"00000000", 23956 => x"00000000", 23957 => x"00000000",
    23958 => x"00000000", 23959 => x"00000000", 23960 => x"00000000",
    23961 => x"00000000", 23962 => x"00000000", 23963 => x"00000000",
    23964 => x"00000000", 23965 => x"00000000", 23966 => x"00000000",
    23967 => x"00000000", 23968 => x"00000000", 23969 => x"00000000",
    23970 => x"00000000", 23971 => x"00000000", 23972 => x"00000000",
    23973 => x"00000000", 23974 => x"00000000", 23975 => x"00000000",
    23976 => x"00000000", 23977 => x"00000000", 23978 => x"00000000",
    23979 => x"00000000", 23980 => x"00000000", 23981 => x"00000000",
    23982 => x"00000000", 23983 => x"00000000", 23984 => x"00000000",
    23985 => x"00000000", 23986 => x"00000000", 23987 => x"00000000",
    23988 => x"00000000", 23989 => x"00000000", 23990 => x"00000000",
    23991 => x"00000000", 23992 => x"00000000", 23993 => x"00000000",
    23994 => x"00000000", 23995 => x"00000000", 23996 => x"00000000",
    23997 => x"00000000", 23998 => x"00000000", 23999 => x"00000000",
    24000 => x"00000000", 24001 => x"00000000", 24002 => x"00000000",
    24003 => x"00000000", 24004 => x"00000000", 24005 => x"00000000",
    24006 => x"00000000", 24007 => x"00000000", 24008 => x"00000000",
    24009 => x"00000000", 24010 => x"00000000", 24011 => x"00000000",
    24012 => x"00000000", 24013 => x"00000000", 24014 => x"00000000",
    24015 => x"00000000", 24016 => x"00000000", 24017 => x"00000000",
    24018 => x"00000000", 24019 => x"00000000", 24020 => x"00000000",
    24021 => x"00000000", 24022 => x"00000000", 24023 => x"00000000",
    24024 => x"00000000", 24025 => x"00000000", 24026 => x"00000000",
    24027 => x"00000000", 24028 => x"00000000", 24029 => x"00000000",
    24030 => x"00000000", 24031 => x"00000000", 24032 => x"00000000",
    24033 => x"00000000", 24034 => x"00000000", 24035 => x"00000000",
    24036 => x"00000000", 24037 => x"00000000", 24038 => x"00000000",
    24039 => x"00000000", 24040 => x"00000000", 24041 => x"00000000",
    24042 => x"00000000", 24043 => x"00000000", 24044 => x"00000000",
    24045 => x"00000000", 24046 => x"00000000", 24047 => x"00000000",
    24048 => x"00000000", 24049 => x"00000000", 24050 => x"00000000",
    24051 => x"00000000", 24052 => x"00000000", 24053 => x"00000000",
    24054 => x"00000000", 24055 => x"00000000", 24056 => x"00000000",
    24057 => x"00000000", 24058 => x"00000000", 24059 => x"00000000",
    24060 => x"00000000", 24061 => x"00000000", 24062 => x"00000000",
    24063 => x"00000000", 24064 => x"00000000", 24065 => x"00000000",
    24066 => x"00000000", 24067 => x"00000000", 24068 => x"00000000",
    24069 => x"00000000", 24070 => x"00000000", 24071 => x"00000000",
    24072 => x"00000000", 24073 => x"00000000", 24074 => x"00000000",
    24075 => x"00000000", 24076 => x"00000000", 24077 => x"00000000",
    24078 => x"00000000", 24079 => x"00000000", 24080 => x"00000000",
    24081 => x"00000000", 24082 => x"00000000", 24083 => x"00000000",
    24084 => x"00000000", 24085 => x"00000000", 24086 => x"00000000",
    24087 => x"00000000", 24088 => x"00000000", 24089 => x"00000000",
    24090 => x"00000000", 24091 => x"00000000", 24092 => x"00000000",
    24093 => x"00000000", 24094 => x"00000000", 24095 => x"00000000",
    24096 => x"00000000", 24097 => x"00000000", 24098 => x"00000000",
    24099 => x"00000000", 24100 => x"00000000", 24101 => x"00000000",
    24102 => x"00000000", 24103 => x"00000000", 24104 => x"00000000",
    24105 => x"00000000", 24106 => x"00000000", 24107 => x"00000000",
    24108 => x"00000000", 24109 => x"00000000", 24110 => x"00000000",
    24111 => x"00000000", 24112 => x"00000000", 24113 => x"00000000",
    24114 => x"00000000", 24115 => x"00000000", 24116 => x"00000000",
    24117 => x"00000000", 24118 => x"00000000", 24119 => x"00000000",
    24120 => x"00000000", 24121 => x"00000000", 24122 => x"00000000",
    24123 => x"00000000", 24124 => x"00000000", 24125 => x"00000000",
    24126 => x"00000000", 24127 => x"00000000", 24128 => x"00000000",
    24129 => x"00000000", 24130 => x"00000000", 24131 => x"00000000",
    24132 => x"00000000", 24133 => x"00000000", 24134 => x"00000000",
    24135 => x"00000000", 24136 => x"00000000", 24137 => x"00000000",
    24138 => x"00000000", 24139 => x"00000000", 24140 => x"00000000",
    24141 => x"00000000", 24142 => x"00000000", 24143 => x"00000000",
    24144 => x"00000000", 24145 => x"00000000", 24146 => x"00000000",
    24147 => x"00000000", 24148 => x"00000000", 24149 => x"00000000",
    24150 => x"00000000", 24151 => x"00000000", 24152 => x"00000000",
    24153 => x"00000000", 24154 => x"00000000", 24155 => x"00000000",
    24156 => x"00000000", 24157 => x"00000000", 24158 => x"00000000",
    24159 => x"00000000", 24160 => x"00000000", 24161 => x"00000000",
    24162 => x"00000000", 24163 => x"00000000", 24164 => x"00000000",
    24165 => x"00000000", 24166 => x"00000000", 24167 => x"00000000",
    24168 => x"00000000", 24169 => x"00000000", 24170 => x"00000000",
    24171 => x"00000000", 24172 => x"00000000", 24173 => x"00000000",
    24174 => x"00000000", 24175 => x"00000000", 24176 => x"00000000",
    24177 => x"00000000", 24178 => x"00000000", 24179 => x"00000000",
    24180 => x"00000000", 24181 => x"00000000", 24182 => x"00000000",
    24183 => x"00000000", 24184 => x"00000000", 24185 => x"00000000",
    24186 => x"00000000", 24187 => x"00000000", 24188 => x"00000000",
    24189 => x"00000000", 24190 => x"00000000", 24191 => x"00000000",
    24192 => x"00000000", 24193 => x"00000000", 24194 => x"00000000",
    24195 => x"00000000", 24196 => x"00000000", 24197 => x"00000000",
    24198 => x"00000000", 24199 => x"00000000", 24200 => x"00000000",
    24201 => x"00000000", 24202 => x"00000000", 24203 => x"00000000",
    24204 => x"00000000", 24205 => x"00000000", 24206 => x"00000000",
    24207 => x"00000000", 24208 => x"00000000", 24209 => x"00000000",
    24210 => x"00000000", 24211 => x"00000000", 24212 => x"00000000",
    24213 => x"00000000", 24214 => x"00000000", 24215 => x"00000000",
    24216 => x"00000000", 24217 => x"00000000", 24218 => x"00000000",
    24219 => x"00000000", 24220 => x"00000000", 24221 => x"00000000",
    24222 => x"00000000", 24223 => x"00000000", 24224 => x"00000000",
    24225 => x"00000000", 24226 => x"00000000", 24227 => x"00000000",
    24228 => x"00000000", 24229 => x"00000000", 24230 => x"00000000",
    24231 => x"00000000", 24232 => x"00000000", 24233 => x"00000000",
    24234 => x"00000000", 24235 => x"00000000", 24236 => x"00000000",
    24237 => x"00000000", 24238 => x"00000000", 24239 => x"00000000",
    24240 => x"00000000", 24241 => x"00000000", 24242 => x"00000000",
    24243 => x"00000000", 24244 => x"00000000", 24245 => x"00000000",
    24246 => x"00000000", 24247 => x"00000000", 24248 => x"00000000",
    24249 => x"00000000", 24250 => x"00000000", 24251 => x"00000000",
    24252 => x"00000000", 24253 => x"00000000", 24254 => x"00000000",
    24255 => x"00000000", 24256 => x"00000000", 24257 => x"00000000",
    24258 => x"00000000", 24259 => x"00000000", 24260 => x"00000000",
    24261 => x"00000000", 24262 => x"00000000", 24263 => x"00000000",
    24264 => x"00000000", 24265 => x"00000000", 24266 => x"00000000",
    24267 => x"00000000", 24268 => x"00000000", 24269 => x"00000000",
    24270 => x"00000000", 24271 => x"00000000", 24272 => x"00000000",
    24273 => x"00000000", 24274 => x"00000000", 24275 => x"00000000",
    24276 => x"00000000", 24277 => x"00000000", 24278 => x"00000000",
    24279 => x"00000000", 24280 => x"00000000", 24281 => x"00000000",
    24282 => x"00000000", 24283 => x"00000000", 24284 => x"00000000",
    24285 => x"00000000", 24286 => x"00000000", 24287 => x"00000000",
    24288 => x"00000000", 24289 => x"00000000", 24290 => x"00000000",
    24291 => x"00000000", 24292 => x"00000000", 24293 => x"00000000",
    24294 => x"00000000", 24295 => x"00000000", 24296 => x"00000000",
    24297 => x"00000000", 24298 => x"00000000", 24299 => x"00000000",
    24300 => x"00000000", 24301 => x"00000000", 24302 => x"00000000",
    24303 => x"00000000", 24304 => x"00000000", 24305 => x"00000000",
    24306 => x"00000000", 24307 => x"00000000", 24308 => x"00000000",
    24309 => x"00000000", 24310 => x"00000000", 24311 => x"00000000",
    24312 => x"00000000", 24313 => x"00000000", 24314 => x"00000000",
    24315 => x"00000000", 24316 => x"00000000", 24317 => x"00000000",
    24318 => x"00000000", 24319 => x"00000000", 24320 => x"00000000",
    24321 => x"00000000", 24322 => x"00000000", 24323 => x"00000000",
    24324 => x"00000000", 24325 => x"00000000", 24326 => x"00000000",
    24327 => x"00000000", 24328 => x"00000000", 24329 => x"00000000",
    24330 => x"00000000", 24331 => x"00000000", 24332 => x"00000000",
    24333 => x"00000000", 24334 => x"00000000", 24335 => x"00000000",
    24336 => x"00000000", 24337 => x"00000000", 24338 => x"00000000",
    24339 => x"00000000", 24340 => x"00000000", 24341 => x"00000000",
    24342 => x"00000000", 24343 => x"00000000", 24344 => x"00000000",
    24345 => x"00000000", 24346 => x"00000000", 24347 => x"00000000",
    24348 => x"00000000", 24349 => x"00000000", 24350 => x"00000000",
    24351 => x"00000000", 24352 => x"00000000", 24353 => x"00000000",
    24354 => x"00000000", 24355 => x"00000000", 24356 => x"00000000",
    24357 => x"00000000", 24358 => x"00000000", 24359 => x"00000000",
    24360 => x"00000000", 24361 => x"00000000", 24362 => x"00000000",
    24363 => x"00000000", 24364 => x"00000000", 24365 => x"00000000",
    24366 => x"00000000", 24367 => x"00000000", 24368 => x"00000000",
    24369 => x"00000000", 24370 => x"00000000", 24371 => x"00000000",
    24372 => x"00000000", 24373 => x"00000000", 24374 => x"00000000",
    24375 => x"00000000", 24376 => x"00000000", 24377 => x"00000000",
    24378 => x"00000000", 24379 => x"00000000", 24380 => x"00000000",
    24381 => x"00000000", 24382 => x"00000000", 24383 => x"00000000",
    24384 => x"00000000", 24385 => x"00000000", 24386 => x"00000000",
    24387 => x"00000000", 24388 => x"00000000", 24389 => x"00000000",
    24390 => x"00000000", 24391 => x"00000000", 24392 => x"00000000",
    24393 => x"00000000", 24394 => x"00000000", 24395 => x"00000000",
    24396 => x"00000000", 24397 => x"00000000", 24398 => x"00000000",
    24399 => x"00000000", 24400 => x"00000000", 24401 => x"00000000",
    24402 => x"00000000", 24403 => x"00000000", 24404 => x"00000000",
    24405 => x"00000000", 24406 => x"00000000", 24407 => x"00000000",
    24408 => x"00000000", 24409 => x"00000000", 24410 => x"00000000",
    24411 => x"00000000", 24412 => x"00000000", 24413 => x"00000000",
    24414 => x"00000000", 24415 => x"00000000", 24416 => x"00000000",
    24417 => x"00000000", 24418 => x"00000000", 24419 => x"00000000",
    24420 => x"00000000", 24421 => x"00000000", 24422 => x"00000000",
    24423 => x"00000000", 24424 => x"00000000", 24425 => x"00000000",
    24426 => x"00000000", 24427 => x"00000000", 24428 => x"00000000",
    24429 => x"00000000", 24430 => x"00000000", 24431 => x"00000000",
    24432 => x"00000000", 24433 => x"00000000", 24434 => x"00000000",
    24435 => x"00000000", 24436 => x"00000000", 24437 => x"00000000",
    24438 => x"00000000", 24439 => x"00000000", 24440 => x"00000000",
    24441 => x"00000000", 24442 => x"00000000", 24443 => x"00000000",
    24444 => x"00000000", 24445 => x"00000000", 24446 => x"00000000",
    24447 => x"00000000", 24448 => x"00000000", 24449 => x"00000000",
    24450 => x"00000000", 24451 => x"00000000", 24452 => x"00000000",
    24453 => x"00000000", 24454 => x"00000000", 24455 => x"00000000",
    24456 => x"00000000", 24457 => x"00000000", 24458 => x"00000000",
    24459 => x"00000000", 24460 => x"00000000", 24461 => x"00000000",
    24462 => x"00000000", 24463 => x"00000000", 24464 => x"00000000",
    24465 => x"00000000", 24466 => x"00000000", 24467 => x"00000000",
    24468 => x"00000000", 24469 => x"00000000", 24470 => x"00000000",
    24471 => x"00000000", 24472 => x"00000000", 24473 => x"00000000",
    24474 => x"00000000", 24475 => x"00000000", 24476 => x"00000000",
    24477 => x"00000000", 24478 => x"00000000", 24479 => x"00000000",
    24480 => x"00000000", 24481 => x"00000000", 24482 => x"00000000",
    24483 => x"00000000", 24484 => x"00000000", 24485 => x"00000000",
    24486 => x"00000000", 24487 => x"00000000", 24488 => x"00000000",
    24489 => x"00000000", 24490 => x"00000000", 24491 => x"00000000",
    24492 => x"00000000", 24493 => x"00000000", 24494 => x"00000000",
    24495 => x"00000000", 24496 => x"00000000", 24497 => x"00000000",
    24498 => x"00000000", 24499 => x"00000000", 24500 => x"00000000",
    24501 => x"00000000", 24502 => x"00000000", 24503 => x"00000000",
    24504 => x"00000000", 24505 => x"00000000", 24506 => x"00000000",
    24507 => x"00000000", 24508 => x"00000000", 24509 => x"00000000",
    24510 => x"00000000", 24511 => x"00000000", 24512 => x"00000000",
    24513 => x"00000000", 24514 => x"00000000", 24515 => x"00000000",
    24516 => x"00000000", 24517 => x"00000000", 24518 => x"00000000",
    24519 => x"00000000", 24520 => x"00000000", 24521 => x"00000000",
    24522 => x"00000000", 24523 => x"00000000", 24524 => x"00000000",
    24525 => x"00000000", 24526 => x"00000000", 24527 => x"00000000",
    24528 => x"00000000", 24529 => x"00000000", 24530 => x"00000000",
    24531 => x"00000000", 24532 => x"00000000", 24533 => x"00000000",
    24534 => x"00000000", 24535 => x"00000000", 24536 => x"00000000",
    24537 => x"00000000", 24538 => x"00000000", 24539 => x"00000000",
    24540 => x"00000000", 24541 => x"00000000", 24542 => x"00000000",
    24543 => x"00000000", 24544 => x"00000000", 24545 => x"00000000",
    24546 => x"00000000", 24547 => x"00000000", 24548 => x"00000000",
    24549 => x"00000000", 24550 => x"00000000", 24551 => x"00000000",
    24552 => x"00000000", 24553 => x"00000000", 24554 => x"00000000",
    24555 => x"00000000", 24556 => x"00000000", 24557 => x"00000000",
    24558 => x"00000000", 24559 => x"00000000", 24560 => x"00000000",
    24561 => x"00000000", 24562 => x"00000000", 24563 => x"00000000",
    24564 => x"00000000", 24565 => x"00000000", 24566 => x"00000000",
    24567 => x"00000000", 24568 => x"00000000", 24569 => x"00000000",
    24570 => x"00000000", 24571 => x"00000000", 24572 => x"00000000",
    24573 => x"00000000", 24574 => x"00000000", 24575 => x"00000000",
    24576 => x"00000000", 24577 => x"00000000", 24578 => x"00000000",
    24579 => x"00000000", 24580 => x"00000000", 24581 => x"00000000",
    24582 => x"00000000", 24583 => x"00000000", 24584 => x"00000000",
    24585 => x"00000000", 24586 => x"00000000", 24587 => x"00000000",
    24588 => x"00000000", 24589 => x"00000000", 24590 => x"00000000",
    24591 => x"00000000", 24592 => x"00000000", 24593 => x"00000000",
    24594 => x"00000000", 24595 => x"00000000", 24596 => x"00000000",
    24597 => x"00000000", 24598 => x"00000000", 24599 => x"00000000",
    24600 => x"00000000", 24601 => x"00000000", 24602 => x"00000000",
    24603 => x"00000000", 24604 => x"00000000", 24605 => x"00000000",
    24606 => x"00000000", 24607 => x"00000000", 24608 => x"00000000",
    24609 => x"00000000", 24610 => x"00000000", 24611 => x"00000000",
    24612 => x"00000000", 24613 => x"00000000", 24614 => x"00000000",
    24615 => x"00000000", 24616 => x"00000000", 24617 => x"00000000",
    24618 => x"00000000", 24619 => x"00000000", 24620 => x"00000000",
    24621 => x"00000000", 24622 => x"00000000", 24623 => x"00000000",
    24624 => x"00000000", 24625 => x"00000000", 24626 => x"00000000",
    24627 => x"00000000", 24628 => x"00000000", 24629 => x"00000000",
    24630 => x"00000000", 24631 => x"00000000", 24632 => x"00000000",
    24633 => x"00000000", 24634 => x"00000000", 24635 => x"00000000",
    24636 => x"00000000", 24637 => x"00000000", 24638 => x"00000000",
    24639 => x"00000000", 24640 => x"00000000", 24641 => x"00000000",
    24642 => x"00000000", 24643 => x"00000000", 24644 => x"00000000",
    24645 => x"00000000", 24646 => x"00000000", 24647 => x"00000000",
    24648 => x"00000000", 24649 => x"00000000", 24650 => x"00000000",
    24651 => x"00000000", 24652 => x"00000000", 24653 => x"00000000",
    24654 => x"00000000", 24655 => x"00000000", 24656 => x"00000000",
    24657 => x"00000000", 24658 => x"00000000", 24659 => x"00000000",
    24660 => x"00000000", 24661 => x"00000000", 24662 => x"00000000",
    24663 => x"00000000", 24664 => x"00000000", 24665 => x"00000000",
    24666 => x"00000000", 24667 => x"00000000", 24668 => x"00000000",
    24669 => x"00000000", 24670 => x"00000000", 24671 => x"00000000",
    24672 => x"00000000", 24673 => x"00000000", 24674 => x"00000000",
    24675 => x"00000000", 24676 => x"00000000", 24677 => x"00000000",
    24678 => x"00000000", 24679 => x"00000000", 24680 => x"00000000",
    24681 => x"00000000", 24682 => x"00000000", 24683 => x"00000000",
    24684 => x"00000000", 24685 => x"00000000", 24686 => x"00000000",
    24687 => x"00000000", 24688 => x"00000000", 24689 => x"00000000",
    24690 => x"00000000", 24691 => x"00000000", 24692 => x"00000000",
    24693 => x"00000000", 24694 => x"00000000", 24695 => x"00000000",
    24696 => x"00000000", 24697 => x"00000000", 24698 => x"00000000",
    24699 => x"00000000", 24700 => x"00000000", 24701 => x"00000000",
    24702 => x"00000000", 24703 => x"00000000", 24704 => x"00000000",
    24705 => x"00000000", 24706 => x"00000000", 24707 => x"00000000",
    24708 => x"00000000", 24709 => x"00000000", 24710 => x"00000000",
    24711 => x"00000000", 24712 => x"00000000", 24713 => x"00000000",
    24714 => x"00000000", 24715 => x"00000000", 24716 => x"00000000",
    24717 => x"00000000", 24718 => x"00000000", 24719 => x"00000000",
    24720 => x"00000000", 24721 => x"00000000", 24722 => x"00000000",
    24723 => x"00000000", 24724 => x"00000000", 24725 => x"00000000",
    24726 => x"00000000", 24727 => x"00000000", 24728 => x"00000000",
    24729 => x"00000000", 24730 => x"00000000", 24731 => x"00000000",
    24732 => x"00000000", 24733 => x"00000000", 24734 => x"00000000",
    24735 => x"00000000", 24736 => x"00000000", 24737 => x"00000000",
    24738 => x"00000000", 24739 => x"00000000", 24740 => x"00000000",
    24741 => x"00000000", 24742 => x"00000000", 24743 => x"00000000",
    24744 => x"00000000", 24745 => x"00000000", 24746 => x"00000000",
    24747 => x"00000000", 24748 => x"00000000", 24749 => x"00000000",
    24750 => x"00000000", 24751 => x"00000000", 24752 => x"00000000",
    24753 => x"00000000", 24754 => x"00000000", 24755 => x"00000000",
    24756 => x"00000000", 24757 => x"00000000", 24758 => x"00000000",
    24759 => x"00000000", 24760 => x"00000000", 24761 => x"00000000",
    24762 => x"00000000", 24763 => x"00000000", 24764 => x"00000000",
    24765 => x"00000000", 24766 => x"00000000", 24767 => x"00000000",
    24768 => x"00000000", 24769 => x"00000000", 24770 => x"00000000",
    24771 => x"00000000", 24772 => x"00000000", 24773 => x"00000000",
    24774 => x"00000000", 24775 => x"00000000", 24776 => x"00000000",
    24777 => x"00000000", 24778 => x"00000000", 24779 => x"00000000",
    24780 => x"00000000", 24781 => x"00000000", 24782 => x"00000000",
    24783 => x"00000000", 24784 => x"00000000", 24785 => x"00000000",
    24786 => x"00000000", 24787 => x"00000000", 24788 => x"00000000",
    24789 => x"00000000", 24790 => x"00000000", 24791 => x"00000000",
    24792 => x"00000000", 24793 => x"00000000", 24794 => x"00000000",
    24795 => x"00000000", 24796 => x"00000000", 24797 => x"00000000",
    24798 => x"00000000", 24799 => x"00000000", 24800 => x"00000000",
    24801 => x"00000000", 24802 => x"00000000", 24803 => x"00000000",
    24804 => x"00000000", 24805 => x"00000000", 24806 => x"00000000",
    24807 => x"00000000", 24808 => x"00000000", 24809 => x"00000000",
    24810 => x"00000000", 24811 => x"00000000", 24812 => x"00000000",
    24813 => x"00000000", 24814 => x"00000000", 24815 => x"00000000",
    24816 => x"00000000", 24817 => x"00000000", 24818 => x"00000000",
    24819 => x"00000000", 24820 => x"00000000", 24821 => x"00000000",
    24822 => x"00000000", 24823 => x"00000000", 24824 => x"00000000",
    24825 => x"00000000", 24826 => x"00000000", 24827 => x"00000000",
    24828 => x"00000000", 24829 => x"00000000", 24830 => x"00000000",
    24831 => x"00000000", 24832 => x"00000000", 24833 => x"00000000",
    24834 => x"00000000", 24835 => x"00000000", 24836 => x"00000000",
    24837 => x"00000000", 24838 => x"00000000", 24839 => x"00000000",
    24840 => x"00000000", 24841 => x"00000000", 24842 => x"00000000",
    24843 => x"00000000", 24844 => x"00000000", 24845 => x"00000000",
    24846 => x"00000000", 24847 => x"00000000", 24848 => x"00000000",
    24849 => x"00000000", 24850 => x"00000000", 24851 => x"00000000",
    24852 => x"00000000", 24853 => x"00000000", 24854 => x"00000000",
    24855 => x"00000000", 24856 => x"00000000", 24857 => x"00000000",
    24858 => x"00000000", 24859 => x"00000000", 24860 => x"00000000",
    24861 => x"00000000", 24862 => x"00000000", 24863 => x"00000000",
    24864 => x"00000000", 24865 => x"00000000", 24866 => x"00000000",
    24867 => x"00000000", 24868 => x"00000000", 24869 => x"00000000",
    24870 => x"00000000", 24871 => x"00000000", 24872 => x"00000000",
    24873 => x"00000000", 24874 => x"00000000", 24875 => x"00000000",
    24876 => x"00000000", 24877 => x"00000000", 24878 => x"00000000",
    24879 => x"00000000", 24880 => x"00000000", 24881 => x"00000000",
    24882 => x"00000000", 24883 => x"00000000", 24884 => x"00000000",
    24885 => x"00000000", 24886 => x"00000000", 24887 => x"00000000",
    24888 => x"00000000", 24889 => x"00000000", 24890 => x"00000000",
    24891 => x"00000000", 24892 => x"00000000", 24893 => x"00000000",
    24894 => x"00000000", 24895 => x"00000000", 24896 => x"00000000",
    24897 => x"00000000", 24898 => x"00000000", 24899 => x"00000000",
    24900 => x"00000000", 24901 => x"00000000", 24902 => x"00000000",
    24903 => x"00000000", 24904 => x"00000000", 24905 => x"00000000",
    24906 => x"00000000", 24907 => x"00000000", 24908 => x"00000000",
    24909 => x"00000000", 24910 => x"00000000", 24911 => x"00000000",
    24912 => x"00000000", 24913 => x"00000000", 24914 => x"00000000",
    24915 => x"00000000", 24916 => x"00000000", 24917 => x"00000000",
    24918 => x"00000000", 24919 => x"00000000", 24920 => x"00000000",
    24921 => x"00000000", 24922 => x"00000000", 24923 => x"00000000",
    24924 => x"00000000", 24925 => x"00000000", 24926 => x"00000000",
    24927 => x"00000000", 24928 => x"00000000", 24929 => x"00000000",
    24930 => x"00000000", 24931 => x"00000000", 24932 => x"00000000",
    24933 => x"00000000", 24934 => x"00000000", 24935 => x"00000000",
    24936 => x"00000000", 24937 => x"00000000", 24938 => x"00000000",
    24939 => x"00000000", 24940 => x"00000000", 24941 => x"00000000",
    24942 => x"00000000", 24943 => x"00000000", 24944 => x"00000000",
    24945 => x"00000000", 24946 => x"00000000", 24947 => x"00000000",
    24948 => x"00000000", 24949 => x"00000000", 24950 => x"00000000",
    24951 => x"00000000", 24952 => x"00000000", 24953 => x"00000000",
    24954 => x"00000000", 24955 => x"00000000", 24956 => x"00000000",
    24957 => x"00000000", 24958 => x"00000000", 24959 => x"00000000",
    24960 => x"00000000", 24961 => x"00000000", 24962 => x"00000000",
    24963 => x"00000000", 24964 => x"00000000", 24965 => x"00000000",
    24966 => x"00000000", 24967 => x"00000000", 24968 => x"00000000",
    24969 => x"00000000", 24970 => x"00000000", 24971 => x"00000000",
    24972 => x"00000000", 24973 => x"00000000", 24974 => x"00000000",
    24975 => x"00000000", 24976 => x"00000000", 24977 => x"00000000",
    24978 => x"00000000", 24979 => x"00000000", 24980 => x"00000000",
    24981 => x"00000000", 24982 => x"00000000", 24983 => x"00000000",
    24984 => x"00000000", 24985 => x"00000000", 24986 => x"00000000",
    24987 => x"00000000", 24988 => x"00000000", 24989 => x"00000000",
    24990 => x"00000000", 24991 => x"00000000", 24992 => x"00000000",
    24993 => x"00000000", 24994 => x"00000000", 24995 => x"00000000",
    24996 => x"00000000", 24997 => x"00000000", 24998 => x"00000000",
    24999 => x"00000000", 25000 => x"00000000", 25001 => x"00000000",
    25002 => x"00000000", 25003 => x"00000000", 25004 => x"00000000",
    25005 => x"00000000", 25006 => x"00000000", 25007 => x"00000000",
    25008 => x"00000000", 25009 => x"00000000", 25010 => x"00000000",
    25011 => x"00000000", 25012 => x"00000000", 25013 => x"00000000",
    25014 => x"00000000", 25015 => x"00000000", 25016 => x"00000000",
    25017 => x"00000000", 25018 => x"00000000", 25019 => x"00000000",
    25020 => x"00000000", 25021 => x"00000000", 25022 => x"00000000",
    25023 => x"00000000", 25024 => x"00000000", 25025 => x"00000000",
    25026 => x"00000000", 25027 => x"00000000", 25028 => x"00000000",
    25029 => x"00000000", 25030 => x"00000000", 25031 => x"00000000",
    25032 => x"00000000", 25033 => x"00000000", 25034 => x"00000000",
    25035 => x"00000000", 25036 => x"00000000", 25037 => x"00000000",
    25038 => x"00000000", 25039 => x"00000000", 25040 => x"00000000",
    25041 => x"00000000", 25042 => x"00000000", 25043 => x"00000000",
    25044 => x"00000000", 25045 => x"00000000", 25046 => x"00000000",
    25047 => x"00000000", 25048 => x"00000000", 25049 => x"00000000",
    25050 => x"00000000", 25051 => x"00000000", 25052 => x"00000000",
    25053 => x"00000000", 25054 => x"00000000", 25055 => x"00000000",
    25056 => x"00000000", 25057 => x"00000000", 25058 => x"00000000",
    25059 => x"00000000", 25060 => x"00000000", 25061 => x"00000000",
    25062 => x"00000000", 25063 => x"00000000", 25064 => x"00000000",
    25065 => x"00000000", 25066 => x"00000000", 25067 => x"00000000",
    25068 => x"00000000", 25069 => x"00000000", 25070 => x"00000000",
    25071 => x"00000000", 25072 => x"00000000", 25073 => x"00000000",
    25074 => x"00000000", 25075 => x"00000000", 25076 => x"00000000",
    25077 => x"00000000", 25078 => x"00000000", 25079 => x"00000000",
    25080 => x"00000000", 25081 => x"00000000", 25082 => x"00000000",
    25083 => x"00000000", 25084 => x"00000000", 25085 => x"00000000",
    25086 => x"00000000", 25087 => x"00000000", 25088 => x"00000000",
    25089 => x"00000000", 25090 => x"00000000", 25091 => x"00000000",
    25092 => x"00000000", 25093 => x"00000000", 25094 => x"00000000",
    25095 => x"00000000", 25096 => x"00000000", 25097 => x"00000000",
    25098 => x"00000000", 25099 => x"00000000", 25100 => x"00000000",
    25101 => x"00000000", 25102 => x"00000000", 25103 => x"00000000",
    25104 => x"00000000", 25105 => x"00000000", 25106 => x"00000000",
    25107 => x"00000000", 25108 => x"00000000", 25109 => x"00000000",
    25110 => x"00000000", 25111 => x"00000000", 25112 => x"00000000",
    25113 => x"00000000", 25114 => x"00000000", 25115 => x"00000000",
    25116 => x"00000000", 25117 => x"00000000", 25118 => x"00000000",
    25119 => x"00000000", 25120 => x"00000000", 25121 => x"00000000",
    25122 => x"00000000", 25123 => x"00000000", 25124 => x"00000000",
    25125 => x"00000000", 25126 => x"00000000", 25127 => x"00000000",
    25128 => x"00000000", 25129 => x"00000000", 25130 => x"00000000",
    25131 => x"00000000", 25132 => x"00000000", 25133 => x"00000000",
    25134 => x"00000000", 25135 => x"00000000", 25136 => x"00000000",
    25137 => x"00000000", 25138 => x"00000000", 25139 => x"00000000",
    25140 => x"00000000", 25141 => x"00000000", 25142 => x"00000000",
    25143 => x"00000000", 25144 => x"00000000", 25145 => x"00000000",
    25146 => x"00000000", 25147 => x"00000000", 25148 => x"00000000",
    25149 => x"00000000", 25150 => x"00000000", 25151 => x"00000000",
    25152 => x"00000000", 25153 => x"00000000", 25154 => x"00000000",
    25155 => x"00000000", 25156 => x"00000000", 25157 => x"00000000",
    25158 => x"00000000", 25159 => x"00000000", 25160 => x"00000000",
    25161 => x"00000000", 25162 => x"00000000", 25163 => x"00000000",
    25164 => x"00000000", 25165 => x"00000000", 25166 => x"00000000",
    25167 => x"00000000", 25168 => x"00000000", 25169 => x"00000000",
    25170 => x"00000000", 25171 => x"00000000", 25172 => x"00000000",
    25173 => x"00000000", 25174 => x"00000000", 25175 => x"00000000",
    25176 => x"00000000", 25177 => x"00000000", 25178 => x"00000000",
    25179 => x"00000000", 25180 => x"00000000", 25181 => x"00000000",
    25182 => x"00000000", 25183 => x"00000000", 25184 => x"00000000",
    25185 => x"00000000", 25186 => x"00000000", 25187 => x"00000000",
    25188 => x"00000000", 25189 => x"00000000", 25190 => x"00000000",
    25191 => x"00000000", 25192 => x"00000000", 25193 => x"00000000",
    25194 => x"00000000", 25195 => x"00000000", 25196 => x"00000000",
    25197 => x"00000000", 25198 => x"00000000", 25199 => x"00000000",
    25200 => x"00000000", 25201 => x"00000000", 25202 => x"00000000",
    25203 => x"00000000", 25204 => x"00000000", 25205 => x"00000000",
    25206 => x"00000000", 25207 => x"00000000", 25208 => x"00000000",
    25209 => x"00000000", 25210 => x"00000000", 25211 => x"00000000",
    25212 => x"00000000", 25213 => x"00000000", 25214 => x"00000000",
    25215 => x"00000000", 25216 => x"00000000", 25217 => x"00000000",
    25218 => x"00000000", 25219 => x"00000000", 25220 => x"00000000",
    25221 => x"00000000", 25222 => x"00000000", 25223 => x"00000000",
    25224 => x"00000000", 25225 => x"00000000", 25226 => x"00000000",
    25227 => x"00000000", 25228 => x"00000000", 25229 => x"00000000",
    25230 => x"00000000", 25231 => x"00000000", 25232 => x"00000000",
    25233 => x"00000000", 25234 => x"00000000", 25235 => x"00000000",
    25236 => x"00000000", 25237 => x"00000000", 25238 => x"00000000",
    25239 => x"00000000", 25240 => x"00000000", 25241 => x"00000000",
    25242 => x"00000000", 25243 => x"00000000", 25244 => x"00000000",
    25245 => x"00000000", 25246 => x"00000000", 25247 => x"00000000",
    25248 => x"00000000", 25249 => x"00000000", 25250 => x"00000000",
    25251 => x"00000000", 25252 => x"00000000", 25253 => x"00000000",
    25254 => x"00000000", 25255 => x"00000000", 25256 => x"00000000",
    25257 => x"00000000", 25258 => x"00000000", 25259 => x"00000000",
    25260 => x"00000000", 25261 => x"00000000", 25262 => x"00000000",
    25263 => x"00000000", 25264 => x"00000000", 25265 => x"00000000",
    25266 => x"00000000", 25267 => x"00000000", 25268 => x"00000000",
    25269 => x"00000000", 25270 => x"00000000", 25271 => x"00000000",
    25272 => x"00000000", 25273 => x"00000000", 25274 => x"00000000",
    25275 => x"00000000", 25276 => x"00000000", 25277 => x"00000000",
    25278 => x"00000000", 25279 => x"00000000", 25280 => x"00000000",
    25281 => x"00000000", 25282 => x"00000000", 25283 => x"00000000",
    25284 => x"00000000", 25285 => x"00000000", 25286 => x"00000000",
    25287 => x"00000000", 25288 => x"00000000", 25289 => x"00000000",
    25290 => x"00000000", 25291 => x"00000000", 25292 => x"00000000",
    25293 => x"00000000", 25294 => x"00000000", 25295 => x"00000000",
    25296 => x"00000000", 25297 => x"00000000", 25298 => x"00000000",
    25299 => x"00000000", 25300 => x"00000000", 25301 => x"00000000",
    25302 => x"00000000", 25303 => x"00000000", 25304 => x"00000000",
    25305 => x"00000000", 25306 => x"00000000", 25307 => x"00000000",
    25308 => x"00000000", 25309 => x"00000000", 25310 => x"00000000",
    25311 => x"00000000", 25312 => x"00000000", 25313 => x"00000000",
    25314 => x"00000000", 25315 => x"00000000", 25316 => x"00000000",
    25317 => x"00000000", 25318 => x"00000000", 25319 => x"00000000",
    25320 => x"00000000", 25321 => x"00000000", 25322 => x"00000000",
    25323 => x"00000000", 25324 => x"00000000", 25325 => x"00000000",
    25326 => x"00000000", 25327 => x"00000000", 25328 => x"00000000",
    25329 => x"00000000", 25330 => x"00000000", 25331 => x"00000000",
    25332 => x"00000000", 25333 => x"00000000", 25334 => x"00000000",
    25335 => x"00000000", 25336 => x"00000000", 25337 => x"00000000",
    25338 => x"00000000", 25339 => x"00000000", 25340 => x"00000000",
    25341 => x"00000000", 25342 => x"00000000", 25343 => x"00000000",
    25344 => x"00000000", 25345 => x"00000000", 25346 => x"00000000",
    25347 => x"00000000", 25348 => x"00000000", 25349 => x"00000000",
    25350 => x"00000000", 25351 => x"00000000", 25352 => x"00000000",
    25353 => x"00000000", 25354 => x"00000000", 25355 => x"00000000",
    25356 => x"00000000", 25357 => x"00000000", 25358 => x"00000000",
    25359 => x"00000000", 25360 => x"00000000", 25361 => x"00000000",
    25362 => x"00000000", 25363 => x"00000000", 25364 => x"00000000",
    25365 => x"00000000", 25366 => x"00000000", 25367 => x"00000000",
    25368 => x"00000000", 25369 => x"00000000", 25370 => x"00000000",
    25371 => x"00000000", 25372 => x"00000000", 25373 => x"00000000",
    25374 => x"00000000", 25375 => x"00000000", 25376 => x"00000000",
    25377 => x"00000000", 25378 => x"00000000", 25379 => x"00000000",
    25380 => x"00000000", 25381 => x"00000000", 25382 => x"00000000",
    25383 => x"00000000", 25384 => x"00000000", 25385 => x"00000000",
    25386 => x"00000000", 25387 => x"00000000", 25388 => x"00000000",
    25389 => x"00000000", 25390 => x"00000000", 25391 => x"00000000",
    25392 => x"00000000", 25393 => x"00000000", 25394 => x"00000000",
    25395 => x"00000000", 25396 => x"00000000", 25397 => x"00000000",
    25398 => x"00000000", 25399 => x"00000000", 25400 => x"00000000",
    25401 => x"00000000", 25402 => x"00000000", 25403 => x"00000000",
    25404 => x"00000000", 25405 => x"00000000", 25406 => x"00000000",
    25407 => x"00000000", 25408 => x"00000000", 25409 => x"00000000",
    25410 => x"00000000", 25411 => x"00000000", 25412 => x"00000000",
    25413 => x"00000000", 25414 => x"00000000", 25415 => x"00000000",
    25416 => x"00000000", 25417 => x"00000000", 25418 => x"00000000",
    25419 => x"00000000", 25420 => x"00000000", 25421 => x"00000000",
    25422 => x"00000000", 25423 => x"00000000", 25424 => x"00000000",
    25425 => x"00000000", 25426 => x"00000000", 25427 => x"00000000",
    25428 => x"00000000", 25429 => x"00000000", 25430 => x"00000000",
    25431 => x"00000000", 25432 => x"00000000", 25433 => x"00000000",
    25434 => x"00000000", 25435 => x"00000000", 25436 => x"00000000",
    25437 => x"00000000", 25438 => x"00000000", 25439 => x"00000000",
    25440 => x"00000000", 25441 => x"00000000", 25442 => x"00000000",
    25443 => x"00000000", 25444 => x"00000000", 25445 => x"00000000",
    25446 => x"00000000", 25447 => x"00000000", 25448 => x"00000000",
    25449 => x"00000000", 25450 => x"00000000", 25451 => x"00000000",
    25452 => x"00000000", 25453 => x"00000000", 25454 => x"00000000",
    25455 => x"00000000", 25456 => x"00000000", 25457 => x"00000000",
    25458 => x"00000000", 25459 => x"00000000", 25460 => x"00000000",
    25461 => x"00000000", 25462 => x"00000000", 25463 => x"00000000",
    25464 => x"00000000", 25465 => x"00000000", 25466 => x"00000000",
    25467 => x"00000000", 25468 => x"00000000", 25469 => x"00000000",
    25470 => x"00000000", 25471 => x"00000000", 25472 => x"00000000",
    25473 => x"00000000", 25474 => x"00000000", 25475 => x"00000000",
    25476 => x"00000000", 25477 => x"00000000", 25478 => x"00000000",
    25479 => x"00000000", 25480 => x"00000000", 25481 => x"00000000",
    25482 => x"00000000", 25483 => x"00000000", 25484 => x"00000000",
    25485 => x"00000000", 25486 => x"00000000", 25487 => x"00000000",
    25488 => x"00000000", 25489 => x"00000000", 25490 => x"00000000",
    25491 => x"00000000", 25492 => x"00000000", 25493 => x"00000000",
    25494 => x"00000000", 25495 => x"00000000", 25496 => x"00000000",
    25497 => x"00000000", 25498 => x"00000000", 25499 => x"00000000",
    25500 => x"00000000", 25501 => x"00000000", 25502 => x"00000000",
    25503 => x"00000000", 25504 => x"00000000", 25505 => x"00000000",
    25506 => x"00000000", 25507 => x"00000000", 25508 => x"00000000",
    25509 => x"00000000", 25510 => x"00000000", 25511 => x"00000000",
    25512 => x"00000000", 25513 => x"00000000", 25514 => x"00000000",
    25515 => x"00000000", 25516 => x"00000000", 25517 => x"00000000",
    25518 => x"00000000", 25519 => x"00000000", 25520 => x"00000000",
    25521 => x"00000000", 25522 => x"00000000", 25523 => x"00000000",
    25524 => x"00000000", 25525 => x"00000000", 25526 => x"00000000",
    25527 => x"00000000", 25528 => x"00000000", 25529 => x"00000000",
    25530 => x"00000000", 25531 => x"00000000", 25532 => x"00000000",
    25533 => x"00000000", 25534 => x"00000000", 25535 => x"00000000",
    25536 => x"00000000", 25537 => x"00000000", 25538 => x"00000000",
    25539 => x"00000000", 25540 => x"00000000", 25541 => x"00000000",
    25542 => x"00000000", 25543 => x"00000000", 25544 => x"00000000",
    25545 => x"00000000", 25546 => x"00000000", 25547 => x"00000000",
    25548 => x"00000000", 25549 => x"00000000", 25550 => x"00000000",
    25551 => x"00000000", 25552 => x"00000000", 25553 => x"00000000",
    25554 => x"00000000", 25555 => x"00000000", 25556 => x"00000000",
    25557 => x"00000000", 25558 => x"00000000", 25559 => x"00000000",
    25560 => x"00000000", 25561 => x"00000000", 25562 => x"00000000",
    25563 => x"00000000", 25564 => x"00000000", 25565 => x"00000000",
    25566 => x"00000000", 25567 => x"00000000", 25568 => x"00000000",
    25569 => x"00000000", 25570 => x"00000000", 25571 => x"00000000",
    25572 => x"00000000", 25573 => x"00000000", 25574 => x"00000000",
    25575 => x"00000000", 25576 => x"00000000", 25577 => x"00000000",
    25578 => x"00000000", 25579 => x"00000000", 25580 => x"00000000",
    25581 => x"00000000", 25582 => x"00000000", 25583 => x"00000000",
    25584 => x"00000000", 25585 => x"00000000", 25586 => x"00000000",
    25587 => x"00000000", 25588 => x"00000000", 25589 => x"00000000",
    25590 => x"00000000", 25591 => x"00000000", 25592 => x"00000000",
    25593 => x"00000000", 25594 => x"00000000", 25595 => x"00000000",
    25596 => x"00000000", 25597 => x"00000000", 25598 => x"00000000",
    25599 => x"00000000", 25600 => x"00000000", 25601 => x"00000000",
    25602 => x"00000000", 25603 => x"00000000", 25604 => x"00000000",
    25605 => x"00000000", 25606 => x"00000000", 25607 => x"00000000",
    25608 => x"00000000", 25609 => x"00000000", 25610 => x"00000000",
    25611 => x"00000000", 25612 => x"00000000", 25613 => x"00000000",
    25614 => x"00000000", 25615 => x"00000000", 25616 => x"00000000",
    25617 => x"00000000", 25618 => x"00000000", 25619 => x"00000000",
    25620 => x"00000000", 25621 => x"00000000", 25622 => x"00000000",
    25623 => x"00000000", 25624 => x"00000000", 25625 => x"00000000",
    25626 => x"00000000", 25627 => x"00000000", 25628 => x"00000000",
    25629 => x"00000000", 25630 => x"00000000", 25631 => x"00000000",
    25632 => x"00000000", 25633 => x"00000000", 25634 => x"00000000",
    25635 => x"00000000", 25636 => x"00000000", 25637 => x"00000000",
    25638 => x"00000000", 25639 => x"00000000", 25640 => x"00000000",
    25641 => x"00000000", 25642 => x"00000000", 25643 => x"00000000",
    25644 => x"00000000", 25645 => x"00000000", 25646 => x"00000000",
    25647 => x"00000000", 25648 => x"00000000", 25649 => x"00000000",
    25650 => x"00000000", 25651 => x"00000000", 25652 => x"00000000",
    25653 => x"00000000", 25654 => x"00000000", 25655 => x"00000000",
    25656 => x"00000000", 25657 => x"00000000", 25658 => x"00000000",
    25659 => x"00000000", 25660 => x"00000000", 25661 => x"00000000",
    25662 => x"00000000", 25663 => x"00000000", 25664 => x"00000000",
    25665 => x"00000000", 25666 => x"00000000", 25667 => x"00000000",
    25668 => x"00000000", 25669 => x"00000000", 25670 => x"00000000",
    25671 => x"00000000", 25672 => x"00000000", 25673 => x"00000000",
    25674 => x"00000000", 25675 => x"00000000", 25676 => x"00000000",
    25677 => x"00000000", 25678 => x"00000000", 25679 => x"00000000",
    25680 => x"00000000", 25681 => x"00000000", 25682 => x"00000000",
    25683 => x"00000000", 25684 => x"00000000", 25685 => x"00000000",
    25686 => x"00000000", 25687 => x"00000000", 25688 => x"00000000",
    25689 => x"00000000", 25690 => x"00000000", 25691 => x"00000000",
    25692 => x"00000000", 25693 => x"00000000", 25694 => x"00000000",
    25695 => x"00000000", 25696 => x"00000000", 25697 => x"00000000",
    25698 => x"00000000", 25699 => x"00000000", 25700 => x"00000000",
    25701 => x"00000000", 25702 => x"00000000", 25703 => x"00000000",
    25704 => x"00000000", 25705 => x"00000000", 25706 => x"00000000",
    25707 => x"00000000", 25708 => x"00000000", 25709 => x"00000000",
    25710 => x"00000000", 25711 => x"00000000", 25712 => x"00000000",
    25713 => x"00000000", 25714 => x"00000000", 25715 => x"00000000",
    25716 => x"00000000", 25717 => x"00000000", 25718 => x"00000000",
    25719 => x"00000000", 25720 => x"00000000", 25721 => x"00000000",
    25722 => x"00000000", 25723 => x"00000000", 25724 => x"00000000",
    25725 => x"00000000", 25726 => x"00000000", 25727 => x"00000000",
    25728 => x"00000000", 25729 => x"00000000", 25730 => x"00000000",
    25731 => x"00000000", 25732 => x"00000000", 25733 => x"00000000",
    25734 => x"00000000", 25735 => x"00000000", 25736 => x"00000000",
    25737 => x"00000000", 25738 => x"00000000", 25739 => x"00000000",
    25740 => x"00000000", 25741 => x"00000000", 25742 => x"00000000",
    25743 => x"00000000", 25744 => x"00000000", 25745 => x"00000000",
    25746 => x"00000000", 25747 => x"00000000", 25748 => x"00000000",
    25749 => x"00000000", 25750 => x"00000000", 25751 => x"00000000",
    25752 => x"00000000", 25753 => x"00000000", 25754 => x"00000000",
    25755 => x"00000000", 25756 => x"00000000", 25757 => x"00000000",
    25758 => x"00000000", 25759 => x"00000000", 25760 => x"00000000",
    25761 => x"00000000", 25762 => x"00000000", 25763 => x"00000000",
    25764 => x"00000000", 25765 => x"00000000", 25766 => x"00000000",
    25767 => x"00000000", 25768 => x"00000000", 25769 => x"00000000",
    25770 => x"00000000", 25771 => x"00000000", 25772 => x"00000000",
    25773 => x"00000000", 25774 => x"00000000", 25775 => x"00000000",
    25776 => x"00000000", 25777 => x"00000000", 25778 => x"00000000",
    25779 => x"00000000", 25780 => x"00000000", 25781 => x"00000000",
    25782 => x"00000000", 25783 => x"00000000", 25784 => x"00000000",
    25785 => x"00000000", 25786 => x"00000000", 25787 => x"00000000",
    25788 => x"00000000", 25789 => x"00000000", 25790 => x"00000000",
    25791 => x"00000000", 25792 => x"00000000", 25793 => x"00000000",
    25794 => x"00000000", 25795 => x"00000000", 25796 => x"00000000",
    25797 => x"00000000", 25798 => x"00000000", 25799 => x"00000000",
    25800 => x"00000000", 25801 => x"00000000", 25802 => x"00000000",
    25803 => x"00000000", 25804 => x"00000000", 25805 => x"00000000",
    25806 => x"00000000", 25807 => x"00000000", 25808 => x"00000000",
    25809 => x"00000000", 25810 => x"00000000", 25811 => x"00000000",
    25812 => x"00000000", 25813 => x"00000000", 25814 => x"00000000",
    25815 => x"00000000", 25816 => x"00000000", 25817 => x"00000000",
    25818 => x"00000000", 25819 => x"00000000", 25820 => x"00000000",
    25821 => x"00000000", 25822 => x"00000000", 25823 => x"00000000",
    25824 => x"00000000", 25825 => x"00000000", 25826 => x"00000000",
    25827 => x"00000000", 25828 => x"00000000", 25829 => x"00000000",
    25830 => x"00000000", 25831 => x"00000000", 25832 => x"00000000",
    25833 => x"00000000", 25834 => x"00000000", 25835 => x"00000000",
    25836 => x"00000000", 25837 => x"00000000", 25838 => x"00000000",
    25839 => x"00000000", 25840 => x"00000000", 25841 => x"00000000",
    25842 => x"00000000", 25843 => x"00000000", 25844 => x"00000000",
    25845 => x"00000000", 25846 => x"00000000", 25847 => x"00000000",
    25848 => x"00000000", 25849 => x"00000000", 25850 => x"00000000",
    25851 => x"00000000", 25852 => x"00000000", 25853 => x"00000000",
    25854 => x"00000000", 25855 => x"00000000", 25856 => x"00000000",
    25857 => x"00000000", 25858 => x"00000000", 25859 => x"00000000",
    25860 => x"00000000", 25861 => x"00000000", 25862 => x"00000000",
    25863 => x"00000000", 25864 => x"00000000", 25865 => x"00000000",
    25866 => x"00000000", 25867 => x"00000000", 25868 => x"00000000",
    25869 => x"00000000", 25870 => x"00000000", 25871 => x"00000000",
    25872 => x"00000000", 25873 => x"00000000", 25874 => x"00000000",
    25875 => x"00000000", 25876 => x"00000000", 25877 => x"00000000",
    25878 => x"00000000", 25879 => x"00000000", 25880 => x"00000000",
    25881 => x"00000000", 25882 => x"00000000", 25883 => x"00000000",
    25884 => x"00000000", 25885 => x"00000000", 25886 => x"00000000",
    25887 => x"00000000", 25888 => x"00000000", 25889 => x"00000000",
    25890 => x"00000000", 25891 => x"00000000", 25892 => x"00000000",
    25893 => x"00000000", 25894 => x"00000000", 25895 => x"00000000",
    25896 => x"00000000", 25897 => x"00000000", 25898 => x"00000000",
    25899 => x"00000000", 25900 => x"00000000", 25901 => x"00000000",
    25902 => x"00000000", 25903 => x"00000000", 25904 => x"00000000",
    25905 => x"00000000", 25906 => x"00000000", 25907 => x"00000000",
    25908 => x"00000000", 25909 => x"00000000", 25910 => x"00000000",
    25911 => x"00000000", 25912 => x"00000000", 25913 => x"00000000",
    25914 => x"00000000", 25915 => x"00000000", 25916 => x"00000000",
    25917 => x"00000000", 25918 => x"00000000", 25919 => x"00000000",
    25920 => x"00000000", 25921 => x"00000000", 25922 => x"00000000",
    25923 => x"00000000", 25924 => x"00000000", 25925 => x"00000000",
    25926 => x"00000000", 25927 => x"00000000", 25928 => x"00000000",
    25929 => x"00000000", 25930 => x"00000000", 25931 => x"00000000",
    25932 => x"00000000", 25933 => x"00000000", 25934 => x"00000000",
    25935 => x"00000000", 25936 => x"00000000", 25937 => x"00000000",
    25938 => x"00000000", 25939 => x"00000000", 25940 => x"00000000",
    25941 => x"00000000", 25942 => x"00000000", 25943 => x"00000000",
    25944 => x"00000000", 25945 => x"00000000", 25946 => x"00000000",
    25947 => x"00000000", 25948 => x"00000000", 25949 => x"00000000",
    25950 => x"00000000", 25951 => x"00000000", 25952 => x"00000000",
    25953 => x"00000000", 25954 => x"00000000", 25955 => x"00000000",
    25956 => x"00000000", 25957 => x"00000000", 25958 => x"00000000",
    25959 => x"00000000", 25960 => x"00000000", 25961 => x"00000000",
    25962 => x"00000000", 25963 => x"00000000", 25964 => x"00000000",
    25965 => x"00000000", 25966 => x"00000000", 25967 => x"00000000",
    25968 => x"00000000", 25969 => x"00000000", 25970 => x"00000000",
    25971 => x"00000000", 25972 => x"00000000", 25973 => x"00000000",
    25974 => x"00000000", 25975 => x"00000000", 25976 => x"00000000",
    25977 => x"00000000", 25978 => x"00000000", 25979 => x"00000000",
    25980 => x"00000000", 25981 => x"00000000", 25982 => x"00000000",
    25983 => x"00000000", 25984 => x"00000000", 25985 => x"00000000",
    25986 => x"00000000", 25987 => x"00000000", 25988 => x"00000000",
    25989 => x"00000000", 25990 => x"00000000", 25991 => x"00000000",
    25992 => x"00000000", 25993 => x"00000000", 25994 => x"00000000",
    25995 => x"00000000", 25996 => x"00000000", 25997 => x"00000000",
    25998 => x"00000000", 25999 => x"00000000", 26000 => x"00000000",
    26001 => x"00000000", 26002 => x"00000000", 26003 => x"00000000",
    26004 => x"00000000", 26005 => x"00000000", 26006 => x"00000000",
    26007 => x"00000000", 26008 => x"00000000", 26009 => x"00000000",
    26010 => x"00000000", 26011 => x"00000000", 26012 => x"00000000",
    26013 => x"00000000", 26014 => x"00000000", 26015 => x"00000000",
    26016 => x"00000000", 26017 => x"00000000", 26018 => x"00000000",
    26019 => x"00000000", 26020 => x"00000000", 26021 => x"00000000",
    26022 => x"00000000", 26023 => x"00000000", 26024 => x"00000000",
    26025 => x"00000000", 26026 => x"00000000", 26027 => x"00000000",
    26028 => x"00000000", 26029 => x"00000000", 26030 => x"00000000",
    26031 => x"00000000", 26032 => x"00000000", 26033 => x"00000000",
    26034 => x"00000000", 26035 => x"00000000", 26036 => x"00000000",
    26037 => x"00000000", 26038 => x"00000000", 26039 => x"00000000",
    26040 => x"00000000", 26041 => x"00000000", 26042 => x"00000000",
    26043 => x"00000000", 26044 => x"00000000", 26045 => x"00000000",
    26046 => x"00000000", 26047 => x"00000000", 26048 => x"00000000",
    26049 => x"00000000", 26050 => x"00000000", 26051 => x"00000000",
    26052 => x"00000000", 26053 => x"00000000", 26054 => x"00000000",
    26055 => x"00000000", 26056 => x"00000000", 26057 => x"00000000",
    26058 => x"00000000", 26059 => x"00000000", 26060 => x"00000000",
    26061 => x"00000000", 26062 => x"00000000", 26063 => x"00000000",
    26064 => x"00000000", 26065 => x"00000000", 26066 => x"00000000",
    26067 => x"00000000", 26068 => x"00000000", 26069 => x"00000000",
    26070 => x"00000000", 26071 => x"00000000", 26072 => x"00000000",
    26073 => x"00000000", 26074 => x"00000000", 26075 => x"00000000",
    26076 => x"00000000", 26077 => x"00000000", 26078 => x"00000000",
    26079 => x"00000000", 26080 => x"00000000", 26081 => x"00000000",
    26082 => x"00000000", 26083 => x"00000000", 26084 => x"00000000",
    26085 => x"00000000", 26086 => x"00000000", 26087 => x"00000000",
    26088 => x"00000000", 26089 => x"00000000", 26090 => x"00000000",
    26091 => x"00000000", 26092 => x"00000000", 26093 => x"00000000",
    26094 => x"00000000", 26095 => x"00000000", 26096 => x"00000000",
    26097 => x"00000000", 26098 => x"00000000", 26099 => x"00000000",
    26100 => x"00000000", 26101 => x"00000000", 26102 => x"00000000",
    26103 => x"00000000", 26104 => x"00000000", 26105 => x"00000000",
    26106 => x"00000000", 26107 => x"00000000", 26108 => x"00000000",
    26109 => x"00000000", 26110 => x"00000000", 26111 => x"00000000",
    26112 => x"00000000", 26113 => x"00000000", 26114 => x"00000000",
    26115 => x"00000000", 26116 => x"00000000", 26117 => x"00000000",
    26118 => x"00000000", 26119 => x"00000000", 26120 => x"00000000",
    26121 => x"00000000", 26122 => x"00000000", 26123 => x"00000000",
    26124 => x"00000000", 26125 => x"00000000", 26126 => x"00000000",
    26127 => x"00000000", 26128 => x"00000000", 26129 => x"00000000",
    26130 => x"00000000", 26131 => x"00000000", 26132 => x"00000000",
    26133 => x"00000000", 26134 => x"00000000", 26135 => x"00000000",
    26136 => x"00000000", 26137 => x"00000000", 26138 => x"00000000",
    26139 => x"00000000", 26140 => x"00000000", 26141 => x"00000000",
    26142 => x"00000000", 26143 => x"00000000", 26144 => x"00000000",
    26145 => x"00000000", 26146 => x"00000000", 26147 => x"00000000",
    26148 => x"00000000", 26149 => x"00000000", 26150 => x"00000000",
    26151 => x"00000000", 26152 => x"00000000", 26153 => x"00000000",
    26154 => x"00000000", 26155 => x"00000000", 26156 => x"00000000",
    26157 => x"00000000", 26158 => x"00000000", 26159 => x"00000000",
    26160 => x"00000000", 26161 => x"00000000", 26162 => x"00000000",
    26163 => x"00000000", 26164 => x"00000000", 26165 => x"00000000",
    26166 => x"00000000", 26167 => x"00000000", 26168 => x"00000000",
    26169 => x"00000000", 26170 => x"00000000", 26171 => x"00000000",
    26172 => x"00000000", 26173 => x"00000000", 26174 => x"00000000",
    26175 => x"00000000", 26176 => x"00000000", 26177 => x"00000000",
    26178 => x"00000000", 26179 => x"00000000", 26180 => x"00000000",
    26181 => x"00000000", 26182 => x"00000000", 26183 => x"00000000",
    26184 => x"00000000", 26185 => x"00000000", 26186 => x"00000000",
    26187 => x"00000000", 26188 => x"00000000", 26189 => x"00000000",
    26190 => x"00000000", 26191 => x"00000000", 26192 => x"00000000",
    26193 => x"00000000", 26194 => x"00000000", 26195 => x"00000000",
    26196 => x"00000000", 26197 => x"00000000", 26198 => x"00000000",
    26199 => x"00000000", 26200 => x"00000000", 26201 => x"00000000",
    26202 => x"00000000", 26203 => x"00000000", 26204 => x"00000000",
    26205 => x"00000000", 26206 => x"00000000", 26207 => x"00000000",
    26208 => x"00000000", 26209 => x"00000000", 26210 => x"00000000",
    26211 => x"00000000", 26212 => x"00000000", 26213 => x"00000000",
    26214 => x"00000000", 26215 => x"00000000", 26216 => x"00000000",
    26217 => x"00000000", 26218 => x"00000000", 26219 => x"00000000",
    26220 => x"00000000", 26221 => x"00000000", 26222 => x"00000000",
    26223 => x"00000000", 26224 => x"00000000", 26225 => x"00000000",
    26226 => x"00000000", 26227 => x"00000000", 26228 => x"00000000",
    26229 => x"00000000", 26230 => x"00000000", 26231 => x"00000000",
    26232 => x"00000000", 26233 => x"00000000", 26234 => x"00000000",
    26235 => x"00000000", 26236 => x"00000000", 26237 => x"00000000",
    26238 => x"00000000", 26239 => x"00000000", 26240 => x"00000000",
    26241 => x"00000000", 26242 => x"00000000", 26243 => x"00000000",
    26244 => x"00000000", 26245 => x"00000000", 26246 => x"00000000",
    26247 => x"00000000", 26248 => x"00000000", 26249 => x"00000000",
    26250 => x"00000000", 26251 => x"00000000", 26252 => x"00000000",
    26253 => x"00000000", 26254 => x"00000000", 26255 => x"00000000",
    26256 => x"00000000", 26257 => x"00000000", 26258 => x"00000000",
    26259 => x"00000000", 26260 => x"00000000", 26261 => x"00000000",
    26262 => x"00000000", 26263 => x"00000000", 26264 => x"00000000",
    26265 => x"00000000", 26266 => x"00000000", 26267 => x"00000000",
    26268 => x"00000000", 26269 => x"00000000", 26270 => x"00000000",
    26271 => x"00000000", 26272 => x"00000000", 26273 => x"00000000",
    26274 => x"00000000", 26275 => x"00000000", 26276 => x"00000000",
    26277 => x"00000000", 26278 => x"00000000", 26279 => x"00000000",
    26280 => x"00000000", 26281 => x"00000000", 26282 => x"00000000",
    26283 => x"00000000", 26284 => x"00000000", 26285 => x"00000000",
    26286 => x"00000000", 26287 => x"00000000", 26288 => x"00000000",
    26289 => x"00000000", 26290 => x"00000000", 26291 => x"00000000",
    26292 => x"00000000", 26293 => x"00000000", 26294 => x"00000000",
    26295 => x"00000000", 26296 => x"00000000", 26297 => x"00000000",
    26298 => x"00000000", 26299 => x"00000000", 26300 => x"00000000",
    26301 => x"00000000", 26302 => x"00000000", 26303 => x"00000000",
    26304 => x"00000000", 26305 => x"00000000", 26306 => x"00000000",
    26307 => x"00000000", 26308 => x"00000000", 26309 => x"00000000",
    26310 => x"00000000", 26311 => x"00000000", 26312 => x"00000000",
    26313 => x"00000000", 26314 => x"00000000", 26315 => x"00000000",
    26316 => x"00000000", 26317 => x"00000000", 26318 => x"00000000",
    26319 => x"00000000", 26320 => x"00000000", 26321 => x"00000000",
    26322 => x"00000000", 26323 => x"00000000", 26324 => x"00000000",
    26325 => x"00000000", 26326 => x"00000000", 26327 => x"00000000",
    26328 => x"00000000", 26329 => x"00000000", 26330 => x"00000000",
    26331 => x"00000000", 26332 => x"00000000", 26333 => x"00000000",
    26334 => x"00000000", 26335 => x"00000000", 26336 => x"00000000",
    26337 => x"00000000", 26338 => x"00000000", 26339 => x"00000000",
    26340 => x"00000000", 26341 => x"00000000", 26342 => x"00000000",
    26343 => x"00000000", 26344 => x"00000000", 26345 => x"00000000",
    26346 => x"00000000", 26347 => x"00000000", 26348 => x"00000000",
    26349 => x"00000000", 26350 => x"00000000", 26351 => x"00000000",
    26352 => x"00000000", 26353 => x"00000000", 26354 => x"00000000",
    26355 => x"00000000", 26356 => x"00000000", 26357 => x"00000000",
    26358 => x"00000000", 26359 => x"00000000", 26360 => x"00000000",
    26361 => x"00000000", 26362 => x"00000000", 26363 => x"00000000",
    26364 => x"00000000", 26365 => x"00000000", 26366 => x"00000000",
    26367 => x"00000000", 26368 => x"00000000", 26369 => x"00000000",
    26370 => x"00000000", 26371 => x"00000000", 26372 => x"00000000",
    26373 => x"00000000", 26374 => x"00000000", 26375 => x"00000000",
    26376 => x"00000000", 26377 => x"00000000", 26378 => x"00000000",
    26379 => x"00000000", 26380 => x"00000000", 26381 => x"00000000",
    26382 => x"00000000", 26383 => x"00000000", 26384 => x"00000000",
    26385 => x"00000000", 26386 => x"00000000", 26387 => x"00000000",
    26388 => x"00000000", 26389 => x"00000000", 26390 => x"00000000",
    26391 => x"00000000", 26392 => x"00000000", 26393 => x"00000000",
    26394 => x"00000000", 26395 => x"00000000", 26396 => x"00000000",
    26397 => x"00000000", 26398 => x"00000000", 26399 => x"00000000",
    26400 => x"00000000", 26401 => x"00000000", 26402 => x"00000000",
    26403 => x"00000000", 26404 => x"00000000", 26405 => x"00000000",
    26406 => x"00000000", 26407 => x"00000000", 26408 => x"00000000",
    26409 => x"00000000", 26410 => x"00000000", 26411 => x"00000000",
    26412 => x"00000000", 26413 => x"00000000", 26414 => x"00000000",
    26415 => x"00000000", 26416 => x"00000000", 26417 => x"00000000",
    26418 => x"00000000", 26419 => x"00000000", 26420 => x"00000000",
    26421 => x"00000000", 26422 => x"00000000", 26423 => x"00000000",
    26424 => x"00000000", 26425 => x"00000000", 26426 => x"00000000",
    26427 => x"00000000", 26428 => x"00000000", 26429 => x"00000000",
    26430 => x"00000000", 26431 => x"00000000", 26432 => x"00000000",
    26433 => x"00000000", 26434 => x"00000000", 26435 => x"00000000",
    26436 => x"00000000", 26437 => x"00000000", 26438 => x"00000000",
    26439 => x"00000000", 26440 => x"00000000", 26441 => x"00000000",
    26442 => x"00000000", 26443 => x"00000000", 26444 => x"00000000",
    26445 => x"00000000", 26446 => x"00000000", 26447 => x"00000000",
    26448 => x"00000000", 26449 => x"00000000", 26450 => x"00000000",
    26451 => x"00000000", 26452 => x"00000000", 26453 => x"00000000",
    26454 => x"00000000", 26455 => x"00000000", 26456 => x"00000000",
    26457 => x"00000000", 26458 => x"00000000", 26459 => x"00000000",
    26460 => x"00000000", 26461 => x"00000000", 26462 => x"00000000",
    26463 => x"00000000", 26464 => x"00000000", 26465 => x"00000000",
    26466 => x"00000000", 26467 => x"00000000", 26468 => x"00000000",
    26469 => x"00000000", 26470 => x"00000000", 26471 => x"00000000",
    26472 => x"00000000", 26473 => x"00000000", 26474 => x"00000000",
    26475 => x"00000000", 26476 => x"00000000", 26477 => x"00000000",
    26478 => x"00000000", 26479 => x"00000000", 26480 => x"00000000",
    26481 => x"00000000", 26482 => x"00000000", 26483 => x"00000000",
    26484 => x"00000000", 26485 => x"00000000", 26486 => x"00000000",
    26487 => x"00000000", 26488 => x"00000000", 26489 => x"00000000",
    26490 => x"00000000", 26491 => x"00000000", 26492 => x"00000000",
    26493 => x"00000000", 26494 => x"00000000", 26495 => x"00000000",
    26496 => x"00000000", 26497 => x"00000000", 26498 => x"00000000",
    26499 => x"00000000", 26500 => x"00000000", 26501 => x"00000000",
    26502 => x"00000000", 26503 => x"00000000", 26504 => x"00000000",
    26505 => x"00000000", 26506 => x"00000000", 26507 => x"00000000",
    26508 => x"00000000", 26509 => x"00000000", 26510 => x"00000000",
    26511 => x"00000000", 26512 => x"00000000", 26513 => x"00000000",
    26514 => x"00000000", 26515 => x"00000000", 26516 => x"00000000",
    26517 => x"00000000", 26518 => x"00000000", 26519 => x"00000000",
    26520 => x"00000000", 26521 => x"00000000", 26522 => x"00000000",
    26523 => x"00000000", 26524 => x"00000000", 26525 => x"00000000",
    26526 => x"00000000", 26527 => x"00000000", 26528 => x"00000000",
    26529 => x"00000000", 26530 => x"00000000", 26531 => x"00000000",
    26532 => x"00000000", 26533 => x"00000000", 26534 => x"00000000",
    26535 => x"00000000", 26536 => x"00000000", 26537 => x"00000000",
    26538 => x"00000000", 26539 => x"00000000", 26540 => x"00000000",
    26541 => x"00000000", 26542 => x"00000000", 26543 => x"00000000",
    26544 => x"00000000", 26545 => x"00000000", 26546 => x"00000000",
    26547 => x"00000000", 26548 => x"00000000", 26549 => x"00000000",
    26550 => x"00000000", 26551 => x"00000000", 26552 => x"00000000",
    26553 => x"00000000", 26554 => x"00000000", 26555 => x"00000000",
    26556 => x"00000000", 26557 => x"00000000", 26558 => x"00000000",
    26559 => x"00000000", 26560 => x"00000000", 26561 => x"00000000",
    26562 => x"00000000", 26563 => x"00000000", 26564 => x"00000000",
    26565 => x"00000000", 26566 => x"00000000", 26567 => x"00000000",
    26568 => x"00000000", 26569 => x"00000000", 26570 => x"00000000",
    26571 => x"00000000", 26572 => x"00000000", 26573 => x"00000000",
    26574 => x"00000000", 26575 => x"00000000", 26576 => x"00000000",
    26577 => x"00000000", 26578 => x"00000000", 26579 => x"00000000",
    26580 => x"00000000", 26581 => x"00000000", 26582 => x"00000000",
    26583 => x"00000000", 26584 => x"00000000", 26585 => x"00000000",
    26586 => x"00000000", 26587 => x"00000000", 26588 => x"00000000",
    26589 => x"00000000", 26590 => x"00000000", 26591 => x"00000000",
    26592 => x"00000000", 26593 => x"00000000", 26594 => x"00000000",
    26595 => x"00000000", 26596 => x"00000000", 26597 => x"00000000",
    26598 => x"00000000", 26599 => x"00000000", 26600 => x"00000000",
    26601 => x"00000000", 26602 => x"00000000", 26603 => x"00000000",
    26604 => x"00000000", 26605 => x"00000000", 26606 => x"00000000",
    26607 => x"00000000", 26608 => x"00000000", 26609 => x"00000000",
    26610 => x"00000000", 26611 => x"00000000", 26612 => x"00000000",
    26613 => x"00000000", 26614 => x"00000000", 26615 => x"00000000",
    26616 => x"00000000", 26617 => x"00000000", 26618 => x"00000000",
    26619 => x"00000000", 26620 => x"00000000", 26621 => x"00000000",
    26622 => x"00000000", 26623 => x"00000000", 26624 => x"00000000",
    26625 => x"00000000", 26626 => x"00000000", 26627 => x"00000000",
    26628 => x"00000000", 26629 => x"00000000", 26630 => x"00000000",
    26631 => x"00000000", 26632 => x"00000000", 26633 => x"00000000",
    26634 => x"00000000", 26635 => x"00000000", 26636 => x"00000000",
    26637 => x"00000000", 26638 => x"00000000", 26639 => x"00000000",
    26640 => x"00000000", 26641 => x"00000000", 26642 => x"00000000",
    26643 => x"00000000", 26644 => x"00000000", 26645 => x"00000000",
    26646 => x"00000000", 26647 => x"00000000", 26648 => x"00000000",
    26649 => x"00000000", 26650 => x"00000000", 26651 => x"00000000",
    26652 => x"00000000", 26653 => x"00000000", 26654 => x"00000000",
    26655 => x"00000000", 26656 => x"00000000", 26657 => x"00000000",
    26658 => x"00000000", 26659 => x"00000000", 26660 => x"00000000",
    26661 => x"00000000", 26662 => x"00000000", 26663 => x"00000000",
    26664 => x"00000000", 26665 => x"00000000", 26666 => x"00000000",
    26667 => x"00000000", 26668 => x"00000000", 26669 => x"00000000",
    26670 => x"00000000", 26671 => x"00000000", 26672 => x"00000000",
    26673 => x"00000000", 26674 => x"00000000", 26675 => x"00000000",
    26676 => x"00000000", 26677 => x"00000000", 26678 => x"00000000",
    26679 => x"00000000", 26680 => x"00000000", 26681 => x"00000000",
    26682 => x"00000000", 26683 => x"00000000", 26684 => x"00000000",
    26685 => x"00000000", 26686 => x"00000000", 26687 => x"00000000",
    26688 => x"00000000", 26689 => x"00000000", 26690 => x"00000000",
    26691 => x"00000000", 26692 => x"00000000", 26693 => x"00000000",
    26694 => x"00000000", 26695 => x"00000000", 26696 => x"00000000",
    26697 => x"00000000", 26698 => x"00000000", 26699 => x"00000000",
    26700 => x"00000000", 26701 => x"00000000", 26702 => x"00000000",
    26703 => x"00000000", 26704 => x"00000000", 26705 => x"00000000",
    26706 => x"00000000", 26707 => x"00000000", 26708 => x"00000000",
    26709 => x"00000000", 26710 => x"00000000", 26711 => x"00000000",
    26712 => x"00000000", 26713 => x"00000000", 26714 => x"00000000",
    26715 => x"00000000", 26716 => x"00000000", 26717 => x"00000000",
    26718 => x"00000000", 26719 => x"00000000", 26720 => x"00000000",
    26721 => x"00000000", 26722 => x"00000000", 26723 => x"00000000",
    26724 => x"00000000", 26725 => x"00000000", 26726 => x"00000000",
    26727 => x"00000000", 26728 => x"00000000", 26729 => x"00000000",
    26730 => x"00000000", 26731 => x"00000000", 26732 => x"00000000",
    26733 => x"00000000", 26734 => x"00000000", 26735 => x"00000000",
    26736 => x"00000000", 26737 => x"00000000", 26738 => x"00000000",
    26739 => x"00000000", 26740 => x"00000000", 26741 => x"00000000",
    26742 => x"00000000", 26743 => x"00000000", 26744 => x"00000000",
    26745 => x"00000000", 26746 => x"00000000", 26747 => x"00000000",
    26748 => x"00000000", 26749 => x"00000000", 26750 => x"00000000",
    26751 => x"00000000", 26752 => x"00000000", 26753 => x"00000000",
    26754 => x"00000000", 26755 => x"00000000", 26756 => x"00000000",
    26757 => x"00000000", 26758 => x"00000000", 26759 => x"00000000",
    26760 => x"00000000", 26761 => x"00000000", 26762 => x"00000000",
    26763 => x"00000000", 26764 => x"00000000", 26765 => x"00000000",
    26766 => x"00000000", 26767 => x"00000000", 26768 => x"00000000",
    26769 => x"00000000", 26770 => x"00000000", 26771 => x"00000000",
    26772 => x"00000000", 26773 => x"00000000", 26774 => x"00000000",
    26775 => x"00000000", 26776 => x"00000000", 26777 => x"00000000",
    26778 => x"00000000", 26779 => x"00000000", 26780 => x"00000000",
    26781 => x"00000000", 26782 => x"00000000", 26783 => x"00000000",
    26784 => x"00000000", 26785 => x"00000000", 26786 => x"00000000",
    26787 => x"00000000", 26788 => x"00000000", 26789 => x"00000000",
    26790 => x"00000000", 26791 => x"00000000", 26792 => x"00000000",
    26793 => x"00000000", 26794 => x"00000000", 26795 => x"00000000",
    26796 => x"00000000", 26797 => x"00000000", 26798 => x"00000000",
    26799 => x"00000000", 26800 => x"00000000", 26801 => x"00000000",
    26802 => x"00000000", 26803 => x"00000000", 26804 => x"00000000",
    26805 => x"00000000", 26806 => x"00000000", 26807 => x"00000000",
    26808 => x"00000000", 26809 => x"00000000", 26810 => x"00000000",
    26811 => x"00000000", 26812 => x"00000000", 26813 => x"00000000",
    26814 => x"00000000", 26815 => x"00000000", 26816 => x"00000000",
    26817 => x"00000000", 26818 => x"00000000", 26819 => x"00000000",
    26820 => x"00000000", 26821 => x"00000000", 26822 => x"00000000",
    26823 => x"00000000", 26824 => x"00000000", 26825 => x"00000000",
    26826 => x"00000000", 26827 => x"00000000", 26828 => x"00000000",
    26829 => x"00000000", 26830 => x"00000000", 26831 => x"00000000",
    26832 => x"00000000", 26833 => x"00000000", 26834 => x"00000000",
    26835 => x"00000000", 26836 => x"00000000", 26837 => x"00000000",
    26838 => x"00000000", 26839 => x"00000000", 26840 => x"00000000",
    26841 => x"00000000", 26842 => x"00000000", 26843 => x"00000000",
    26844 => x"00000000", 26845 => x"00000000", 26846 => x"00000000",
    26847 => x"00000000", 26848 => x"00000000", 26849 => x"00000000",
    26850 => x"00000000", 26851 => x"00000000", 26852 => x"00000000",
    26853 => x"00000000", 26854 => x"00000000", 26855 => x"00000000",
    26856 => x"00000000", 26857 => x"00000000", 26858 => x"00000000",
    26859 => x"00000000", 26860 => x"00000000", 26861 => x"00000000",
    26862 => x"00000000", 26863 => x"00000000", 26864 => x"00000000",
    26865 => x"00000000", 26866 => x"00000000", 26867 => x"00000000",
    26868 => x"00000000", 26869 => x"00000000", 26870 => x"00000000",
    26871 => x"00000000", 26872 => x"00000000", 26873 => x"00000000",
    26874 => x"00000000", 26875 => x"00000000", 26876 => x"00000000",
    26877 => x"00000000", 26878 => x"00000000", 26879 => x"00000000",
    26880 => x"00000000", 26881 => x"00000000", 26882 => x"00000000",
    26883 => x"00000000", 26884 => x"00000000", 26885 => x"00000000",
    26886 => x"00000000", 26887 => x"00000000", 26888 => x"00000000",
    26889 => x"00000000", 26890 => x"00000000", 26891 => x"00000000",
    26892 => x"00000000", 26893 => x"00000000", 26894 => x"00000000",
    26895 => x"00000000", 26896 => x"00000000", 26897 => x"00000000",
    26898 => x"00000000", 26899 => x"00000000", 26900 => x"00000000",
    26901 => x"00000000", 26902 => x"00000000", 26903 => x"00000000",
    26904 => x"00000000", 26905 => x"00000000", 26906 => x"00000000",
    26907 => x"00000000", 26908 => x"00000000", 26909 => x"00000000",
    26910 => x"00000000", 26911 => x"00000000", 26912 => x"00000000",
    26913 => x"00000000", 26914 => x"00000000", 26915 => x"00000000",
    26916 => x"00000000", 26917 => x"00000000", 26918 => x"00000000",
    26919 => x"00000000", 26920 => x"00000000", 26921 => x"00000000",
    26922 => x"00000000", 26923 => x"00000000", 26924 => x"00000000",
    26925 => x"00000000", 26926 => x"00000000", 26927 => x"00000000",
    26928 => x"00000000", 26929 => x"00000000", 26930 => x"00000000",
    26931 => x"00000000", 26932 => x"00000000", 26933 => x"00000000",
    26934 => x"00000000", 26935 => x"00000000", 26936 => x"00000000",
    26937 => x"00000000", 26938 => x"00000000", 26939 => x"00000000",
    26940 => x"00000000", 26941 => x"00000000", 26942 => x"00000000",
    26943 => x"00000000", 26944 => x"00000000", 26945 => x"00000000",
    26946 => x"00000000", 26947 => x"00000000", 26948 => x"00000000",
    26949 => x"00000000", 26950 => x"00000000", 26951 => x"00000000",
    26952 => x"00000000", 26953 => x"00000000", 26954 => x"00000000",
    26955 => x"00000000", 26956 => x"00000000", 26957 => x"00000000",
    26958 => x"00000000", 26959 => x"00000000", 26960 => x"00000000",
    26961 => x"00000000", 26962 => x"00000000", 26963 => x"00000000",
    26964 => x"00000000", 26965 => x"00000000", 26966 => x"00000000",
    26967 => x"00000000", 26968 => x"00000000", 26969 => x"00000000",
    26970 => x"00000000", 26971 => x"00000000", 26972 => x"00000000",
    26973 => x"00000000", 26974 => x"00000000", 26975 => x"00000000",
    26976 => x"00000000", 26977 => x"00000000", 26978 => x"00000000",
    26979 => x"00000000", 26980 => x"00000000", 26981 => x"00000000",
    26982 => x"00000000", 26983 => x"00000000", 26984 => x"00000000",
    26985 => x"00000000", 26986 => x"00000000", 26987 => x"00000000",
    26988 => x"00000000", 26989 => x"00000000", 26990 => x"00000000",
    26991 => x"00000000", 26992 => x"00000000", 26993 => x"00000000",
    26994 => x"00000000", 26995 => x"00000000", 26996 => x"00000000",
    26997 => x"00000000", 26998 => x"00000000", 26999 => x"00000000",
    27000 => x"00000000", 27001 => x"00000000", 27002 => x"00000000",
    27003 => x"00000000", 27004 => x"00000000", 27005 => x"00000000",
    27006 => x"00000000", 27007 => x"00000000", 27008 => x"00000000",
    27009 => x"00000000", 27010 => x"00000000", 27011 => x"00000000",
    27012 => x"00000000", 27013 => x"00000000", 27014 => x"00000000",
    27015 => x"00000000", 27016 => x"00000000", 27017 => x"00000000",
    27018 => x"00000000", 27019 => x"00000000", 27020 => x"00000000",
    27021 => x"00000000", 27022 => x"00000000", 27023 => x"00000000",
    27024 => x"00000000", 27025 => x"00000000", 27026 => x"00000000",
    27027 => x"00000000", 27028 => x"00000000", 27029 => x"00000000",
    27030 => x"00000000", 27031 => x"00000000", 27032 => x"00000000",
    27033 => x"00000000", 27034 => x"00000000", 27035 => x"00000000",
    27036 => x"00000000", 27037 => x"00000000", 27038 => x"00000000",
    27039 => x"00000000", 27040 => x"00000000", 27041 => x"00000000",
    27042 => x"00000000", 27043 => x"00000000", 27044 => x"00000000",
    27045 => x"00000000", 27046 => x"00000000", 27047 => x"00000000",
    27048 => x"00000000", 27049 => x"00000000", 27050 => x"00000000",
    27051 => x"00000000", 27052 => x"00000000", 27053 => x"00000000",
    27054 => x"00000000", 27055 => x"00000000", 27056 => x"00000000",
    27057 => x"00000000", 27058 => x"00000000", 27059 => x"00000000",
    27060 => x"00000000", 27061 => x"00000000", 27062 => x"00000000",
    27063 => x"00000000", 27064 => x"00000000", 27065 => x"00000000",
    27066 => x"00000000", 27067 => x"00000000", 27068 => x"00000000",
    27069 => x"00000000", 27070 => x"00000000", 27071 => x"00000000",
    27072 => x"00000000", 27073 => x"00000000", 27074 => x"00000000",
    27075 => x"00000000", 27076 => x"00000000", 27077 => x"00000000",
    27078 => x"00000000", 27079 => x"00000000", 27080 => x"00000000",
    27081 => x"00000000", 27082 => x"00000000", 27083 => x"00000000",
    27084 => x"00000000", 27085 => x"00000000", 27086 => x"00000000",
    27087 => x"00000000", 27088 => x"00000000", 27089 => x"00000000",
    27090 => x"00000000", 27091 => x"00000000", 27092 => x"00000000",
    27093 => x"00000000", 27094 => x"00000000", 27095 => x"00000000",
    27096 => x"00000000", 27097 => x"00000000", 27098 => x"00000000",
    27099 => x"00000000", 27100 => x"00000000", 27101 => x"00000000",
    27102 => x"00000000", 27103 => x"00000000", 27104 => x"00000000",
    27105 => x"00000000", 27106 => x"00000000", 27107 => x"00000000",
    27108 => x"00000000", 27109 => x"00000000", 27110 => x"00000000",
    27111 => x"00000000", 27112 => x"00000000", 27113 => x"00000000",
    27114 => x"00000000", 27115 => x"00000000", 27116 => x"00000000",
    27117 => x"00000000", 27118 => x"00000000", 27119 => x"00000000",
    27120 => x"00000000", 27121 => x"00000000", 27122 => x"00000000",
    27123 => x"00000000", 27124 => x"00000000", 27125 => x"00000000",
    27126 => x"00000000", 27127 => x"00000000", 27128 => x"00000000",
    27129 => x"00000000", 27130 => x"00000000", 27131 => x"00000000",
    27132 => x"00000000", 27133 => x"00000000", 27134 => x"00000000",
    27135 => x"00000000", 27136 => x"00000000", 27137 => x"00000000",
    27138 => x"00000000", 27139 => x"00000000", 27140 => x"00000000",
    27141 => x"00000000", 27142 => x"00000000", 27143 => x"00000000",
    27144 => x"00000000", 27145 => x"00000000", 27146 => x"00000000",
    27147 => x"00000000", 27148 => x"00000000", 27149 => x"00000000",
    27150 => x"00000000", 27151 => x"00000000", 27152 => x"00000000",
    27153 => x"00000000", 27154 => x"00000000", 27155 => x"00000000",
    27156 => x"00000000", 27157 => x"00000000", 27158 => x"00000000",
    27159 => x"00000000", 27160 => x"00000000", 27161 => x"00000000",
    27162 => x"00000000", 27163 => x"00000000", 27164 => x"00000000",
    27165 => x"00000000", 27166 => x"00000000", 27167 => x"00000000",
    27168 => x"00000000", 27169 => x"00000000", 27170 => x"00000000",
    27171 => x"00000000", 27172 => x"00000000", 27173 => x"00000000",
    27174 => x"00000000", 27175 => x"00000000", 27176 => x"00000000",
    27177 => x"00000000", 27178 => x"00000000", 27179 => x"00000000",
    27180 => x"00000000", 27181 => x"00000000", 27182 => x"00000000",
    27183 => x"00000000", 27184 => x"00000000", 27185 => x"00000000",
    27186 => x"00000000", 27187 => x"00000000", 27188 => x"00000000",
    27189 => x"00000000", 27190 => x"00000000", 27191 => x"00000000",
    27192 => x"00000000", 27193 => x"00000000", 27194 => x"00000000",
    27195 => x"00000000", 27196 => x"00000000", 27197 => x"00000000",
    27198 => x"00000000", 27199 => x"00000000", 27200 => x"00000000",
    27201 => x"00000000", 27202 => x"00000000", 27203 => x"00000000",
    27204 => x"00000000", 27205 => x"00000000", 27206 => x"00000000",
    27207 => x"00000000", 27208 => x"00000000", 27209 => x"00000000",
    27210 => x"00000000", 27211 => x"00000000", 27212 => x"00000000",
    27213 => x"00000000", 27214 => x"00000000", 27215 => x"00000000",
    27216 => x"00000000", 27217 => x"00000000", 27218 => x"00000000",
    27219 => x"00000000", 27220 => x"00000000", 27221 => x"00000000",
    27222 => x"00000000", 27223 => x"00000000", 27224 => x"00000000",
    27225 => x"00000000", 27226 => x"00000000", 27227 => x"00000000",
    27228 => x"00000000", 27229 => x"00000000", 27230 => x"00000000",
    27231 => x"00000000", 27232 => x"00000000", 27233 => x"00000000",
    27234 => x"00000000", 27235 => x"00000000", 27236 => x"00000000",
    27237 => x"00000000", 27238 => x"00000000", 27239 => x"00000000",
    27240 => x"00000000", 27241 => x"00000000", 27242 => x"00000000",
    27243 => x"00000000", 27244 => x"00000000", 27245 => x"00000000",
    27246 => x"00000000", 27247 => x"00000000", 27248 => x"00000000",
    27249 => x"00000000", 27250 => x"00000000", 27251 => x"00000000",
    27252 => x"00000000", 27253 => x"00000000", 27254 => x"00000000",
    27255 => x"00000000", 27256 => x"00000000", 27257 => x"00000000",
    27258 => x"00000000", 27259 => x"00000000", 27260 => x"00000000",
    27261 => x"00000000", 27262 => x"00000000", 27263 => x"00000000",
    27264 => x"00000000", 27265 => x"00000000", 27266 => x"00000000",
    27267 => x"00000000", 27268 => x"00000000", 27269 => x"00000000",
    27270 => x"00000000", 27271 => x"00000000", 27272 => x"00000000",
    27273 => x"00000000", 27274 => x"00000000", 27275 => x"00000000",
    27276 => x"00000000", 27277 => x"00000000", 27278 => x"00000000",
    27279 => x"00000000", 27280 => x"00000000", 27281 => x"00000000",
    27282 => x"00000000", 27283 => x"00000000", 27284 => x"00000000",
    27285 => x"00000000", 27286 => x"00000000", 27287 => x"00000000",
    27288 => x"00000000", 27289 => x"00000000", 27290 => x"00000000",
    27291 => x"00000000", 27292 => x"00000000", 27293 => x"00000000",
    27294 => x"00000000", 27295 => x"00000000", 27296 => x"00000000",
    27297 => x"00000000", 27298 => x"00000000", 27299 => x"00000000",
    27300 => x"00000000", 27301 => x"00000000", 27302 => x"00000000",
    27303 => x"00000000", 27304 => x"00000000", 27305 => x"00000000",
    27306 => x"00000000", 27307 => x"00000000", 27308 => x"00000000",
    27309 => x"00000000", 27310 => x"00000000", 27311 => x"00000000",
    27312 => x"00000000", 27313 => x"00000000", 27314 => x"00000000",
    27315 => x"00000000", 27316 => x"00000000", 27317 => x"00000000",
    27318 => x"00000000", 27319 => x"00000000", 27320 => x"00000000",
    27321 => x"00000000", 27322 => x"00000000", 27323 => x"00000000",
    27324 => x"00000000", 27325 => x"00000000", 27326 => x"00000000",
    27327 => x"00000000", 27328 => x"00000000", 27329 => x"00000000",
    27330 => x"00000000", 27331 => x"00000000", 27332 => x"00000000",
    27333 => x"00000000", 27334 => x"00000000", 27335 => x"00000000",
    27336 => x"00000000", 27337 => x"00000000", 27338 => x"00000000",
    27339 => x"00000000", 27340 => x"00000000", 27341 => x"00000000",
    27342 => x"00000000", 27343 => x"00000000", 27344 => x"00000000",
    27345 => x"00000000", 27346 => x"00000000", 27347 => x"00000000",
    27348 => x"00000000", 27349 => x"00000000", 27350 => x"00000000",
    27351 => x"00000000", 27352 => x"00000000", 27353 => x"00000000",
    27354 => x"00000000", 27355 => x"00000000", 27356 => x"00000000",
    27357 => x"00000000", 27358 => x"00000000", 27359 => x"00000000",
    27360 => x"00000000", 27361 => x"00000000", 27362 => x"00000000",
    27363 => x"00000000", 27364 => x"00000000", 27365 => x"00000000",
    27366 => x"00000000", 27367 => x"00000000", 27368 => x"00000000",
    27369 => x"00000000", 27370 => x"00000000", 27371 => x"00000000",
    27372 => x"00000000", 27373 => x"00000000", 27374 => x"00000000",
    27375 => x"00000000", 27376 => x"00000000", 27377 => x"00000000",
    27378 => x"00000000", 27379 => x"00000000", 27380 => x"00000000",
    27381 => x"00000000", 27382 => x"00000000", 27383 => x"00000000",
    27384 => x"00000000", 27385 => x"00000000", 27386 => x"00000000",
    27387 => x"00000000", 27388 => x"00000000", 27389 => x"00000000",
    27390 => x"00000000", 27391 => x"00000000", 27392 => x"00000000",
    27393 => x"00000000", 27394 => x"00000000", 27395 => x"00000000",
    27396 => x"00000000", 27397 => x"00000000", 27398 => x"00000000",
    27399 => x"00000000", 27400 => x"00000000", 27401 => x"00000000",
    27402 => x"00000000", 27403 => x"00000000", 27404 => x"00000000",
    27405 => x"00000000", 27406 => x"00000000", 27407 => x"00000000",
    27408 => x"00000000", 27409 => x"00000000", 27410 => x"00000000",
    27411 => x"00000000", 27412 => x"00000000", 27413 => x"00000000",
    27414 => x"00000000", 27415 => x"00000000", 27416 => x"00000000",
    27417 => x"00000000", 27418 => x"00000000", 27419 => x"00000000",
    27420 => x"00000000", 27421 => x"00000000", 27422 => x"00000000",
    27423 => x"00000000", 27424 => x"00000000", 27425 => x"00000000",
    27426 => x"00000000", 27427 => x"00000000", 27428 => x"00000000",
    27429 => x"00000000", 27430 => x"00000000", 27431 => x"00000000",
    27432 => x"00000000", 27433 => x"00000000", 27434 => x"00000000",
    27435 => x"00000000", 27436 => x"00000000", 27437 => x"00000000",
    27438 => x"00000000", 27439 => x"00000000", 27440 => x"00000000",
    27441 => x"00000000", 27442 => x"00000000", 27443 => x"00000000",
    27444 => x"00000000", 27445 => x"00000000", 27446 => x"00000000",
    27447 => x"00000000", 27448 => x"00000000", 27449 => x"00000000",
    27450 => x"00000000", 27451 => x"00000000", 27452 => x"00000000",
    27453 => x"00000000", 27454 => x"00000000", 27455 => x"00000000",
    27456 => x"00000000", 27457 => x"00000000", 27458 => x"00000000",
    27459 => x"00000000", 27460 => x"00000000", 27461 => x"00000000",
    27462 => x"00000000", 27463 => x"00000000", 27464 => x"00000000",
    27465 => x"00000000", 27466 => x"00000000", 27467 => x"00000000",
    27468 => x"00000000", 27469 => x"00000000", 27470 => x"00000000",
    27471 => x"00000000", 27472 => x"00000000", 27473 => x"00000000",
    27474 => x"00000000", 27475 => x"00000000", 27476 => x"00000000",
    27477 => x"00000000", 27478 => x"00000000", 27479 => x"00000000",
    27480 => x"00000000", 27481 => x"00000000", 27482 => x"00000000",
    27483 => x"00000000", 27484 => x"00000000", 27485 => x"00000000",
    27486 => x"00000000", 27487 => x"00000000", 27488 => x"00000000",
    27489 => x"00000000", 27490 => x"00000000", 27491 => x"00000000",
    27492 => x"00000000", 27493 => x"00000000", 27494 => x"00000000",
    27495 => x"00000000", 27496 => x"00000000", 27497 => x"00000000",
    27498 => x"00000000", 27499 => x"00000000", 27500 => x"00000000",
    27501 => x"00000000", 27502 => x"00000000", 27503 => x"00000000",
    27504 => x"00000000", 27505 => x"00000000", 27506 => x"00000000",
    27507 => x"00000000", 27508 => x"00000000", 27509 => x"00000000",
    27510 => x"00000000", 27511 => x"00000000", 27512 => x"00000000",
    27513 => x"00000000", 27514 => x"00000000", 27515 => x"00000000",
    27516 => x"00000000", 27517 => x"00000000", 27518 => x"00000000",
    27519 => x"00000000", 27520 => x"00000000", 27521 => x"00000000",
    27522 => x"00000000", 27523 => x"00000000", 27524 => x"00000000",
    27525 => x"00000000", 27526 => x"00000000", 27527 => x"00000000",
    27528 => x"00000000", 27529 => x"00000000", 27530 => x"00000000",
    27531 => x"00000000", 27532 => x"00000000", 27533 => x"00000000",
    27534 => x"00000000", 27535 => x"00000000", 27536 => x"00000000",
    27537 => x"00000000", 27538 => x"00000000", 27539 => x"00000000",
    27540 => x"00000000", 27541 => x"00000000", 27542 => x"00000000",
    27543 => x"00000000", 27544 => x"00000000", 27545 => x"00000000",
    27546 => x"00000000", 27547 => x"00000000", 27548 => x"00000000",
    27549 => x"00000000", 27550 => x"00000000", 27551 => x"00000000",
    27552 => x"00000000", 27553 => x"00000000", 27554 => x"00000000",
    27555 => x"00000000", 27556 => x"00000000", 27557 => x"00000000",
    27558 => x"00000000", 27559 => x"00000000", 27560 => x"00000000",
    27561 => x"00000000", 27562 => x"00000000", 27563 => x"00000000",
    27564 => x"00000000", 27565 => x"00000000", 27566 => x"00000000",
    27567 => x"00000000", 27568 => x"00000000", 27569 => x"00000000",
    27570 => x"00000000", 27571 => x"00000000", 27572 => x"00000000",
    27573 => x"00000000", 27574 => x"00000000", 27575 => x"00000000",
    27576 => x"00000000", 27577 => x"00000000", 27578 => x"00000000",
    27579 => x"00000000", 27580 => x"00000000", 27581 => x"00000000",
    27582 => x"00000000", 27583 => x"00000000", 27584 => x"00000000",
    27585 => x"00000000", 27586 => x"00000000", 27587 => x"00000000",
    27588 => x"00000000", 27589 => x"00000000", 27590 => x"00000000",
    27591 => x"00000000", 27592 => x"00000000", 27593 => x"00000000",
    27594 => x"00000000", 27595 => x"00000000", 27596 => x"00000000",
    27597 => x"00000000", 27598 => x"00000000", 27599 => x"00000000",
    27600 => x"00000000", 27601 => x"00000000", 27602 => x"00000000",
    27603 => x"00000000", 27604 => x"00000000", 27605 => x"00000000",
    27606 => x"00000000", 27607 => x"00000000", 27608 => x"00000000",
    27609 => x"00000000", 27610 => x"00000000", 27611 => x"00000000",
    27612 => x"00000000", 27613 => x"00000000", 27614 => x"00000000",
    27615 => x"00000000", 27616 => x"00000000", 27617 => x"00000000",
    27618 => x"00000000", 27619 => x"00000000", 27620 => x"00000000",
    27621 => x"00000000", 27622 => x"00000000", 27623 => x"00000000",
    27624 => x"00000000", 27625 => x"00000000", 27626 => x"00000000",
    27627 => x"00000000", 27628 => x"00000000", 27629 => x"00000000",
    27630 => x"00000000", 27631 => x"00000000", 27632 => x"00000000",
    27633 => x"00000000", 27634 => x"00000000", 27635 => x"00000000",
    27636 => x"00000000", 27637 => x"00000000", 27638 => x"00000000",
    27639 => x"00000000", 27640 => x"00000000", 27641 => x"00000000",
    27642 => x"00000000", 27643 => x"00000000", 27644 => x"00000000",
    27645 => x"00000000", 27646 => x"00000000", 27647 => x"00000000",
    27648 => x"00000000", 27649 => x"00000000", 27650 => x"00000000",
    27651 => x"00000000", 27652 => x"00000000", 27653 => x"00000000",
    27654 => x"00000000", 27655 => x"00000000", 27656 => x"00000000",
    27657 => x"00000000", 27658 => x"00000000", 27659 => x"00000000",
    27660 => x"00000000", 27661 => x"00000000", 27662 => x"00000000",
    27663 => x"00000000", 27664 => x"00000000", 27665 => x"00000000",
    27666 => x"00000000", 27667 => x"00000000", 27668 => x"00000000",
    27669 => x"00000000", 27670 => x"00000000", 27671 => x"00000000",
    27672 => x"00000000", 27673 => x"00000000", 27674 => x"00000000",
    27675 => x"00000000", 27676 => x"00000000", 27677 => x"00000000",
    27678 => x"00000000", 27679 => x"00000000", 27680 => x"00000000",
    27681 => x"00000000", 27682 => x"00000000", 27683 => x"00000000",
    27684 => x"00000000", 27685 => x"00000000", 27686 => x"00000000",
    27687 => x"00000000", 27688 => x"00000000", 27689 => x"00000000",
    27690 => x"00000000", 27691 => x"00000000", 27692 => x"00000000",
    27693 => x"00000000", 27694 => x"00000000", 27695 => x"00000000",
    27696 => x"00000000", 27697 => x"00000000", 27698 => x"00000000",
    27699 => x"00000000", 27700 => x"00000000", 27701 => x"00000000",
    27702 => x"00000000", 27703 => x"00000000", 27704 => x"00000000",
    27705 => x"00000000", 27706 => x"00000000", 27707 => x"00000000",
    27708 => x"00000000", 27709 => x"00000000", 27710 => x"00000000",
    27711 => x"00000000", 27712 => x"00000000", 27713 => x"00000000",
    27714 => x"00000000", 27715 => x"00000000", 27716 => x"00000000",
    27717 => x"00000000", 27718 => x"00000000", 27719 => x"00000000",
    27720 => x"00000000", 27721 => x"00000000", 27722 => x"00000000",
    27723 => x"00000000", 27724 => x"00000000", 27725 => x"00000000",
    27726 => x"00000000", 27727 => x"00000000", 27728 => x"00000000",
    27729 => x"00000000", 27730 => x"00000000", 27731 => x"00000000",
    27732 => x"00000000", 27733 => x"00000000", 27734 => x"00000000",
    27735 => x"00000000", 27736 => x"00000000", 27737 => x"00000000",
    27738 => x"00000000", 27739 => x"00000000", 27740 => x"00000000",
    27741 => x"00000000", 27742 => x"00000000", 27743 => x"00000000",
    27744 => x"00000000", 27745 => x"00000000", 27746 => x"00000000",
    27747 => x"00000000", 27748 => x"00000000", 27749 => x"00000000",
    27750 => x"00000000", 27751 => x"00000000", 27752 => x"00000000",
    27753 => x"00000000", 27754 => x"00000000", 27755 => x"00000000",
    27756 => x"00000000", 27757 => x"00000000", 27758 => x"00000000",
    27759 => x"00000000", 27760 => x"00000000", 27761 => x"00000000",
    27762 => x"00000000", 27763 => x"00000000", 27764 => x"00000000",
    27765 => x"00000000", 27766 => x"00000000", 27767 => x"00000000",
    27768 => x"00000000", 27769 => x"00000000", 27770 => x"00000000",
    27771 => x"00000000", 27772 => x"00000000", 27773 => x"00000000",
    27774 => x"00000000", 27775 => x"00000000", 27776 => x"00000000",
    27777 => x"00000000", 27778 => x"00000000", 27779 => x"00000000",
    27780 => x"00000000", 27781 => x"00000000", 27782 => x"00000000",
    27783 => x"00000000", 27784 => x"00000000", 27785 => x"00000000",
    27786 => x"00000000", 27787 => x"00000000", 27788 => x"00000000",
    27789 => x"00000000", 27790 => x"00000000", 27791 => x"00000000",
    27792 => x"00000000", 27793 => x"00000000", 27794 => x"00000000",
    27795 => x"00000000", 27796 => x"00000000", 27797 => x"00000000",
    27798 => x"00000000", 27799 => x"00000000", 27800 => x"00000000",
    27801 => x"00000000", 27802 => x"00000000", 27803 => x"00000000",
    27804 => x"00000000", 27805 => x"00000000", 27806 => x"00000000",
    27807 => x"00000000", 27808 => x"00000000", 27809 => x"00000000",
    27810 => x"00000000", 27811 => x"00000000", 27812 => x"00000000",
    27813 => x"00000000", 27814 => x"00000000", 27815 => x"00000000",
    27816 => x"00000000", 27817 => x"00000000", 27818 => x"00000000",
    27819 => x"00000000", 27820 => x"00000000", 27821 => x"00000000",
    27822 => x"00000000", 27823 => x"00000000", 27824 => x"00000000",
    27825 => x"00000000", 27826 => x"00000000", 27827 => x"00000000",
    27828 => x"00000000", 27829 => x"00000000", 27830 => x"00000000",
    27831 => x"00000000", 27832 => x"00000000", 27833 => x"00000000",
    27834 => x"00000000", 27835 => x"00000000", 27836 => x"00000000",
    27837 => x"00000000", 27838 => x"00000000", 27839 => x"00000000",
    27840 => x"00000000", 27841 => x"00000000", 27842 => x"00000000",
    27843 => x"00000000", 27844 => x"00000000", 27845 => x"00000000",
    27846 => x"00000000", 27847 => x"00000000", 27848 => x"00000000",
    27849 => x"00000000", 27850 => x"00000000", 27851 => x"00000000",
    27852 => x"00000000", 27853 => x"00000000", 27854 => x"00000000",
    27855 => x"00000000", 27856 => x"00000000", 27857 => x"00000000",
    27858 => x"00000000", 27859 => x"00000000", 27860 => x"00000000",
    27861 => x"00000000", 27862 => x"00000000", 27863 => x"00000000",
    27864 => x"00000000", 27865 => x"00000000", 27866 => x"00000000",
    27867 => x"00000000", 27868 => x"00000000", 27869 => x"00000000",
    27870 => x"00000000", 27871 => x"00000000", 27872 => x"00000000",
    27873 => x"00000000", 27874 => x"00000000", 27875 => x"00000000",
    27876 => x"00000000", 27877 => x"00000000", 27878 => x"00000000",
    27879 => x"00000000", 27880 => x"00000000", 27881 => x"00000000",
    27882 => x"00000000", 27883 => x"00000000", 27884 => x"00000000",
    27885 => x"00000000", 27886 => x"00000000", 27887 => x"00000000",
    27888 => x"00000000", 27889 => x"00000000", 27890 => x"00000000",
    27891 => x"00000000", 27892 => x"00000000", 27893 => x"00000000",
    27894 => x"00000000", 27895 => x"00000000", 27896 => x"00000000",
    27897 => x"00000000", 27898 => x"00000000", 27899 => x"00000000",
    27900 => x"00000000", 27901 => x"00000000", 27902 => x"00000000",
    27903 => x"00000000", 27904 => x"00000000", 27905 => x"00000000",
    27906 => x"00000000", 27907 => x"00000000", 27908 => x"00000000",
    27909 => x"00000000", 27910 => x"00000000", 27911 => x"00000000",
    27912 => x"00000000", 27913 => x"00000000", 27914 => x"00000000",
    27915 => x"00000000", 27916 => x"00000000", 27917 => x"00000000",
    27918 => x"00000000", 27919 => x"00000000", 27920 => x"00000000",
    27921 => x"00000000", 27922 => x"00000000", 27923 => x"00000000",
    27924 => x"00000000", 27925 => x"00000000", 27926 => x"00000000",
    27927 => x"00000000", 27928 => x"00000000", 27929 => x"00000000",
    27930 => x"00000000", 27931 => x"00000000", 27932 => x"00000000",
    27933 => x"00000000", 27934 => x"00000000", 27935 => x"00000000",
    27936 => x"00000000", 27937 => x"00000000", 27938 => x"00000000",
    27939 => x"00000000", 27940 => x"00000000", 27941 => x"00000000",
    27942 => x"00000000", 27943 => x"00000000", 27944 => x"00000000",
    27945 => x"00000000", 27946 => x"00000000", 27947 => x"00000000",
    27948 => x"00000000", 27949 => x"00000000", 27950 => x"00000000",
    27951 => x"00000000", 27952 => x"00000000", 27953 => x"00000000",
    27954 => x"00000000", 27955 => x"00000000", 27956 => x"00000000",
    27957 => x"00000000", 27958 => x"00000000", 27959 => x"00000000",
    27960 => x"00000000", 27961 => x"00000000", 27962 => x"00000000",
    27963 => x"00000000", 27964 => x"00000000", 27965 => x"00000000",
    27966 => x"00000000", 27967 => x"00000000", 27968 => x"00000000",
    27969 => x"00000000", 27970 => x"00000000", 27971 => x"00000000",
    27972 => x"00000000", 27973 => x"00000000", 27974 => x"00000000",
    27975 => x"00000000", 27976 => x"00000000", 27977 => x"00000000",
    27978 => x"00000000", 27979 => x"00000000", 27980 => x"00000000",
    27981 => x"00000000", 27982 => x"00000000", 27983 => x"00000000",
    27984 => x"00000000", 27985 => x"00000000", 27986 => x"00000000",
    27987 => x"00000000", 27988 => x"00000000", 27989 => x"00000000",
    27990 => x"00000000", 27991 => x"00000000", 27992 => x"00000000",
    27993 => x"00000000", 27994 => x"00000000", 27995 => x"00000000",
    27996 => x"00000000", 27997 => x"00000000", 27998 => x"00000000",
    27999 => x"00000000", 28000 => x"00000000", 28001 => x"00000000",
    28002 => x"00000000", 28003 => x"00000000", 28004 => x"00000000",
    28005 => x"00000000", 28006 => x"00000000", 28007 => x"00000000",
    28008 => x"00000000", 28009 => x"00000000", 28010 => x"00000000",
    28011 => x"00000000", 28012 => x"00000000", 28013 => x"00000000",
    28014 => x"00000000", 28015 => x"00000000", 28016 => x"00000000",
    28017 => x"00000000", 28018 => x"00000000", 28019 => x"00000000",
    28020 => x"00000000", 28021 => x"00000000", 28022 => x"00000000",
    28023 => x"00000000", 28024 => x"00000000", 28025 => x"00000000",
    28026 => x"00000000", 28027 => x"00000000", 28028 => x"00000000",
    28029 => x"00000000", 28030 => x"00000000", 28031 => x"00000000",
    28032 => x"00000000", 28033 => x"00000000", 28034 => x"00000000",
    28035 => x"00000000", 28036 => x"00000000", 28037 => x"00000000",
    28038 => x"00000000", 28039 => x"00000000", 28040 => x"00000000",
    28041 => x"00000000", 28042 => x"00000000", 28043 => x"00000000",
    28044 => x"00000000", 28045 => x"00000000", 28046 => x"00000000",
    28047 => x"00000000", 28048 => x"00000000", 28049 => x"00000000",
    28050 => x"00000000", 28051 => x"00000000", 28052 => x"00000000",
    28053 => x"00000000", 28054 => x"00000000", 28055 => x"00000000",
    28056 => x"00000000", 28057 => x"00000000", 28058 => x"00000000",
    28059 => x"00000000", 28060 => x"00000000", 28061 => x"00000000",
    28062 => x"00000000", 28063 => x"00000000", 28064 => x"00000000",
    28065 => x"00000000", 28066 => x"00000000", 28067 => x"00000000",
    28068 => x"00000000", 28069 => x"00000000", 28070 => x"00000000",
    28071 => x"00000000", 28072 => x"00000000", 28073 => x"00000000",
    28074 => x"00000000", 28075 => x"00000000", 28076 => x"00000000",
    28077 => x"00000000", 28078 => x"00000000", 28079 => x"00000000",
    28080 => x"00000000", 28081 => x"00000000", 28082 => x"00000000",
    28083 => x"00000000", 28084 => x"00000000", 28085 => x"00000000",
    28086 => x"00000000", 28087 => x"00000000", 28088 => x"00000000",
    28089 => x"00000000", 28090 => x"00000000", 28091 => x"00000000",
    28092 => x"00000000", 28093 => x"00000000", 28094 => x"00000000",
    28095 => x"00000000", 28096 => x"00000000", 28097 => x"00000000",
    28098 => x"00000000", 28099 => x"00000000", 28100 => x"00000000",
    28101 => x"00000000", 28102 => x"00000000", 28103 => x"00000000",
    28104 => x"00000000", 28105 => x"00000000", 28106 => x"00000000",
    28107 => x"00000000", 28108 => x"00000000", 28109 => x"00000000",
    28110 => x"00000000", 28111 => x"00000000", 28112 => x"00000000",
    28113 => x"00000000", 28114 => x"00000000", 28115 => x"00000000",
    28116 => x"00000000", 28117 => x"00000000", 28118 => x"00000000",
    28119 => x"00000000", 28120 => x"00000000", 28121 => x"00000000",
    28122 => x"00000000", 28123 => x"00000000", 28124 => x"00000000",
    28125 => x"00000000", 28126 => x"00000000", 28127 => x"00000000",
    28128 => x"00000000", 28129 => x"00000000", 28130 => x"00000000",
    28131 => x"00000000", 28132 => x"00000000", 28133 => x"00000000",
    28134 => x"00000000", 28135 => x"00000000", 28136 => x"00000000",
    28137 => x"00000000", 28138 => x"00000000", 28139 => x"00000000",
    28140 => x"00000000", 28141 => x"00000000", 28142 => x"00000000",
    28143 => x"00000000", 28144 => x"00000000", 28145 => x"00000000",
    28146 => x"00000000", 28147 => x"00000000", 28148 => x"00000000",
    28149 => x"00000000", 28150 => x"00000000", 28151 => x"00000000",
    28152 => x"00000000", 28153 => x"00000000", 28154 => x"00000000",
    28155 => x"00000000", 28156 => x"00000000", 28157 => x"00000000",
    28158 => x"00000000", 28159 => x"00000000", 28160 => x"00000000",
    28161 => x"00000000", 28162 => x"00000000", 28163 => x"00000000",
    28164 => x"00000000", 28165 => x"00000000", 28166 => x"00000000",
    28167 => x"00000000", 28168 => x"00000000", 28169 => x"00000000",
    28170 => x"00000000", 28171 => x"00000000", 28172 => x"00000000",
    28173 => x"00000000", 28174 => x"00000000", 28175 => x"00000000",
    28176 => x"00000000", 28177 => x"00000000", 28178 => x"00000000",
    28179 => x"00000000", 28180 => x"00000000", 28181 => x"00000000",
    28182 => x"00000000", 28183 => x"00000000", 28184 => x"00000000",
    28185 => x"00000000", 28186 => x"00000000", 28187 => x"00000000",
    28188 => x"00000000", 28189 => x"00000000", 28190 => x"00000000",
    28191 => x"00000000", 28192 => x"00000000", 28193 => x"00000000",
    28194 => x"00000000", 28195 => x"00000000", 28196 => x"00000000",
    28197 => x"00000000", 28198 => x"00000000", 28199 => x"00000000",
    28200 => x"00000000", 28201 => x"00000000", 28202 => x"00000000",
    28203 => x"00000000", 28204 => x"00000000", 28205 => x"00000000",
    28206 => x"00000000", 28207 => x"00000000", 28208 => x"00000000",
    28209 => x"00000000", 28210 => x"00000000", 28211 => x"00000000",
    28212 => x"00000000", 28213 => x"00000000", 28214 => x"00000000",
    28215 => x"00000000", 28216 => x"00000000", 28217 => x"00000000",
    28218 => x"00000000", 28219 => x"00000000", 28220 => x"00000000",
    28221 => x"00000000", 28222 => x"00000000", 28223 => x"00000000",
    28224 => x"00000000", 28225 => x"00000000", 28226 => x"00000000",
    28227 => x"00000000", 28228 => x"00000000", 28229 => x"00000000",
    28230 => x"00000000", 28231 => x"00000000", 28232 => x"00000000",
    28233 => x"00000000", 28234 => x"00000000", 28235 => x"00000000",
    28236 => x"00000000", 28237 => x"00000000", 28238 => x"00000000",
    28239 => x"00000000", 28240 => x"00000000", 28241 => x"00000000",
    28242 => x"00000000", 28243 => x"00000000", 28244 => x"00000000",
    28245 => x"00000000", 28246 => x"00000000", 28247 => x"00000000",
    28248 => x"00000000", 28249 => x"00000000", 28250 => x"00000000",
    28251 => x"00000000", 28252 => x"00000000", 28253 => x"00000000",
    28254 => x"00000000", 28255 => x"00000000", 28256 => x"00000000",
    28257 => x"00000000", 28258 => x"00000000", 28259 => x"00000000",
    28260 => x"00000000", 28261 => x"00000000", 28262 => x"00000000",
    28263 => x"00000000", 28264 => x"00000000", 28265 => x"00000000",
    28266 => x"00000000", 28267 => x"00000000", 28268 => x"00000000",
    28269 => x"00000000", 28270 => x"00000000", 28271 => x"00000000",
    28272 => x"00000000", 28273 => x"00000000", 28274 => x"00000000",
    28275 => x"00000000", 28276 => x"00000000", 28277 => x"00000000",
    28278 => x"00000000", 28279 => x"00000000", 28280 => x"00000000",
    28281 => x"00000000", 28282 => x"00000000", 28283 => x"00000000",
    28284 => x"00000000", 28285 => x"00000000", 28286 => x"00000000",
    28287 => x"00000000", 28288 => x"00000000", 28289 => x"00000000",
    28290 => x"00000000", 28291 => x"00000000", 28292 => x"00000000",
    28293 => x"00000000", 28294 => x"00000000", 28295 => x"00000000",
    28296 => x"00000000", 28297 => x"00000000", 28298 => x"00000000",
    28299 => x"00000000", 28300 => x"00000000", 28301 => x"00000000",
    28302 => x"00000000", 28303 => x"00000000", 28304 => x"00000000",
    28305 => x"00000000", 28306 => x"00000000", 28307 => x"00000000",
    28308 => x"00000000", 28309 => x"00000000", 28310 => x"00000000",
    28311 => x"00000000", 28312 => x"00000000", 28313 => x"00000000",
    28314 => x"00000000", 28315 => x"00000000", 28316 => x"00000000",
    28317 => x"00000000", 28318 => x"00000000", 28319 => x"00000000",
    28320 => x"00000000", 28321 => x"00000000", 28322 => x"00000000",
    28323 => x"00000000", 28324 => x"00000000", 28325 => x"00000000",
    28326 => x"00000000", 28327 => x"00000000", 28328 => x"00000000",
    28329 => x"00000000", 28330 => x"00000000", 28331 => x"00000000",
    28332 => x"00000000", 28333 => x"00000000", 28334 => x"00000000",
    28335 => x"00000000", 28336 => x"00000000", 28337 => x"00000000",
    28338 => x"00000000", 28339 => x"00000000", 28340 => x"00000000",
    28341 => x"00000000", 28342 => x"00000000", 28343 => x"00000000",
    28344 => x"00000000", 28345 => x"00000000", 28346 => x"00000000",
    28347 => x"00000000", 28348 => x"00000000", 28349 => x"00000000",
    28350 => x"00000000", 28351 => x"00000000", 28352 => x"00000000",
    28353 => x"00000000", 28354 => x"00000000", 28355 => x"00000000",
    28356 => x"00000000", 28357 => x"00000000", 28358 => x"00000000",
    28359 => x"00000000", 28360 => x"00000000", 28361 => x"00000000",
    28362 => x"00000000", 28363 => x"00000000", 28364 => x"00000000",
    28365 => x"00000000", 28366 => x"00000000", 28367 => x"00000000",
    28368 => x"00000000", 28369 => x"00000000", 28370 => x"00000000",
    28371 => x"00000000", 28372 => x"00000000", 28373 => x"00000000",
    28374 => x"00000000", 28375 => x"00000000", 28376 => x"00000000",
    28377 => x"00000000", 28378 => x"00000000", 28379 => x"00000000",
    28380 => x"00000000", 28381 => x"00000000", 28382 => x"00000000",
    28383 => x"00000000", 28384 => x"00000000", 28385 => x"00000000",
    28386 => x"00000000", 28387 => x"00000000", 28388 => x"00000000",
    28389 => x"00000000", 28390 => x"00000000", 28391 => x"00000000",
    28392 => x"00000000", 28393 => x"00000000", 28394 => x"00000000",
    28395 => x"00000000", 28396 => x"00000000", 28397 => x"00000000",
    28398 => x"00000000", 28399 => x"00000000", 28400 => x"00000000",
    28401 => x"00000000", 28402 => x"00000000", 28403 => x"00000000",
    28404 => x"00000000", 28405 => x"00000000", 28406 => x"00000000",
    28407 => x"00000000", 28408 => x"00000000", 28409 => x"00000000",
    28410 => x"00000000", 28411 => x"00000000", 28412 => x"00000000",
    28413 => x"00000000", 28414 => x"00000000", 28415 => x"00000000",
    28416 => x"00000000", 28417 => x"00000000", 28418 => x"00000000",
    28419 => x"00000000", 28420 => x"00000000", 28421 => x"00000000",
    28422 => x"00000000", 28423 => x"00000000", 28424 => x"00000000",
    28425 => x"00000000", 28426 => x"00000000", 28427 => x"00000000",
    28428 => x"00000000", 28429 => x"00000000", 28430 => x"00000000",
    28431 => x"00000000", 28432 => x"00000000", 28433 => x"00000000",
    28434 => x"00000000", 28435 => x"00000000", 28436 => x"00000000",
    28437 => x"00000000", 28438 => x"00000000", 28439 => x"00000000",
    28440 => x"00000000", 28441 => x"00000000", 28442 => x"00000000",
    28443 => x"00000000", 28444 => x"00000000", 28445 => x"00000000",
    28446 => x"00000000", 28447 => x"00000000", 28448 => x"00000000",
    28449 => x"00000000", 28450 => x"00000000", 28451 => x"00000000",
    28452 => x"00000000", 28453 => x"00000000", 28454 => x"00000000",
    28455 => x"00000000", 28456 => x"00000000", 28457 => x"00000000",
    28458 => x"00000000", 28459 => x"00000000", 28460 => x"00000000",
    28461 => x"00000000", 28462 => x"00000000", 28463 => x"00000000",
    28464 => x"00000000", 28465 => x"00000000", 28466 => x"00000000",
    28467 => x"00000000", 28468 => x"00000000", 28469 => x"00000000",
    28470 => x"00000000", 28471 => x"00000000", 28472 => x"00000000",
    28473 => x"00000000", 28474 => x"00000000", 28475 => x"00000000",
    28476 => x"00000000", 28477 => x"00000000", 28478 => x"00000000",
    28479 => x"00000000", 28480 => x"00000000", 28481 => x"00000000",
    28482 => x"00000000", 28483 => x"00000000", 28484 => x"00000000",
    28485 => x"00000000", 28486 => x"00000000", 28487 => x"00000000",
    28488 => x"00000000", 28489 => x"00000000", 28490 => x"00000000",
    28491 => x"00000000", 28492 => x"00000000", 28493 => x"00000000",
    28494 => x"00000000", 28495 => x"00000000", 28496 => x"00000000",
    28497 => x"00000000", 28498 => x"00000000", 28499 => x"00000000",
    28500 => x"00000000", 28501 => x"00000000", 28502 => x"00000000",
    28503 => x"00000000", 28504 => x"00000000", 28505 => x"00000000",
    28506 => x"00000000", 28507 => x"00000000", 28508 => x"00000000",
    28509 => x"00000000", 28510 => x"00000000", 28511 => x"00000000",
    28512 => x"00000000", 28513 => x"00000000", 28514 => x"00000000",
    28515 => x"00000000", 28516 => x"00000000", 28517 => x"00000000",
    28518 => x"00000000", 28519 => x"00000000", 28520 => x"00000000",
    28521 => x"00000000", 28522 => x"00000000", 28523 => x"00000000",
    28524 => x"00000000", 28525 => x"00000000", 28526 => x"00000000",
    28527 => x"00000000", 28528 => x"00000000", 28529 => x"00000000",
    28530 => x"00000000", 28531 => x"00000000", 28532 => x"00000000",
    28533 => x"00000000", 28534 => x"00000000", 28535 => x"00000000",
    28536 => x"00000000", 28537 => x"00000000", 28538 => x"00000000",
    28539 => x"00000000", 28540 => x"00000000", 28541 => x"00000000",
    28542 => x"00000000", 28543 => x"00000000", 28544 => x"00000000",
    28545 => x"00000000", 28546 => x"00000000", 28547 => x"00000000",
    28548 => x"00000000", 28549 => x"00000000", 28550 => x"00000000",
    28551 => x"00000000", 28552 => x"00000000", 28553 => x"00000000",
    28554 => x"00000000", 28555 => x"00000000", 28556 => x"00000000",
    28557 => x"00000000", 28558 => x"00000000", 28559 => x"00000000",
    28560 => x"00000000", 28561 => x"00000000", 28562 => x"00000000",
    28563 => x"00000000", 28564 => x"00000000", 28565 => x"00000000",
    28566 => x"00000000", 28567 => x"00000000", 28568 => x"00000000",
    28569 => x"00000000", 28570 => x"00000000", 28571 => x"00000000",
    28572 => x"00000000", 28573 => x"00000000", 28574 => x"00000000",
    28575 => x"00000000", 28576 => x"00000000", 28577 => x"00000000",
    28578 => x"00000000", 28579 => x"00000000", 28580 => x"00000000",
    28581 => x"00000000", 28582 => x"00000000", 28583 => x"00000000",
    28584 => x"00000000", 28585 => x"00000000", 28586 => x"00000000",
    28587 => x"00000000", 28588 => x"00000000", 28589 => x"00000000",
    28590 => x"00000000", 28591 => x"00000000", 28592 => x"00000000",
    28593 => x"00000000", 28594 => x"00000000", 28595 => x"00000000",
    28596 => x"00000000", 28597 => x"00000000", 28598 => x"00000000",
    28599 => x"00000000", 28600 => x"00000000", 28601 => x"00000000",
    28602 => x"00000000", 28603 => x"00000000", 28604 => x"00000000",
    28605 => x"00000000", 28606 => x"00000000", 28607 => x"00000000",
    28608 => x"00000000", 28609 => x"00000000", 28610 => x"00000000",
    28611 => x"00000000", 28612 => x"00000000", 28613 => x"00000000",
    28614 => x"00000000", 28615 => x"00000000", 28616 => x"00000000",
    28617 => x"00000000", 28618 => x"00000000", 28619 => x"00000000",
    28620 => x"00000000", 28621 => x"00000000", 28622 => x"00000000",
    28623 => x"00000000", 28624 => x"00000000", 28625 => x"00000000",
    28626 => x"00000000", 28627 => x"00000000", 28628 => x"00000000",
    28629 => x"00000000", 28630 => x"00000000", 28631 => x"00000000",
    28632 => x"00000000", 28633 => x"00000000", 28634 => x"00000000",
    28635 => x"00000000", 28636 => x"00000000", 28637 => x"00000000",
    28638 => x"00000000", 28639 => x"00000000", 28640 => x"00000000",
    28641 => x"00000000", 28642 => x"00000000", 28643 => x"00000000",
    28644 => x"00000000", 28645 => x"00000000", 28646 => x"00000000",
    28647 => x"00000000", 28648 => x"00000000", 28649 => x"00000000",
    28650 => x"00000000", 28651 => x"00000000", 28652 => x"00000000",
    28653 => x"00000000", 28654 => x"00000000", 28655 => x"00000000",
    28656 => x"00000000", 28657 => x"00000000", 28658 => x"00000000",
    28659 => x"00000000", 28660 => x"00000000", 28661 => x"00000000",
    28662 => x"00000000", 28663 => x"00000000", 28664 => x"00000000",
    28665 => x"00000000", 28666 => x"00000000", 28667 => x"00000000",
    28668 => x"00000000", 28669 => x"00000000", 28670 => x"00000000",
    28671 => x"00000000", 28672 => x"00000000", 28673 => x"00000000",
    28674 => x"00000000", 28675 => x"00000000", 28676 => x"00000000",
    28677 => x"00000000", 28678 => x"00000000", 28679 => x"00000000",
    28680 => x"00000000", 28681 => x"00000000", 28682 => x"00000000",
    28683 => x"00000000", 28684 => x"00000000", 28685 => x"00000000",
    28686 => x"00000000", 28687 => x"00000000", 28688 => x"00000000",
    28689 => x"00000000", 28690 => x"00000000", 28691 => x"00000000",
    28692 => x"00000000", 28693 => x"00000000", 28694 => x"00000000",
    28695 => x"00000000", 28696 => x"00000000", 28697 => x"00000000",
    28698 => x"00000000", 28699 => x"00000000", 28700 => x"00000000",
    28701 => x"00000000", 28702 => x"00000000", 28703 => x"00000000",
    28704 => x"00000000", 28705 => x"00000000", 28706 => x"00000000",
    28707 => x"00000000", 28708 => x"00000000", 28709 => x"00000000",
    28710 => x"00000000", 28711 => x"00000000", 28712 => x"00000000",
    28713 => x"00000000", 28714 => x"00000000", 28715 => x"00000000",
    28716 => x"00000000", 28717 => x"00000000", 28718 => x"00000000",
    28719 => x"00000000", 28720 => x"00000000", 28721 => x"00000000",
    28722 => x"00000000", 28723 => x"00000000", 28724 => x"00000000",
    28725 => x"00000000", 28726 => x"00000000", 28727 => x"00000000",
    28728 => x"00000000", 28729 => x"00000000", 28730 => x"00000000",
    28731 => x"00000000", 28732 => x"00000000", 28733 => x"00000000",
    28734 => x"00000000", 28735 => x"00000000", 28736 => x"00000000",
    28737 => x"00000000", 28738 => x"00000000", 28739 => x"00000000",
    28740 => x"00000000", 28741 => x"00000000", 28742 => x"00000000",
    28743 => x"00000000", 28744 => x"00000000", 28745 => x"00000000",
    28746 => x"00000000", 28747 => x"00000000", 28748 => x"00000000",
    28749 => x"00000000", 28750 => x"00000000", 28751 => x"00000000",
    28752 => x"00000000", 28753 => x"00000000", 28754 => x"00000000",
    28755 => x"00000000", 28756 => x"00000000", 28757 => x"00000000",
    28758 => x"00000000", 28759 => x"00000000", 28760 => x"00000000",
    28761 => x"00000000", 28762 => x"00000000", 28763 => x"00000000",
    28764 => x"00000000", 28765 => x"00000000", 28766 => x"00000000",
    28767 => x"00000000", 28768 => x"00000000", 28769 => x"00000000",
    28770 => x"00000000", 28771 => x"00000000", 28772 => x"00000000",
    28773 => x"00000000", 28774 => x"00000000", 28775 => x"00000000",
    28776 => x"00000000", 28777 => x"00000000", 28778 => x"00000000",
    28779 => x"00000000", 28780 => x"00000000", 28781 => x"00000000",
    28782 => x"00000000", 28783 => x"00000000", 28784 => x"00000000",
    28785 => x"00000000", 28786 => x"00000000", 28787 => x"00000000",
    28788 => x"00000000", 28789 => x"00000000", 28790 => x"00000000",
    28791 => x"00000000", 28792 => x"00000000", 28793 => x"00000000",
    28794 => x"00000000", 28795 => x"00000000", 28796 => x"00000000",
    28797 => x"00000000", 28798 => x"00000000", 28799 => x"00000000",
    28800 => x"00000000", 28801 => x"00000000", 28802 => x"00000000",
    28803 => x"00000000", 28804 => x"00000000", 28805 => x"00000000",
    28806 => x"00000000", 28807 => x"00000000", 28808 => x"00000000",
    28809 => x"00000000", 28810 => x"00000000", 28811 => x"00000000",
    28812 => x"00000000", 28813 => x"00000000", 28814 => x"00000000",
    28815 => x"00000000", 28816 => x"00000000", 28817 => x"00000000",
    28818 => x"00000000", 28819 => x"00000000", 28820 => x"00000000",
    28821 => x"00000000", 28822 => x"00000000", 28823 => x"00000000",
    28824 => x"00000000", 28825 => x"00000000", 28826 => x"00000000",
    28827 => x"00000000", 28828 => x"00000000", 28829 => x"00000000",
    28830 => x"00000000", 28831 => x"00000000", 28832 => x"00000000",
    28833 => x"00000000", 28834 => x"00000000", 28835 => x"00000000",
    28836 => x"00000000", 28837 => x"00000000", 28838 => x"00000000",
    28839 => x"00000000", 28840 => x"00000000", 28841 => x"00000000",
    28842 => x"00000000", 28843 => x"00000000", 28844 => x"00000000",
    28845 => x"00000000", 28846 => x"00000000", 28847 => x"00000000",
    28848 => x"00000000", 28849 => x"00000000", 28850 => x"00000000",
    28851 => x"00000000", 28852 => x"00000000", 28853 => x"00000000",
    28854 => x"00000000", 28855 => x"00000000", 28856 => x"00000000",
    28857 => x"00000000", 28858 => x"00000000", 28859 => x"00000000",
    28860 => x"00000000", 28861 => x"00000000", 28862 => x"00000000",
    28863 => x"00000000", 28864 => x"00000000", 28865 => x"00000000",
    28866 => x"00000000", 28867 => x"00000000", 28868 => x"00000000",
    28869 => x"00000000", 28870 => x"00000000", 28871 => x"00000000",
    28872 => x"00000000", 28873 => x"00000000", 28874 => x"00000000",
    28875 => x"00000000", 28876 => x"00000000", 28877 => x"00000000",
    28878 => x"00000000", 28879 => x"00000000", 28880 => x"00000000",
    28881 => x"00000000", 28882 => x"00000000", 28883 => x"00000000",
    28884 => x"00000000", 28885 => x"00000000", 28886 => x"00000000",
    28887 => x"00000000", 28888 => x"00000000", 28889 => x"00000000",
    28890 => x"00000000", 28891 => x"00000000", 28892 => x"00000000",
    28893 => x"00000000", 28894 => x"00000000", 28895 => x"00000000",
    28896 => x"00000000", 28897 => x"00000000", 28898 => x"00000000",
    28899 => x"00000000", 28900 => x"00000000", 28901 => x"00000000",
    28902 => x"00000000", 28903 => x"00000000", 28904 => x"00000000",
    28905 => x"00000000", 28906 => x"00000000", 28907 => x"00000000",
    28908 => x"00000000", 28909 => x"00000000", 28910 => x"00000000",
    28911 => x"00000000", 28912 => x"00000000", 28913 => x"00000000",
    28914 => x"00000000", 28915 => x"00000000", 28916 => x"00000000",
    28917 => x"00000000", 28918 => x"00000000", 28919 => x"00000000",
    28920 => x"00000000", 28921 => x"00000000", 28922 => x"00000000",
    28923 => x"00000000", 28924 => x"00000000", 28925 => x"00000000",
    28926 => x"00000000", 28927 => x"00000000", 28928 => x"00000000",
    28929 => x"00000000", 28930 => x"00000000", 28931 => x"00000000",
    28932 => x"00000000", 28933 => x"00000000", 28934 => x"00000000",
    28935 => x"00000000", 28936 => x"00000000", 28937 => x"00000000",
    28938 => x"00000000", 28939 => x"00000000", 28940 => x"00000000",
    28941 => x"00000000", 28942 => x"00000000", 28943 => x"00000000",
    28944 => x"00000000", 28945 => x"00000000", 28946 => x"00000000",
    28947 => x"00000000", 28948 => x"00000000", 28949 => x"00000000",
    28950 => x"00000000", 28951 => x"00000000", 28952 => x"00000000",
    28953 => x"00000000", 28954 => x"00000000", 28955 => x"00000000",
    28956 => x"00000000", 28957 => x"00000000", 28958 => x"00000000",
    28959 => x"00000000", 28960 => x"00000000", 28961 => x"00000000",
    28962 => x"00000000", 28963 => x"00000000", 28964 => x"00000000",
    28965 => x"00000000", 28966 => x"00000000", 28967 => x"00000000",
    28968 => x"00000000", 28969 => x"00000000", 28970 => x"00000000",
    28971 => x"00000000", 28972 => x"00000000", 28973 => x"00000000",
    28974 => x"00000000", 28975 => x"00000000", 28976 => x"00000000",
    28977 => x"00000000", 28978 => x"00000000", 28979 => x"00000000",
    28980 => x"00000000", 28981 => x"00000000", 28982 => x"00000000",
    28983 => x"00000000", 28984 => x"00000000", 28985 => x"00000000",
    28986 => x"00000000", 28987 => x"00000000", 28988 => x"00000000",
    28989 => x"00000000", 28990 => x"00000000", 28991 => x"00000000",
    28992 => x"00000000", 28993 => x"00000000", 28994 => x"00000000",
    28995 => x"00000000", 28996 => x"00000000", 28997 => x"00000000",
    28998 => x"00000000", 28999 => x"00000000", 29000 => x"00000000",
    29001 => x"00000000", 29002 => x"00000000", 29003 => x"00000000",
    29004 => x"00000000", 29005 => x"00000000", 29006 => x"00000000",
    29007 => x"00000000", 29008 => x"00000000", 29009 => x"00000000",
    29010 => x"00000000", 29011 => x"00000000", 29012 => x"00000000",
    29013 => x"00000000", 29014 => x"00000000", 29015 => x"00000000",
    29016 => x"00000000", 29017 => x"00000000", 29018 => x"00000000",
    29019 => x"00000000", 29020 => x"00000000", 29021 => x"00000000",
    29022 => x"00000000", 29023 => x"00000000", 29024 => x"00000000",
    29025 => x"00000000", 29026 => x"00000000", 29027 => x"00000000",
    29028 => x"00000000", 29029 => x"00000000", 29030 => x"00000000",
    29031 => x"00000000", 29032 => x"00000000", 29033 => x"00000000",
    29034 => x"00000000", 29035 => x"00000000", 29036 => x"00000000",
    29037 => x"00000000", 29038 => x"00000000", 29039 => x"00000000",
    29040 => x"00000000", 29041 => x"00000000", 29042 => x"00000000",
    29043 => x"00000000", 29044 => x"00000000", 29045 => x"00000000",
    29046 => x"00000000", 29047 => x"00000000", 29048 => x"00000000",
    29049 => x"00000000", 29050 => x"00000000", 29051 => x"00000000",
    29052 => x"00000000", 29053 => x"00000000", 29054 => x"00000000",
    29055 => x"00000000", 29056 => x"00000000", 29057 => x"00000000",
    29058 => x"00000000", 29059 => x"00000000", 29060 => x"00000000",
    29061 => x"00000000", 29062 => x"00000000", 29063 => x"00000000",
    29064 => x"00000000", 29065 => x"00000000", 29066 => x"00000000",
    29067 => x"00000000", 29068 => x"00000000", 29069 => x"00000000",
    29070 => x"00000000", 29071 => x"00000000", 29072 => x"00000000",
    29073 => x"00000000", 29074 => x"00000000", 29075 => x"00000000",
    29076 => x"00000000", 29077 => x"00000000", 29078 => x"00000000",
    29079 => x"00000000", 29080 => x"00000000", 29081 => x"00000000",
    29082 => x"00000000", 29083 => x"00000000", 29084 => x"00000000",
    29085 => x"00000000", 29086 => x"00000000", 29087 => x"00000000",
    29088 => x"00000000", 29089 => x"00000000", 29090 => x"00000000",
    29091 => x"00000000", 29092 => x"00000000", 29093 => x"00000000",
    29094 => x"00000000", 29095 => x"00000000", 29096 => x"00000000",
    29097 => x"00000000", 29098 => x"00000000", 29099 => x"00000000",
    29100 => x"00000000", 29101 => x"00000000", 29102 => x"00000000",
    29103 => x"00000000", 29104 => x"00000000", 29105 => x"00000000",
    29106 => x"00000000", 29107 => x"00000000", 29108 => x"00000000",
    29109 => x"00000000", 29110 => x"00000000", 29111 => x"00000000",
    29112 => x"00000000", 29113 => x"00000000", 29114 => x"00000000",
    29115 => x"00000000", 29116 => x"00000000", 29117 => x"00000000",
    29118 => x"00000000", 29119 => x"00000000", 29120 => x"00000000",
    29121 => x"00000000", 29122 => x"00000000", 29123 => x"00000000",
    29124 => x"00000000", 29125 => x"00000000", 29126 => x"00000000",
    29127 => x"00000000", 29128 => x"00000000", 29129 => x"00000000",
    29130 => x"00000000", 29131 => x"00000000", 29132 => x"00000000",
    29133 => x"00000000", 29134 => x"00000000", 29135 => x"00000000",
    29136 => x"00000000", 29137 => x"00000000", 29138 => x"00000000",
    29139 => x"00000000", 29140 => x"00000000", 29141 => x"00000000",
    29142 => x"00000000", 29143 => x"00000000", 29144 => x"00000000",
    29145 => x"00000000", 29146 => x"00000000", 29147 => x"00000000",
    29148 => x"00000000", 29149 => x"00000000", 29150 => x"00000000",
    29151 => x"00000000", 29152 => x"00000000", 29153 => x"00000000",
    29154 => x"00000000", 29155 => x"00000000", 29156 => x"00000000",
    29157 => x"00000000", 29158 => x"00000000", 29159 => x"00000000",
    29160 => x"00000000", 29161 => x"00000000", 29162 => x"00000000",
    29163 => x"00000000", 29164 => x"00000000", 29165 => x"00000000",
    29166 => x"00000000", 29167 => x"00000000", 29168 => x"00000000",
    29169 => x"00000000", 29170 => x"00000000", 29171 => x"00000000",
    29172 => x"00000000", 29173 => x"00000000", 29174 => x"00000000",
    29175 => x"00000000", 29176 => x"00000000", 29177 => x"00000000",
    29178 => x"00000000", 29179 => x"00000000", 29180 => x"00000000",
    29181 => x"00000000", 29182 => x"00000000", 29183 => x"00000000",
    29184 => x"00000000", 29185 => x"00000000", 29186 => x"00000000",
    29187 => x"00000000", 29188 => x"00000000", 29189 => x"00000000",
    29190 => x"00000000", 29191 => x"00000000", 29192 => x"00000000",
    29193 => x"00000000", 29194 => x"00000000", 29195 => x"00000000",
    29196 => x"00000000", 29197 => x"00000000", 29198 => x"00000000",
    29199 => x"00000000", 29200 => x"00000000", 29201 => x"00000000",
    29202 => x"00000000", 29203 => x"00000000", 29204 => x"00000000",
    29205 => x"00000000", 29206 => x"00000000", 29207 => x"00000000",
    29208 => x"00000000", 29209 => x"00000000", 29210 => x"00000000",
    29211 => x"00000000", 29212 => x"00000000", 29213 => x"00000000",
    29214 => x"00000000", 29215 => x"00000000", 29216 => x"00000000",
    29217 => x"00000000", 29218 => x"00000000", 29219 => x"00000000",
    29220 => x"00000000", 29221 => x"00000000", 29222 => x"00000000",
    29223 => x"00000000", 29224 => x"00000000", 29225 => x"00000000",
    29226 => x"00000000", 29227 => x"00000000", 29228 => x"00000000",
    29229 => x"00000000", 29230 => x"00000000", 29231 => x"00000000",
    29232 => x"00000000", 29233 => x"00000000", 29234 => x"00000000",
    29235 => x"00000000", 29236 => x"00000000", 29237 => x"00000000",
    29238 => x"00000000", 29239 => x"00000000", 29240 => x"00000000",
    29241 => x"00000000", 29242 => x"00000000", 29243 => x"00000000",
    29244 => x"00000000", 29245 => x"00000000", 29246 => x"00000000",
    29247 => x"00000000", 29248 => x"00000000", 29249 => x"00000000",
    29250 => x"00000000", 29251 => x"00000000", 29252 => x"00000000",
    29253 => x"00000000", 29254 => x"00000000", 29255 => x"00000000",
    29256 => x"00000000", 29257 => x"00000000", 29258 => x"00000000",
    29259 => x"00000000", 29260 => x"00000000", 29261 => x"00000000",
    29262 => x"00000000", 29263 => x"00000000", 29264 => x"00000000",
    29265 => x"00000000", 29266 => x"00000000", 29267 => x"00000000",
    29268 => x"00000000", 29269 => x"00000000", 29270 => x"00000000",
    29271 => x"00000000", 29272 => x"00000000", 29273 => x"00000000",
    29274 => x"00000000", 29275 => x"00000000", 29276 => x"00000000",
    29277 => x"00000000", 29278 => x"00000000", 29279 => x"00000000",
    29280 => x"00000000", 29281 => x"00000000", 29282 => x"00000000",
    29283 => x"00000000", 29284 => x"00000000", 29285 => x"00000000",
    29286 => x"00000000", 29287 => x"00000000", 29288 => x"00000000",
    29289 => x"00000000", 29290 => x"00000000", 29291 => x"00000000",
    29292 => x"00000000", 29293 => x"00000000", 29294 => x"00000000",
    29295 => x"00000000", 29296 => x"00000000", 29297 => x"00000000",
    29298 => x"00000000", 29299 => x"00000000", 29300 => x"00000000",
    29301 => x"00000000", 29302 => x"00000000", 29303 => x"00000000",
    29304 => x"00000000", 29305 => x"00000000", 29306 => x"00000000",
    29307 => x"00000000", 29308 => x"00000000", 29309 => x"00000000",
    29310 => x"00000000", 29311 => x"00000000", 29312 => x"00000000",
    29313 => x"00000000", 29314 => x"00000000", 29315 => x"00000000",
    29316 => x"00000000", 29317 => x"00000000", 29318 => x"00000000",
    29319 => x"00000000", 29320 => x"00000000", 29321 => x"00000000",
    29322 => x"00000000", 29323 => x"00000000", 29324 => x"00000000",
    29325 => x"00000000", 29326 => x"00000000", 29327 => x"00000000",
    29328 => x"00000000", 29329 => x"00000000", 29330 => x"00000000",
    29331 => x"00000000", 29332 => x"00000000", 29333 => x"00000000",
    29334 => x"00000000", 29335 => x"00000000", 29336 => x"00000000",
    29337 => x"00000000", 29338 => x"00000000", 29339 => x"00000000",
    29340 => x"00000000", 29341 => x"00000000", 29342 => x"00000000",
    29343 => x"00000000", 29344 => x"00000000", 29345 => x"00000000",
    29346 => x"00000000", 29347 => x"00000000", 29348 => x"00000000",
    29349 => x"00000000", 29350 => x"00000000", 29351 => x"00000000",
    29352 => x"00000000", 29353 => x"00000000", 29354 => x"00000000",
    29355 => x"00000000", 29356 => x"00000000", 29357 => x"00000000",
    29358 => x"00000000", 29359 => x"00000000", 29360 => x"00000000",
    29361 => x"00000000", 29362 => x"00000000", 29363 => x"00000000",
    29364 => x"00000000", 29365 => x"00000000", 29366 => x"00000000",
    29367 => x"00000000", 29368 => x"00000000", 29369 => x"00000000",
    29370 => x"00000000", 29371 => x"00000000", 29372 => x"00000000",
    29373 => x"00000000", 29374 => x"00000000", 29375 => x"00000000",
    29376 => x"00000000", 29377 => x"00000000", 29378 => x"00000000",
    29379 => x"00000000", 29380 => x"00000000", 29381 => x"00000000",
    29382 => x"00000000", 29383 => x"00000000", 29384 => x"00000000",
    29385 => x"00000000", 29386 => x"00000000", 29387 => x"00000000",
    29388 => x"00000000", 29389 => x"00000000", 29390 => x"00000000",
    29391 => x"00000000", 29392 => x"00000000", 29393 => x"00000000",
    29394 => x"00000000", 29395 => x"00000000", 29396 => x"00000000",
    29397 => x"00000000", 29398 => x"00000000", 29399 => x"00000000",
    29400 => x"00000000", 29401 => x"00000000", 29402 => x"00000000",
    29403 => x"00000000", 29404 => x"00000000", 29405 => x"00000000",
    29406 => x"00000000", 29407 => x"00000000", 29408 => x"00000000",
    29409 => x"00000000", 29410 => x"00000000", 29411 => x"00000000",
    29412 => x"00000000", 29413 => x"00000000", 29414 => x"00000000",
    29415 => x"00000000", 29416 => x"00000000", 29417 => x"00000000",
    29418 => x"00000000", 29419 => x"00000000", 29420 => x"00000000",
    29421 => x"00000000", 29422 => x"00000000", 29423 => x"00000000",
    29424 => x"00000000", 29425 => x"00000000", 29426 => x"00000000",
    29427 => x"00000000", 29428 => x"00000000", 29429 => x"00000000",
    29430 => x"00000000", 29431 => x"00000000", 29432 => x"00000000",
    29433 => x"00000000", 29434 => x"00000000", 29435 => x"00000000",
    29436 => x"00000000", 29437 => x"00000000", 29438 => x"00000000",
    29439 => x"00000000", 29440 => x"00000000", 29441 => x"00000000",
    29442 => x"00000000", 29443 => x"00000000", 29444 => x"00000000",
    29445 => x"00000000", 29446 => x"00000000", 29447 => x"00000000",
    29448 => x"00000000", 29449 => x"00000000", 29450 => x"00000000",
    29451 => x"00000000", 29452 => x"00000000", 29453 => x"00000000",
    29454 => x"00000000", 29455 => x"00000000", 29456 => x"00000000",
    29457 => x"00000000", 29458 => x"00000000", 29459 => x"00000000",
    29460 => x"00000000", 29461 => x"00000000", 29462 => x"00000000",
    29463 => x"00000000", 29464 => x"00000000", 29465 => x"00000000",
    29466 => x"00000000", 29467 => x"00000000", 29468 => x"00000000",
    29469 => x"00000000", 29470 => x"00000000", 29471 => x"00000000",
    29472 => x"00000000", 29473 => x"00000000", 29474 => x"00000000",
    29475 => x"00000000", 29476 => x"00000000", 29477 => x"00000000",
    29478 => x"00000000", 29479 => x"00000000", 29480 => x"00000000",
    29481 => x"00000000", 29482 => x"00000000", 29483 => x"00000000",
    29484 => x"00000000", 29485 => x"00000000", 29486 => x"00000000",
    29487 => x"00000000", 29488 => x"00000000", 29489 => x"00000000",
    29490 => x"00000000", 29491 => x"00000000", 29492 => x"00000000",
    29493 => x"00000000", 29494 => x"00000000", 29495 => x"00000000",
    29496 => x"00000000", 29497 => x"00000000", 29498 => x"00000000",
    29499 => x"00000000", 29500 => x"00000000", 29501 => x"00000000",
    29502 => x"00000000", 29503 => x"00000000", 29504 => x"00000000",
    29505 => x"00000000", 29506 => x"00000000", 29507 => x"00000000",
    29508 => x"00000000", 29509 => x"00000000", 29510 => x"00000000",
    29511 => x"00000000", 29512 => x"00000000", 29513 => x"00000000",
    29514 => x"00000000", 29515 => x"00000000", 29516 => x"00000000",
    29517 => x"00000000", 29518 => x"00000000", 29519 => x"00000000",
    29520 => x"00000000", 29521 => x"00000000", 29522 => x"00000000",
    29523 => x"00000000", 29524 => x"00000000", 29525 => x"00000000",
    29526 => x"00000000", 29527 => x"00000000", 29528 => x"00000000",
    29529 => x"00000000", 29530 => x"00000000", 29531 => x"00000000",
    29532 => x"00000000", 29533 => x"00000000", 29534 => x"00000000",
    29535 => x"00000000", 29536 => x"00000000", 29537 => x"00000000",
    29538 => x"00000000", 29539 => x"00000000", 29540 => x"00000000",
    29541 => x"00000000", 29542 => x"00000000", 29543 => x"00000000",
    29544 => x"00000000", 29545 => x"00000000", 29546 => x"00000000",
    29547 => x"00000000", 29548 => x"00000000", 29549 => x"00000000",
    29550 => x"00000000", 29551 => x"00000000", 29552 => x"00000000",
    29553 => x"00000000", 29554 => x"00000000", 29555 => x"00000000",
    29556 => x"00000000", 29557 => x"00000000", 29558 => x"00000000",
    29559 => x"00000000", 29560 => x"00000000", 29561 => x"00000000",
    29562 => x"00000000", 29563 => x"00000000", 29564 => x"00000000",
    29565 => x"00000000", 29566 => x"00000000", 29567 => x"00000000",
    29568 => x"00000000", 29569 => x"00000000", 29570 => x"00000000",
    29571 => x"00000000", 29572 => x"00000000", 29573 => x"00000000",
    29574 => x"00000000", 29575 => x"00000000", 29576 => x"00000000",
    29577 => x"00000000", 29578 => x"00000000", 29579 => x"00000000",
    29580 => x"00000000", 29581 => x"00000000", 29582 => x"00000000",
    29583 => x"00000000", 29584 => x"00000000", 29585 => x"00000000",
    29586 => x"00000000", 29587 => x"00000000", 29588 => x"00000000",
    29589 => x"00000000", 29590 => x"00000000", 29591 => x"00000000",
    29592 => x"00000000", 29593 => x"00000000", 29594 => x"00000000",
    29595 => x"00000000", 29596 => x"00000000", 29597 => x"00000000",
    29598 => x"00000000", 29599 => x"00000000", 29600 => x"00000000",
    29601 => x"00000000", 29602 => x"00000000", 29603 => x"00000000",
    29604 => x"00000000", 29605 => x"00000000", 29606 => x"00000000",
    29607 => x"00000000", 29608 => x"00000000", 29609 => x"00000000",
    29610 => x"00000000", 29611 => x"00000000", 29612 => x"00000000",
    29613 => x"00000000", 29614 => x"00000000", 29615 => x"00000000",
    29616 => x"00000000", 29617 => x"00000000", 29618 => x"00000000",
    29619 => x"00000000", 29620 => x"00000000", 29621 => x"00000000",
    29622 => x"00000000", 29623 => x"00000000", 29624 => x"00000000",
    29625 => x"00000000", 29626 => x"00000000", 29627 => x"00000000",
    29628 => x"00000000", 29629 => x"00000000", 29630 => x"00000000",
    29631 => x"00000000", 29632 => x"00000000", 29633 => x"00000000",
    29634 => x"00000000", 29635 => x"00000000", 29636 => x"00000000",
    29637 => x"00000000", 29638 => x"00000000", 29639 => x"00000000",
    29640 => x"00000000", 29641 => x"00000000", 29642 => x"00000000",
    29643 => x"00000000", 29644 => x"00000000", 29645 => x"00000000",
    29646 => x"00000000", 29647 => x"00000000", 29648 => x"00000000",
    29649 => x"00000000", 29650 => x"00000000", 29651 => x"00000000",
    29652 => x"00000000", 29653 => x"00000000", 29654 => x"00000000",
    29655 => x"00000000", 29656 => x"00000000", 29657 => x"00000000",
    29658 => x"00000000", 29659 => x"00000000", 29660 => x"00000000",
    29661 => x"00000000", 29662 => x"00000000", 29663 => x"00000000",
    29664 => x"00000000", 29665 => x"00000000", 29666 => x"00000000",
    29667 => x"00000000", 29668 => x"00000000", 29669 => x"00000000",
    29670 => x"00000000", 29671 => x"00000000", 29672 => x"00000000",
    29673 => x"00000000", 29674 => x"00000000", 29675 => x"00000000",
    29676 => x"00000000", 29677 => x"00000000", 29678 => x"00000000",
    29679 => x"00000000", 29680 => x"00000000", 29681 => x"00000000",
    29682 => x"00000000", 29683 => x"00000000", 29684 => x"00000000",
    29685 => x"00000000", 29686 => x"00000000", 29687 => x"00000000",
    29688 => x"00000000", 29689 => x"00000000", 29690 => x"00000000",
    29691 => x"00000000", 29692 => x"00000000", 29693 => x"00000000",
    29694 => x"00000000", 29695 => x"00000000", 29696 => x"00000000",
    29697 => x"00000000", 29698 => x"00000000", 29699 => x"00000000",
    29700 => x"00000000", 29701 => x"00000000", 29702 => x"00000000",
    29703 => x"00000000", 29704 => x"00000000", 29705 => x"00000000",
    29706 => x"00000000", 29707 => x"00000000", 29708 => x"00000000",
    29709 => x"00000000", 29710 => x"00000000", 29711 => x"00000000",
    29712 => x"00000000", 29713 => x"00000000", 29714 => x"00000000",
    29715 => x"00000000", 29716 => x"00000000", 29717 => x"00000000",
    29718 => x"00000000", 29719 => x"00000000", 29720 => x"00000000",
    29721 => x"00000000", 29722 => x"00000000", 29723 => x"00000000",
    29724 => x"00000000", 29725 => x"00000000", 29726 => x"00000000",
    29727 => x"00000000", 29728 => x"00000000", 29729 => x"00000000",
    29730 => x"00000000", 29731 => x"00000000", 29732 => x"00000000",
    29733 => x"00000000", 29734 => x"00000000", 29735 => x"00000000",
    29736 => x"00000000", 29737 => x"00000000", 29738 => x"00000000",
    29739 => x"00000000", 29740 => x"00000000", 29741 => x"00000000",
    29742 => x"00000000", 29743 => x"00000000", 29744 => x"00000000",
    29745 => x"00000000", 29746 => x"00000000", 29747 => x"00000000",
    29748 => x"00000000", 29749 => x"00000000", 29750 => x"00000000",
    29751 => x"00000000", 29752 => x"00000000", 29753 => x"00000000",
    29754 => x"00000000", 29755 => x"00000000", 29756 => x"00000000",
    29757 => x"00000000", 29758 => x"00000000", 29759 => x"00000000",
    29760 => x"00000000", 29761 => x"00000000", 29762 => x"00000000",
    29763 => x"00000000", 29764 => x"00000000", 29765 => x"00000000",
    29766 => x"00000000", 29767 => x"00000000", 29768 => x"00000000",
    29769 => x"00000000", 29770 => x"00000000", 29771 => x"00000000",
    29772 => x"00000000", 29773 => x"00000000", 29774 => x"00000000",
    29775 => x"00000000", 29776 => x"00000000", 29777 => x"00000000",
    29778 => x"00000000", 29779 => x"00000000", 29780 => x"00000000",
    29781 => x"00000000", 29782 => x"00000000", 29783 => x"00000000",
    29784 => x"00000000", 29785 => x"00000000", 29786 => x"00000000",
    29787 => x"00000000", 29788 => x"00000000", 29789 => x"00000000",
    29790 => x"00000000", 29791 => x"00000000", 29792 => x"00000000",
    29793 => x"00000000", 29794 => x"00000000", 29795 => x"00000000",
    29796 => x"00000000", 29797 => x"00000000", 29798 => x"00000000",
    29799 => x"00000000", 29800 => x"00000000", 29801 => x"00000000",
    29802 => x"00000000", 29803 => x"00000000", 29804 => x"00000000",
    29805 => x"00000000", 29806 => x"00000000", 29807 => x"00000000",
    29808 => x"00000000", 29809 => x"00000000", 29810 => x"00000000",
    29811 => x"00000000", 29812 => x"00000000", 29813 => x"00000000",
    29814 => x"00000000", 29815 => x"00000000", 29816 => x"00000000",
    29817 => x"00000000", 29818 => x"00000000", 29819 => x"00000000",
    29820 => x"00000000", 29821 => x"00000000", 29822 => x"00000000",
    29823 => x"00000000", 29824 => x"00000000", 29825 => x"00000000",
    29826 => x"00000000", 29827 => x"00000000", 29828 => x"00000000",
    29829 => x"00000000", 29830 => x"00000000", 29831 => x"00000000",
    29832 => x"00000000", 29833 => x"00000000", 29834 => x"00000000",
    29835 => x"00000000", 29836 => x"00000000", 29837 => x"00000000",
    29838 => x"00000000", 29839 => x"00000000", 29840 => x"00000000",
    29841 => x"00000000", 29842 => x"00000000", 29843 => x"00000000",
    29844 => x"00000000", 29845 => x"00000000", 29846 => x"00000000",
    29847 => x"00000000", 29848 => x"00000000", 29849 => x"00000000",
    29850 => x"00000000", 29851 => x"00000000", 29852 => x"00000000",
    29853 => x"00000000", 29854 => x"00000000", 29855 => x"00000000",
    29856 => x"00000000", 29857 => x"00000000", 29858 => x"00000000",
    29859 => x"00000000", 29860 => x"00000000", 29861 => x"00000000",
    29862 => x"00000000", 29863 => x"00000000", 29864 => x"00000000",
    29865 => x"00000000", 29866 => x"00000000", 29867 => x"00000000",
    29868 => x"00000000", 29869 => x"00000000", 29870 => x"00000000",
    29871 => x"00000000", 29872 => x"00000000", 29873 => x"00000000",
    29874 => x"00000000", 29875 => x"00000000", 29876 => x"00000000",
    29877 => x"00000000", 29878 => x"00000000", 29879 => x"00000000",
    29880 => x"00000000", 29881 => x"00000000", 29882 => x"00000000",
    29883 => x"00000000", 29884 => x"00000000", 29885 => x"00000000",
    29886 => x"00000000", 29887 => x"00000000", 29888 => x"00000000",
    29889 => x"00000000", 29890 => x"00000000", 29891 => x"00000000",
    29892 => x"00000000", 29893 => x"00000000", 29894 => x"00000000",
    29895 => x"00000000", 29896 => x"00000000", 29897 => x"00000000",
    29898 => x"00000000", 29899 => x"00000000", 29900 => x"00000000",
    29901 => x"00000000", 29902 => x"00000000", 29903 => x"00000000",
    29904 => x"00000000", 29905 => x"00000000", 29906 => x"00000000",
    29907 => x"00000000", 29908 => x"00000000", 29909 => x"00000000",
    29910 => x"00000000", 29911 => x"00000000", 29912 => x"00000000",
    29913 => x"00000000", 29914 => x"00000000", 29915 => x"00000000",
    29916 => x"00000000", 29917 => x"00000000", 29918 => x"00000000",
    29919 => x"00000000", 29920 => x"00000000", 29921 => x"00000000",
    29922 => x"00000000", 29923 => x"00000000", 29924 => x"00000000",
    29925 => x"00000000", 29926 => x"00000000", 29927 => x"00000000",
    29928 => x"00000000", 29929 => x"00000000", 29930 => x"00000000",
    29931 => x"00000000", 29932 => x"00000000", 29933 => x"00000000",
    29934 => x"00000000", 29935 => x"00000000", 29936 => x"00000000",
    29937 => x"00000000", 29938 => x"00000000", 29939 => x"00000000",
    29940 => x"00000000", 29941 => x"00000000", 29942 => x"00000000",
    29943 => x"00000000", 29944 => x"00000000", 29945 => x"00000000",
    29946 => x"00000000", 29947 => x"00000000", 29948 => x"00000000",
    29949 => x"00000000", 29950 => x"00000000", 29951 => x"00000000",
    29952 => x"00000000", 29953 => x"00000000", 29954 => x"00000000",
    29955 => x"00000000", 29956 => x"00000000", 29957 => x"00000000",
    29958 => x"00000000", 29959 => x"00000000", 29960 => x"00000000",
    29961 => x"00000000", 29962 => x"00000000", 29963 => x"00000000",
    29964 => x"00000000", 29965 => x"00000000", 29966 => x"00000000",
    29967 => x"00000000", 29968 => x"00000000", 29969 => x"00000000",
    29970 => x"00000000", 29971 => x"00000000", 29972 => x"00000000",
    29973 => x"00000000", 29974 => x"00000000", 29975 => x"00000000",
    29976 => x"00000000", 29977 => x"00000000", 29978 => x"00000000",
    29979 => x"00000000", 29980 => x"00000000", 29981 => x"00000000",
    29982 => x"00000000", 29983 => x"00000000", 29984 => x"00000000",
    29985 => x"00000000", 29986 => x"00000000", 29987 => x"00000000",
    29988 => x"00000000", 29989 => x"00000000", 29990 => x"00000000",
    29991 => x"00000000", 29992 => x"00000000", 29993 => x"00000000",
    29994 => x"00000000", 29995 => x"00000000", 29996 => x"00000000",
    29997 => x"00000000", 29998 => x"00000000", 29999 => x"00000000",
    30000 => x"00000000", 30001 => x"00000000", 30002 => x"00000000",
    30003 => x"00000000", 30004 => x"00000000", 30005 => x"00000000",
    30006 => x"00000000", 30007 => x"00000000", 30008 => x"00000000",
    30009 => x"00000000", 30010 => x"00000000", 30011 => x"00000000",
    30012 => x"00000000", 30013 => x"00000000", 30014 => x"00000000",
    30015 => x"00000000", 30016 => x"00000000", 30017 => x"00000000",
    30018 => x"00000000", 30019 => x"00000000", 30020 => x"00000000",
    30021 => x"00000000", 30022 => x"00000000", 30023 => x"00000000",
    30024 => x"00000000", 30025 => x"00000000", 30026 => x"00000000",
    30027 => x"00000000", 30028 => x"00000000", 30029 => x"00000000",
    30030 => x"00000000", 30031 => x"00000000", 30032 => x"00000000",
    30033 => x"00000000", 30034 => x"00000000", 30035 => x"00000000",
    30036 => x"00000000", 30037 => x"00000000", 30038 => x"00000000",
    30039 => x"00000000", 30040 => x"00000000", 30041 => x"00000000",
    30042 => x"00000000", 30043 => x"00000000", 30044 => x"00000000",
    30045 => x"00000000", 30046 => x"00000000", 30047 => x"00000000",
    30048 => x"00000000", 30049 => x"00000000", 30050 => x"00000000",
    30051 => x"00000000", 30052 => x"00000000", 30053 => x"00000000",
    30054 => x"00000000", 30055 => x"00000000", 30056 => x"00000000",
    30057 => x"00000000", 30058 => x"00000000", 30059 => x"00000000",
    30060 => x"00000000", 30061 => x"00000000", 30062 => x"00000000",
    30063 => x"00000000", 30064 => x"00000000", 30065 => x"00000000",
    30066 => x"00000000", 30067 => x"00000000", 30068 => x"00000000",
    30069 => x"00000000", 30070 => x"00000000", 30071 => x"00000000",
    30072 => x"00000000", 30073 => x"00000000", 30074 => x"00000000",
    30075 => x"00000000", 30076 => x"00000000", 30077 => x"00000000",
    30078 => x"00000000", 30079 => x"00000000", 30080 => x"00000000",
    30081 => x"00000000", 30082 => x"00000000", 30083 => x"00000000",
    30084 => x"00000000", 30085 => x"00000000", 30086 => x"00000000",
    30087 => x"00000000", 30088 => x"00000000", 30089 => x"00000000",
    30090 => x"00000000", 30091 => x"00000000", 30092 => x"00000000",
    30093 => x"00000000", 30094 => x"00000000", 30095 => x"00000000",
    30096 => x"00000000", 30097 => x"00000000", 30098 => x"00000000",
    30099 => x"00000000", 30100 => x"00000000", 30101 => x"00000000",
    30102 => x"00000000", 30103 => x"00000000", 30104 => x"00000000",
    30105 => x"00000000", 30106 => x"00000000", 30107 => x"00000000",
    30108 => x"00000000", 30109 => x"00000000", 30110 => x"00000000",
    30111 => x"00000000", 30112 => x"00000000", 30113 => x"00000000",
    30114 => x"00000000", 30115 => x"00000000", 30116 => x"00000000",
    30117 => x"00000000", 30118 => x"00000000", 30119 => x"00000000",
    30120 => x"00000000", 30121 => x"00000000", 30122 => x"00000000",
    30123 => x"00000000", 30124 => x"00000000", 30125 => x"00000000",
    30126 => x"00000000", 30127 => x"00000000", 30128 => x"00000000",
    30129 => x"00000000", 30130 => x"00000000", 30131 => x"00000000",
    30132 => x"00000000", 30133 => x"00000000", 30134 => x"00000000",
    30135 => x"00000000", 30136 => x"00000000", 30137 => x"00000000",
    30138 => x"00000000", 30139 => x"00000000", 30140 => x"00000000",
    30141 => x"00000000", 30142 => x"00000000", 30143 => x"00000000",
    30144 => x"00000000", 30145 => x"00000000", 30146 => x"00000000",
    30147 => x"00000000", 30148 => x"00000000", 30149 => x"00000000",
    30150 => x"00000000", 30151 => x"00000000", 30152 => x"00000000",
    30153 => x"00000000", 30154 => x"00000000", 30155 => x"00000000",
    30156 => x"00000000", 30157 => x"00000000", 30158 => x"00000000",
    30159 => x"00000000", 30160 => x"00000000", 30161 => x"00000000",
    30162 => x"00000000", 30163 => x"00000000", 30164 => x"00000000",
    30165 => x"00000000", 30166 => x"00000000", 30167 => x"00000000",
    30168 => x"00000000", 30169 => x"00000000", 30170 => x"00000000",
    30171 => x"00000000", 30172 => x"00000000", 30173 => x"00000000",
    30174 => x"00000000", 30175 => x"00000000", 30176 => x"00000000",
    30177 => x"00000000", 30178 => x"00000000", 30179 => x"00000000",
    30180 => x"00000000", 30181 => x"00000000", 30182 => x"00000000",
    30183 => x"00000000", 30184 => x"00000000", 30185 => x"00000000",
    30186 => x"00000000", 30187 => x"00000000", 30188 => x"00000000",
    30189 => x"00000000", 30190 => x"00000000", 30191 => x"00000000",
    30192 => x"00000000", 30193 => x"00000000", 30194 => x"00000000",
    30195 => x"00000000", 30196 => x"00000000", 30197 => x"00000000",
    30198 => x"00000000", 30199 => x"00000000", 30200 => x"00000000",
    30201 => x"00000000", 30202 => x"00000000", 30203 => x"00000000",
    30204 => x"00000000", 30205 => x"00000000", 30206 => x"00000000",
    30207 => x"00000000", 30208 => x"00000000", 30209 => x"00000000",
    30210 => x"00000000", 30211 => x"00000000", 30212 => x"00000000",
    30213 => x"00000000", 30214 => x"00000000", 30215 => x"00000000",
    30216 => x"00000000", 30217 => x"00000000", 30218 => x"00000000",
    30219 => x"00000000", 30220 => x"00000000", 30221 => x"00000000",
    30222 => x"00000000", 30223 => x"00000000", 30224 => x"00000000",
    30225 => x"00000000", 30226 => x"00000000", 30227 => x"00000000",
    30228 => x"00000000", 30229 => x"00000000", 30230 => x"00000000",
    30231 => x"00000000", 30232 => x"00000000", 30233 => x"00000000",
    30234 => x"00000000", 30235 => x"00000000", 30236 => x"00000000",
    30237 => x"00000000", 30238 => x"00000000", 30239 => x"00000000",
    30240 => x"00000000", 30241 => x"00000000", 30242 => x"00000000",
    30243 => x"00000000", 30244 => x"00000000", 30245 => x"00000000",
    30246 => x"00000000", 30247 => x"00000000", 30248 => x"00000000",
    30249 => x"00000000", 30250 => x"00000000", 30251 => x"00000000",
    30252 => x"00000000", 30253 => x"00000000", 30254 => x"00000000",
    30255 => x"00000000", 30256 => x"00000000", 30257 => x"00000000",
    30258 => x"00000000", 30259 => x"00000000", 30260 => x"00000000",
    30261 => x"00000000", 30262 => x"00000000", 30263 => x"00000000",
    30264 => x"00000000", 30265 => x"00000000", 30266 => x"00000000",
    30267 => x"00000000", 30268 => x"00000000", 30269 => x"00000000",
    30270 => x"00000000", 30271 => x"00000000", 30272 => x"00000000",
    30273 => x"00000000", 30274 => x"00000000", 30275 => x"00000000",
    30276 => x"00000000", 30277 => x"00000000", 30278 => x"00000000",
    30279 => x"00000000", 30280 => x"00000000", 30281 => x"00000000",
    30282 => x"00000000", 30283 => x"00000000", 30284 => x"00000000",
    30285 => x"00000000", 30286 => x"00000000", 30287 => x"00000000",
    30288 => x"00000000", 30289 => x"00000000", 30290 => x"00000000",
    30291 => x"00000000", 30292 => x"00000000", 30293 => x"00000000",
    30294 => x"00000000", 30295 => x"00000000", 30296 => x"00000000",
    30297 => x"00000000", 30298 => x"00000000", 30299 => x"00000000",
    30300 => x"00000000", 30301 => x"00000000", 30302 => x"00000000",
    30303 => x"00000000", 30304 => x"00000000", 30305 => x"00000000",
    30306 => x"00000000", 30307 => x"00000000", 30308 => x"00000000",
    30309 => x"00000000", 30310 => x"00000000", 30311 => x"00000000",
    30312 => x"00000000", 30313 => x"00000000", 30314 => x"00000000",
    30315 => x"00000000", 30316 => x"00000000", 30317 => x"00000000",
    30318 => x"00000000", 30319 => x"00000000", 30320 => x"00000000",
    30321 => x"00000000", 30322 => x"00000000", 30323 => x"00000000",
    30324 => x"00000000", 30325 => x"00000000", 30326 => x"00000000",
    30327 => x"00000000", 30328 => x"00000000", 30329 => x"00000000",
    30330 => x"00000000", 30331 => x"00000000", 30332 => x"00000000",
    30333 => x"00000000", 30334 => x"00000000", 30335 => x"00000000",
    30336 => x"00000000", 30337 => x"00000000", 30338 => x"00000000",
    30339 => x"00000000", 30340 => x"00000000", 30341 => x"00000000",
    30342 => x"00000000", 30343 => x"00000000", 30344 => x"00000000",
    30345 => x"00000000", 30346 => x"00000000", 30347 => x"00000000",
    30348 => x"00000000", 30349 => x"00000000", 30350 => x"00000000",
    30351 => x"00000000", 30352 => x"00000000", 30353 => x"00000000",
    30354 => x"00000000", 30355 => x"00000000", 30356 => x"00000000",
    30357 => x"00000000", 30358 => x"00000000", 30359 => x"00000000",
    30360 => x"00000000", 30361 => x"00000000", 30362 => x"00000000",
    30363 => x"00000000", 30364 => x"00000000", 30365 => x"00000000",
    30366 => x"00000000", 30367 => x"00000000", 30368 => x"00000000",
    30369 => x"00000000", 30370 => x"00000000", 30371 => x"00000000",
    30372 => x"00000000", 30373 => x"00000000", 30374 => x"00000000",
    30375 => x"00000000", 30376 => x"00000000", 30377 => x"00000000",
    30378 => x"00000000", 30379 => x"00000000", 30380 => x"00000000",
    30381 => x"00000000", 30382 => x"00000000", 30383 => x"00000000",
    30384 => x"00000000", 30385 => x"00000000", 30386 => x"00000000",
    30387 => x"00000000", 30388 => x"00000000", 30389 => x"00000000",
    30390 => x"00000000", 30391 => x"00000000", 30392 => x"00000000",
    30393 => x"00000000", 30394 => x"00000000", 30395 => x"00000000",
    30396 => x"00000000", 30397 => x"00000000", 30398 => x"00000000",
    30399 => x"00000000", 30400 => x"00000000", 30401 => x"00000000",
    30402 => x"00000000", 30403 => x"00000000", 30404 => x"00000000",
    30405 => x"00000000", 30406 => x"00000000", 30407 => x"00000000",
    30408 => x"00000000", 30409 => x"00000000", 30410 => x"00000000",
    30411 => x"00000000", 30412 => x"00000000", 30413 => x"00000000",
    30414 => x"00000000", 30415 => x"00000000", 30416 => x"00000000",
    30417 => x"00000000", 30418 => x"00000000", 30419 => x"00000000",
    30420 => x"00000000", 30421 => x"00000000", 30422 => x"00000000",
    30423 => x"00000000", 30424 => x"00000000", 30425 => x"00000000",
    30426 => x"00000000", 30427 => x"00000000", 30428 => x"00000000",
    30429 => x"00000000", 30430 => x"00000000", 30431 => x"00000000",
    30432 => x"00000000", 30433 => x"00000000", 30434 => x"00000000",
    30435 => x"00000000", 30436 => x"00000000", 30437 => x"00000000",
    30438 => x"00000000", 30439 => x"00000000", 30440 => x"00000000",
    30441 => x"00000000", 30442 => x"00000000", 30443 => x"00000000",
    30444 => x"00000000", 30445 => x"00000000", 30446 => x"00000000",
    30447 => x"00000000", 30448 => x"00000000", 30449 => x"00000000",
    30450 => x"00000000", 30451 => x"00000000", 30452 => x"00000000",
    30453 => x"00000000", 30454 => x"00000000", 30455 => x"00000000",
    30456 => x"00000000", 30457 => x"00000000", 30458 => x"00000000",
    30459 => x"00000000", 30460 => x"00000000", 30461 => x"00000000",
    30462 => x"00000000", 30463 => x"00000000", 30464 => x"00000000",
    30465 => x"00000000", 30466 => x"00000000", 30467 => x"00000000",
    30468 => x"00000000", 30469 => x"00000000", 30470 => x"00000000",
    30471 => x"00000000", 30472 => x"00000000", 30473 => x"00000000",
    30474 => x"00000000", 30475 => x"00000000", 30476 => x"00000000",
    30477 => x"00000000", 30478 => x"00000000", 30479 => x"00000000",
    30480 => x"00000000", 30481 => x"00000000", 30482 => x"00000000",
    30483 => x"00000000", 30484 => x"00000000", 30485 => x"00000000",
    30486 => x"00000000", 30487 => x"00000000", 30488 => x"00000000",
    30489 => x"00000000", 30490 => x"00000000", 30491 => x"00000000",
    30492 => x"00000000", 30493 => x"00000000", 30494 => x"00000000",
    30495 => x"00000000", 30496 => x"00000000", 30497 => x"00000000",
    30498 => x"00000000", 30499 => x"00000000", 30500 => x"00000000",
    30501 => x"00000000", 30502 => x"00000000", 30503 => x"00000000",
    30504 => x"00000000", 30505 => x"00000000", 30506 => x"00000000",
    30507 => x"00000000", 30508 => x"00000000", 30509 => x"00000000",
    30510 => x"00000000", 30511 => x"00000000", 30512 => x"00000000",
    30513 => x"00000000", 30514 => x"00000000", 30515 => x"00000000",
    30516 => x"00000000", 30517 => x"00000000", 30518 => x"00000000",
    30519 => x"00000000", 30520 => x"00000000", 30521 => x"00000000",
    30522 => x"00000000", 30523 => x"00000000", 30524 => x"00000000",
    30525 => x"00000000", 30526 => x"00000000", 30527 => x"00000000",
    30528 => x"00000000", 30529 => x"00000000", 30530 => x"00000000",
    30531 => x"00000000", 30532 => x"00000000", 30533 => x"00000000",
    30534 => x"00000000", 30535 => x"00000000", 30536 => x"00000000",
    30537 => x"00000000", 30538 => x"00000000", 30539 => x"00000000",
    30540 => x"00000000", 30541 => x"00000000", 30542 => x"00000000",
    30543 => x"00000000", 30544 => x"00000000", 30545 => x"00000000",
    30546 => x"00000000", 30547 => x"00000000", 30548 => x"00000000",
    30549 => x"00000000", 30550 => x"00000000", 30551 => x"00000000",
    30552 => x"00000000", 30553 => x"00000000", 30554 => x"00000000",
    30555 => x"00000000", 30556 => x"00000000", 30557 => x"00000000",
    30558 => x"00000000", 30559 => x"00000000", 30560 => x"00000000",
    30561 => x"00000000", 30562 => x"00000000", 30563 => x"00000000",
    30564 => x"00000000", 30565 => x"00000000", 30566 => x"00000000",
    30567 => x"00000000", 30568 => x"00000000", 30569 => x"00000000",
    30570 => x"00000000", 30571 => x"00000000", 30572 => x"00000000",
    30573 => x"00000000", 30574 => x"00000000", 30575 => x"00000000",
    30576 => x"00000000", 30577 => x"00000000", 30578 => x"00000000",
    30579 => x"00000000", 30580 => x"00000000", 30581 => x"00000000",
    30582 => x"00000000", 30583 => x"00000000", 30584 => x"00000000",
    30585 => x"00000000", 30586 => x"00000000", 30587 => x"00000000",
    30588 => x"00000000", 30589 => x"00000000", 30590 => x"00000000",
    30591 => x"00000000", 30592 => x"00000000", 30593 => x"00000000",
    30594 => x"00000000", 30595 => x"00000000", 30596 => x"00000000",
    30597 => x"00000000", 30598 => x"00000000", 30599 => x"00000000",
    30600 => x"00000000", 30601 => x"00000000", 30602 => x"00000000",
    30603 => x"00000000", 30604 => x"00000000", 30605 => x"00000000",
    30606 => x"00000000", 30607 => x"00000000", 30608 => x"00000000",
    30609 => x"00000000", 30610 => x"00000000", 30611 => x"00000000",
    30612 => x"00000000", 30613 => x"00000000", 30614 => x"00000000",
    30615 => x"00000000", 30616 => x"00000000", 30617 => x"00000000",
    30618 => x"00000000", 30619 => x"00000000", 30620 => x"00000000",
    30621 => x"00000000", 30622 => x"00000000", 30623 => x"00000000",
    30624 => x"00000000", 30625 => x"00000000", 30626 => x"00000000",
    30627 => x"00000000", 30628 => x"00000000", 30629 => x"00000000",
    30630 => x"00000000", 30631 => x"00000000", 30632 => x"00000000",
    30633 => x"00000000", 30634 => x"00000000", 30635 => x"00000000",
    30636 => x"00000000", 30637 => x"00000000", 30638 => x"00000000",
    30639 => x"00000000", 30640 => x"00000000", 30641 => x"00000000",
    30642 => x"00000000", 30643 => x"00000000", 30644 => x"00000000",
    30645 => x"00000000", 30646 => x"00000000", 30647 => x"00000000",
    30648 => x"00000000", 30649 => x"00000000", 30650 => x"00000000",
    30651 => x"00000000", 30652 => x"00000000", 30653 => x"00000000",
    30654 => x"00000000", 30655 => x"00000000", 30656 => x"00000000",
    30657 => x"00000000", 30658 => x"00000000", 30659 => x"00000000",
    30660 => x"00000000", 30661 => x"00000000", 30662 => x"00000000",
    30663 => x"00000000", 30664 => x"00000000", 30665 => x"00000000",
    30666 => x"00000000", 30667 => x"00000000", 30668 => x"00000000",
    30669 => x"00000000", 30670 => x"00000000", 30671 => x"00000000",
    30672 => x"00000000", 30673 => x"00000000", 30674 => x"00000000",
    30675 => x"00000000", 30676 => x"00000000", 30677 => x"00000000",
    30678 => x"00000000", 30679 => x"00000000", 30680 => x"00000000",
    30681 => x"00000000", 30682 => x"00000000", 30683 => x"00000000",
    30684 => x"00000000", 30685 => x"00000000", 30686 => x"00000000",
    30687 => x"00000000", 30688 => x"00000000", 30689 => x"00000000",
    30690 => x"00000000", 30691 => x"00000000", 30692 => x"00000000",
    30693 => x"00000000", 30694 => x"00000000", 30695 => x"00000000",
    30696 => x"00000000", 30697 => x"00000000", 30698 => x"00000000",
    30699 => x"00000000", 30700 => x"00000000", 30701 => x"00000000",
    30702 => x"00000000", 30703 => x"00000000", 30704 => x"00000000",
    30705 => x"00000000", 30706 => x"00000000", 30707 => x"00000000",
    30708 => x"00000000", 30709 => x"00000000", 30710 => x"00000000",
    30711 => x"00000000", 30712 => x"00000000", 30713 => x"00000000",
    30714 => x"00000000", 30715 => x"00000000", 30716 => x"00000000",
    30717 => x"00000000", 30718 => x"00000000", 30719 => x"00000000",
    30720 => x"00000000", 30721 => x"00000000", 30722 => x"00000000",
    30723 => x"00000000", 30724 => x"00000000", 30725 => x"00000000",
    30726 => x"00000000", 30727 => x"00000000", 30728 => x"00000000",
    30729 => x"00000000", 30730 => x"00000000", 30731 => x"00000000",
    30732 => x"00000000", 30733 => x"00000000", 30734 => x"00000000",
    30735 => x"00000000", 30736 => x"00000000", 30737 => x"00000000",
    30738 => x"00000000", 30739 => x"00000000", 30740 => x"00000000",
    30741 => x"00000000", 30742 => x"00000000", 30743 => x"00000000",
    30744 => x"00000000", 30745 => x"00000000", 30746 => x"00000000",
    30747 => x"00000000", 30748 => x"00000000", 30749 => x"00000000",
    30750 => x"00000000", 30751 => x"00000000", 30752 => x"00000000",
    30753 => x"00000000", 30754 => x"00000000", 30755 => x"00000000",
    30756 => x"00000000", 30757 => x"00000000", 30758 => x"00000000",
    30759 => x"00000000", 30760 => x"00000000", 30761 => x"00000000",
    30762 => x"00000000", 30763 => x"00000000", 30764 => x"00000000",
    30765 => x"00000000", 30766 => x"00000000", 30767 => x"00000000",
    30768 => x"00000000", 30769 => x"00000000", 30770 => x"00000000",
    30771 => x"00000000", 30772 => x"00000000", 30773 => x"00000000",
    30774 => x"00000000", 30775 => x"00000000", 30776 => x"00000000",
    30777 => x"00000000", 30778 => x"00000000", 30779 => x"00000000",
    30780 => x"00000000", 30781 => x"00000000", 30782 => x"00000000",
    30783 => x"00000000", 30784 => x"00000000", 30785 => x"00000000",
    30786 => x"00000000", 30787 => x"00000000", 30788 => x"00000000",
    30789 => x"00000000", 30790 => x"00000000", 30791 => x"00000000",
    30792 => x"00000000", 30793 => x"00000000", 30794 => x"00000000",
    30795 => x"00000000", 30796 => x"00000000", 30797 => x"00000000",
    30798 => x"00000000", 30799 => x"00000000", 30800 => x"00000000",
    30801 => x"00000000", 30802 => x"00000000", 30803 => x"00000000",
    30804 => x"00000000", 30805 => x"00000000", 30806 => x"00000000",
    30807 => x"00000000", 30808 => x"00000000", 30809 => x"00000000",
    30810 => x"00000000", 30811 => x"00000000", 30812 => x"00000000",
    30813 => x"00000000", 30814 => x"00000000", 30815 => x"00000000",
    30816 => x"00000000", 30817 => x"00000000", 30818 => x"00000000",
    30819 => x"00000000", 30820 => x"00000000", 30821 => x"00000000",
    30822 => x"00000000", 30823 => x"00000000", 30824 => x"00000000",
    30825 => x"00000000", 30826 => x"00000000", 30827 => x"00000000",
    30828 => x"00000000", 30829 => x"00000000", 30830 => x"00000000",
    30831 => x"00000000", 30832 => x"00000000", 30833 => x"00000000",
    30834 => x"00000000", 30835 => x"00000000", 30836 => x"00000000",
    30837 => x"00000000", 30838 => x"00000000", 30839 => x"00000000",
    30840 => x"00000000", 30841 => x"00000000", 30842 => x"00000000",
    30843 => x"00000000", 30844 => x"00000000", 30845 => x"00000000",
    30846 => x"00000000", 30847 => x"00000000", 30848 => x"00000000",
    30849 => x"00000000", 30850 => x"00000000", 30851 => x"00000000",
    30852 => x"00000000", 30853 => x"00000000", 30854 => x"00000000",
    30855 => x"00000000", 30856 => x"00000000", 30857 => x"00000000",
    30858 => x"00000000", 30859 => x"00000000", 30860 => x"00000000",
    30861 => x"00000000", 30862 => x"00000000", 30863 => x"00000000",
    30864 => x"00000000", 30865 => x"00000000", 30866 => x"00000000",
    30867 => x"00000000", 30868 => x"00000000", 30869 => x"00000000",
    30870 => x"00000000", 30871 => x"00000000", 30872 => x"00000000",
    30873 => x"00000000", 30874 => x"00000000", 30875 => x"00000000",
    30876 => x"00000000", 30877 => x"00000000", 30878 => x"00000000",
    30879 => x"00000000", 30880 => x"00000000", 30881 => x"00000000",
    30882 => x"00000000", 30883 => x"00000000", 30884 => x"00000000",
    30885 => x"00000000", 30886 => x"00000000", 30887 => x"00000000",
    30888 => x"00000000", 30889 => x"00000000", 30890 => x"00000000",
    30891 => x"00000000", 30892 => x"00000000", 30893 => x"00000000",
    30894 => x"00000000", 30895 => x"00000000", 30896 => x"00000000",
    30897 => x"00000000", 30898 => x"00000000", 30899 => x"00000000",
    30900 => x"00000000", 30901 => x"00000000", 30902 => x"00000000",
    30903 => x"00000000", 30904 => x"00000000", 30905 => x"00000000",
    30906 => x"00000000", 30907 => x"00000000", 30908 => x"00000000",
    30909 => x"00000000", 30910 => x"00000000", 30911 => x"00000000",
    30912 => x"00000000", 30913 => x"00000000", 30914 => x"00000000",
    30915 => x"00000000", 30916 => x"00000000", 30917 => x"00000000",
    30918 => x"00000000", 30919 => x"00000000", 30920 => x"00000000",
    30921 => x"00000000", 30922 => x"00000000", 30923 => x"00000000",
    30924 => x"00000000", 30925 => x"00000000", 30926 => x"00000000",
    30927 => x"00000000", 30928 => x"00000000", 30929 => x"00000000",
    30930 => x"00000000", 30931 => x"00000000", 30932 => x"00000000",
    30933 => x"00000000", 30934 => x"00000000", 30935 => x"00000000",
    30936 => x"00000000", 30937 => x"00000000", 30938 => x"00000000",
    30939 => x"00000000", 30940 => x"00000000", 30941 => x"00000000",
    30942 => x"00000000", 30943 => x"00000000", 30944 => x"00000000",
    30945 => x"00000000", 30946 => x"00000000", 30947 => x"00000000",
    30948 => x"00000000", 30949 => x"00000000", 30950 => x"00000000",
    30951 => x"00000000", 30952 => x"00000000", 30953 => x"00000000",
    30954 => x"00000000", 30955 => x"00000000", 30956 => x"00000000",
    30957 => x"00000000", 30958 => x"00000000", 30959 => x"00000000",
    30960 => x"00000000", 30961 => x"00000000", 30962 => x"00000000",
    30963 => x"00000000", 30964 => x"00000000", 30965 => x"00000000",
    30966 => x"00000000", 30967 => x"00000000", 30968 => x"00000000",
    30969 => x"00000000", 30970 => x"00000000", 30971 => x"00000000",
    30972 => x"00000000", 30973 => x"00000000", 30974 => x"00000000",
    30975 => x"00000000", 30976 => x"00000000", 30977 => x"00000000",
    30978 => x"00000000", 30979 => x"00000000", 30980 => x"00000000",
    30981 => x"00000000", 30982 => x"00000000", 30983 => x"00000000",
    30984 => x"00000000", 30985 => x"00000000", 30986 => x"00000000",
    30987 => x"00000000", 30988 => x"00000000", 30989 => x"00000000",
    30990 => x"00000000", 30991 => x"00000000", 30992 => x"00000000",
    30993 => x"00000000", 30994 => x"00000000", 30995 => x"00000000",
    30996 => x"00000000", 30997 => x"00000000", 30998 => x"00000000",
    30999 => x"00000000", 31000 => x"00000000", 31001 => x"00000000",
    31002 => x"00000000", 31003 => x"00000000", 31004 => x"00000000",
    31005 => x"00000000", 31006 => x"00000000", 31007 => x"00000000",
    31008 => x"00000000", 31009 => x"00000000", 31010 => x"00000000",
    31011 => x"00000000", 31012 => x"00000000", 31013 => x"00000000",
    31014 => x"00000000", 31015 => x"00000000", 31016 => x"00000000",
    31017 => x"00000000", 31018 => x"00000000", 31019 => x"00000000",
    31020 => x"00000000", 31021 => x"00000000", 31022 => x"00000000",
    31023 => x"00000000", 31024 => x"00000000", 31025 => x"00000000",
    31026 => x"00000000", 31027 => x"00000000", 31028 => x"00000000",
    31029 => x"00000000", 31030 => x"00000000", 31031 => x"00000000",
    31032 => x"00000000", 31033 => x"00000000", 31034 => x"00000000",
    31035 => x"00000000", 31036 => x"00000000", 31037 => x"00000000",
    31038 => x"00000000", 31039 => x"00000000", 31040 => x"00000000",
    31041 => x"00000000", 31042 => x"00000000", 31043 => x"00000000",
    31044 => x"00000000", 31045 => x"00000000", 31046 => x"00000000",
    31047 => x"00000000", 31048 => x"00000000", 31049 => x"00000000",
    31050 => x"00000000", 31051 => x"00000000", 31052 => x"00000000",
    31053 => x"00000000", 31054 => x"00000000", 31055 => x"00000000",
    31056 => x"00000000", 31057 => x"00000000", 31058 => x"00000000",
    31059 => x"00000000", 31060 => x"00000000", 31061 => x"00000000",
    31062 => x"00000000", 31063 => x"00000000", 31064 => x"00000000",
    31065 => x"00000000", 31066 => x"00000000", 31067 => x"00000000",
    31068 => x"00000000", 31069 => x"00000000", 31070 => x"00000000",
    31071 => x"00000000", 31072 => x"00000000", 31073 => x"00000000",
    31074 => x"00000000", 31075 => x"00000000", 31076 => x"00000000",
    31077 => x"00000000", 31078 => x"00000000", 31079 => x"00000000",
    31080 => x"00000000", 31081 => x"00000000", 31082 => x"00000000",
    31083 => x"00000000", 31084 => x"00000000", 31085 => x"00000000",
    31086 => x"00000000", 31087 => x"00000000", 31088 => x"00000000",
    31089 => x"00000000", 31090 => x"00000000", 31091 => x"00000000",
    31092 => x"00000000", 31093 => x"00000000", 31094 => x"00000000",
    31095 => x"00000000", 31096 => x"00000000", 31097 => x"00000000",
    31098 => x"00000000", 31099 => x"00000000", 31100 => x"00000000",
    31101 => x"00000000", 31102 => x"00000000", 31103 => x"00000000",
    31104 => x"00000000", 31105 => x"00000000", 31106 => x"00000000",
    31107 => x"00000000", 31108 => x"00000000", 31109 => x"00000000",
    31110 => x"00000000", 31111 => x"00000000", 31112 => x"00000000",
    31113 => x"00000000", 31114 => x"00000000", 31115 => x"00000000",
    31116 => x"00000000", 31117 => x"00000000", 31118 => x"00000000",
    31119 => x"00000000", 31120 => x"00000000", 31121 => x"00000000",
    31122 => x"00000000", 31123 => x"00000000", 31124 => x"00000000",
    31125 => x"00000000", 31126 => x"00000000", 31127 => x"00000000",
    31128 => x"00000000", 31129 => x"00000000", 31130 => x"00000000",
    31131 => x"00000000", 31132 => x"00000000", 31133 => x"00000000",
    31134 => x"00000000", 31135 => x"00000000", 31136 => x"00000000",
    31137 => x"00000000", 31138 => x"00000000", 31139 => x"00000000",
    31140 => x"00000000", 31141 => x"00000000", 31142 => x"00000000",
    31143 => x"00000000", 31144 => x"00000000", 31145 => x"00000000",
    31146 => x"00000000", 31147 => x"00000000", 31148 => x"00000000",
    31149 => x"00000000", 31150 => x"00000000", 31151 => x"00000000",
    31152 => x"00000000", 31153 => x"00000000", 31154 => x"00000000",
    31155 => x"00000000", 31156 => x"00000000", 31157 => x"00000000",
    31158 => x"00000000", 31159 => x"00000000", 31160 => x"00000000",
    31161 => x"00000000", 31162 => x"00000000", 31163 => x"00000000",
    31164 => x"00000000", 31165 => x"00000000", 31166 => x"00000000",
    31167 => x"00000000", 31168 => x"00000000", 31169 => x"00000000",
    31170 => x"00000000", 31171 => x"00000000", 31172 => x"00000000",
    31173 => x"00000000", 31174 => x"00000000", 31175 => x"00000000",
    31176 => x"00000000", 31177 => x"00000000", 31178 => x"00000000",
    31179 => x"00000000", 31180 => x"00000000", 31181 => x"00000000",
    31182 => x"00000000", 31183 => x"00000000", 31184 => x"00000000",
    31185 => x"00000000", 31186 => x"00000000", 31187 => x"00000000",
    31188 => x"00000000", 31189 => x"00000000", 31190 => x"00000000",
    31191 => x"00000000", 31192 => x"00000000", 31193 => x"00000000",
    31194 => x"00000000", 31195 => x"00000000", 31196 => x"00000000",
    31197 => x"00000000", 31198 => x"00000000", 31199 => x"00000000",
    31200 => x"00000000", 31201 => x"00000000", 31202 => x"00000000",
    31203 => x"00000000", 31204 => x"00000000", 31205 => x"00000000",
    31206 => x"00000000", 31207 => x"00000000", 31208 => x"00000000",
    31209 => x"00000000", 31210 => x"00000000", 31211 => x"00000000",
    31212 => x"00000000", 31213 => x"00000000", 31214 => x"00000000",
    31215 => x"00000000", 31216 => x"00000000", 31217 => x"00000000",
    31218 => x"00000000", 31219 => x"00000000", 31220 => x"00000000",
    31221 => x"00000000", 31222 => x"00000000", 31223 => x"00000000",
    31224 => x"00000000", 31225 => x"00000000", 31226 => x"00000000",
    31227 => x"00000000", 31228 => x"00000000", 31229 => x"00000000",
    31230 => x"00000000", 31231 => x"00000000", 31232 => x"00000000",
    31233 => x"00000000", 31234 => x"00000000", 31235 => x"00000000",
    31236 => x"00000000", 31237 => x"00000000", 31238 => x"00000000",
    31239 => x"00000000", 31240 => x"00000000", 31241 => x"00000000",
    31242 => x"00000000", 31243 => x"00000000", 31244 => x"00000000",
    31245 => x"00000000", 31246 => x"00000000", 31247 => x"00000000",
    31248 => x"00000000", 31249 => x"00000000", 31250 => x"00000000",
    31251 => x"00000000", 31252 => x"00000000", 31253 => x"00000000",
    31254 => x"00000000", 31255 => x"00000000", 31256 => x"00000000",
    31257 => x"00000000", 31258 => x"00000000", 31259 => x"00000000",
    31260 => x"00000000", 31261 => x"00000000", 31262 => x"00000000",
    31263 => x"00000000", 31264 => x"00000000", 31265 => x"00000000",
    31266 => x"00000000", 31267 => x"00000000", 31268 => x"00000000",
    31269 => x"00000000", 31270 => x"00000000", 31271 => x"00000000",
    31272 => x"00000000", 31273 => x"00000000", 31274 => x"00000000",
    31275 => x"00000000", 31276 => x"00000000", 31277 => x"00000000",
    31278 => x"00000000", 31279 => x"00000000", 31280 => x"00000000",
    31281 => x"00000000", 31282 => x"00000000", 31283 => x"00000000",
    31284 => x"00000000", 31285 => x"00000000", 31286 => x"00000000",
    31287 => x"00000000", 31288 => x"00000000", 31289 => x"00000000",
    31290 => x"00000000", 31291 => x"00000000", 31292 => x"00000000",
    31293 => x"00000000", 31294 => x"00000000", 31295 => x"00000000",
    31296 => x"00000000", 31297 => x"00000000", 31298 => x"00000000",
    31299 => x"00000000", 31300 => x"00000000", 31301 => x"00000000",
    31302 => x"00000000", 31303 => x"00000000", 31304 => x"00000000",
    31305 => x"00000000", 31306 => x"00000000", 31307 => x"00000000",
    31308 => x"00000000", 31309 => x"00000000", 31310 => x"00000000",
    31311 => x"00000000", 31312 => x"00000000", 31313 => x"00000000",
    31314 => x"00000000", 31315 => x"00000000", 31316 => x"00000000",
    31317 => x"00000000", 31318 => x"00000000", 31319 => x"00000000",
    31320 => x"00000000", 31321 => x"00000000", 31322 => x"00000000",
    31323 => x"00000000", 31324 => x"00000000", 31325 => x"00000000",
    31326 => x"00000000", 31327 => x"00000000", 31328 => x"00000000",
    31329 => x"00000000", 31330 => x"00000000", 31331 => x"00000000",
    31332 => x"00000000", 31333 => x"00000000", 31334 => x"00000000",
    31335 => x"00000000", 31336 => x"00000000", 31337 => x"00000000",
    31338 => x"00000000", 31339 => x"00000000", 31340 => x"00000000",
    31341 => x"00000000", 31342 => x"00000000", 31343 => x"00000000",
    31344 => x"00000000", 31345 => x"00000000", 31346 => x"00000000",
    31347 => x"00000000", 31348 => x"00000000", 31349 => x"00000000",
    31350 => x"00000000", 31351 => x"00000000", 31352 => x"00000000",
    31353 => x"00000000", 31354 => x"00000000", 31355 => x"00000000",
    31356 => x"00000000", 31357 => x"00000000", 31358 => x"00000000",
    31359 => x"00000000", 31360 => x"00000000", 31361 => x"00000000",
    31362 => x"00000000", 31363 => x"00000000", 31364 => x"00000000",
    31365 => x"00000000", 31366 => x"00000000", 31367 => x"00000000",
    31368 => x"00000000", 31369 => x"00000000", 31370 => x"00000000",
    31371 => x"00000000", 31372 => x"00000000", 31373 => x"00000000",
    31374 => x"00000000", 31375 => x"00000000", 31376 => x"00000000",
    31377 => x"00000000", 31378 => x"00000000", 31379 => x"00000000",
    31380 => x"00000000", 31381 => x"00000000", 31382 => x"00000000",
    31383 => x"00000000", 31384 => x"00000000", 31385 => x"00000000",
    31386 => x"00000000", 31387 => x"00000000", 31388 => x"00000000",
    31389 => x"00000000", 31390 => x"00000000", 31391 => x"00000000",
    31392 => x"00000000", 31393 => x"00000000", 31394 => x"00000000",
    31395 => x"00000000", 31396 => x"00000000", 31397 => x"00000000",
    31398 => x"00000000", 31399 => x"00000000", 31400 => x"00000000",
    31401 => x"00000000", 31402 => x"00000000", 31403 => x"00000000",
    31404 => x"00000000", 31405 => x"00000000", 31406 => x"00000000",
    31407 => x"00000000", 31408 => x"00000000", 31409 => x"00000000",
    31410 => x"00000000", 31411 => x"00000000", 31412 => x"00000000",
    31413 => x"00000000", 31414 => x"00000000", 31415 => x"00000000",
    31416 => x"00000000", 31417 => x"00000000", 31418 => x"00000000",
    31419 => x"00000000", 31420 => x"00000000", 31421 => x"00000000",
    31422 => x"00000000", 31423 => x"00000000", 31424 => x"00000000",
    31425 => x"00000000", 31426 => x"00000000", 31427 => x"00000000",
    31428 => x"00000000", 31429 => x"00000000", 31430 => x"00000000",
    31431 => x"00000000", 31432 => x"00000000", 31433 => x"00000000",
    31434 => x"00000000", 31435 => x"00000000", 31436 => x"00000000",
    31437 => x"00000000", 31438 => x"00000000", 31439 => x"00000000",
    31440 => x"00000000", 31441 => x"00000000", 31442 => x"00000000",
    31443 => x"00000000", 31444 => x"00000000", 31445 => x"00000000",
    31446 => x"00000000", 31447 => x"00000000", 31448 => x"00000000",
    31449 => x"00000000", 31450 => x"00000000", 31451 => x"00000000",
    31452 => x"00000000", 31453 => x"00000000", 31454 => x"00000000",
    31455 => x"00000000", 31456 => x"00000000", 31457 => x"00000000",
    31458 => x"00000000", 31459 => x"00000000", 31460 => x"00000000",
    31461 => x"00000000", 31462 => x"00000000", 31463 => x"00000000",
    31464 => x"00000000", 31465 => x"00000000", 31466 => x"00000000",
    31467 => x"00000000", 31468 => x"00000000", 31469 => x"00000000",
    31470 => x"00000000", 31471 => x"00000000", 31472 => x"00000000",
    31473 => x"00000000", 31474 => x"00000000", 31475 => x"00000000",
    31476 => x"00000000", 31477 => x"00000000", 31478 => x"00000000",
    31479 => x"00000000", 31480 => x"00000000", 31481 => x"00000000",
    31482 => x"00000000", 31483 => x"00000000", 31484 => x"00000000",
    31485 => x"00000000", 31486 => x"00000000", 31487 => x"00000000",
    31488 => x"00000000", 31489 => x"00000000", 31490 => x"00000000",
    31491 => x"00000000", 31492 => x"00000000", 31493 => x"00000000",
    31494 => x"00000000", 31495 => x"00000000", 31496 => x"00000000",
    31497 => x"00000000", 31498 => x"00000000", 31499 => x"00000000",
    31500 => x"00000000", 31501 => x"00000000", 31502 => x"00000000",
    31503 => x"00000000", 31504 => x"00000000", 31505 => x"00000000",
    31506 => x"00000000", 31507 => x"00000000", 31508 => x"00000000",
    31509 => x"00000000", 31510 => x"00000000", 31511 => x"00000000",
    31512 => x"00000000", 31513 => x"00000000", 31514 => x"00000000",
    31515 => x"00000000", 31516 => x"00000000", 31517 => x"00000000",
    31518 => x"00000000", 31519 => x"00000000", 31520 => x"00000000",
    31521 => x"00000000", 31522 => x"00000000", 31523 => x"00000000",
    31524 => x"00000000", 31525 => x"00000000", 31526 => x"00000000",
    31527 => x"00000000", 31528 => x"00000000", 31529 => x"00000000",
    31530 => x"00000000", 31531 => x"00000000", 31532 => x"00000000",
    31533 => x"00000000", 31534 => x"00000000", 31535 => x"00000000",
    31536 => x"00000000", 31537 => x"00000000", 31538 => x"00000000",
    31539 => x"00000000", 31540 => x"00000000", 31541 => x"00000000",
    31542 => x"00000000", 31543 => x"00000000", 31544 => x"00000000",
    31545 => x"00000000", 31546 => x"00000000", 31547 => x"00000000",
    31548 => x"00000000", 31549 => x"00000000", 31550 => x"00000000",
    31551 => x"00000000", 31552 => x"00000000", 31553 => x"00000000",
    31554 => x"00000000", 31555 => x"00000000", 31556 => x"00000000",
    31557 => x"00000000", 31558 => x"00000000", 31559 => x"00000000",
    31560 => x"00000000", 31561 => x"00000000", 31562 => x"00000000",
    31563 => x"00000000", 31564 => x"00000000", 31565 => x"00000000",
    31566 => x"00000000", 31567 => x"00000000", 31568 => x"00000000",
    31569 => x"00000000", 31570 => x"00000000", 31571 => x"00000000",
    31572 => x"00000000", 31573 => x"00000000", 31574 => x"00000000",
    31575 => x"00000000", 31576 => x"00000000", 31577 => x"00000000",
    31578 => x"00000000", 31579 => x"00000000", 31580 => x"00000000",
    31581 => x"00000000", 31582 => x"00000000", 31583 => x"00000000",
    31584 => x"00000000", 31585 => x"00000000", 31586 => x"00000000",
    31587 => x"00000000", 31588 => x"00000000", 31589 => x"00000000",
    31590 => x"00000000", 31591 => x"00000000", 31592 => x"00000000",
    31593 => x"00000000", 31594 => x"00000000", 31595 => x"00000000",
    31596 => x"00000000", 31597 => x"00000000", 31598 => x"00000000",
    31599 => x"00000000", 31600 => x"00000000", 31601 => x"00000000",
    31602 => x"00000000", 31603 => x"00000000", 31604 => x"00000000",
    31605 => x"00000000", 31606 => x"00000000", 31607 => x"00000000",
    31608 => x"00000000", 31609 => x"00000000", 31610 => x"00000000",
    31611 => x"00000000", 31612 => x"00000000", 31613 => x"00000000",
    31614 => x"00000000", 31615 => x"00000000", 31616 => x"00000000",
    31617 => x"00000000", 31618 => x"00000000", 31619 => x"00000000",
    31620 => x"00000000", 31621 => x"00000000", 31622 => x"00000000",
    31623 => x"00000000", 31624 => x"00000000", 31625 => x"00000000",
    31626 => x"00000000", 31627 => x"00000000", 31628 => x"00000000",
    31629 => x"00000000", 31630 => x"00000000", 31631 => x"00000000",
    31632 => x"00000000", 31633 => x"00000000", 31634 => x"00000000",
    31635 => x"00000000", 31636 => x"00000000", 31637 => x"00000000",
    31638 => x"00000000", 31639 => x"00000000", 31640 => x"00000000",
    31641 => x"00000000", 31642 => x"00000000", 31643 => x"00000000",
    31644 => x"00000000", 31645 => x"00000000", 31646 => x"00000000",
    31647 => x"00000000", 31648 => x"00000000", 31649 => x"00000000",
    31650 => x"00000000", 31651 => x"00000000", 31652 => x"00000000",
    31653 => x"00000000", 31654 => x"00000000", 31655 => x"00000000",
    31656 => x"00000000", 31657 => x"00000000", 31658 => x"00000000",
    31659 => x"00000000", 31660 => x"00000000", 31661 => x"00000000",
    31662 => x"00000000", 31663 => x"00000000", 31664 => x"00000000",
    31665 => x"00000000", 31666 => x"00000000", 31667 => x"00000000",
    31668 => x"00000000", 31669 => x"00000000", 31670 => x"00000000",
    31671 => x"00000000", 31672 => x"00000000", 31673 => x"00000000",
    31674 => x"00000000", 31675 => x"00000000", 31676 => x"00000000",
    31677 => x"00000000", 31678 => x"00000000", 31679 => x"00000000",
    31680 => x"00000000", 31681 => x"00000000", 31682 => x"00000000",
    31683 => x"00000000", 31684 => x"00000000", 31685 => x"00000000",
    31686 => x"00000000", 31687 => x"00000000", 31688 => x"00000000",
    31689 => x"00000000", 31690 => x"00000000", 31691 => x"00000000",
    31692 => x"00000000", 31693 => x"00000000", 31694 => x"00000000",
    31695 => x"00000000", 31696 => x"00000000", 31697 => x"00000000",
    31698 => x"00000000", 31699 => x"00000000", 31700 => x"00000000",
    31701 => x"00000000", 31702 => x"00000000", 31703 => x"00000000",
    31704 => x"00000000", 31705 => x"00000000", 31706 => x"00000000",
    31707 => x"00000000", 31708 => x"00000000", 31709 => x"00000000",
    31710 => x"00000000", 31711 => x"00000000", 31712 => x"00000000",
    31713 => x"00000000", 31714 => x"00000000", 31715 => x"00000000",
    31716 => x"00000000", 31717 => x"00000000", 31718 => x"00000000",
    31719 => x"00000000", 31720 => x"00000000", 31721 => x"00000000",
    31722 => x"00000000", 31723 => x"00000000", 31724 => x"00000000",
    31725 => x"00000000", 31726 => x"00000000", 31727 => x"00000000",
    31728 => x"00000000", 31729 => x"00000000", 31730 => x"00000000",
    31731 => x"00000000", 31732 => x"00000000", 31733 => x"00000000",
    31734 => x"00000000", 31735 => x"00000000", 31736 => x"00000000",
    31737 => x"00000000", 31738 => x"00000000", 31739 => x"00000000",
    31740 => x"00000000", 31741 => x"00000000", 31742 => x"00000000",
    31743 => x"00000000", 31744 => x"00000000", 31745 => x"00000000",
    31746 => x"00000000", 31747 => x"00000000", 31748 => x"00000000",
    31749 => x"00000000", 31750 => x"00000000", 31751 => x"00000000",
    31752 => x"00000000", 31753 => x"00000000", 31754 => x"00000000",
    31755 => x"00000000", 31756 => x"00000000", 31757 => x"00000000",
    31758 => x"00000000", 31759 => x"00000000", 31760 => x"00000000",
    31761 => x"00000000", 31762 => x"00000000", 31763 => x"00000000",
    31764 => x"00000000", 31765 => x"00000000", 31766 => x"00000000",
    31767 => x"00000000", 31768 => x"00000000", 31769 => x"00000000",
    31770 => x"00000000", 31771 => x"00000000", 31772 => x"00000000",
    31773 => x"00000000", 31774 => x"00000000", 31775 => x"00000000",
    31776 => x"00000000", 31777 => x"00000000", 31778 => x"00000000",
    31779 => x"00000000", 31780 => x"00000000", 31781 => x"00000000",
    31782 => x"00000000", 31783 => x"00000000", 31784 => x"00000000",
    31785 => x"00000000", 31786 => x"00000000", 31787 => x"00000000",
    31788 => x"00000000", 31789 => x"00000000", 31790 => x"00000000",
    31791 => x"00000000", 31792 => x"00000000", 31793 => x"00000000",
    31794 => x"00000000", 31795 => x"00000000", 31796 => x"00000000",
    31797 => x"00000000", 31798 => x"00000000", 31799 => x"00000000",
    31800 => x"00000000", 31801 => x"00000000", 31802 => x"00000000",
    31803 => x"00000000", 31804 => x"00000000", 31805 => x"00000000",
    31806 => x"00000000", 31807 => x"00000000", 31808 => x"00000000",
    31809 => x"00000000", 31810 => x"00000000", 31811 => x"00000000",
    31812 => x"00000000", 31813 => x"00000000", 31814 => x"00000000",
    31815 => x"00000000", 31816 => x"00000000", 31817 => x"00000000",
    31818 => x"00000000", 31819 => x"00000000", 31820 => x"00000000",
    31821 => x"00000000", 31822 => x"00000000", 31823 => x"00000000",
    31824 => x"00000000", 31825 => x"00000000", 31826 => x"00000000",
    31827 => x"00000000", 31828 => x"00000000", 31829 => x"00000000",
    31830 => x"00000000", 31831 => x"00000000", 31832 => x"00000000",
    31833 => x"00000000", 31834 => x"00000000", 31835 => x"00000000",
    31836 => x"00000000", 31837 => x"00000000", 31838 => x"00000000",
    31839 => x"00000000", 31840 => x"00000000", 31841 => x"00000000",
    31842 => x"00000000", 31843 => x"00000000", 31844 => x"00000000",
    31845 => x"00000000", 31846 => x"00000000", 31847 => x"00000000",
    31848 => x"00000000", 31849 => x"00000000", 31850 => x"00000000",
    31851 => x"00000000", 31852 => x"00000000", 31853 => x"00000000",
    31854 => x"00000000", 31855 => x"00000000", 31856 => x"00000000",
    31857 => x"00000000", 31858 => x"00000000", 31859 => x"00000000",
    31860 => x"00000000", 31861 => x"00000000", 31862 => x"00000000",
    31863 => x"00000000", 31864 => x"00000000", 31865 => x"00000000",
    31866 => x"00000000", 31867 => x"00000000", 31868 => x"00000000",
    31869 => x"00000000", 31870 => x"00000000", 31871 => x"00000000",
    31872 => x"00000000", 31873 => x"00000000", 31874 => x"00000000",
    31875 => x"00000000", 31876 => x"00000000", 31877 => x"00000000",
    31878 => x"00000000", 31879 => x"00000000", 31880 => x"00000000",
    31881 => x"00000000", 31882 => x"00000000", 31883 => x"00000000",
    31884 => x"00000000", 31885 => x"00000000", 31886 => x"00000000",
    31887 => x"00000000", 31888 => x"00000000", 31889 => x"00000000",
    31890 => x"00000000", 31891 => x"00000000", 31892 => x"00000000",
    31893 => x"00000000", 31894 => x"00000000", 31895 => x"00000000",
    31896 => x"00000000", 31897 => x"00000000", 31898 => x"00000000",
    31899 => x"00000000", 31900 => x"00000000", 31901 => x"00000000",
    31902 => x"00000000", 31903 => x"00000000", 31904 => x"00000000",
    31905 => x"00000000", 31906 => x"00000000", 31907 => x"00000000",
    31908 => x"00000000", 31909 => x"00000000", 31910 => x"00000000",
    31911 => x"00000000", 31912 => x"00000000", 31913 => x"00000000",
    31914 => x"00000000", 31915 => x"00000000", 31916 => x"00000000",
    31917 => x"00000000", 31918 => x"00000000", 31919 => x"00000000",
    31920 => x"00000000", 31921 => x"00000000", 31922 => x"00000000",
    31923 => x"00000000", 31924 => x"00000000", 31925 => x"00000000",
    31926 => x"00000000", 31927 => x"00000000", 31928 => x"00000000",
    31929 => x"00000000", 31930 => x"00000000", 31931 => x"00000000",
    31932 => x"00000000", 31933 => x"00000000", 31934 => x"00000000",
    31935 => x"00000000", 31936 => x"00000000", 31937 => x"00000000",
    31938 => x"00000000", 31939 => x"00000000", 31940 => x"00000000",
    31941 => x"00000000", 31942 => x"00000000", 31943 => x"00000000",
    31944 => x"00000000", 31945 => x"00000000", 31946 => x"00000000",
    31947 => x"00000000", 31948 => x"00000000", 31949 => x"00000000",
    31950 => x"00000000", 31951 => x"00000000", 31952 => x"00000000",
    31953 => x"00000000", 31954 => x"00000000", 31955 => x"00000000",
    31956 => x"00000000", 31957 => x"00000000", 31958 => x"00000000",
    31959 => x"00000000", 31960 => x"00000000", 31961 => x"00000000",
    31962 => x"00000000", 31963 => x"00000000", 31964 => x"00000000",
    31965 => x"00000000", 31966 => x"00000000", 31967 => x"00000000",
    31968 => x"00000000", 31969 => x"00000000", 31970 => x"00000000",
    31971 => x"00000000", 31972 => x"00000000", 31973 => x"00000000",
    31974 => x"00000000", 31975 => x"00000000", 31976 => x"00000000",
    31977 => x"00000000", 31978 => x"00000000", 31979 => x"00000000",
    31980 => x"00000000", 31981 => x"00000000", 31982 => x"00000000",
    31983 => x"00000000", 31984 => x"00000000", 31985 => x"00000000",
    31986 => x"00000000", 31987 => x"00000000", 31988 => x"00000000",
    31989 => x"00000000", 31990 => x"00000000", 31991 => x"00000000",
    31992 => x"00000000", 31993 => x"00000000", 31994 => x"00000000",
    31995 => x"00000000", 31996 => x"00000000", 31997 => x"00000000",
    31998 => x"00000000", 31999 => x"00000000", 32000 => x"00000000",
    32001 => x"00000000", 32002 => x"00000000", 32003 => x"00000000",
    32004 => x"00000000", 32005 => x"00000000", 32006 => x"00000000",
    32007 => x"00000000", 32008 => x"00000000", 32009 => x"00000000",
    32010 => x"00000000", 32011 => x"00000000", 32012 => x"00000000",
    32013 => x"00000000", 32014 => x"00000000", 32015 => x"00000000",
    32016 => x"00000000", 32017 => x"00000000", 32018 => x"00000000",
    32019 => x"00000000", 32020 => x"00000000", 32021 => x"00000000",
    32022 => x"00000000", 32023 => x"00000000", 32024 => x"00000000",
    32025 => x"00000000", 32026 => x"00000000", 32027 => x"00000000",
    32028 => x"00000000", 32029 => x"00000000", 32030 => x"00000000",
    32031 => x"00000000", 32032 => x"00000000", 32033 => x"00000000",
    32034 => x"00000000", 32035 => x"00000000", 32036 => x"00000000",
    32037 => x"00000000", 32038 => x"00000000", 32039 => x"00000000",
    32040 => x"00000000", 32041 => x"00000000", 32042 => x"00000000",
    32043 => x"00000000", 32044 => x"00000000", 32045 => x"00000000",
    32046 => x"00000000", 32047 => x"00000000", 32048 => x"00000000",
    32049 => x"00000000", 32050 => x"00000000", 32051 => x"00000000",
    32052 => x"00000000", 32053 => x"00000000", 32054 => x"00000000",
    32055 => x"00000000", 32056 => x"00000000", 32057 => x"00000000",
    32058 => x"00000000", 32059 => x"00000000", 32060 => x"00000000",
    32061 => x"00000000", 32062 => x"00000000", 32063 => x"00000000",
    32064 => x"00000000", 32065 => x"00000000", 32066 => x"00000000",
    32067 => x"00000000", 32068 => x"00000000", 32069 => x"00000000",
    32070 => x"00000000", 32071 => x"00000000", 32072 => x"00000000",
    32073 => x"00000000", 32074 => x"00000000", 32075 => x"00000000",
    32076 => x"00000000", 32077 => x"00000000", 32078 => x"00000000",
    32079 => x"00000000", 32080 => x"00000000", 32081 => x"00000000",
    32082 => x"00000000", 32083 => x"00000000", 32084 => x"00000000",
    32085 => x"00000000", 32086 => x"00000000", 32087 => x"00000000",
    32088 => x"00000000", 32089 => x"00000000", 32090 => x"00000000",
    32091 => x"00000000", 32092 => x"00000000", 32093 => x"00000000",
    32094 => x"00000000", 32095 => x"00000000", 32096 => x"00000000",
    32097 => x"00000000", 32098 => x"00000000", 32099 => x"00000000",
    32100 => x"00000000", 32101 => x"00000000", 32102 => x"00000000",
    32103 => x"00000000", 32104 => x"00000000", 32105 => x"00000000",
    32106 => x"00000000", 32107 => x"00000000", 32108 => x"00000000",
    32109 => x"00000000", 32110 => x"00000000", 32111 => x"00000000",
    32112 => x"00000000", 32113 => x"00000000", 32114 => x"00000000",
    32115 => x"00000000", 32116 => x"00000000", 32117 => x"00000000",
    32118 => x"00000000", 32119 => x"00000000", 32120 => x"00000000",
    32121 => x"00000000", 32122 => x"00000000", 32123 => x"00000000",
    32124 => x"00000000", 32125 => x"00000000", 32126 => x"00000000",
    32127 => x"00000000", 32128 => x"00000000", 32129 => x"00000000",
    32130 => x"00000000", 32131 => x"00000000", 32132 => x"00000000",
    32133 => x"00000000", 32134 => x"00000000", 32135 => x"00000000",
    32136 => x"00000000", 32137 => x"00000000", 32138 => x"00000000",
    32139 => x"00000000", 32140 => x"00000000", 32141 => x"00000000",
    32142 => x"00000000", 32143 => x"00000000", 32144 => x"00000000",
    32145 => x"00000000", 32146 => x"00000000", 32147 => x"00000000",
    32148 => x"00000000", 32149 => x"00000000", 32150 => x"00000000",
    32151 => x"00000000", 32152 => x"00000000", 32153 => x"00000000",
    32154 => x"00000000", 32155 => x"00000000", 32156 => x"00000000",
    32157 => x"00000000", 32158 => x"00000000", 32159 => x"00000000",
    32160 => x"00000000", 32161 => x"00000000", 32162 => x"00000000",
    32163 => x"00000000", 32164 => x"00000000", 32165 => x"00000000",
    32166 => x"00000000", 32167 => x"00000000", 32168 => x"00000000",
    32169 => x"00000000", 32170 => x"00000000", 32171 => x"00000000",
    32172 => x"00000000", 32173 => x"00000000", 32174 => x"00000000",
    32175 => x"00000000", 32176 => x"00000000", 32177 => x"00000000",
    32178 => x"00000000", 32179 => x"00000000", 32180 => x"00000000",
    32181 => x"00000000", 32182 => x"00000000", 32183 => x"00000000",
    32184 => x"00000000", 32185 => x"00000000", 32186 => x"00000000",
    32187 => x"00000000", 32188 => x"00000000", 32189 => x"00000000",
    32190 => x"00000000", 32191 => x"00000000", 32192 => x"00000000",
    32193 => x"00000000", 32194 => x"00000000", 32195 => x"00000000",
    32196 => x"00000000", 32197 => x"00000000", 32198 => x"00000000",
    32199 => x"00000000", 32200 => x"00000000", 32201 => x"00000000",
    32202 => x"00000000", 32203 => x"00000000", 32204 => x"00000000",
    32205 => x"00000000", 32206 => x"00000000", 32207 => x"00000000",
    32208 => x"00000000", 32209 => x"00000000", 32210 => x"00000000",
    32211 => x"00000000", 32212 => x"00000000", 32213 => x"00000000",
    32214 => x"00000000", 32215 => x"00000000", 32216 => x"00000000",
    32217 => x"00000000", 32218 => x"00000000", 32219 => x"00000000",
    32220 => x"00000000", 32221 => x"00000000", 32222 => x"00000000",
    32223 => x"00000000", 32224 => x"00000000", 32225 => x"00000000",
    32226 => x"00000000", 32227 => x"00000000", 32228 => x"00000000",
    32229 => x"00000000", 32230 => x"00000000", 32231 => x"00000000",
    32232 => x"00000000", 32233 => x"00000000", 32234 => x"00000000",
    32235 => x"00000000", 32236 => x"00000000", 32237 => x"00000000",
    32238 => x"00000000", 32239 => x"00000000", 32240 => x"00000000",
    32241 => x"00000000", 32242 => x"00000000", 32243 => x"00000000",
    32244 => x"00000000", 32245 => x"00000000", 32246 => x"00000000",
    32247 => x"00000000", 32248 => x"00000000", 32249 => x"00000000",
    32250 => x"00000000", 32251 => x"00000000", 32252 => x"00000000",
    32253 => x"00000000", 32254 => x"00000000", 32255 => x"00000000",
    32256 => x"00000000", 32257 => x"00000000", 32258 => x"00000000",
    32259 => x"00000000", 32260 => x"00000000", 32261 => x"00000000",
    32262 => x"00000000", 32263 => x"00000000", 32264 => x"00000000",
    32265 => x"00000000", 32266 => x"00000000", 32267 => x"00000000",
    32268 => x"00000000", 32269 => x"00000000", 32270 => x"00000000",
    32271 => x"00000000", 32272 => x"00000000", 32273 => x"00000000",
    32274 => x"00000000", 32275 => x"00000000", 32276 => x"00000000",
    32277 => x"00000000", 32278 => x"00000000", 32279 => x"00000000",
    32280 => x"00000000", 32281 => x"00000000", 32282 => x"00000000",
    32283 => x"00000000", 32284 => x"00000000", 32285 => x"00000000",
    32286 => x"00000000", 32287 => x"00000000", 32288 => x"00000000",
    32289 => x"00000000", 32290 => x"00000000", 32291 => x"00000000",
    32292 => x"00000000", 32293 => x"00000000", 32294 => x"00000000",
    32295 => x"00000000", 32296 => x"00000000", 32297 => x"00000000",
    32298 => x"00000000", 32299 => x"00000000", 32300 => x"00000000",
    32301 => x"00000000", 32302 => x"00000000", 32303 => x"00000000",
    32304 => x"00000000", 32305 => x"00000000", 32306 => x"00000000",
    32307 => x"00000000", 32308 => x"00000000", 32309 => x"00000000",
    32310 => x"00000000", 32311 => x"00000000", 32312 => x"00000000",
    32313 => x"00000000", 32314 => x"00000000", 32315 => x"00000000",
    32316 => x"00000000", 32317 => x"00000000", 32318 => x"00000000",
    32319 => x"00000000", 32320 => x"00000000", 32321 => x"00000000",
    32322 => x"00000000", 32323 => x"00000000", 32324 => x"00000000",
    32325 => x"00000000", 32326 => x"00000000", 32327 => x"00000000",
    32328 => x"00000000", 32329 => x"00000000", 32330 => x"00000000",
    32331 => x"00000000", 32332 => x"00000000", 32333 => x"00000000",
    32334 => x"00000000", 32335 => x"00000000", 32336 => x"00000000",
    32337 => x"00000000", 32338 => x"00000000", 32339 => x"00000000",
    32340 => x"00000000", 32341 => x"00000000", 32342 => x"00000000",
    32343 => x"00000000", 32344 => x"00000000", 32345 => x"00000000",
    32346 => x"00000000", 32347 => x"00000000", 32348 => x"00000000",
    32349 => x"00000000", 32350 => x"00000000", 32351 => x"00000000",
    32352 => x"00000000", 32353 => x"00000000", 32354 => x"00000000",
    32355 => x"00000000", 32356 => x"00000000", 32357 => x"00000000",
    32358 => x"00000000", 32359 => x"00000000", 32360 => x"00000000",
    32361 => x"00000000", 32362 => x"00000000", 32363 => x"00000000",
    32364 => x"00000000", 32365 => x"00000000", 32366 => x"00000000",
    32367 => x"00000000", 32368 => x"00000000", 32369 => x"00000000",
    32370 => x"00000000", 32371 => x"00000000", 32372 => x"00000000",
    32373 => x"00000000", 32374 => x"00000000", 32375 => x"00000000",
    32376 => x"00000000", 32377 => x"00000000", 32378 => x"00000000",
    32379 => x"00000000", 32380 => x"00000000", 32381 => x"00000000",
    32382 => x"00000000", 32383 => x"00000000", 32384 => x"00000000",
    32385 => x"00000000", 32386 => x"00000000", 32387 => x"00000000",
    32388 => x"00000000", 32389 => x"00000000", 32390 => x"00000000",
    32391 => x"00000000", 32392 => x"00000000", 32393 => x"00000000",
    32394 => x"00000000", 32395 => x"00000000", 32396 => x"00000000",
    32397 => x"00000000", 32398 => x"00000000", 32399 => x"00000000",
    32400 => x"00000000", 32401 => x"00000000", 32402 => x"00000000",
    32403 => x"00000000", 32404 => x"00000000", 32405 => x"00000000",
    32406 => x"00000000", 32407 => x"00000000", 32408 => x"00000000",
    32409 => x"00000000", 32410 => x"00000000", 32411 => x"00000000",
    32412 => x"00000000", 32413 => x"00000000", 32414 => x"00000000",
    32415 => x"00000000", 32416 => x"00000000", 32417 => x"00000000",
    32418 => x"00000000", 32419 => x"00000000", 32420 => x"00000000",
    32421 => x"00000000", 32422 => x"00000000", 32423 => x"00000000",
    32424 => x"00000000", 32425 => x"00000000", 32426 => x"00000000",
    32427 => x"00000000", 32428 => x"00000000", 32429 => x"00000000",
    32430 => x"00000000", 32431 => x"00000000", 32432 => x"00000000",
    32433 => x"00000000", 32434 => x"00000000", 32435 => x"00000000",
    32436 => x"00000000", 32437 => x"00000000", 32438 => x"00000000",
    32439 => x"00000000", 32440 => x"00000000", 32441 => x"00000000",
    32442 => x"00000000", 32443 => x"00000000", 32444 => x"00000000",
    32445 => x"00000000", 32446 => x"00000000", 32447 => x"00000000",
    32448 => x"00000000", 32449 => x"00000000", 32450 => x"00000000",
    32451 => x"00000000", 32452 => x"00000000", 32453 => x"00000000",
    32454 => x"00000000", 32455 => x"00000000", 32456 => x"00000000",
    32457 => x"00000000", 32458 => x"00000000", 32459 => x"00000000",
    32460 => x"00000000", 32461 => x"00000000", 32462 => x"00000000",
    32463 => x"00000000", 32464 => x"00000000", 32465 => x"00000000",
    32466 => x"00000000", 32467 => x"00000000", 32468 => x"00000000",
    32469 => x"00000000", 32470 => x"00000000", 32471 => x"00000000",
    32472 => x"00000000", 32473 => x"00000000", 32474 => x"00000000",
    32475 => x"00000000", 32476 => x"00000000", 32477 => x"00000000",
    32478 => x"00000000", 32479 => x"00000000", 32480 => x"00000000",
    32481 => x"00000000", 32482 => x"00000000", 32483 => x"00000000",
    32484 => x"00000000", 32485 => x"00000000", 32486 => x"00000000",
    32487 => x"00000000", 32488 => x"00000000", 32489 => x"00000000",
    32490 => x"00000000", 32491 => x"00000000", 32492 => x"00000000",
    32493 => x"00000000", 32494 => x"00000000", 32495 => x"00000000",
    32496 => x"00000000", 32497 => x"00000000", 32498 => x"00000000",
    32499 => x"00000000", 32500 => x"00000000", 32501 => x"00000000",
    32502 => x"00000000", 32503 => x"00000000", 32504 => x"00000000",
    32505 => x"00000000", 32506 => x"00000000", 32507 => x"00000000",
    32508 => x"00000000", 32509 => x"00000000", 32510 => x"00000000",
    32511 => x"00000000", 32512 => x"00000000", 32513 => x"00000000",
    32514 => x"00000000", 32515 => x"00000000", 32516 => x"00000000",
    32517 => x"00000000", 32518 => x"00000000", 32519 => x"00000000",
    32520 => x"00000000", 32521 => x"00000000", 32522 => x"00000000",
    32523 => x"00000000", 32524 => x"00000000", 32525 => x"00000000",
    32526 => x"00000000", 32527 => x"00000000", 32528 => x"00000000",
    32529 => x"00000000", 32530 => x"00000000", 32531 => x"00000000",
    32532 => x"00000000", 32533 => x"00000000", 32534 => x"00000000",
    32535 => x"00000000", 32536 => x"00000000", 32537 => x"00000000",
    32538 => x"00000000", 32539 => x"00000000", 32540 => x"00000000",
    32541 => x"00000000", 32542 => x"00000000", 32543 => x"00000000",
    32544 => x"00000000", 32545 => x"00000000", 32546 => x"00000000",
    32547 => x"00000000", 32548 => x"00000000", 32549 => x"00000000",
    32550 => x"00000000", 32551 => x"00000000", 32552 => x"00000000",
    32553 => x"00000000", 32554 => x"00000000", 32555 => x"00000000",
    32556 => x"00000000", 32557 => x"00000000", 32558 => x"00000000",
    32559 => x"00000000", 32560 => x"00000000", 32561 => x"00000000",
    32562 => x"00000000", 32563 => x"00000000", 32564 => x"00000000",
    32565 => x"00000000", 32566 => x"00000000", 32567 => x"00000000",
    32568 => x"00000000", 32569 => x"00000000", 32570 => x"00000000",
    32571 => x"00000000", 32572 => x"00000000", 32573 => x"00000000",
    32574 => x"00000000", 32575 => x"00000000", 32576 => x"00000000",
    32577 => x"00000000", 32578 => x"00000000", 32579 => x"00000000",
    32580 => x"00000000", 32581 => x"00000000", 32582 => x"00000000",
    32583 => x"00000000", 32584 => x"00000000", 32585 => x"00000000",
    32586 => x"00000000", 32587 => x"00000000", 32588 => x"00000000",
    32589 => x"00000000", 32590 => x"00000000", 32591 => x"00000000",
    32592 => x"00000000", 32593 => x"00000000", 32594 => x"00000000",
    32595 => x"00000000", 32596 => x"00000000", 32597 => x"00000000",
    32598 => x"00000000", 32599 => x"00000000", 32600 => x"00000000",
    32601 => x"00000000", 32602 => x"00000000", 32603 => x"00000000",
    32604 => x"00000000", 32605 => x"00000000", 32606 => x"00000000",
    32607 => x"00000000", 32608 => x"00000000", 32609 => x"00000000",
    32610 => x"00000000", 32611 => x"00000000", 32612 => x"00000000",
    32613 => x"00000000", 32614 => x"00000000", 32615 => x"00000000",
    32616 => x"00000000", 32617 => x"00000000", 32618 => x"00000000",
    32619 => x"00000000", 32620 => x"00000000", 32621 => x"00000000",
    32622 => x"00000000", 32623 => x"00000000", 32624 => x"00000000",
    32625 => x"00000000", 32626 => x"00000000", 32627 => x"00000000",
    32628 => x"00000000", 32629 => x"00000000", 32630 => x"00000000",
    32631 => x"00000000", 32632 => x"00000000", 32633 => x"00000000",
    32634 => x"00000000", 32635 => x"00000000", 32636 => x"00000000",
    32637 => x"00000000", 32638 => x"00000000", 32639 => x"00000000",
    32640 => x"00000000", 32641 => x"00000000", 32642 => x"00000000",
    32643 => x"00000000", 32644 => x"00000000", 32645 => x"00000000",
    32646 => x"00000000", 32647 => x"00000000", 32648 => x"00000000",
    32649 => x"00000000", 32650 => x"00000000", 32651 => x"00000000",
    32652 => x"00000000", 32653 => x"00000000", 32654 => x"00000000",
    32655 => x"00000000", 32656 => x"00000000", 32657 => x"00000000",
    32658 => x"00000000", 32659 => x"00000000", 32660 => x"00000000",
    32661 => x"00000000", 32662 => x"00000000", 32663 => x"00000000",
    32664 => x"00000000", 32665 => x"00000000", 32666 => x"00000000",
    32667 => x"00000000", 32668 => x"00000000", 32669 => x"00000000",
    32670 => x"00000000", 32671 => x"00000000", 32672 => x"00000000",
    32673 => x"00000000", 32674 => x"00000000", 32675 => x"00000000",
    32676 => x"00000000", 32677 => x"00000000", 32678 => x"00000000",
    32679 => x"00000000", 32680 => x"00000000", 32681 => x"00000000",
    32682 => x"00000000", 32683 => x"00000000", 32684 => x"00000000",
    32685 => x"00000000", 32686 => x"00000000", 32687 => x"00000000",
    32688 => x"00000000", 32689 => x"00000000", 32690 => x"00000000",
    32691 => x"00000000", 32692 => x"00000000", 32693 => x"00000000",
    32694 => x"00000000", 32695 => x"00000000", 32696 => x"00000000",
    32697 => x"00000000", 32698 => x"00000000", 32699 => x"00000000",
    32700 => x"00000000", 32701 => x"00000000", 32702 => x"00000000",
    32703 => x"00000000", 32704 => x"00000000", 32705 => x"00000000",
    32706 => x"00000000", 32707 => x"00000000", 32708 => x"00000000",
    32709 => x"00000000", 32710 => x"00000000", 32711 => x"00000000",
    32712 => x"00000000", 32713 => x"00000000", 32714 => x"00000000",
    32715 => x"00000000", 32716 => x"00000000", 32717 => x"00000000",
    32718 => x"00000000", 32719 => x"00000000", 32720 => x"00000000",
    32721 => x"00000000", 32722 => x"00000000", 32723 => x"00000000",
    32724 => x"00000000", 32725 => x"00000000", 32726 => x"00000000",
    32727 => x"00000000", 32728 => x"00000000", 32729 => x"00000000",
    32730 => x"00000000", 32731 => x"00000000", 32732 => x"00000000",
    32733 => x"00000000", 32734 => x"00000000", 32735 => x"00000000",
    32736 => x"00000000", 32737 => x"00000000", 32738 => x"00000000",
    32739 => x"00000000", 32740 => x"00000000", 32741 => x"00000000",
    32742 => x"00000000", 32743 => x"00000000", 32744 => x"00000000",
    32745 => x"00000000", 32746 => x"00000000", 32747 => x"00000000",
    32748 => x"00000000", 32749 => x"00000000", 32750 => x"00000000",
    32751 => x"00000000", 32752 => x"00000000", 32753 => x"00000000",
    32754 => x"00000000", 32755 => x"00000000", 32756 => x"00000000",
    32757 => x"00000000", 32758 => x"00000000", 32759 => x"00000000",
    32760 => x"00000000", 32761 => x"00000000", 32762 => x"00000000",
    32763 => x"00000000", 32764 => x"00000000", 32765 => x"00000000",
    32766 => x"00000000", 32767 => x"00000000");
end wrc_bin_pkg;

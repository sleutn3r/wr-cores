// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Shs5826zkrmCRZnjjbJKw+xc3r2c94GdTDYwJD1tIc/SYjvnNcesn5YT9AMbwhVu
QzgyOV/9nge2DLajat8N2gdgrXenizoX3WxnGVDVW0ZvCWqPD8XtmwSFcgvpqp4F
HtQxzctDz11GU2LmqMNij4TCjqx/ouJYRm76gvwXVnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 18016)
3FzOS2yEGOb5Ccqtg2UnlSaLEuVrelietpmwiiT1d+Fvt6ycVIZOdQHqoBXzsHIn
uTJBSYleIT/Wajd36f+XDrL3TKUMr5WUZ+v3FoOtJCpN02C1CUevBvhbb0UpDg7N
zAGVq+MzB/kgE1uIgSURk1nJwLHo8LgRf1c3W+Tcxmm8e0qaMRucp8ZEKu6UNMAR
TUYbZk978GFVN7MYYtT7uFALbyC6FSiulRR5JGJdBcDbTsBRMxPrE6ZgamuFGNyH
ihBNThNyqhC+hIcszvn5JbvMIkf8JDK+BD7OClf8lzodzgRtlAEHqBc/Vf0ekn9Z
GwvVnCIA+VGKCnnCFiwhbMB/wGmiZ11CVdqPuiA00txU6+r1vdc4PW3e3qPVmREa
rLsCm2NY+v8n9MCaK+L4pyb/7TkMsrZVJzF2+Q4GrOgx0PvNslKLTrs+6YjSOtB2
6U2Mj1PoBoxjwAV24poXv4bGJRQVZ027Jm5EWB0sh+7iqXN9jqAW6vVcfbigWO5g
O5DRIIgfHla0z4GiIy2ltL3SzhsaxEpNYjV/heVtQqhro3vmGbgz/yIL2XSuCe6E
ZnRtiGgDsRzsXcnkxYRdwdUAflHBbhHzjRRqmxlOK9Kn+3uSiCa4M4x4jcvSpFNY
DaYnqvMR8cnl7qHn8rX1UKZQXB+Zl5BuqN4RvDILBb12hn85vRHBxQ2XTOpMpE8n
AC9qF6LdJZ0R2BIzYjK5czmm1FcXDbLe6ZQ60VNO9TaaIuL/2umq/xnepCL4eNRK
YgUtjpfymMyzLsPyb47MhqMFcrO1ytJOptdBT0RSMz1YToXJLp1fc7C+4y0DbASc
1l70s/ux+MuAXgkT3KUnVAjwezEm4+D7h+pPJz9ixOD+m2nSae7HZhf6EXxuUKWs
xMFT1Y2g36x5ZKs5TDxRxAQBVYSdYxkD8HKqU1NZeanS7INw0sdpwa4kKjJ2IuU+
7JSI+Yi3nH18UIUyfqYPK/nI0KBYxIgaJBppW7kUf1h++oTkjnVHGG8JaK93i0+W
cgVUmZ79WfBGnJfGRSV6DsOnum8qehgw7EWI4049tcIdLI4SQoFmdqp41a7oviNa
Yy1LI6GRUSVUVBFHSNjFhGi3phC0sWtrtwqxpvIieiS9RXTK171ndRySTuzuSAYy
r+68AfAs/6HK+aR1Jm7GAIap7wBLvmym2ZC6vxNAGKiQonjlvNiVLXZSKjrPUDXr
bdPQv4IX06AZeRGdH1AYrCfte+DT5aHX/DtCsg56iz7RuxArQdjdSHLt/HcMDbKG
CQq5fzdZsDTni0yvhN43dI+gFHqxwsOnF19BFBSnKxtXnGVWJJLGBlTBI7/Gbyrm
dpf1unxapk6MZFn7gg+OKxeXVl/zHz75/UKEuf3ZPUJYSCKrHohV7EBz4JvZaGaZ
YcUBh6XNNMwKFJqJo8nBggQbSk2ENDt9+xLafnJ60JahrvNq3eLM+rjMDdIIpyZx
w78rqanLnZG/90XIOEGTR/5DVo6mPAmMTcmmxmhDMqYd8MlQOr/G+4w2e2FXChTu
++DHY2YsCzcp9W0AuogjnmSqZzGb7ExyM1lE7qpaPpBGYp7FGNRZAyjEcmIMt0H9
uKOwdJzauucczHY1DeXKZ/z2wSN3F1YJaJQf9GmE/FoEgVV+0yITbmny1JgiL65J
30E8653UhZdEzPULloA1iyRjaMTPtyRckhB/dqAW6Qfhxus+Itz5xkoj8NGPpYaH
V2O0sYvUBUM9sGaNOBSaMW5btvzN7dr3G2jVF4SXgAx8o+C2ayDkLA0oOdcJqWZx
+bosur+v4lljDdxWyMt2jaV8NKImA4BktkCaJTTFRuJdyPfPHSOKi7YMqxC9d6Oc
9+RzGCS5nxydpNQOk0dYrImpOWFE1Ek/NQyXP81G5t636nNdddjYKGipqf78rttd
R5k76AKPAEV2W/TGQf6jIkGSQRiTZJGbmVuR+56y3sEP8wPG8kJsHityHriOCtx9
pDOkeui6P7aQ18JkSi9SANWwYzQMAiMyy8YBLQ37AKTGSZQTFZ27/KmZqBbEavJE
2eV+7ERbu434nvzwnnp8hFVpIy21IX9u0IYYicwiH/1YpWvavTflzzNO42WDfsP6
xMVRiQOT7ehXKzdyubcrzMQxUHTVN5qpsxxxhKSwAVYDy9IcjUnAfanguvT9gJxj
gKpCyAc91bNK7hjY4VSLuN23aBtYZkyitLYrrflMZtqWk938wIZ+Gaue7Rdch4tq
vL/c+aD7f2+enwbrVb5QTo73LWUAuwjLs+5owTokZsW7mdqwK087x9VnV/onkqQc
dkO3eR7Iwjokm7VSVwF4rGxdf9iiTsXQNpjg4bKa2Q08+rVDcZUfU6o8qSL4vPms
DVkeWxdE8ucFXHH/ZqYlWRlnwBK9i8xS4p2EYpXp8vaO0xcoFpYK6nrZ0Nl6ckw7
HZEpWarMkip/0+QH2KBGowupavTkUj4YbSYUZqDTN8pQU606Ym/rjPNGXO3mk+Vo
nnWhZjxYWTCkmGVUwv1mAu80Q4EYvs2hviS3Q8UK21QO3Dj9ySNt01lUcsducBAl
p8m3DxFkPevqJ6qidyO9oslJWiO/Yt8QpX4sSLP7tS3L4K7wPdaWygiM50pdWjmv
RyBpZDJeUkMRjNcCGYRqlLo4DQTbypJxe5CBxo/N7twCOAXIi9NZtYKFZ8Xvmrnf
EqAV/Asxo1JvCtnEME3I1aAkA6zfwMV7LaFyB13Y/dU36uiv9W7zo+5iTd1Y0o17
tE4RNX8j9ikGISZhq037fbd92EBJR3VhjESt8y+NoBifqrvLBqoi8IZxOmK2CSBZ
Sc5BX7KcyuWU0J6A8GmbnukkaLRO92Y3HVrkQPfU3DtQp596J/ZDssSGUDgB6iY6
vD8QRlOWee1E4xIUXwc7NsWpB7xTGoGw5W2opBYir8e9BVjUxAVFvxm6mOVWp6u5
xXSOPEUw35ZYQNBjI2EmNvE1r9JupY1PPf3m0Recp0jg62dRlFKMBkOrmZUCyHTW
Zlzb4TFl7UugEwUnkNYGaDITxoh+Ho30cz9FzfvZFqthhyVLYzc/6yheC3m9AvGF
53MUNCStT7E7HefsnlZM+Y3XeLPUx0FjhHZY0NIgqOCSl75wtZgVe4Ob89kOBNEP
L5oZxJCiAjyNrS4aGg+1hWnawGNYK0Btbc9iGqIgUfN+8TjW43aXLHwzcHzBhVPR
RiLYk2O2uy1OxQmbMOGBKzVncP65OUrau+gy5hu/wjsA1mlEYwGodLt/z6JlHdMM
7LyyDeRkEodPMlJd3slJbdDqpYZyf16EBbV/kXj4DvL1FiuqB7lFHAl1TWppWN5E
SuYRP3nAA3mpzCXBlYc48Zu/Y/bQnPc+qsYDDxtaxupTxxezvhMk52qTnfuS2A+9
NbGVmBC5wFNIODFeUbpl3JEzbvyrZrDQbsGaSCnl9LgkdSCQ9gHBq6rGO4I5Xm+v
kLYJmrw3oZZvBfyBG3XM+csLwA0euoiCaHMB22+9/y7xblwMQUAQIdjk5Wc8GcwF
Y5h8W6DzXdLtiYQ7ON8FA88iMbemf7Cu9IfD8Sjpiv9oJfo0DCOOD5P7Y1XqthD6
4eUaD/2V6EjQb2wHyyS+dbCB340vn96Qv3t85A0NSfZavcl93oXCo09lhIjXMfDl
4Q5rG7vo076SmVtu1vJ/MaltABRdeG52VMkgycxKxHzXKNtI7+HE+9aGlCxcg+Ls
xAeRE1J+4QOuR9x9kL0W5PXwhJHBDnWIk8azg+hq4HvL3sbnCaIHfHp6J+8G3FKU
V63Je+ZcIQXS9ZFFg9dJvlrBfaCUL3sR0p6FOUI553zibXJk0BfnOr2O35+SIbX1
AMSadJfKuO7pQw4O7hZQOSMQK9Sylcn1rYlx16Nn3FYDrkgY+Yg437O5Pv1QkUO9
eSRBHIKQDZVVrbwMHLplV1VFecXhkqrVZ2CNsGSOoFHDmC61X05epqQG9bW9hFU2
hKsESg7pjioXVOgbNFT1m9BFNVBBw75VEFTYNgDP2h+IG+rLy8lDaAp3FFaDeOfn
qtJqnLkCRHMjJKMePn/gluSosvl8JH0DIujrcRkt2fl29tDOLSEyP9dcqWuJ/90U
lbtbfVtJnebyh4OK+EgwMt+DT+eU9u9gF7rfJc7GWpMOeehNn5GvHSRH97oqvt3I
9EdR6lVXZ917TEqUff+KnQ2XjfEw7k2JBbuN2DXoXzAQD8/IyvjhHu6g4ckcx5Vb
Zf+8QjcodCaFuQisQX2ViuKSBynRWOKxF3qELaLky05I56EhSkvVYndYb36CsPab
GZT7EvxJ5sMYeSgs2EL1Dcz6MFSXpvlSnLx6aKSrzzLMkF42NluEbKwRz8EOypVg
vJJ6wInf3E5rTj//wO+8TcyxGblFp85jR8YA15NLa8Z17DJ3pqYIMTCGugdAsJMu
vF/Q6gudHKt5Kr2lIEa5xuqEiTFEXB6aflkYHjGkrQ6fJ0U2TiiATU9YNQ+pwZe8
LlDhNvnm/3NYvxy+kFxsXi3r2NW9Vdzb2NzQbJjdod6FPXyJA6ZCFI9LhK5v5tsO
OFj6/3X4rtQ4VXpTvPbJw16/QPaBy/G7i3PzQnMw+kIfKPx6EjffxwK32gkR+ab7
ffgtHz5wFbcLMJQ4TvgiT4vCS1aehFCyFnaHeOfuxZ/X1xcpZE9F6//yMns6hq3u
zPSLtYnYmJJ6gfNaLiNYLggx+B0jaIlgmCdT8gXO4viS3ey2+uFT9KaQMrViPAX3
Aoae+yDoMNFue/HaAgj0quI8MNqXn29GdC0B00a3TWp9MeY2/wzSLGC5sKFHV5iS
1toYXLmzDo7t2V75T2okTf+WMXcx2doZ/bDNJ/G7L7QL6iVmHvi3TNxHIiTnoxE8
ROJyyhKbUK+r2T5bJHZ6P1AdsoJyEtJFReEah+BD2xygpMcNCqQNrUn5wn9F4PVP
IjKROBVYzy/IfPskswgR9eSEQR7XksU1JAlzHU/e9OPgGCQUaWw4Dys9prANiWQL
xXr/1RXci3KJNiyICrmO2bpP13/xdWYNOjzqT43LaumSjKp1Hyxz/T7GjjA+Z1Nc
Bfjzx4vZuc9hodBH9Fr588bzo5zOmjKku3bijynnHdhdG6fwgYL83tyHT/W7WYZV
20YjQwfRRQMA9Hs4TA4KwaHNRhY78C+7QhwjBe2fqXUouo/meUUh8DdjUKLrXGE4
uRkblUIqR8+7VrZ7lkr/7bCQrAnRdHocvZW413TTuMu1SlzQxGbGAWi6cdi/HXoA
Wv2c41lpikDQL5t8XlU0wVIoUZDuskwpjdj8O6yFrMjBrjyO9vsdfTpXZ4ffY0rv
ogjZc1v24A/67WCIRtfzbOxDx7dHj643YYM56a3N4k+VhnQmap4Yht417d2KDIVz
tBNscltHq88BC6vwtMM+5wgDejruUoLzs7QHYWLXOt7pIYLbRL4Xu7ovRSdx698U
C47dRQt4Gmuy5KlViTi5zQqRCZ84sCgKKvoUtRBBxSf6+KDbqCfXfIasqQbJtpvs
wG3pmgMaa9ODW/LSz3sRSRe9RRqSnfN9Ze8ILd+hOwYtwuH0q0LWCYCCTWm1fgUv
uAosH/kWmYmuWJ9afwGsnkSZx2rBTzK96kS5UOFqVjUE/05SeBU05/OCEFllN6Kn
ZOkOep2VNUfMnWIutWzsDBA4IXtNrjMm1GAoba4gZC5rr0sxmk7SuLUarKTuBolt
ulbNXM06Qsdt6NOJ7lry8uQfDnoKBdmOnYeOabOvUVtmx/bbkWc8xybtlgkdjbFm
IWizzJJNiY4vcPwDVFdbzLhsa9+A110XflZrJ4aNvk94mza4sAM5vB/hSNPZH201
RXi4NgtGxyopPr2FhO0z7r3P/wQcE5i6hyxW+CCFZ3a1uY7hahcnTXJSWQgUTlxs
Pm3e11FgSWDINt3+HyFpBuKgM9mmMv8xF8bVFtg8xjPni+wUmLR5zVUED/D3p3BW
WjgChUeVPCjSJzLyVIX7IUk/LQU25WC2KpgCQNGhVCc9IQyoHQ7ySgLZZK4Z+uIK
RddUKro7QPpchISSB8RIClyS12KbbgqedH7E+Yl8GcCD0upt0bRNalTiyTFnkdjl
nP8FfSTBJ0xWfQu3S2Qt3aJV38Y1Z+4eZVd6XFkYKIAQrAhiKwhPfSusMB4w4k2Y
TA0PJJFl2Z18c6b02mZBFLC/y78r43wRavETKqjtL4zFvr/BIVwxVxgJjrTF6ED3
Q7txqPPaBzHwSwcD2ISdx4KJWsGGqnqwnB12Fap/8N+IloWSu9c4VyBNK3/mYm4T
IPKc18gx7w3QhXklIPKv7IysDyXk/Rr5oyGpnSZaHyMZX8oOI47e6mzbzypUxlk6
jOJjTtxdjMjwnUGKvbhLi0q7wigTxfnOWATcd+lim6RpoAa4RuPZFeZd6L1onXO3
B+klbiMq40pB6NHATEC4+gyQhtVspTBTYnSMUouPKdXdiyr2k8WwuJ16EQi0IuRx
yNv6zfPyzH2szVvo4OE9Ejk1EeH4bKFW4alOlxU4X0mKA//r9VCKUGUkA0NG/U6E
pokjCT5OKRAZYz9Jk7eHNbKXAcC+83FFIpVHR9UflSCq/2l/54zcv+VMbD0SGqql
pNpoHfjqpfKostgJmSkKB5O16ti7dvANTJWrTYft7fMqUiuJyG4cK/DjuwPI7o5S
3XhBOQm3yaTkhmYwCUcroEET1Bnd0Yo3UrOo7pijnoJVFZzTf/9yF5VYJPGls16m
g8/DKF/WxxkU/UrvJhAr2umNxoOIfm9/SNdgIxVlPx9aROSS3kCFiw6Ss39a215f
yA0mJOeSBVGnNCraiUGxW0HttqZGHQNkVLYqzdNeXK74lx01Sp6b8x4FEKLdW4pn
DCOMBr3M5q4zxCZ0GqgKzeM2gDMtZwo4hWxmjDFQALdfTnWpSty/s7br/oEV1qbh
Qu0UdOv142drCL40PxqG7xPEa4dJcJfMjnyNJO+2qNtJoGViPwPkPcn2nGEfNSBf
OerpDAAKS+lr850AS+PugSvO73kGdhYjT898Dxv2VtKBXPAY6of0Oc8rU82m6WHQ
q8IanT+3AEougtQptiOv9osyuL78IYzlwby8mHrajUlwM0AdM0oAbl2JOXmo3Dyx
6Qc5SyOWFJ9xA2Ud9frlSKA3FFRkRwG8wxXP+eyxRNGuyfoLOMCMEIk0h/u10s6W
CKEn5SllPQ2ocxGMiTSMMR0O3FwAw4TnUXAO4ogHJbxxdZlogzhzRwGnjxJfYMrs
3wuGYmI9PpXqAB5xcWY50uibbheYf/lclU45HBuTiEFj8UUr7AjKngacw2BtCizQ
COK7wOZLqaLSLXyIxnlgz/ZPt0WzxOXuJi8fVjlcZnu7Uh4lnr5CKAg/p3Qyt3KL
7LUQ/mWwhXWXrIXQmQnm87cXoh5YL96eKzIZy40+CXGb8AtJGxdBJsZwtu0WPmDm
XTx15C9S43RObmeyBA/sGu82I4teCZ+g2QjzO90sK3z6pc/8Ln4rnv2UmIm4C/kH
4Yf7DeNy5sXbmCEa7ZfwMg+2uyLVwMu7KwlqWuyDU9tWRthQzCKJl7djQ3Prhv/3
acDgJdOI7x89aR0IkM/E0LG+mOYehQbxGqqpXnp+xZX1C1CAB+3J7FtH4JhFT8Mk
0FEibAeo0UZB/O2uIkO1ubdS1vrkrKOnnoSgvXIGHeOUuuDGu+rG7gQCSenS4dnF
cxTjFXZT1FfdSZaV/nhNDiY2RdNwNZWGYT8oDVcL2d4ApxOYErZiSvAsVEcSFh3y
bwaW3ur9bNJ5wTttR/UjJ3EyJV8uyQwKLtAcCr0ynKkgr4F/T4ddDnRZeinZOIMT
jK3gGdMXSmqWa4DHkzB7pZY/wdX7J+snU4jIdwSniaDWuvR7lbpqhDG+OpHJZG1m
fZH0ehJ03hgROQSd1jR2F3C9rWmdVVLGgVD8FV9gReIiMeEbGXope2TkDPhaQlGk
w5gW0kkY8ogVUgmIh2gHXGrA4wQ7wwP8rujQj20tIxM/lqix3LWQw9gqZ/Lh+0jQ
t+eoy0/jnigwn+oavu0c6+XGLA7XGTK1Pbj9GhxCqysfu/VmWvamuVPIkqPAJVjz
namAk6zAkIwMWm03BfV8Y7Lu84uPEePEZozjCNh4IOOKzC4xyV4u5EEUGaa/Jpw7
1mdXZLWMgvC33sZn7K3NoblIcOITqnRWyg6NiJR4I0pghmVS3Q3a7ZH2hlQgXExz
pxmzMobzzoSh9P9HKzQ/IJbq6TN+psKiuWnDRqLvyWgLpijBHDisNiwRk887RsQl
aPtxYgamQ3LRBj416xdtuFH6KDCXvihRvXnolfdQheaH6J7+GQnZ6B14kpaWif9g
3x++SnQ30isTCpO1ANXjOyLPyX+eB09SdS96V1PzSnuxQ6G8rmZJMH6XnONNI89k
2JjJy/9PUVgFo8FkpODGoHanS89eUty1sbBnFnTOu1PLI6EqeE8GVDMaUvIgJfFb
+sMiQzBLENx2KuJVhKC3eNYBcrPhOAKMmhUSdHQXNN9BPLQovSROj3dStZ4kWPmT
KoBbZhSo9vxGkNCjQ7pRZgBsgZyt7YfkbPPAZAh4SGxGekCOmQGP682iWSaZWBJu
f3BKmYA/wm9G1XrfF3+sUcCkYoJ9ar/WRVDeukAvlxnyshRux/r3mB238j8839oE
NmXLOzkBDk5zooQi3xftPpAWP14fElXbL1DMWKL31NF+JC9primz3iFMMA3NmSra
iCvNAZa4YAkNQsyvUImKqPv2WpE54nQvK5If5W7kmALKGsgzrUH2JY/AiiCG9lcn
az02HZow+KXuvqAtVS9+t+KE0E+ignmkdJQwVP5jKEYeDSkVFlzMMZM1/5wn/aEg
WF/hdVbhreodZAKQPHo+CyOh/50jnc3DRDkblyFl/vjmwMhr5c81f2VW5omstLhZ
YlOelqkuPZZulpSZchxMg7GihRkZwai9Silk8gHGDk4K3EDq4HoysmUMsHiQqV8G
1dJBFZYW8JtPxv2JIGr1Nosz78iKQECGVGOKLZwOMFT174K3bOU/ew1pKi7Y3KE8
BSMfLNErms57ecjoYDy/wiql/Hg0tNoR46XaHaL09YTbsrkXdj1mrqsS60pPsjxu
O6hNgVqPJxz1+BCKi/QLL1Y1DcLPaIid1G0d6hO8Gj6q2yjyV3HMhiQPxkb9tCF7
RJcw6QEuGIyAry2Z6IPTDlQeaTo5llVlTM9lXttNxqCqRibTEbBogElrYx4/IJTN
b9/MybEfhLe/14zOlz30WHN0Jh/a806/bMF9aNsOZUxs5ZSZ4cemccVppTmGR7kK
xH5LstZgJci80l3A8A3JyDIDxxZqaQnCJAVbOUYHmiqxtczELF0CWxOZqxH7Uens
20UflD+gxD/BM/yMgexuObz2oNWZM9ZWhEqAPlidGI0rhSRGDssVflmA2IINI/RV
mDJeWs5XFdcKyPzpiy8nsyxsCqufJleRZFULArVJbgTJ2ra1avLW3XDcwkcyQDC5
oDBaNdpBoBs9D7iJDkHk0VkJuOMFqHZc0ph4auVcvL41fnGtkqApk7b/1e5NHSwF
NmWt9TNfXU33IYgFLAeEynvkNNzYdRWiTUFuaC5baPCNMLGxxf4IazIupbsXXzJr
JDds2LdXFMbdQI9jN5QXXG4As6D+XsTL/e7nHmBjiEc0CwQEQzL0IeNX2sRnAlP4
+9Gp9Dkd9obS51i0GOmkBTo36jA0mihaDtt5N7NPjoOiqphPoZ9eRRaa9cMRnbtb
oJANVzKrcm4jtxRT/bg80oc4Ujklk2P2oWoKoDSbguvtK2Je6vtm0eUQZxyRSHib
XMy4riw+K4bob/N5jmSv7k2ucUqECNb8c7VTQomW0LRT0J6MY+gSKCHjjZXQ0cwh
n9npMm+iLTQScSuUWRIDmKniGi995GxGdHoNqZPlBoK2u3y5j/kU8KqvgQ9A26iJ
UFPA7NTyRGLTK+LXzLcwrVgcJxyAIXTAwWVrYNWEKyDTn5b5IwN1DjLMLpt4TjAP
pVdDU+gjeahYa7EwZZt9iwo0IN5Ts8hc0qxLfDesy+NxyeYJJJmVug6r7XlGN/s4
bO++htnsKw1uzutv0cVbi7BK38eurRxClML2Ig5ac8EiQv7PCwNQLd5EzN+e5Ftq
erEW/SbXLeGVrfJ2bafUoIj9umhKFTebZ2kTtZ8ygK/OqK41b8r3N/pAV6mhZt7E
p5IaOGNufhBiBGf6beWvKL7CT+qiwm7C2Wvxu8FNlIjv/da7xjTCLCJ7W3Zpkq6p
m61+gS6cw3lOBKJqjOcxNbKpyQ5tqw7YZiA8+f+HwvALTqfA8ytFU2v2FmfeZgYx
eT4BiCmjN7LwIsJ6YdLrbghppKcfZY5QKzInO8NUjQbZgNJrSVBS7nTiPBBS4IAD
0iZCngoopym20c0+WQ9QJgXU8rlTc/uF1vHqtw7M6+Fe+/OoynN6CNRaoy3oQvWX
CTMx1f+CkHCKaP/heg4J/px32HmA4/P2NnlTJtfdkLnjWE0OV+GibwYjwk5giPDz
bEh7Mv0mBhzS+O2sGkAoVXs2ZVAkZfl7r0PbKxISK47Am8ZXhmVnQEkab+hcnyGz
Xot9CSHS7xU+IENniCTxya3D/fBkjc3f9qicMdSUOG6g8R3To3p0J2m6VgUyn609
sgzRAJX2mqj/5BMe7nSRWuqW2Tl1W3VeyT5R02UNhNaW9bYX1cZyEjZqwPQ2L7+0
/4vSxaPJZWpZx5QEQzBBHPbbgXGwF9MAs+d+N4Hk23DulfBMk8yUrJXiGTh1lVp8
Qcwqhwpe/q5K7Zear+/TqVRqK57aQ1bM+MrdKj6cZdY/Za4xreziitJZiCaczP70
xFARyKoHZgX3UkOVPMte5R4Kc1Jhhuier7gqoHVv3Q9XPdvHe/pK3qyRREvmn4sE
TGgy2rk4iQi+lDnQGmTjhgahuVr34jOsVZrLuNn8jsSgatOnTsXqcqJpTSdKnNCq
K7ou1cK6iwv8WeumXR2D43eeNfxcP8NjlFy9A3hfjnYz1xru8rw6rJMDgivPabex
EfzRuqIkyfE4QtOnYVzJ0aXbsvhvJbScO83wtxKlPhvZ1IYaCEgvF9ZUUGHRTkCH
WT7wcQgMeGeXwaneaEU+JdyoqMliEgfvK3s1XAK/GqCtBU+EOB0Xdjo0F9NND02n
lsbS78jO+MYdJX6kdyUO5EA9Umj9pHohm0Zkj+HRymIBuhDHlcZCa6hqFbwrFDa4
Nfw1F8hDQAfeDzAN+5O8Sr2vcsMhqBY8Ed4IPRC5fcxi63JAhKztHnh7QNWf6/E1
3qRaOsUIa5jddF3Tfm0aZ3+VgvxllyKrpOZvASK998FBKXvxR9rkQUy1xHLxe6GG
0WfF9fvu6mHEI6/eMJlSlJaFMIki31EQ1XEKvH886yDOxIXkSDaTOzhTuob8fQ+N
UBUm2ICJ4VYE5ZU08i2K9kDoPs8IvtWXoi8wL2BNw9eqJnOe25XaixRJiQiVYbQY
O7WdTt5ai0CbdB//1oinT4Ru2Sc/5VIPh0qfhb6cmfm7tvOEwHuxBoWOL0vL+ZXL
Hus5VMmDpj1UsKM1/qhkXJS7YUAv70/6Xyidroxd6OiySIT6JfFzOMLXoKUyZUoA
NKa3fVDFLupTtpZemzRdnmxugXWISn3t7x0QItej6GVS2YpofAEmhpBG6vPQVJ8b
bXVeVqOGG4No2+lHzO2ibybqmLpyrcBOuG65zBC458TuKcmlcwTgAgZU3HxJSeG3
fZP/wLRE9bceKx5yKIFgewamVlxB11C7mqFl4NmZalMuCSo1t9jok0NKFyUeuQtT
g8umuZ5VkaSaDvGZ97IQS4cde2Ob56HB8IyeiT++GWWPAuEBKX7wLu6GU4nvID5p
B8b4Q1WegC7c2K2JYfdP6zpOe5F+CGhcr8EZEqnEP6B4Bsm+GRlazd+XnBN3OPg2
yysfVoNNhYfyAhptohM/TOEN/aEMze/wfhtvBnUxiQ2xzZTi7G7rQ6YXIGl4Jx0W
tYylDdGJgZ6umtRrd0TpLtbR+JPKyYxInVng2eDhJ0n6pHOLusfnGUvrcbVAcok+
OP4J/CGkex7cCzDk8EaGiSiJyB4NUc5i55v8VoLs6hUQ2vheT4LUJ7VjhtZVmA8G
mmlXLVK6a8Y4+gHZ7pH7UpmaoTM7WEnHLqEjpZS9wzGBA7yoUdzawJ0pZEdRDY6K
fr+n3OAhaHE/BUQtuVn9/IIVzJ8g8whr9wBJtZHab1yUWPLufM96bBWuAfn52BOr
WSCbQfb2HYPy4FtAlNrudQxGWGyKXqJOIlOXF+7jNWkZjsC9H1GqZoinBb+Ruw2f
sH7ynrF2/rniwck+IgPe3lNQaEE7VVDo6HJrkzeTIE4rTsjle38wAUsBRAfbsGgc
nlDYU6+QcPUVhJGBcBTDJIcmvi989SOy+wQa4UrLyCKgVc4TD3TpRHD30IFIEvSj
eAXF9qh/w9WdVXF8sqTjYQyfxbo15uZv7jXK2n2JQZ0yrTDEELiGL3BZbLoWGnhd
QCmZrr0kl8xp1X8no/2ijngr80ssR8RHGTvT2D+MMNNx7t5R7d+PrzsVfRHs86qL
zl2d7pB8Uh+3mJ5dUhf/+X/SAtccd7sxh2sv/ETG9/FzFzQEvRCLlDgVFBPS7KLW
Tim8O6XAYlTrxKIsyKBMlzgAuwloOxoJ6PaZ/JIcjzE0/Dpm+rCU85C/rYHiuR/Q
MspsDTD1G8LuQkYgnJH6lLjcS9JFXzvDqjr5O73Nayw51lX+0MlIGND77RSSR09y
SSJieMP8mTWsTvt/6tT5lEPUiUuriF42bt06TPtCbPWPmyLYmZ/5wxa9JTwT2IJK
M0PJjIrdMV1SQpzLuyRnEAAsBHqP0pq6TvBArWx0bQKjpFGE8tqggRKklBLtH+VC
LVxQzsk/31t/ohypJirI7SlSzMLsIPlIKpIUR06H5xqOwfU7gg2vhJTMNkAVYamv
3QXrPiQ1FrcsGkviE68+3rkrtFgPgMvI5GF6MOYfrH9HXB5X3ZhFrSs4d+Bk3+lS
sqhb79psV0PlDEHteZVOSiYxtGwYK8AHILW26m9B8eedJKCHNcwMG5Zd/hivSVq5
iBAthji+G4VZkPuHTT5THh7PbZkk/E7mQ+RsfKP2K0tKSN5pUzq1DAISrR5comX3
ehsSBJIR/8i3TqDD5GB7nF3qZT18U2v7To7Xnwju/otDMjD/7S8g+8izVdLGJszB
GMJzCxW2OfXxS8ZuFYKppGlbqrJQXerIIbbkcj1v8fLBWu3jRFQ2Bl6PTnFo7CuZ
+jHwaVJVi7c/PyStBB1CJi2tMUB/iyMkKhMGlkplv0w04jC1HTPzfRCi0ZUQRhfo
w5/DQq9bTl2lyzGYgdTt8SGs3lvCiQRLVzavUMWa4eAAH+R570AFw6OPCF3CBtVV
PeNMJ5XHwyQOu3GpRmLd8tT3YG6POIqNFec531TJFOpj1mTm4XiO4mlUTsndPCLq
ZCCdng7YJ8K82ZMU9WsBxK3D+UFg/mpod/ywH4+8wG0yfkZEk+weMriE/0aQ0cZl
tjf6pX1+YJlMcMh5BnjUyRZYRb6QhSKXyE58A38b5dvxz1eXYICtneCSmKzuKb5j
F3LoGZM30kHxGs3Gr/oyP0fiodrL05rJNEQNsav3cSGIXRNNJujPsgsNGs6t4toU
nNPjWW1HNx8UOv0CX+eAuqXNGvUSRAXJkkh8d6pkKBAz94JsHm0Nj5wDW4epAIYV
J5zLagf7y9hP/8oGF94LrxuHX+HKqxhOPMA8qQItRt9QDOwFFSLe+8aw0MLa4frX
yWCeJlJ9KW+JHK+JzpiXZYgCvVnaXurWgunF96SXjRNYlKyZySqPe9wJuc+WS6Fp
ttoUkdpsOFVQwwFeETJt7U7jeoVGfOlhdPemrRjgIdzVLQQXiOVPWC2vkjQgzr9R
++pJ1+b4DS3YTFE2KsLLDl+z0HFwNPps6SaiS5wfuez6gmN+5J3/NGqqVfNyaUNi
abZC9CKXP88HtCyNCwoJ3UJgOqZy6qYUXcIh1r+K46mLmgeazTqZrpbtiHOfJjWU
wqlVBmEX6p99yBpXbvNOKHuiwL8A+Tzu+iBskuM6wq7ZnpVilc77u8D2o+AxNngd
mkk/G/1/+TJMHTsSBIzchWcGOpyv4xIfsSPyDFBTFlvLwvjeZAd2lXvYK01T2Lr5
Y4isbt4gkexiUaOFr4QYpCLY69wHs+wuwVsEpLmyCXSEZiBtrNbKwuoBg/xmetvi
fkckkNqS2go1E+h+9Sco137Tl2amk8hBkeFOv/SiFwazaf+2e871VOSWhMfDgrU/
XabdtMBtwamWETnuJhsvei/bz3yUkH3jjir/BUTeox7EtkfZy/00dwQgiAXl92ax
E4MoIq0W3dKOlZSIeNhl0qcR3EBkrIqn4VCdDhHRSmUxpEou39tscFctYFfBfnEo
y3ytSCfCY6rDffaA3O+aDhvxDbHeJE4pFWlBbm208zCjI3yC//ZmB9bDtcKmc9i+
yDOHoF8+zbPUfb+ya0nTOdwVaNBITdWNim70AtN00k0TB8uUxzuT3xBKvSyTDqg1
/4FWOuQSN19NFSaBD7gMzuLTbVryiDbxx3j4nd/Nc4SbSLrWXbhWIof/pwszMyNX
wtv2D4JLzvLBRHf/JTNgq2sNukkAIWAaKM0Y7ILipbi3Y4+I8Zk9BigFtq1XvgQ6
xU0bh7G73xKf+eE9ksM5e5/STYNl4W8aWBlpBZ8r+Qzusi5pPirRQO/MLEa9SaTc
FpZshayp0aX4bemnIrMeE1F+HcnC6L9/qQxeCf921nTcuPn2kSLi30jpFOtWNRuj
PfVoS6t7D4uvHAoAPT3obKpVjTVUwQAh3HmEC7si7QD9xHeEWZgLtOl2E3HHwIni
YyGg4RDWWVYl29wl1cFKybOdOAfusBdxQo+q5WrL1k8rdGkVpjACdXZ/UJ8FL9R4
uRDaNiNuBhpHqVK+gvntZljhaWJzPDqxIxsj8XTybndpELjLoZ07G8xV52NBRCHO
mEewSjQ5nsuDiuUJYWaobkIhNNiqIbLvWGIfrp8J+SwSqB9FKLvkjDoX2Pvdg0W+
dtcwnj1Jb7zNm88NaQIneIBucPSK6GVVlVbUINmvVuNPB5XjFCDzbUk2f3OET/t1
popzr95tucv8qMQAfIq5DXfcS5Xz/7GScPM5tg9J0Cr1VfQiui2w8cDNDJIPIK36
EopXDgMREz1lL78sVXzqBObSiOwAEMB/HLJmv1sgsORUrdKx68TK9nMnXN2VXKH0
FowCBniZadW7mJs1g78rQNb0Zl6/NpbyNGCNcYSsnmVjnCbrm5jIH/BAsIsUUQad
XuI0vOC/AGEiuXUjsCx3BYrgw1nZi2gXhjtpCQijHr9TeWJFSfpfLZtdZL8DkwKq
JaUvPhWgSrAcu8n9GaKJ1k7KgCyOBMLvqxqe3aQ0GllFIGj1rknkNb7/p4AlBG+H
sCW6agIRGHL6IvoHetrdn8cw1jc4ao9BRmsVaxBGG/enEZa/IEStmrH2asHR5B14
bE2QoyW/6hO/y/mcXRVNafF8Z7PqpSkVaDL9igoqaPAMZLvWnR6YvDDNwy50y1mu
PhTBBHyunzivswDorYcz+21J7O7HG2k3ZV4U+QO14W7epD6iJyb5Osha8kNby+LN
eprd5Myw2Xh0FPPIR8D6ngTQNsk44MRF1Nfjhh18DeTyLhFy3s/xdgbZHvjzM0K4
u0Y2O4FSThiTideww1Ppyzrp/Nv9nZBwhAS86vXbcHIHcqjID/fCVyt4PL8tTyN2
HVqmikF41qLb1ODS4cSJ7SbdCfMa6ibOxAu2FlpYi7SfW0mr+DT/4SFFag1cY5hl
PVHpxViNZO3+ohQZB0kIfthqKgeQHRLc7wB8qY/Li6Wztkk9R7K1KzI9qeEN3bfQ
hgvtNvL/IBC+OvtItfhlzTYMZXBREbILfNDudPt/sDLzxut2/8RaFBCjGbRYorzf
eMQOw3JcjbF1KjIWfktFa+KvB8m2JSjIv/bvz5FbzDmLd+iavQ8T1hifqb7EKMJ/
GJIE5gy31bksQ1f04cFUJhJf6NqUG/ZV5NxJObjsugBxYoM7Fg4pbjd8s53yo31u
uY9ReecJX9mhdHUFv+blChzN8k8JVKobEQRU+uzgIdeoYa9kFJnPOdjeQn7tnKSb
/vANwHH9aZ7vhRU8iaYY5SvLsQ8ScS34HUhu3fJ8zkVi0YMhorkdfpfQBo7ZAQXo
JCqAWEcI9AChycKdKQFcwliQhm2dlYnaeyCAdYkYUxhNTf+8XLqz0QfkxDxmjiI8
29fXzG4WJqHFf7YRpZHvxspZt7XiN1oNe5ecfnz0+82s7+QZXM4x4DJSrnYJhkUK
c2XnGi1Y9dTgwJut12DXl9DSf+lKcApcS4KulblS3GFS1X+pxTKRc5NCIVK93YOR
k1aimJWLf0mjT6B+HU5FRAI4Xw5vWaSnU017GhQ2s2OfaJbfMyYiEmf/yMvfQGwK
yY2jAB9KvZjuyduO6vrZRfhDkTi+ybpDbTdjfaln33utQBEAW16qnxZSbWZqW8s1
OEU6K6Mlw60iYIs3F2d70GS2FMuSHLMdm16XK/nWUZRIgxNu5+EcJIJiVDdBbQUx
TSd1mVyl6qfeOfzY/GprwSq9fbcuE6dBpWsnBfuAB6tVrFfTJshCpgBk0mJeODDT
l6cE6xh4zCmO6YSk6VxyBnTWFbe3ATcM4vk/OnB6q9HrFqys8sEy3rX/IZDUqIVK
sbeRXhY1GxLEhHTEjlZ/JBrg/ZMrDQ3qUAV2XmVWQ0SWZc8IXR+YHaJmR+MJAW94
ItqNfZKU6il68ZpbSyz/z7/5g15jdTpNDEaqOrtueoyy2Fzd/CwODEZx3tUQdJ3t
65tqkUgYgnEtYsq4I0J2+8eTg05Xlbq+M6K3R2YiHO+dyx6ZbqjsgDHqb63I/S24
1ZiA5Jd41Wf+VCabMIdkB80RiP4qWj3EAObHOv+BnKcGPnN/0x6jL4zB0utjmgxB
ux+9cCf/7NRvBLmdecKxB8TyZpMj4EixQa7lxGhiVwrIVRHSXvE/LRK+WVR1clWC
/hdS65dBWtKK+briqqBFC6xXXRO4LAI5Qq14QQdKNdKdBziwK2Lj5tb5/ltt33NO
RSbfZNu+p2d7nJTOOvKTTb4KBGP5a1u65xjk267xZR59mQ/jbEOyop0tukLvVCHa
bWqOUgTNMkzJ/cYCvSdtFo9BiUdq26WVX0yaRSwHyz7U+QzAeYDY+t5WhbI8fXii
HOCl7v7MfINay1FxTLx+NQwPqwbELL2ZE/GlqrJksHYl3OQRLEtT4Opg5S+fWKDI
qgxzuW7BL1C+F4GvftubiuhsNcSNJfhMfmOFjARHWUDgB/222zrvMWw9Nhoj+cjf
zfkywZCwG1D67xhcKC9WrGKEI9DSf7n5azjgzKeAu5bCPXAbgpn0Pj+AQ1Sizt+C
RlV0GnsE+g6248n++bvWQZDyJrEPAfTboHwCamBAle5dE+G3EdV/IltkgsDU+63C
/tjyfjf3DwrZfGfUY+2Ulq2IKFgKkrzYVRmd2NNhcqwGg9fNIUDHpktMfxl3CbOt
GZi7+m+luzSJFBgkXhBwxfOvx6WmUiwTBZz2mySHPst7jiVyDNn0iE0uHBhAa7c1
MHoMQrH1qo9dfXBW35R7OBQVXRo7MtI3ZwyhBAL8MRMVuNh5UvmzWxtIX6HcrroQ
bbcr2DQeuYbp7nLUW7bJ+wVPJWCPJ5xcbiB4JV/7d4W2yx6Prx4LjRPgGdg1ogft
C7iKHEBS6GVkwa2EeOpsyKkFZU8RNY3GE0WuqwJU1duOgu3N4QOIpgC6r8iwMrZU
po/IS9g6g1kuBDjnWNPWE6Vb1C1hSNhlX6r735l0cVQxugI3EwTW2wwfOrXRtq2z
XdbOi2iPl8qTkZeYLPc1YUaFnIZ52rAy9Ibx+HlyBmkSZHJrC/VCs7gfDDkHYXVf
B5hpLnSNAEvwN9w7E5YnaY4hr9GJnBCGMhNUrJy1/PQapUUKHjrgrfUwFvH0JE9h
IhABpKuSnjq7gzSsoIyXB7oagJDLSPKLGDVF3RnCPyX6MLnF/am7BLAXn6XmtQn/
6QMq3ly7KKgE949gObqJodcydB7Kh9IVRR7xU5wTcA96kM1MOzrlm32jZRXS6XzW
o7hOQUfjkFwOHTBQpH+nSL0n/bdR6gPnBq7IssBImXGF/Lfb1P/TaJfFjxdKIOF3
Wjnw7zhw9Vi0EIT3tzKD0scbrmrMbG7DgkUGPcTbC1NQoyrTCHX+Q/BP+mhJN7r0
KeFqtqkNO5FnkUxEdn49CIDo85/s/sFCBK/X2MQQY8tEe3B+WwUO2go9hRHSbRKw
gUZD/Wf8Xzqr9tj3KUulpxDU6j49oVG/0VpAVaPkVXYLp2IKntbbZb8iSoIC8oNb
WO932uYOMJp6NnZWZ5Hapw6cw6nzQ2nA2YqwbLxK08yXlN+X9JVJXaSC4m2rsp+K
korXn42v730mxPcH3s2Rmb/JbHwy+SxFkiGHw5nyhbPn+5sAXm54wH7mn/gumF+r
UIzlFUtKnGpxXw8hXOEcjx5z/fuYbx+VwArlXJPF6uq7yv7a4HkhM/z6xG95ZuKE
3/Q/qw3w0BsrGV5ldHsdL7fflUPWKCIKCUlQeo2yE9iqvY+5ITHLbT3VU/Qc80cL
IPci1lMxu77rWQ3yEE0COUbPQljHUdS0A09cgpPADAAbhklsnO0gKUcJOYg8frS/
C4bjqnpAbruOX2FjZXwIXFDd7EhZrA1+Eo/eVKWSED8pUu36cCvCeePDnGRW4nEO
g1RFC/2YY//OiJLTRCAFUUvBiXWRlRQf07l1l338128pyAP0DLM0oUHRjjqibbuk
YCSZk9WV7Jq7ZQlp6bPzsjCIdNM2DEWJ9dTg1tGoE1d/0HNOUE2fPYYG0Ukd2zeq
1ZDbFn+YOuWZqmxIRasU3ZizbcjXisq+snnD3vYoMTAUdgeZiAMIlYi4nIYiS2K3
/9hhlyjUYSlKhriFLtBA/LWDm5KGRydEH5PtPu63GRXoMhhUeg/Mqwv9RhxlGFYr
UTHWLLcfAr5z4rFKq+4ezVYhT+U0YkOrZldm5WZMmWnshYcFK6seCYa8bPC95DN1
z5Lo9Z9CT7z77/mEUlO/CPUOR5MGoT+JyZvsdr3xuhkjYdsOtw5BAlV/m2QMB29/
WiwluGkydWApJms9Np968v+zluV6PAi99ME28Z2Mr8X0CJv2hCpl7BkAmpvj9Vpy
XWVpT/pKR5vvAWk7yZ8EyU7P9OhQGWgSO8mlM3a2lgHjVGPdKHo84fjDwueIFhWp
/B/YtMMzorNKPOaKxx1MzpiIYlo6JqonCnWby0Piu9wZl9PeCFWPiZeWONrVyz9w
3tj3MhvRhcurTY6D8SgJZeRdEJuZVtTEHiHCLarfGDjULHVZFYfYWkS3ry9dRBXi
UoSPNo3oPVynYNzurT+uumhMsScgBt/9cgypPwjjh3n0j0hahxgfK0wcjjJyZjSR
L/9/mz6WuQ8uYHMYhZnVJxLqnHfNdp8WZSWU1D3bUKsW62dWc0kkAtNri2yDT9KN
EB5PIeQRymeNwwssUd7gg6cUEE8SZx3/vj4crTTLP1tQ4aK+vaRieWG0tnBq8Xf5
0LQHytpDMKiINvl0kPfA5B0UvCnHfq6Vt4QZPRWuHzJXiSGrHf6Xc9h+fFmYdfTE
I/AClBX5e558FHu1sVf5NeAkEhrpMQXVYThJlxqNqFm2XKEm31CqO4kxg3fVJ62h
OUku3sXqQc4rLrWP1TuFY5+aT+2o7mUsZuZSQlwJA0SezIolYWQkBFld1AFP2NSi
ZTxpdoZ+dVvfLulf1AOeW7Nm6ZNiHkLZvDXr8kMVPB+j5sgbqNCH0YXBSpBgJ31I
jFuEclZfRDIYJjcSyp4kYABFd6HrzcF3pP8vmlz5NN4/ZKy/TVMBqAD/kJz3DV/5
mDFbbKOgfwX5t9elmgke5uN3msRMl1/NqQ54AMJ54Fpk3NnHytBfxdQy0Dqr1m1i
EwypNrwqXZoJbgksVq6ge2VJDJHaHaIoBKLN5qLDbCc2RvQ5q4Mpi8SFV/jcjfOG
4u5MubGPmj2cbgokskj8nd6zcKrdcUID0fW9ztqr0Qbvd/T2n3ZmOtvcCmh7c8Gg
0JFaIUQ8WD5vJo6tRVfuQeqzGZoHQYBpwbQ4W5b/e4qMxBxf+ievjXhxMcRi2iM0
q9W+jqhK2GSCaDJcLcW+wWiG9ao2cw2JcgLLG+aOh+Kc/xKaQ4W4xncltHVOvC66
thAKcA7GFPde2TGRpPWJ86nQmOOtFljje80EaNj7ZJhyvqD05XKJSGaUTBHrr4GR
S22gDd225G6I93/t/2eegGbzfC4mSrF3HHaGIv8MmlfezJo/oIiYFHW5u2+anyEg
ZvnUtzvwGMc7zzmE7Zd5vz0Z1petNNMzOS6HT6IfSG710B3GwkTWcbYkxOgl7Rwt
lOG6Lppuk1qqsUHyRf02PR+yWA4L3G1fWFScGACXuirAReZ8OgrOapGzjfmd0DUo
HZyi/+UQN2Ngnff6BY1QbUEiuMGiRK3dhljnM8DRS9ht666bqtUzmArMAqPbMy7i
C1JCPDf4tkvuDiJsI+0+w54qmcY5xASlKoeu67RavUqZIvGNbqnlAvksnPtDgqmL
VJD2ituuDeObzV+tGJ2uyarta3ZQoEqyUFE8Vf6/LMUNz+BGvCxPx24NW7HmceQV
s1XckIOidI2JUs9e+xnERJVUTvlJW8jptRvWT7/fBNuFZHAWGZGmyPwd2urbg7SD
UmxglADyatvHxHEAP4wY0Up/G1E/IY2WgzuznC17R7kHr6QvmLkj2oJGo2n91Wgw
XJ+A1lLBRNrwoqJgiF1EHTe1m7Sp7aJB68j40Cw8id7avlIuZCbyopyOQZekBLG6
8YUvhKQhQe6l4blYvXpSANKsDPdgJPmCmncxTjygV5ehqe4U/YOHO59ZOWrk/lOk
iBp0koBJ3V8SVLQNsFVrKTtMb1p5Dm2uLrP3tpVNRfdDc8OQtiHFDY8hEaqKbc+o
ZPBjUrKgM+409tJ3JVcxcLcIjT3DkUfWgMrVvS4dve/qNga6bb/iKPmytYcf2iVp
ep+HG0oEVjIRTOuczK/EKLabkT5Qg9HyyFvgKvqL61hFCmeENRFxkg5d7S14FzBF
gRaYiyulvyFeXqrKxYeXLT0dA1IJPPLSb6laDuL9bALIaOiTUIaatqD0uZBpSP5o
iWL/5jgnXjyYP5A+CIfG4hMAeFU0/G2sZp2V/zPizU+y01MjaD8X+vYVnbu6Dy2b
fSNt873jLyloa+pjQs7A2oYUlgMIejnB3oa7flHuJvQ6WJ5FBs0BLZmpzuqcT/la
XcTR2z41yQa9Y0MLPTLwfOmAdO/V0eWTy4mDbIZGt3aIMrLOUHNusGJ7ZwcWYjSU
hmII/tQOhT51aD5xAvmRALQ6wSlnhahoeBOl0i8ps9MPBGIyLoqPg5jQufGkRM7T
3fODjCDrOMPod17hEiXQnC1ZzI2e/I+K9BBswnAFU5UW+i6PXRl21hb/Nhht0r4p
7y5Y3syMoLFprW0nLzEfiM7s5Z3tQY0NyEmf1Ri5g/hg4J0Qv+iWuM4Vr+xAqmPI
UUJ3KGTwG3T6b1hn3UAVZvFRwbrcbDupyoJjgDUiqvZVfS0hGppCQ00alEszPx0W
+Bq71mjZ5jwrEcwbt9xdkr48frEIBG4i3oHDKkSG5CCcMKcSHfLk8NqSbbDYuOUK
+SbMa2S+GGL7YnGDp/12MVv5+rdV9w3Jdh3nl0dzAxEVBpZfWaxq+fCHL1pJU9W8
y/BVNmXv7En9oJ4W945gTodfCMc1PwTVWn75WauYIDRVXJek7KpQ7q9vRBICatNl
cFx1imm69VAPMKkER/xnVvv58dOn+D6WE89VcqGI+Yo30LcUFCdtQw1Z36r/B5dV
3TEofWNZMo5x9zTxNFNmgYMDQ1pz0ycgzy9Z4UaESLQguTYjJyWHfrl2OZGiF+Rm
+0azE66rM9Eca2SxUnvQFW6/1LK16TY/wYKKGLCSw2dr5gIgstrUt65rVcJGKNRF
E7VjgVzMp+3OJxYjCXbDQXUQEmxyMVZnXOgYyz6aerDV75bDQSiHYRW3S7atLnQR
5VEHHxx/YSCrRnLfDA7przWLjwEh/N6/baAC9paJ5Z5EjnuFk7Y+eSUEonEJhv/t
MzkuDfB++3GBLInz3NKqoCrZzaUuNZBVRTimDhToL/78LAmwDnxoQkeZMPyIbqy5
FQB7TiHJjuKvHHgRGL2MH0jynwhNCGy0iwXIHIyRoslQWzrZgNCI/3XIqQkysW4b
je2YCqrtQscOIG4RGQS6o+GhWQ55wD5iFqZOmRI4Tc8UBUR4Wq/pMojMial1BUwS
UJADdlyzrzAuw1kkjdus4LfRo8NgHIh4hY/RpsBKD550mwvwLwog8oEGme4Uqai2
Gj734MvgQ06K5rXu2i/DCJ7yUi9AyHzrB7wXdm5wfw0DbG0lzFbN1oz7N5flLUce
r7gfCdJ9hOFe+87BiaraPdj2CMAh4swt5HVENt9Jep1wfEK4raLAe3aKZKdSfx8l
Ww4cDZi1yGfc/lQqriKTT//ZkVoE+buSAN9yMXrdzpT1MXXgbAm302i6j0pPA32g
aJ1WArh9sD9kcYZEC2AbNRu7zY3aVQblZxsrcIccu2HKQGXaQYVEXqBApRBS6EMV
qyIk1GoXzrnbgrloMVvmBd+AZC5dX626/kC4z40aqC1Vp1IjO+ffptqdC+scj5Gs
zHCSXtotySDZGQw87pyLBSXqaipGC/Z9cC9DytWWhasYJFrDkGdYbZCOWYPY3izA
qNFfRBqCOiLt1FjnYPhdKjIE+EVGZNWYCqZHUrMtiOcHgrJcCRdMt8VUIunWXsxD
ee3J15EVLSDgzUFmKcddnERgA89sMxyDdApfjwbinEMIYt41A3z4Vdl7DHTg1H4+
auLKHYxh4Q4/ziN2Xw0XTGVJcVLX+JhS0HTKhlL9MXlH62sm/+S5FqK36llzcITa
5Wm9e3SJvfWf5k0IhBG/QlTMHewwERNtsvSJpqdP3yIFHTdGBfurdV/9UW+me6uu
ajjHGXS0+L8HMsLlaf/t/TL/wOGdAl0FOTAzVsrbTFch6e3xr/0Jvevizw/bkYVj
+F9ZzNrP3JZXcOYmt38UfyJ9sm5hRXMHihJFtx6metvzNjBo57otnOwV/finZlLk
v50ae3VJY7W4evciUIn2I1OwbxrN1+jICPHgCS9Ab9wcS4YOayvuayeLLwiB/T9w
A6WwhyzWCjIVksLky0uJhLPC6bbYm62Uk1XUonjz+px2vr7ZxjxCt6fc4s4Ft0B9
FhJkj3CJ1QugvneuAC0bjHUzFv6/ffeKqoD5LIJhkP86bTauImnj5DdLb8oEXFto
ksarz6+f1fjE/XvSnynDLCwYu7d6fk1J2uIAzhSWqq36H7dDOb5hZ7X/uKa0NXjF
cB9Ia1EjnzuQS7Ovf/x5srg+IsfaZqiwsBLVq0afhcrmuyogx0ce6ZS/ONd7m8Co
1ari+CSGV2fWPmVhX5GDI9efTqUs6cy2x44oBqQ+HFNUgUg00WmN98PZ8txjr2pj
240oIdMOTAFUNh01ki0648EWK42+7RcqkZ2aQr51M81JCrpUBKX0PKCSWasIJK+M
fDWp6LrhhhNKPwG13ec2PzFD6yPwdU9LBqEwYrT5ywC0Fs7m+wAd1z9cHOPBFE8m
vZ/AcG5MQ9Pk+trXD1oOztk/af70l6NWilxxhVry6K5qFxjGUSN6uYQ/8xC96GsP
/erXo4dtAxuMRGn+Ok6x+v07S0DXBU/ZRnuSaxQATtJzOWlNfvP+otb4HyeEVpFD
4UDkl0lWltQOxtskfyGqIaipTLfLTMuiZEDBF23ixpAdGBkGYGoWboFuUSn4AZ8x
z8DSnPJneqyPRSZM3Yf41IqUFLDdQCzS+uCJ3a6xy43Pg8sWZkV5A+j33QqhRKi5
LySj2IbY1SIsApX0+1e5A0ncLcH/Gmc0XvmkpjyWnnbK74EftVt2M+sQfYt4T66c
j85qwM4g4Mc61qKxsPTjHA==
`pragma protect end_protected

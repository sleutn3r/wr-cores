// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HEmbODtJbFsd32Ki9B2KbMS7dAi5btQ5WhFN7PYHRyMk73DBIlbLIJ1NvMoA+a2B
G7CL0IrpjTfMl4MnYV3VA0cKRCR+wgTZKCXol0S3eni+Sd4EQ6BJaSLidvA2Yu5w
JQffZ7CjQ+BerFKBWIGloNNsVQR8/5uomrY4BckdUOc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15376)
ofaBpfIIK5tXGcjh2H5wd2toEWDE450e0UwYDIvt4bgyxmbYARMhTvXQ/VisUnov
RE8yDIb/LNXVRiOC73Aei5We+V6cPBic5PSj4E9VQBU4ykkspi6uV95Aokq4bdgm
UMxodZOrmOi1XPsPbwHc7sjDuVKFYIl1DhNn7prrJRnzP0R7XeOAMkm4qfRU29iq
JHSj3poXSXcFdADPSnq6CoiN+iP6i3HPrdduNmZBSbkmvLmYePmfEuc9hT6BOUGw
6QSAUxxbixM64AP5PQ1Zwnx7PmapqN9IMYhaUJFvYTxhmO/whyybWjTv7VaWjbtx
7PfkRyQzXhreS+x27BdwimvV2AHBGRz89pKB2nHjXcAnX76x36BKtYEflVb+G3p+
04WLi+6JMQIa96GQQL9qGvuWs+JSSQCAGIoSjmdnyv/VlfORH+R92wl84OMgntTI
qtkYSBEvxp46YdQa7J2iluqvMpT2UzwGda7BaPTY5PiEhOGq2MTq1DFWW1twkoEd
/fmrUdya9JDWRqvOD5TDPRC4FkArropYK9fWVY3sPyeLZ3lGJ8SJYaSEsWLgrLJs
gImji2eFdEWSp9wJ7PpjD1TPJK/R4X74/l5CE7tP2yBzJYIoobrkQIlzyq//Kn51
uyyTlwIBDjQJ6+BkLSmt0pZfjEKyJsE1Y3lbCQ46WZCeHwTE0CLymboLVxwXVZaV
MMhG1nshYR0+QjVKSKu2+FFLxrx1ysujaaf1pNXPEKaCFG/7jvvzLneoc8CsatGa
VW47CKoBxAWK4qdN/iPdGstavT9qfj19Wl9YXeBQtCsJdQVpcPte46P/e+jxhdy0
fBo8/ojz8IbklK59HFFohEoy39B8sHZ4dIjh8BPk1qJO9FGyrU9blOeC5oE7xP14
KvxWHrVO28uBCFUorChI6xM4ZZM5SD6npqYyp1c9GaKlcmd/fToK8rWKR1YJhInz
4tYDqSXoaf/UmppxcBTzo5inmtiSiytwri0FJjjasi3yzCqf39LLwQ8KiZlCGYsU
+bvAu4mdFMzcp6t5lktWtN0Le3GwqaONh/aY/9maB0EJnb8Gt9jTDqbXe5Ng5P19
6+dFc6v/lNjwogICe2aPlB9y/iM/oQaaEwJN7C7cjdWkVDrjRkI0k+76yzy62RTB
BT2zIr9alU/Nh3oyf1JrjYK0owdgnHfIM+k4xLxBayfcLn2xu672mQWQA9fPWaFX
mbykRAPPytlQX8IOt45x2JKfkDKOTHOL/s9AcnNeIwxKHryDVA4w/RkG3vFq/wac
0pRhAPRPiPtGuPFvYmWRjPWXMo3HL3xIo1qDDgy7QRp9AAnmdQ8AhdB/w7Gu3Cnm
PDuabte7aWQaI44SLPvW90H52ZMmTq4QxPIT+jy5MT4Zm86JE5uEDbjHCsYqgq1F
iFJD8zy88bBZROFPJHP+dVlCsYIp1+Z4RWpwP+chzB422LlGquFvyVKeBp1Vc5zR
vG8z9zAwE+uf/NVdPVtDlhcnM6Osf4K29tdag9tmWFRko/uqGX7kpDS1dHHLqdjt
7S18jUhmcR2vjeR8xCkGUsK+vM50jZDJuaCY9ecyCvXD1Z030zq/tOwKxCjiT9q1
jT2h1ivAtMp206cK8EGSPZ12VbEJwgPZG5ttyvI2r9WI3mRoGxzDzOqINW6YY+78
M47pM83cKp0z/SIR8LGY/vumQ+kjm35aI8L2V5FuF9thOZvEjOroZKpHqwnpwVNH
mDlHB8JR622MoMdKc6L+BmA5E9z08WI/rlr8MjZyW777qMpwEqVKfIN2rKVYT7RI
xlFgXJ9O+tv5T8ATJE1eD6DcwGch7JK9RqC3HP4cIeaWPRFwmY6A0WTWZyPzjeab
w/WqmSFyItxamZeLQyZkQPzo0O+q4wZpsmWYahLfsL9RcC24Z2gDf1Sk2OSL7jwi
432XdkDVeceRl/S7zsv38W4kqhJ9d6dqlG+bzvQCR4SeB36sHARVPUFPgv2keiG5
aR2ol2ouvhoaiS7er4Qx0izh+mErBNPHEhRGq/2P4lFffA9b4ZID31x0vsPke3oc
6tvLw++4nhk2RklGX1Q/ApXrb4yNWrxiD44URcCzURxKIg0ShZluuB9uFThF8Skp
6l8ln4o5YA+iE+9cwwaAj9nbIpKSt85Awqv7NS7j55Uni3e6b42unilIFLW6YHl+
nUU+vt4XeuCyfpWa2gVed+Mmad2jHWxsABx7Q+sfibQ47kLHHEOT3jQNZzTK2WyK
4Bv0BJqyZSJ12csmxB272gUOlTHbLmsGoTr+2RypHT48R6gMCyaV1kgyPYsGZS0e
mufttgBDF0uzqYv5Js3L8nOXD1LfgZj+6Dq6HVDwdyoM5jl12bsQ2zQLZ3vyvfjD
zjils2m1YVxdD7CXxkMK1FHcnpOQTlheDmjU+JIzo4NTOr14kqtGE//O1lSyqmfc
td9q2NZZSpydvxQfEiw6dPJionoSD7pODwaBdlEbwMyvM7pCS9WPXErE/2RdrCmM
B4dF5kY25bIpk91oOQvd3n2HpDc5z+KFYSwvtW4UGN1f7Dws8FdxwZZGEiBLcGY4
5+Ny3TZ6YR03MoB/iTLqrYGUiYnbCh9bes/mvpOT+6PqxPU+9VdsqDLx+pvXEo4I
2PMfkFSR34TNJjp04ZEIvmtgM+/UZH4H4HaLGbEVQl6eIfEylcuFCFonIyKa982T
j7GV/Zd8Jq2uM2HjDx03uVuPe2evBulDYyfMikWWj1ybBoGyHtAdbsZvs4vF0HDm
g8dgN+ZDEXivOdHdCslweJJscbRTkpwwuBnDisK+BOqYuF3qkW8RGCJYy9VBFFuP
+Uw+f1gUxONp81V1RhR/1NJIldXDSl45/9GSkkfXiKYhCXSds96KU5rBeMvccal+
q/DJPpupkOpiGc5OEwV7Yq7rXh64jJ6udj8wAm056LjpnaTIdndOcpfogtV6fUda
uh9ZcmtRGnUUy41mP2rHz352N37h2+JAIazIj4rOvbY0fZj8gJSs7wl4QAtrMIuH
3Na4iMP3eXVAmKdclNlugzg9Ng77BmhCNw7OiqHM1WV4dKqnTv9cMwIY7/Jqlco3
7oHADRtGdzUAQrBTNdpZ2k+OHepP7gvda92aW1uHHbf3EqkKl1oBTPNQnwj1NGJA
GiMC89TRlEFf98R5SCnk3uhVm+7vylVk5LlRgue4HJFtFdcQGlie3anoYZXNUhXt
YBznCW+SiQrC7lcwVWa2W3QwoqmE/aXL3g+aC4zxHnGAJ66ihPX/pW/fCU68p6tY
l1cw+MEVIEcCy/7kVUT64mExzKxVdxlKOs6BuuDnjDV1pVyMmTSuf7d7XT20JseE
XvKSpysAItX7n8S4HFDgIgJmY3axlq/8rVMOCb/lwdcg1tooNmhDM8qoUtZENDGV
uXrdsVqQBQTDRji3G1f5Lpw+kZWqN6lTPpJgBoeu02fa6JnEjFDloQqwH8gwIbcV
6W4c3RB8uNoAn5vUkCASnmAE4UtZZKYWju5JQdyi6fZ7uZbqCbA6yHGUi71ZlGfs
XaXKGg9nGncyJzSuQbUv0kjjcCgeMgWdc5kIjv9Lyj+G9ub0wd8FrPoh8nJWe1PU
Et3vYARoNVODVikTHJXHi2ZVlRO2WE28TX+ANAzG9M70yrOxSU5bCpilmDinm1EV
TiMbcul/Ugm4dDBZzbYSeheLyADmTL/sOeC+4dUnpgEipEAA5da8HbwmV4WRseSu
58O2eQ7p+Z2PUkAYoN2Kt4r9LNgSmjFFuQQSJCmPep4yMJ+a+JA6il6z1qEpJN3q
zsolV5ZeTGouuk/nKvMV65ZP/PdtGW2QO0tmlRV6+e595UgcMaijozO2oBu4eurJ
60WZWnfQ00yGu8LaEoifY0OUBqfcJEiHFtqiPamq9T4OffEPm/EY3iwLsde2zCsK
RQb5z6fxJNW2KCxqZbNquB44xO2f108p6sPUmrEhNKDJICI8eXsGv6qsT1IDLhZp
9dD1vqjjddbFDxfwJSJ7yAkxDColCaHOO6omkZQH+QcAWwggfaG/vvHaJZSOijUx
you6YoLM2kliQetTLjlYTYLeIOtzFA6uHwVhVhaeB0KjwHdl0BarY0xOswdglL0r
3BIJbdCUMdaPlCZfTYF3SFKIsC3LZxXA5AJ7zWKTtqiaQ1/ZATfzokicj3FHy2IK
q+DZocC1z8kSN6BgMzdR2rGg96Y/7V/Iy909HgrmxDObt75tJ8Yf6RW5yD/VsX6b
zGWzihQuFHmCmvtWhAjlUMPUMAv97dmMO8piOF/D1R0t5I/Y9pVI3NU7Rh31ZmIL
XsIYWCF+y5tZr/yvtwtT12yqVKlxN9dYrxEGTWTu9Y0876enpXJ0JIIGpLpM4kOE
gCO8PafKqYrPL48JycFrwZ9e0y8QkgCRVVhGSBHNbnt0/3DdQt8fzUrvtUb7c9rc
mTlcInYqCLgPcxXzlwgVO+0ipd3nyXnrAf/PYkx6faGZulMxIlgqJAoqAso6oi/e
Ma1wLe7NDKDBNXKoGk6qNEkrQ8MulovnXu8GU3yT/xQb6kpP4RJNzorjnv7N3FP0
tdxTXJckyOi4K1dNf8CQZR9WZlVKXmoMpvLuPRl7dWd6mdZVFOxRFFLAHa7S62RY
Bn9kL+3XHrv8X7vaNeQVWk6qRx5GT+ImnJfkQQApDmjLosSjAnEyrRZiDqHa01fv
d0e45HXQNEyaPpzD8DH+M6vSbkHhoulxvPuwotQMKqZAUO0Orj8H6vE8iX5cj1Sx
oyy5QCBJIBzLOz0sauuaiczGRlxw2k9hwiNahwDANMM0azH7X7T6NyVNjTN2f+5+
WmZwwBXU6zaPm7x9bXVr9NGA5/ijgIWzZSmKmMpIes98LNLLsDgpOn/t35YKMlUL
8WlnucYMnz/ipMh7HYOm7l3YfdwHDurSoQj6OfIrcTJiu0FAI19tgt0el3e+idLa
ImV+qpcx/LOkzU/P72C9VAU0c8B/3QGOHIzFlY3DVr52RwUckeIP6K+/jG1wbD+O
+B6TY4cmErbl4c2pN6h00kRUBWCtOsiatSvfkOm4C7ZCiqf34ftIVumcAO1RvGWj
/55MEucP2RkAdqSRMkW75CXkhHa9tj4pYE2nrwCIWKSdYTjsr0K6zIW/lysyqSnv
10M5KHVDuBHVUEXnhszER1wbSpKYkkKDEPP8dSM7s8ed+ChtNwucuGacnPgP+rTQ
+irGdKyJySm50UP4+WGv/CXaSn6xdNjWaghZ5GVkC/XmWqyIltZ9FeYh7sWlW1X3
VIVHp/D2LsbBzKkIJpEGl3M8F739tzk+OhiYQY+fpsLt0AovmhJCM16jO6GYbcuq
4zGx0lw4PQWg5pSeaybWWjPLOrk+xDBstyl9qk3rPMdiv17ELip8WKdPwvonBv4P
pGzYzsjJmNm3JNe13Iumcj3/h0R9zNJnn/CwiE5JO/3/KLRnTftVuoyn5Cj9ArYq
BZd+NqUh4QOq5nFQr6IZ8zxkg46BRzFZsSahe+zJJ7LNMTIml6ywjrgrLsChXIZU
KL2L0+h2v0WZyAsLftUxuDtFY+GjQ6r3fyyQieP6QhrjBLqu3Bk9+TOGHw7Rmazx
7D1Mi3pdx9a39RwlfjZ3WaUgIU9hqn/c72+Awxsn4xK+wXyKtpBf9tqUIRp73YFx
7Qo1IayOeAfAMKh/WKN49XyzixkLxZVhxOmmM9wH3ML3n9EdfNdngtqtY4PaUaxG
sFa2MO+apM9atxD4/d8Jv6dthFIBNxJd5BhxwJEl66R2GFqliTX0ke6EW5HostCx
X299zdhesfpWNO0tPjnGS/16QXsc6l5x+AYtabDFtvyl06QcuglOPYpS2qXXec1v
iBwuZM4pUi2ELKp3KkOD0JghGxqcKSqbBzbcpxQdoyBvJehegVptsiKGmgrl3M6Z
wfRSp28FkNT5wSEyBiZewguIl4EmQfRYeji7N5kE+Cm+Us3f5+FYC5M3sT84cgMM
+pQ/dLSDKvQtDXU0Xv48+FAWHnLRDVShxj1d202/NMj+/Fr088k72hL7iEB8s7dQ
DP4sGK9921I3r5aNDLZ+lghy9VmaNPFw47F3k//ZstRp1a4CDmexUVOYsaE5F6Vd
/Y+4zAGkjuTTbVaVb9WoKneD1Y5Xas93JlRB7q+PubIgIq8fonI38dT+Fe5MZYiJ
RQZ6MXSx+QF5bxVuAUyfzM/6r98s7dH5q5zum6bCvnr21okLM7Dk/lG1ube8Vl5b
c1beW6+++w+EN3LHEdxEqWy2eS7wFEf4BSGLPEzRV+ju3tqgsqwIY0XbJ4KEYaF8
mnHplzB+3h1pWZVBB/3DUJuj0H6KPFXp9O10MNMetOOnbNwj5aBz6yVrveIehS12
A9EvOL/wzauNQB8dReZjOH9tzrGtzRCjwMbH5s1chOrBAwSDZXREBBPd84m52w4m
ctCoJCIMEDosFcoBRWnfSgzEIv4rPooguLyZKQG1wdMnsovdFLTRjHIZoT9LNeWM
n9p9e8+wifgulO7AJuDT5ehQnSD0ELbebGc333nTkpeAwt/Ca78C3YpQEJ58NFDY
1htslQg/1k/E3mLzWyeB9cxttCk9rKTS8lkiL4Z/NDDZnJIdOUwe06OwuuA+MyUB
JMeTxarleW2pryUnjGO40sHNEitLPo+mQ/FDI04VnmQ61ahr0ewF50Cu0tCiE/1c
HD4TTPIk5Pdk7/rNGcrH0+6lSUTNcEGZvPJjq38VwKPicsj98AGfYTtAt2IBIeK0
Z0Gtppq9M7dSvAl7jxIwvLkx643iQCausOOrAsr6KC2Mg2Zy9L+XIkt+aOOKV27L
5wTCPxTVtMYXLiMpBvWamZqEwLJJZ002WB2PCl0qld5sollVeXDPPv3h7XgQSnDG
mGZsbOia4HFjakf0yErxVSBwfD2EgfJJzRiTA4yMmI2xKvZEefgiBH54MUxra835
FFxrdyHnXNZrR6eoQmkR1DFkt/TueWr2gax7adtELTGHntAR9f8QZvumeCrQdELo
gFqni6In69Au3t5l2PRHZP/ez3MxuxeoZyfFM1dg0sk+fnPOXoFSub5M4lNCIzOT
pClD8ABp1DOPOXRqJtewLn7SyHnhPSQCAwbh6/254K2CYmCdEy0VYs54gavgFBJo
YdnWVKxncKCHK1TVJt83fNvtDehQlfbpJ41jHyPZ9C603ud05fKuCVlRLFJvlqND
302ODHvbM2g7BIMplhx8bEo/QOEfaUSDXJX6UJPHOhhtEeudGYVJySWQBcc6aP1y
1YcDY79jVC9ee+HbZY3JeAZt41Nj8Quwy6QD4E4tbcD1ilpKRYblLd9mQquVVrn8
0kGIjvmw7M1nrK6i9a9rVd2WSHMVyqx446H0MSUSYXTQot9Rot7M/3xD6dB9drYK
fnqk41sa0cSt8d5brtSuPQm5ALh7OUUDpzS1vOUBct+zXaHglTtdsRZuz1B2DuSE
AmPFyVVTucsz4/14f2qAlPnfWGuxULG7d5CXwa0040Cuth9FDVgdxRLB8N8Clzmd
FQwgF2lslkeFPOItCgAw5EkrO/GOkxA+PzYnx0qwKhWG5W2nFsJ1cWYYuyDjKgaC
nQUYmXnvVt3jRIA5o0QjuXD9kJCTIr8oEhSJWq1cIZus2v0jUCN/+pVnh7oMAwTI
ZRpWykVOXNQ8Vx/aDUt/GLbX3h86RegP3uLxNyziOUrWekojMFpYsDucfffpQtel
82wqIKz4UsPyfEEfC7R+iIwXjgaEkNXN1viuECkAtx4z9qSVNrJyRpDRoPoNkCpl
43OcSr1474G4DcObMjd2PgNHG8r/dgesepJYfzoa40OSZdBsm4RLN4y017MfZIRN
aa2acDaC7v19MAtO1MSgcavNQKlXwTbd3vesTwS7n+Gc3JrTP3Vjhw0l21gmdl5R
MJHxPEm9hhgCvEbTijufRuoGFKM5dwfHsVI7X2KH7lM9dS93a/roKDy7Oa5GS/gn
mJTcBwRPmH6BVWugZ03axXSQeyN6AG7ImBEJ0s3Iv5CtSaPGAr3oCfolflpTLhvR
8zr0Be6hwZsnyWRe1cf4P3Fb3A9H4t1JZ852ROMMyaWYCu1bsq5JCNJmxTotIBHl
ulFAxCmIjcD7zYUGuNj2h4W2SJn2cOvQiPJ4m3HzpgP7HR19caMQjqlq3tUGnaih
Ljuc/kVp2VWeb9KFO+VzmiOlHM9HOmohXpcA4G6M4gHZ6q9bkSBXjRBlS50i2Rjt
TUJkZgF7d7R91lEdOfFZ0+uwCLEftEaRXZTkHJymJrp5A9FxURiAHqivnrrizTEI
f+bUP3Daled8sHyBezsOcMBxiqd7jyA36+8iiZoFOj4+cXmk3MgTmVKIAei+HcXF
7Nxr+Dk1zDSghf8vh+RM+mItC6IkwYoQ6Iwe7540ixAx/2VkH4xjgG5CT3+XyUyf
W3f0Y9L/Mkc6YXLPxLhCCm3nP3icPcFMs6roVLfLtuDGkTpk8keL2tm4NANfnY8/
0ykOaSc/DDpcMnrmshhpGB/5NXzAk8mGt++UWXQZSK7Y3g5jno25h20sToQ/mYaU
ltjVxWMPbdRERxKlEBadKwfSNrWKpgwYndSi3SeaQ0O+mBU7V9kmkaZbnOh7zK5g
ynyJyDRn8hdBBaiWYr68NPXkTuKrTFUYvKYdND+njinVXicLB92OIzTmao8usd6m
mDJI2wcuDrHTEyxWNfbPr4MooCAlZSs2euWEgL6ddoJaMsIsevHJPsPR6ZM8BPCa
eUtOW+Wui40HPc4eDm5NEEttnNu0gXcyaT596pduI+uYjnybA/BGc4gTxh2RRBrG
wVc6Foywj3mf2l7HcPLUT8hCzlkYvzidftkKts8PW6kz02+rijT4dteUQdRJB+pS
3PkokO+TpPUmGmyUcFABI1QDFxIj86sR2vUph+nvXXhVCE/v1xZD1SyLIAaLkGB9
XN/nlq/pgonz/WpZAstRhQxqmWUvKOxdliiPESvQwL33tzPDqaVy8s/X4Ea7DX0R
+Ds0CnUrK3lVi5iGRkofvGmkql0LCVGTURM87Q0dda+dggOxxySHDDdh/FuHv2SW
o1SKQ+ShHVbdsCcCKrKp65v87fP8TSpPNdkm3JI1cI6pxakcuA+MkkqLU3jGEkwK
b6/f+KqrYUNruSffgCYllQtT/f9bNG64Yuiwexn+atjQLI78qG6Ph7T3vjPLYGb5
zzvnlxLh2OMSq2tpw558SZ4RvdJIhjPuIkzGF5sCwjU+Wj9DtkSN8esgB8xV81EO
8Ix5JNtmpcVAxtrb3z0+IvJKNxT8haFTSUvPWOLLFKD4cV5rXMvQmgMFW+odF1V/
hSaMqcuyOim220IbIyQE5xxDrfTnoolvr+8DcEsZUXw6SODU2nK50gSFJ88Ajibq
4uUXsqvMEJmbhsb/MSsEsNsJYVhqbMtZOzA+LDLTXs1q3duKs+vLpl1Q3BM7c3cZ
NbMIlXdjZuEO/tC/oVY8eTT66eDo0ZUzLZ1RLJlf9rEEvypRR7dlkLfSROhBRHFA
S1p6oTW6jecN8rcKDpVRlqnv6GOrUPd6Ji39ECYkbqWhjeHe2fKzV0emBPgNAKsF
xqYbzP4LHN/jrhbAN8eLYrSXJU2aMyhXRcsnwCnRiqPmTINH4VpPI0I2aVlCKw/v
In2DOB++s11avVXMmVRxa46nXkJLHGahev5zD6rtZJhnlNBhUxstu4IEKKxNUceU
YoRyDPVIOeWM0R1gedQ1yxG4hIzDMbI5rFycmLMqWLQWX2z61iCNp+1W1CapYxxb
2DzRqlntakngu65LRoxlFT9m+7j/IaqJpoXDiCJpskqcyYEZEsbQqDkprX2YDYR0
wcIzY2FJdfh06nlauah56cfMr/M+pflsdXh4sowAfZ7ASTmecEhfCwnivhHSJ2+v
IYuGO1+Qu9yHjrkAsxc65Ic75x2Zp5v3mtQ8uRqH5wTZoP1f0FGH3hzW9Ppi7HGk
oT5GU7DJEHGiCjK8nT7K+y4k4MH6+sqCH3GCZ0jeG122bCI4vVvYZMWi1dsi3djd
i6B4xtShy6Pf0tiY1nr7mhdS6r1MCqjSzfBJC43iZqoYExXzh4iSHSImuRBG5HFE
64N8gp3RgSz9m9G/cfVZx2OjkKRX6Z3r+0gmRS3/RO3/FRGnYtQQTB7acPYx23Gz
PVcXUsnLUgCWb/hbuFs3UQSwur+LKxA/E7AgnNW9nmdWxwshhYkQDnL6tbrhvtOj
QdHJUYb61GChX13hX9hn72jualTd0tVrHD8CcT1qkE1GC/5yd62N/Q/8rzYEoMB+
PMouKw23avqg3WKKVGVLnVbUI5QujxMiRNMwfq2ApkNuUZTM8WQ5HkXH/VgdZx54
yuL1tMgKQ0K2ppO6vpALH9cnfVJCBSMAjzb14uNk0lOR+21tiqFzBbzjlvuABUIZ
CPHclywlHO0xM4oi6bs9P1/hIqxkS2/l/whSzRjXEtmdnpaMRGmeWyMyfhp85Ntx
BdiHO57MG5cjwS1IF+4ShpvlJvpB9yn1Cd77x38dUtHJwY3NWTXhzNtmhUs4CNca
l4vHUUeRxU5wMbWGWrm5JaZtmcJ1/s96Q/sp67ighCYe4eTfi3yaoB59ZGtB9h++
JrwFo9JPu+Qw/BxNXqJzCmQg9uvJeGLOEzp/DlDNHcOlBemvrEYksxXIFBY+tsrM
W+YE9HF9hSLh9Nv71/2yJMYklTbmrfxbMGJjeY/FNRHSn+gMeWEddIZBWj7MLJsD
IYwGxTrypPWGlpvbn0ru63OxOhj0rQ8ft6FlgWjC9Yjc9L5IM97KnN0thqsd/Xl1
tmgjJOcIgxyTDXOFEzwp7j8QNrHllNTvx2rpgSckqK2T2EyZdeUEldXpduIz2WSU
XqiAf2pxDrS9TN/9MC8HcLjdHa9IDPBasKfUOu8DlwDhZT1B6BvUFOALQVwqyVXP
H9To6N5hOWFgFkrR3UkzuPSKu4TF92Ci+QFbGHZ28l9eD0MIKWeTLs3AwdYOC3mv
wt8wXIDb1qGeyPRvHW1uvRpfXHwxbhtvD87MDXrty31JxNHGyuU3JO6k7+rvaEF5
QMP0FXqrKIx1makUg9hGox9PnK5TAtgf0T6g/lf1WV1/OYuPXl/1ZSt2i5sI6Gjk
UzpoNx40uoOG8e+Hc1t2aXJEgtLl8+SNc1GIqknJZdPe820jnVjRSv0r2k8TkhZp
owLzj7rJylGDqZLfSjMEamQqYLFqrWP3JBxKauvcP9Mgo1k8kD1a2b8O2DrGhGiN
yiyZ2pY7OrtfV0GHqfhEej8ZUI03luwhcNbgUvu/ZdPGCb496R4Z7ftq7f98y8fH
R4GzOaKR9D5W8k9IJZl/lTsJGzonERp+die2+FNsNti1jXZ5/KRk9gv6AHtx+LRr
uUpPC/YJGFc1JtlasSzEncyEJ6nhylXXcU9wlZR5gdgNi/Ee5DgreKGnDIvmfVJT
pv0zDScFP7TdyBYYKjNGjF7pj8uRIa2wyyjL54oSyXp/N1+8AEF80iG+xLuHDcsr
7cB4MAlxLvWnQxTmhXVHjYlwrYHbKbyec6yaAEOwrYnt8s+Isokw4ma/Ijgo0mRR
pTpo3ib/XhqTkGELVzkp4S9jbf8iYOWYkT/7XDqgRLFzE+P+nj8vp5AQ9Vxk8QdO
ChvCzWdbunI1+H6ousBtll9LbVh78XpQ38/NKJ2LbfiIhfIwVyThTSNbpp9zYMNV
7ux8DjACSdC1Z41nSLydmkd2nEcnpsSVzoNj1GLe3qiPWw3GqXq8S4kXa8OnpO5j
SqdWd5sowwYVkH85iq62N01shBd1TlIZhxLT00VxanqXrgHwcx2tPHHNZN9FGEBL
K3UDIfeBW5ZsL0/sLDgB4PrEatLkugz2eHCP6qM2EomzFCOMd9krKtXNRfQTEJtt
aOJ1/yX1m5GbCUzBgrPS/Ub1PjHLmM9FyrWRIby/0uGGviGV+Vyl9QDDRmygL9pC
jKMA+bnJlQIGv82xsznyTyF6mk2gtK/HiIQALuiwOAV6hPf8RVJCgA71O5/iPx1s
T3O/UCKZSEMEsRmLXl51/jergoxBXXmN6MmTr48hCQMzwToQhgyvj5tli/2iOy2N
fBL6ihYJNtLngnvI68MjPKNGHO2OLH4t+RzYS9b4b6M3S/OUbGOmyB7jHUxCwxFV
zhOCl7YLH56ypvcsN9oJWFuChZpR/YOElAZgbujs5NDB1ZPYCC0aqTujKu3TOOc9
VjgGgeU4AprlIyeR4njE0Elg5DsC2k1bJ81cn61eVvnKYGd8zlXAL/88Fm4+VVrt
4Srng6B1BlBaLzPyVnwZNT0MCc+kx8SzWcGFH6XQ/9I4AvTWzzAn/QkA3Pr9cx4F
8rQqinLHE9QuqT7qv/nfEL1uH8xCSOY/8IuYburNMyE7GghJb4Oz31gTdCfvEnzX
vnJlq5EZU0yc8MJ9Fc30xhO+Sw6hiSVfpUEIBBD8UFkGNdXjbPyy1KMFKFE7IHGH
vC/pELFKYtls1PqqiCIi+XlCkG6x5zly3L5BxwE95kD2hptqKuvEePQzcUWIP6V2
u0BuOcHbtv9QUtyjqEJDMZLjw9a12pQHWprEyLoXztcnTq4MIV6OZziamQ/Uv0c2
Z/PMxg3A+Yo3iZ2ytICM+Ladf9RGvfDi6kDNmW9v70BuayI84DnmE/MVHpxGgGnB
nX3wynHnNUWUibI5D2RBxDEq3LJ2iEv7rMoCeQ86zn1pGK1kjjRNBd8GUo62tBAQ
1p5T2OD1r3UFeEiW5SvQCj+jwd2bzYWxxUYzsaLBY7Q9uTK0RSEzqLGHt93Q4KZP
+to1I/oboZPrB7nXRoXHu5KaC3xeav115STSwXE+PUcmHM2L+8UII8GXSYpPThTa
uewxuOXZgmELTmzntUqKkkiHgs2bqvWZKUsumoJ/+2kQxOV1VpXO39RC5OMlRuK/
hUJS5aR8CC6AjnaZyTWstVp1M6tqohU905/mnUmTR355GsqDmbpiwHwfSIoaTHXj
jkppy95SsUX0bXEHZshCuYOkgFZswG16EMPyxHiOVHrJxPhopXdP1SCA7ye/rjvc
slEjkPs1IGE6f7u30sEOCK1PqB16x+FrPzwMb1/0H93nXYsGUycmZmca5q/s/yMi
A7gf+E8YsHmOUZ2SS15My+997Cvn/3zWhUYjxZB41Sw4hviKqbb14paoo58toQnY
PNhfQj+2FCTnv4oi3vDPQ2vTRR0C8LZnTbmEp2u5k3jMSkSbmzpIRWhSVwPL03Jk
Sa54/IPzdWqaa/XezysDhSZxC30ZXkVg3IT+MgoWPis6//bPWxTAtNrO5WpWsW2Y
w7qu2hTSVuXfupieqVGsWubr4GN9BnHHC3PrAzgLBqxIUCYoZj0kA/x1xzxJR6lT
WcsZ1s6CE/B/0pqr8TjSicgG5ptY0EoUUZfw+SGNPfUNw80q1qAQjnIfEBr4rLzL
suRtsIkOSv/U9QdTRJKnzNwQMJQTvPneAGyQOujUwY3cquj4PKt9cQv/mgp5gE4N
HI49Q9yDcAE//dS+9NNaPgqoL+870y5255RxpRZf8O3Qwq+YBF++4pHbb8DosrMt
pyhysbYSGcL/5Tp1XA2Pb6Oc1ZMwZaIgdi62sLSycYC25RDQl2cCkaxvd4XSnLev
geGgnz5ugQa7vXYPRNyqVC9AqlqCyaNpFsAasqavAiiczH1hWrvN2eA1FdHDLGii
04Y+mNwFWP+b0tzD0fhL3WSX8L9sdBmPYTavtBRxVsXFTY3CLhSKQ1OwtDpopCnc
sp1FDiL85zlj1D74OY+0tgC0KGdr7lEWWSLTlGAVZb9LCwY4+6NecxT5F0CmOV4b
bAlWuGHAPlwnK765Xs8es5lQU/zCmhTPv137MIOL/phDUChlVHyxLDzNZMCVy5ok
D1/tYU6Ip/S+cWZjDE4GKC5UdIbcjJfHXgN5w5k4fln72V5pbjH7d7eGvW271IkL
/GDoDmNCeLdp5Rp+3AZGZGf4pLelmspRmbkCrh+Xw3eCBkVa9Rr70D6SNm2ccCoU
g4BYX0EH7jq5qpAi1nUk/6M6JZk6+RxxnT5Cw6RdCrwzXUWAxQf4jxjP6yVvZQSD
1+jkR7MA9YTNgxvkfhmdtH6El3tmIVWuoWSUS4UqmX78eX8ycWdgnwSGydke3/st
WaOLJuMMD0Xh7EvnTle2uvgRzwu9VThCyE4P5jjKnMqr++R3/PHEbRraB6uxWrTh
CRWfRhbq4TDlBpYFXNNeqBkAIxk8AhBt0ZtuxAgOPol4ROF4mV6zgpt1NatTmatS
I8wMjdoChTSYN7T7ju9H3aWb8DbqiPoEufh9SirP4yl4SYJs3bggNnqvPGd9D4rL
JORcJAHHPAIMiUaJD7hO6IdDURBxKB+NfFPNgDVudZa6oBwYXKu1u/M/OnBIysE4
YvaA4RybJsgs5b5atUYrnN/20npNy5sZq7kPxPNuzH3EKBcQaEbkduDQnxPLGSQe
QsZ4FnvY9EiSF4nUonIoqH0qrfk1qfr+ICc30ArW19g3j6ig3viZPPlhvaeIr8xC
2ErbQcmU3AfmCr15T3Dec2SO7Awe0OAfS96gqYUaLxYsXXLmSKKfju/2Ikqfrt9Z
t803D1bIXgjJmsS3Z31PivCIVKXqomsiRH3jRMgdHUreQrPX3ImGygR45GaEEtd9
t/O48Fv/IKArn1/jU80QeflVw6kH5rGkbmuhlYqQtg1gnTjy1RDRdA61B80C/dkJ
e5jETVJc8KWK1O3EUTcFlbly7eC4vaMiX546VddP6TGlr6MNePxuiVymyR0v9w6e
CNGQzj4+ls65m0XmTiKct2c+2G5Gl1lRPatbIV4EY4k+2kkiSkYGPWh+AEG57qkZ
2elnCRbVkrtX3KCrpLn0hQdDFhv1UkQ5LLNJWljmZdqqObKTmVBuwcTHGpH8rZ6/
YWD+N1casGwqwWTvajvsTcxky8BrzSgfZgkMtqDZLRJYuJSlphilhv7HrDn/dhco
lSz6qT29o/H5tmLPO7t7AJYRF3V2kFL7BdDM6niU/YCoEYigb0Bn0NgMbezBeBsY
PqxSToSj0Prq6igCOncjEQj9utXiIfMS3IWM5J+EWAb9PDNtyezBh8bmMKkg5PNf
eJgu2YXsRPokDQElg0hfW4jEFhkv+kftXSh9WV0bUt8COxQSgNduXvbiErlmroB9
dBP/y3L3HzMED15q0wmVJ3OM42txzGWttdvYknNQ025uyTjTMpnXfTT3zUk2r5uP
bR6GLQ9b+iKEikRP0ZMPHvQTY6JKpjlMgQbVbJNsuXS1hGCreCZT/BKseilhLAeK
nrUaN79Vu46J5IBmrWznNRAWo0gSOXHAv4T1SS6q0YVeWu+FxrxIPiEWn8cZDFXV
vFO2oq462/vZrpBhpGobA5ud54NSQKE7VcNkSKflnjdPCFwaro1r3CVxM7A20V7D
5PBzZl7RnYkKGZflvT48xypvxvJP4j8fX2RwFOfH9k4BKLZUepcQbF4ikXV5YvVi
tobnvIjmoKttZH9JFvihGmeMGMrtzie32qAiPc/2ACaB2AoLhjTqsSz1HxjgKUNb
7rN95a9cKLL/46uCV6n/CYEpRjqzVBgViem1Plbs3qA6GSY0ZDg83J+qhZP/9uDj
KVxyqJtEUdyD9k8V4xZZHdnf4xEQH8/OaRmXB9IOYzmlPgkhRcB9wwo5udGa6ynP
a5RpN4NQHxjhrGr+FcrmP5KTNp/8zwlEzcAQc7iXFS95EojSWUNyb6pgGvOuG9bK
0z68+Q8mgNYGivvoy9m3PNaIDG00TDwirdGXd0A+mzvZGt0qVKZ79YWMWa/qOVTC
PIBLKnlufOXXsZSXtPLIIBepDfZKUyxPou8HiKxmiU0puhqMO7jkCYxERIkMClmo
7RcCFSV0pp8EZe98WqQCzcAhsm30Ise8aVzPht9xkHoQrOmSGjLwuiZXleq/9cw1
exdsj1sbpsR35L0+EAsC9pM0CSOM4/RBnz0SCCgNMxvdXlMJ8H/L+2qHOPA6tPIi
vlZQ9eEJALeQCYqe8btlHcPokrNox4hQ+ucnpOaA12hc2o8RZzsukoa/De9c+B4x
AF9Vp6niA9Vv1mO9DNpgDyJMxI0oWOVeUybuRcs0u6RQaejq+tNaUqiAAGPJHXDK
IO/xaOxUMOHKlM6R5EF060eEAGSSg5PVG+RfCOOhpgqcQ1uM0/9FiT2R79icslKm
H/SjeR9M5dnJtN7N25hU59HrxyK7OxmKkuDR7sbYl8oVZggo0/tZ/bUNmaX4BdGx
9QjGqckgCyRSeBOOweI3GARU6TGc8PbSgISJJ2STO5KY1quo74Z8im6TnfIvh+ZA
ow7/D2fBsS5x26NH/M4B7Tl4CZO7iTYhb5JTzLLRU4uRgpQaZ+tHGLWl9eRzsojE
5A0VuLSChsdS3Wj1h3rdQrcDGg5eaEG1vW67yaecjJpKeVSnUQZhaQnN6ZNyVsJ0
/07E7NqndN38/OqvbLCcOevbe5sccIgegVuDslehy1Xooed0yLXMvE/TyWjj0no0
i7VqHyzPhIkkh0QnFRU9216JHjZzKDA/GT/pOOl+sw8o90y+hKq6WdlzsCXI5x40
0zm2L2s1pjGWbR0vuGqOoX+YFmW6zpNDRQHcBpUPhhGO9ulwwlQVIQwcXSM00waj
BIA7bAimWg62GUjdzl4UDxkt+y90dYdmBzzVGVGBT5W3Sb8+wwpyTD2z7eVmqCys
+IDVD2E7lVSsGnlkXqdABt60Iz+Wm2PBt7rKRl0XIZ1n3Z8MG5BveJOijzr32ws6
nNtEZpavJfzeo3OQ5Mc8B8wP0kSTNGZKWJz/iDBSNsrX+clJ/k3brsts6XA+jU+f
j0u52outkYsrzTF6eFvmQgGUeQGVa8JMFvawxdw1VFwBeck0nZkQkxVd1pWJPSeb
G0IXnKG7c78EpawmQ1SDhzkdXzeWwMbNxLdcPvGBCqfj6ojkXd068lVI2BV77Vku
+onTJfvx9owNdwRe5juZKtOFMdC7xsLR4d2hSiTHNy0r29wSH+KflsUZ2cPceoYv
WHqMmbGxYaqzhqWvyAKy3PSUFqs0D/ckBRQV2hQ1EVnVcFVJIwwSY5xSo6Oqxp1y
yS/KpsrlIzdgtPpHViCBool1zJDcOy8BCG9JMkqc/cUqAmL4Zc+z4wM9j0sXqOgd
ElO/CYOqu6vTTmgSAf5ALosC8KEsd3AgBMrLoESiWMXplPWkGh7h+z2lAfNUCt+u
dF24rm/NEK/ar8n2Ylg5vhL35FlC784KuSQtb6nuGI3VwykVpTNee9LFZxmEWxks
49VwJXpqeAjRfTiD7S165PGGQwE03G46uOpEDWB8+YeTg7sv5Uj30t3a7yUJcEjz
Wtrv8naL+Al8wnGs4k0YUM4x4Dwuzu0vMAYkcOs3JhXajwLUcML1vSXaD0rUhZ2b
0UF8BPLIj5DL++DOjOKwG57hQefUXcGAIOeWN8hqsG2Ru8Kkr+X9zLGrEUGFb4E9
FtcXlzQEOSXb+g/J0i/+lOzQ9JlH+c/uGZzFexX93SjMYGIJUpEfRdn/YvcuoMjX
ZL4ShjazXgFFxDEnRWpALrPziCTZEP9OjxtUjJPWfjHzbIdfy84nZeJGYYmQqA10
aWZOiO8STW3o5838VQoPV1hcoryUlzrAZB+lL9SSdCLZs5D7wsZO8LJTTURgfq5a
YwhffZ2K+gdbxniBKYmCUn4f5Z7FlHJuQ7dKQomfaLi1ERUNj8A0gcrgIzZRQDQw
G4w4jP+PaQ/3kMExVsVnwIgWbV0nwOR4Txpl+TDjrSIMPi6nfziXhVBeU86Gt8mR
cXDjw0wdIx5u85cQspz9xXhsHZDRRSEv1YsbnyOaHp8holvGeQqYuCdf9drw5edq
msUqsaftIQd+CRt9oi463c083FsplB6rQsK9fnf3b9pL9Xzx+oRZDbjnKReyCvdr
7c+G4WUMq7gXTCxQod1wsyWDkFIoyTtsfsvySLZY4Sk7tWtmwD3476KnyaAixGJP
cnvmD8Nyf1Z0fHSsd6T46Q8XaCKqXJktoxzXdnEKaJ4w3Rs8XA+8rcA0XajuZbwG
FG+bbEeJNBI+EUM5/a05z3N0eVu8XdP9Z6lz25XVCTzUFTKIyKlb9H8IsxwZUOzX
gPJSmjuJhT5cBh95oFLfXez7uguF7ZIuBXOhfeUe92GZDdreH3uNXRrShYwgrkEz
1MPu1B01DsH1HZOijt7kV1S2MomDAnIVAigali/JMFsqBIM36PaHAszNG6jNt74P
8Y5Nw3OR3WrskIXuFbzZ/ENCF6px3MoNsQFznqpIjXtpbopwavx6vLOKMQyTr8KA
dN6nWoz/s14mpIvksuPAYG5NB66BHlFVj45+Goi+8DP2D9pkPDci8GAGiiwN0csS
QlVtoLHr+Jq70k2M5oBUrxxd5Q9MeZKw1fRnEA16R+wC8DP6OkuQAkWZfeMHQsEQ
UsdUkFg9iU9ZLC3eIrZd29lSJLtx6ieDKBNFK+YzD08JbHf71+a08I2qITc7KvMB
UbRTdS9fCrvIqn9uISg4iXYe4ZPsS02E3HJa5R5Kq+EQEIpJDjEoSQ6z/uuC55/I
LpRKXxeU8kHRT2oMT9JJHcOXiCxXK8NHGVXAuxeCxDFI7fCg2YqvGD+8e5cqyRC5
wiCFUjsjZywVcivP1q0dBm5iI45sD74epA0eiUuJQT8qKFoDiLDaLdEAaNtVJvls
gRYO5VQoleaa+A0RwWP5D8iIwqsGZr2VskylyhycCYwDkAFAPd8gUpFoNgjSs2tD
27mhSaiX3lO7DZx0FH7W+hyqqyfqmrOgMydkw2JFF6azRBfX/avDqNs2UbzspR+t
LigBIRgau1v/5vxU8K81CMFGpdAaQOY4n6yuzKlok9k5Q+9z/8PcDQEKhK0Weu9D
aboLIxlvzaZFqBxBydOGQpcBVnvG91BihWwEQdny71XMxE+Y4tpgAF4e8lROf/WO
TT4cJ2Vk+7KemKVp1prbe51gjb0tQZtZFr1FVtRFnvdNSyrJnAoM097CLcKaU9Km
d2gDER2AwUSXLRInfRxW7xcpbpYsYcyKVTrfC5jXt1Rx9tJp7pf+Bdxd1YM2Cehq
6PDOSI9hG3TnmkFDDAnzki+VBh9HUOWx5v/MYlzp6zE+FVdvwodR4a/Iibh+rOhA
yKxI9Xa34oN0rxfM/dZyko8M13AvMJOXUkYnQxwQJUKz/2K8mlJZzA1Gt3mFyrts
IMsxhytROl/Z5mazDVasM9oJkgEOtbFB25Sl/UfUUR2TG30685OHWOU3H+6MNHfy
jU6iFqDLSduwZk0ErcGviI0cLib9a7hnMYps0SlUSqWXxuVisJScrZ9QmIhjyFQU
YaCpVe5MO/+4PsxnWvO6CTXYWtQ8jvtmWHcPIm8gYzCFfJjTib68zEuV1abRU5W7
U45e4hAMj04k+O2lBK03l6R4VqclGMd1k7wbVYqLH3Op8MQYv/1Y3644XIpkZRTE
REqtnzVdvNCxdGEf0d8c8H+b37c5LCQ5zdVNfQzZ4vv3lg+V76rTNvmkFf9uWqHq
ba/o5q65N6UrY/lHhyUXN89hMn6eg8/f1snTCE5yO2YjFaeR3EG8/YruKwDJxWGQ
9d0IVKKwBUZRT/CWG8vGetdxilrZ4y82rYMwbF8Oj/95cLbdDrjxjs+FKNK9VvHw
h3x74Msx0U6+r/tMwTNB0EZQq1PNHBvzOr95yV9dCNEfdM6pAoS30JwsZv/Cz25Z
p6l7CflE/0luHzbOSeaQ7yUsVsqmELsjhNmmK7o9zidUBBKqVfDT5rgNqTfu9g7k
+sr7HwG/D6/MdVyOkF9iNWlJXdR29Nl4iBIKEB4vn0AIm56CPcVMY97HbNyYhHc1
obFuYhCecXynuXH+06MSXivaNC9r9dHnmIKc8hozp8ng/lbTB1mhgakg26nd3Z22
UCIHuL1C1klI7RAUSCpA6Pq+Z68F4osVURuAfpyz7BSg3JWHujK9F6ebNHVoDRZ6
WoOlJRD6CGF0/tlYTTish8ltCaj8oBZZ8wA3mac1MTkp86B20iaiuzFuyiOO+aCB
GZR/xLJ+gDEUMTEcDqWUIHXQ6HDKV31nvjKiKCwkfQxSOUhPi35wfxNjKsvTLGEv
A/OPyySyOFQL0hJhuE5KB2A2Q7ptLQ0Ohp6L2DWkqjmp+JQbdpfJIFc2iVVtRyo5
U+beWChslKHX3d3Lm/3q7k6/aBp6YgvUzSRuYvFuKXOH1sR5be+TfG2iyzB9mAZA
UUvPYWMcNCRjswHqi9310+fz1gwv6N2ZkQCCYaULmZBflby1ry60lpqpf5cTozty
Phf5tM5aU1FESy6flp1N1PBvdBxrOf7AfWT/gbt5//HvQhLy2Vk13YymUy+R2ICB
LKl9MqWOlBgNwiKDMmTsDSDLc4dH1hdpTwwy3CTriZ0vuBiUch5OG1iaefVZNmvA
c+GuGL5kXsLq9uYxTkwJPfXVKN35k2e9xCWOkHUEnFGtXuVCTQUB8vBJ3awyABYd
rrxBDgg5iFRVwNTR+oHRG/iRyali62hPtnN8VAD6Qm/Qzbawug/BX5uWwvIqC4N4
AfLk6WLbb1luj4+mX8jAYA==
`pragma protect end_protected

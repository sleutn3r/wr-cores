-------------------------------------------------------------------------------
-- Title      : Digital Pattern Generator
-- Project    : White Rabbit generator
-------------------------------------------------------------------------------
-- File       : PatternGeneratorModule.vhd
-- Author     : Peter Schakel
-- Company    : KVI
-- Created    : 2012-08-14
-- Last update: 2012-09-28
-- Platform   : FPGA-generic
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description:
--
-- Outputs a user configurable digital pattern on a trigger signal
-- The Pattern is written sequentially to a memory block with the Wishbone Bus.
-- After an external trigger this pattern is read back and set on the output.
-- This is done on the White Rabbit 125 MHz clock.
-- The Whishbone Bus addresses are described in the wb_PatternGenerator documentation.
-- 
-- 
-- Generics
--     g_nrofoutputs : number of parallel bits for the pattern
--     g_patterndepthbits : number of bits used for momory addresses: 2^g_patterndepthbits defines number of words in pattern
--
-- Inputs
--     clk_sys_i : 125MHz Whishbone bus clock
--     rst_n_i : reset: low active
--     gpio_slave_i : Record with Whishbone Bus signals
--     wr_clock_i : White Rabbit 125MHz clock
--     trigger_i : Trigger to start the pattern
--
-- Outputs
--     gpio_slave_o : Record with Whishbone Bus signals
--     pattern_o : Pattern output
--
-- Components
--     wb_PatternGenerator : module with interface to Wishbone bus, generated by wbgen2
--     PatternGenerator : Pattern generator
--     posedge_to_pulse : Makes one pulse from a rising edge in a different clock domain
--
--
-------------------------------------------------------------------------------
-- Copyright (c) 2012 KVI / Peter Schakel
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all ;
use ieee.std_logic_arith.all ;

library work;
use work.genram_pkg.all;
use work.wishbone_pkg.all;

entity PatternGeneratorModule is
	generic(
		g_nrofoutputs      : integer := 32;
		g_patterndepthbits : integer := 7;
		g_periodbits       : integer := 16
	);
	port(
		clk_sys_i                              : in std_logic;
		rst_n_i                                : in std_logic;
		gpio_slave_i                           : in t_wishbone_slave_in;
		gpio_slave_o                           : out t_wishbone_slave_out;
		wr_clock_i                             : in std_logic;
		trigger_i                              : in std_logic;
		pattern_o                              : out std_logic_vector(g_nrofoutputs-1 downto 0)
    );
end PatternGeneratorModule;

architecture struct of PatternGeneratorModule is

component wb_PatternGenerator is
  port (
-- 
    rst_n_i                                  : in     std_logic;
-- 
    wb_clk_i                                 : in     std_logic;
-- 
    wb_addr_i                                : in     std_logic_vector(1 downto 0);
-- 
    wb_data_i                                : in     std_logic_vector(31 downto 0);
-- 
    wb_data_o                                : out    std_logic_vector(31 downto 0);
-- 
    wb_cyc_i                                 : in     std_logic;
-- 
    wb_sel_i                                 : in     std_logic_vector(3 downto 0);
-- 
    wb_stb_i                                 : in     std_logic;
-- 
    wb_we_i                                  : in     std_logic;
-- 
    wb_ack_o                                 : out    std_logic;
-- Ports for PASS_THROUGH field: 'data_in' in reg: 'Pattern data input '
    wbpattern_data_in_o                      : out    std_logic_vector(31 downto 0);
    wbpattern_data_in_wr_o                   : out    std_logic;
-- Port for std_logic_vector field: 'period' in reg: 'Pattern period time'
    wbpattern_period_period_o                : out    std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'Enable' in reg: 'Pattern control'
    wbpattern_control_enable_o               : out    std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Load pattern' in reg: 'Pattern control'
    wbpattern_control_load_o                 : out    std_logic_vector(0 downto 0);
-- Ports for PASS_THROUGH field: 'Stop pattern' in reg: 'Pattern control'
    wbpattern_control_stop_o                 : out    std_logic_vector(0 downto 0);
    wbpattern_control_stop_wr_o              : out    std_logic;
-- Ports for PASS_THROUGH field: 'Soft trigger' in reg: 'Pattern control'
    wbpattern_control_softtrigger_o          : out    std_logic_vector(0 downto 0);
    wbpattern_control_softtrigger_wr_o       : out    std_logic;
-- Port for std_logic_vector field: 'Pattern busy' in reg: 'Pattern Status'
    wbpattern_status_pattern_busy_i          : in     std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Not used' in reg: 'Pattern Status'
    wbpattern_status_reserved_i              : in     std_logic_vector(14 downto 0);
-- Port for std_logic_vector field: 'Pattern width' in reg: 'Pattern Status'
    wbpattern_status_width_i                 : in     std_logic_vector(7 downto 0);
-- Port for std_logic_vector field: 'Bits for pattern memory depth' in reg: 'Pattern Status'
    wbpattern_status_depthbits_i             : in     std_logic_vector(7 downto 0)
  );
end component;

component PatternGenerator is
  generic(
    g_nrofoutputs : integer := 32;
    g_patterndepthbits : integer := 7;
	g_periodbits : integer := 16);
  port(
	whiterabbit_clock_i                      : in  std_logic;
	wishbone_clock_i                         : in  std_logic;
	reset_i                                  : in  std_logic;
	data_i                                   : in  std_logic_vector(g_nrofoutputs-1 downto 0);
	data_write_i                             : in  std_logic;
	period_i                                 : in  std_logic_vector(g_periodbits-1 downto 0);
	data_enable_i                            : in  std_logic;
	enable_i                                 : in  std_logic;
	start_i                                  : in  std_logic;
	force_start_i                            : in  std_logic;
	busy_o                                   : out std_logic;
	pattern_o                                : out std_logic_vector(g_nrofoutputs-1 downto 0));
end component;

component posedge_to_pulse is
	port (
		clock_in                               : in  std_logic;
		clock_out                              : in  std_logic;
		en_clk                                 : in  std_logic;
		signal_in                              : in  std_logic;
		pulse                                  : out std_logic
	);
end component;

signal wbpattern_data_s                      : std_logic_vector(31 downto 0);
signal wbpattern_data_wr_s                   : std_logic;
signal wbpattern_period_period_s             : std_logic_vector(31 downto 0);
signal wbpattern_control_enable_s            : std_logic_vector(0 downto 0);
signal wbpattern_control_load_s              : std_logic_vector(0 downto 0);
signal wbpattern_control_stop_s              : std_logic_vector(0 downto 0);
signal wbpattern_control_stop_wr_s           : std_logic;
signal wbpattern_control_stop0_s             : std_logic;
signal wbpattern_control_stop_sync_s         : std_logic;
signal wbpattern_control_softtrigger_s       : std_logic_vector(0 downto 0);
signal wbpattern_control_softtrigger_wr_s    : std_logic;
signal wbpattern_control_softtrigger0_s      : std_logic;
signal wbpattern_control_softtrigger_sync_s  : std_logic;
signal wbpattern_status_pattern_busy_s       : std_logic_vector(0 downto 0);

signal patterngen_reset_s                    : std_logic;
signal wbpattern_softtrigger_wr_sync_s       : std_logic;
signal pattern_busy_s                        : std_logic;

  
  
	
	
begin

		
		
wb_PatternGenerator1: wb_PatternGenerator port map(
    rst_n_i => rst_n_i,
    wb_clk_i => clk_sys_i,
    wb_addr_i => gpio_slave_i.adr(3 downto 2),
    wb_data_i => gpio_slave_i.dat,
    wb_data_o => gpio_slave_o.dat,
    wb_cyc_i => gpio_slave_i.cyc,
    wb_sel_i => gpio_slave_i.sel,
    wb_stb_i => gpio_slave_i.stb,
    wb_we_i => gpio_slave_i.we,
    wb_ack_o => gpio_slave_o.ack ,
    wbpattern_data_in_o => wbpattern_data_s,
    wbpattern_data_in_wr_o => wbpattern_data_wr_s,
	 wbpattern_period_period_o => wbpattern_period_period_s,
    wbpattern_control_enable_o => wbpattern_control_enable_s,
    wbpattern_control_load_o => wbpattern_control_load_s,
    wbpattern_control_stop_o => wbpattern_control_stop_s,
	 wbpattern_control_stop_wr_o => wbpattern_control_stop_wr_s,
    wbpattern_control_softtrigger_o => wbpattern_control_softtrigger_s,
    wbpattern_control_softtrigger_wr_o => wbpattern_control_softtrigger_wr_s,
    wbpattern_status_pattern_busy_i => wbpattern_status_pattern_busy_s,
    wbpattern_status_reserved_i => (others => '0'),
    wbpattern_status_width_i => conv_std_logic_vector(g_nrofoutputs,8),
    wbpattern_status_depthbits_i => conv_std_logic_vector(g_patterndepthbits,8)
  );

wbpattern_control_stop0_s <= '1' when wbpattern_control_stop_s(0)='1' and wbpattern_control_stop_wr_s='1' else '0';
sync_stop: posedge_to_pulse port map(
	clock_in => clk_sys_i,
	clock_out => wr_clock_i,
	en_clk => '1',
	signal_in => wbpattern_control_stop0_s,
	pulse => wbpattern_control_stop_sync_s);
patterngen_reset_s <= '1' when (rst_n_i='0') or (wbpattern_control_stop_sync_s='1') else '0';
	
wbpattern_control_softtrigger0_s <= '1' when wbpattern_control_softtrigger_s(0)='1' and wbpattern_control_softtrigger_wr_s='1' else '0';
sync_start: posedge_to_pulse port map(
	clock_in => clk_sys_i,
	clock_out => wr_clock_i,
	en_clk => '1',
	signal_in => wbpattern_control_softtrigger0_s,
	pulse => wbpattern_control_softtrigger_sync_s);

PatternGenerator1: PatternGenerator 
  generic map(
    g_nrofoutputs => g_nrofoutputs,
    g_patterndepthbits => g_nrofoutputs,
	 g_periodbits => g_periodbits)
  port map(
    whiterabbit_clock_i => wr_clock_i,
    wishbone_clock_i => clk_sys_i,
    reset_i => patterngen_reset_s,
    data_i => wbpattern_data_s(g_nrofoutputs-1 downto 0),
    data_write_i => wbpattern_data_wr_s,
	 period_i => wbpattern_period_period_s(g_periodbits-1 downto 0),
    data_enable_i => wbpattern_control_load_s(0),
    enable_i => wbpattern_control_enable_s(0),
    start_i => trigger_i,
    force_start_i => wbpattern_control_softtrigger_sync_s,
    busy_o => pattern_busy_s,
    pattern_o => pattern_o);
	 
process(clk_sys_i) -- synchronise to prevent busy_o to be dtermined as clock signal
begin
	if rising_edge(clk_sys_i) then
		wbpattern_status_pattern_busy_s(0) <= pattern_busy_s;
	end if;
end process;
  
end struct;


// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IEZWab19M98iUGZlsWa5nvowK+j2mXqtkBVW6Dp/aJfOJd+bkm3tMrfV/tYfySeS
SJocpQUQMU9j0m80TBhfGxttzicyzNkTmiZVgoEFaOVrb6NcAP+YDLiQAbuOpT4Q
Hbkocr6kxTVsO6zLRcPbg46WqBxJW/6IVilPbs9tR0c=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
S4K83UlgWjU7hwrtb5DmwcUNplt9Hydozh/Eypsnl3tYpWEghw5DlsWt7TlZHa4Q
GyChr7V/wS9UbvZCYGUnKEoVAhrSkhCfIpCN2v8mpfh45OYkwccuBoSAlMYl0a1F
g/bD6KnX9phJwwKNgsj2xIpuYYo0eiBEoeDjVNPXT9jI7NOCkn3N7E8sYqKghtHB
aaQE65dXiQ5wcokD/KY92Kpec3AbAFeUJ0si7UF9n2g6yzkeNGnMe17tB8EDKGHo
ohGn4Ov8O880p0F2f9ZWZI68SPhWxZBEyYFiximxnh+kjqtwgZMHeEiiQ8XWTiTE
pG1YY0W0kgMMC0tlR00lL/jVYyahZaeQqZWCJglg1BFHB0t1eGisJ+qSG2Tgf0NO
PAGWu4pMDWnEu+pXjFbCgGH/oRr9BTVcD4kCLZYFQzqokcIMZ487I6/On+qL2/KL
5V1/z44U+j2wf3ARB29WdZ5owJ9V9nbrJss5SVpIM3vpjXh0xTyAql/h7zldQ40X
Hw/9dGkK+zQlhc6wTm6vN1a3KXp6gDbRYElsevSzpay9I5X8/JzrPEc9EwvKo7Nz
zFbIGyl5Yin+vzFUMtQJP3KL2nvPnpgBOvvhz3QkRE4AkVdKvushoD939XtjVhCk
KGFcJE95C6zEg7sb5ysQUvG29yr9XxY2YDztQHtid1msyQmxcbqz7Sli2pPlVvxa
3CTnv3XGbDZ+DjFLZU6cp7zp9yI2lFfyz1BT4lEnH3rHHOghhYVhRTwp25h49NcD
QtqGP4kbbWG3FGcgg0yGpRLSiVeFYAyPpUVu5riMLgnrZIg5yNyIunAqpwd0ba0t
RNphySZlNH7sY6PnSFCyIeDis09O4LM9vKjiCIDogZ8Jbd9nJSrId9OyK/Z5y2rb
VFGMg6wgcnLpuAojmoUTPbXEMPqoirdyxFlHMYtpE6A1B8BejHoSC6Bh57qKkuKY
1ByMWfTHRUNX22TkSG3761puZddXoRZ6rjbnNjrA+I5XkekXCOTxsiHmzLRhkKPI
2pzjB7fbopP/i4kgy+NtK/0F4BhOsDNJVD3I2CYmyw6hqHqlvyMY68pAXXrPlBai
k088+NrEsFqbXIOK+DZPJ3ZdTaV/4jcLG6BVp+846TLzqDKkE2IjVzBhJf327MSH
s00jfEdxkWLok3V7n8HdMfRUGAfC/FWOPI1ltyXpcjSetrV6tl00Zp8dOvVNnPAu
woST7eaBOf6RpazlKL017r8iOCsziTz1dmjqOv3MO4PwkJaeoMIUZza5nejRPJ+F
eYrVI+9dw3j4LAbozy2wOtwVFll7XwsF3kZPwB3GNNfy9JZj/X0UW9bx+kpt3zMh
iuF95kqvb9TdE2xzYDw1GadvQ9TvCHd+j/4TxGW8vgjiY2IpVNuUROBUDu8rKyX5
FzVWBBCGconK2EKH9Ekh/UoH5EVS5wYA127nqGmoH1QpKrBQpb6nyXSbm5VSfWRC
80FSq3mkJXDwPjH4lvK6/99QtZn3mqfNibS8e2AizLLVIGq5XFS3kuYZMwdQGMK5
egKufRGnTLsS6QxU56V+3c3C9co/QXoO8eKxTjQgVpbp8pCe0vLs9MNvWFrmVnz3
/dTY9dQgbTPzmrJKlTPTq3TUW3tks3Qn+5+j+9kk4rGPPt/ofo5+nzwPDhmupgKj
f8sWrCBaP48rDMUKkY2B8tmieEVIywSFhclOYqaTgMBTf9jQQQMl37b9KASi81y+
xT7h01uLDz2R0KPuIIyCv3xsiIDT/o2TbWVVqCzQeI0gvLsLjqIvZH8rycUGK8ec
bXtlZpUxH2tydfIAssm/jizpFZnz0Reo983C2wfArE+82U9BetwpGAboqrOkfiiS
O9FEdjYr85BOUWwaodbv4g46KvUemcz1la7reesl0qN2MBphFuGtiODMlkSJbTmB
mhWgOODSbf5EQxP81Hk5xbIeEzxtjzcjvyYNYIoPs2NoxRnoujYPevmUuWGZ+isb
t5e3sgoigiqn6Ca3+J4htdQoovY/IM2S3q7ZovahEbXRjUlaXSRp7KfOcKN/FGlY
T03YwtISP22zj8HmNIxgQWZ90K2uWGw81izqBRmwKg48IhRej+bOPG/qQ1D/WMP9
TvAt5kzeoN9bBBTPDpNMFgiPWi/4GHOoQX1JjCYgSDJZ+9Koq/v6AfVdI24ylGs8
nIu8h5DkNCOpy5WXhXIA7zzrHo3x+/fpaIzPRBKg7337J+/ELWJQFaWeIzARoxQk
AOBuJdBrfvGRZ+jERVkjXlmfUBQQ6B0Se7vawFjEAOzYTTzZTr1dn7g9ncnFChPW
4eyHhKnd56rM0FRWe2mejAad6kgKbLsZeUlukPj1katC0JoQsRXX+OD8Y3HodAki
yVkMnuO2iIumnuXStGAvnh9afQVUCD9lEOwZnbrEl/y5IeIvv3PluQxglFG4vBY+
4VRfYKnqLoEJ8OWbT3Y4ViYDahyAJiCitDJrzpNuQ9V2ZQVFTULtr/aNUfsVy7nQ
6JXdrGVwP3pFK2HUdL0bHCyx+R7ex6t5JPd6QNo5a+8nxOx5TR5BxueuEGCQSSWo
YtZsjallIrGm4CX8FMIB1JETCjzq/DSkYgngytuxZgboVp8KMfRmsudAeHDUuu6V
m26R24KDDIR5guB0zGKddiG+GybW8zDXu8AdgD1F0p28Q591f5oqmeGQe9dzAidA
G88HA4BRdWG30vzMY0ziFUH45Xu5d7YQZ4EpOQhKc0leog7Ec8b+ykgBVMm/zKIK
5Uv6aMYIS+AJpx0qEyaw6ZFMGMQ9KAiu2yNRPHOUh2W0G1rXUoL/y3kdToJqkvBa
T+gSQLwh9i7kerTLldBu5BHnPDdrmYwJk646pxjY3Ta5mx150/hCXwW4yrGTLePL
FYQFH7a9JnfKYaCstkjEaw==
`pragma protect end_protected

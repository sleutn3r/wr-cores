// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:45 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TBgwFgm1tKJwc6XmxEgWAfxOIK2c8OJAIBe2agtWRyDnmC3j7wo68dMJPDc+Jbjl
QVMG3j3H7TdobfTvzHY0uABJXZpSPywQMpytwvpq+aMQb9MgvBsa1KSkCMeu6lEb
0eupKO86jHC6iQeZFzoCpqMRGrbuVveo6LtOzO9/63Q=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21472)
1yLSsLZZKoUD6G/pN/uJxDxYYKpikCFgFGVn/pt/2jQ/6m2Gzg1s0svNwM6POQzX
/mmmrltgbn4Snp5KRD2h8em7dHp2sf1TYwqrR9KljBMWwXzaKZm2SG5N/Js29HBg
II1aMItrbiCvDEykhmdCtmC/EYVsK0mi/R/No/YOHTpbBrdt7mfke5E5Ae2AjA64
DSzQa+XfitgxQF22X6a3u2dxnVHSgwbGCDHsBhtvgs5xgDoetDFbX4E3YupJrfKj
is4y5wBZEizlEWVKJeAD5wZ1C69zKMS4WQ//7XgN5h1IIhG8+3rhIFFnA1+8qmpb
tVLMaRAaGTGnV7SaySinpmiaXPgXwZLUQ4T7WQ3FNMfUCoIQY0snbgETl4RKZl/a
zIzuun/hafMVqTvJ1tQGUmvelmr6FWqxaA+QrTu/+hFqmkzoSu4czCTfv00nbGMs
8B6Z8s7Yesy9bb2+PC5FaeR+Hk1qqkm4tKeuYDjVme8o+KyVHZjsOhpYKfCBaMWN
1BffHhxnz++1+k1SL72nzXyg1VWgrOYUSTrhKnRux0YhJy13O2t/Aai8jk1j5Vvi
y+Xt+TLUxRoBkzV6BgYKVjszAYWRhJO1fa6R6r60kAYUaInsUvZHm0A64hgLGrwG
XlCiGPUT8Ah9z2pdG+YTFW8Sh/BFADIxiGrwDyyoZr4BMrEPRjfk3ERaCiP0raR0
XCxVJG7aENfufdDDbBSASqaCTKyDoZOym73SxGB8lgtzdFd5bJ/5zUpRHkvA/ld9
NsIu1ZGlt3zb/afSTrpr21y29veHyiAKr7qRdC2uDw6+K4FN3PHaX8ZKX8gfzJf6
m0mgIpodmBlVXeDzZ81nEUuYz6W1m2ocC0PNmmjeZSZZapOtMJqV741ZUMkjgtLG
xQUplDnp4hCAYomv4bOQTb3xj2qd6YZgL5f0/PIw4oKAYEW5QTHUhoqGsQI3Q2wJ
nQrjJbSpveE8Mk+7W+d1DSXicOa2fKZY5lnLDMZCmLxrTjmVINjHE10IYtD0/8RS
qzWiNlP9osH+9sa7a2Xdygnh28rUSGtKNVPFIIug8AIXb7peVuaG0WzttITlwCer
mo8iUwGM8d1U46QGf6Aqky0I9gjSgjbmMulk1BsOawgfkbIovQ6QgQz/Jeej8ZMa
jHL68/bUTTuaTtjGdVemqVBIkbA4PfJruV9Y8ChfMCq7zl8BUsSWNRZSup28Efo2
I5CmkHCm38i7mrp1oHAM6xd/aKlQWTi56Uj9MEEzdvE23O/7SVGU9QmpYmBKop5t
kaRdKej3X/45MhisSKxiCRMirz8GavHta1VcdZvh2rUFEQvnoWtrQxkNjRoGRglu
VJYPHSiri7RstoqAk0mc2u3G1fDAs6mGUDhjV3ohHegrLGI1BkP+/ZZtry+liXFk
WCpiJ8kmjt+PFOsFwsVrD30A68Ag7wSROzsnALHKfUZtkuWjnPTDLVZUQY1zCw8M
uarnzzL9qgUiWvaeP8S3982mw+cJ64tsa1SOPpoFdHiCh4qGADsF3GKzLxLCXrr7
bV/Efjak01dV7K8hi4Q7dGVUoXwkJC7LBTNbiS9x2dZa/8jux9Z9nWxdmASBZi1e
KzJyL0dzrPezi9BaGBJguEcMhSc4AVM0GZCzHv9x9EzMwN8GloOU8rl4ZiIc7jGD
gd9WV/xLHHqF6Y9OedvXkOUMxGZJnBJXiD8/CL/s64tQxnXoRm88vOAPmRMDd0fz
tnVpep49JHnV8UxXXbvFRGCMN4XUR83n5tEk2gZYHGIscAzAgHTKbcuoDSwpN4MU
RkORD/scKMAHy2B+muDnYESi+OKiCFpb2mbuoCZOU2YALakSXbgHjmhxHYKBNNoL
eYZvE4YSC55ZXAssUni+loUPHQ7pSKuaPvDOAcRjgteFQGP4pIypo4eQQSbskjB8
Dk4Qo4W9e8qep1ZbquLeZCdhhGvUvK1JP2F/ZTj1sKhmjZGZjFHkaU3+k575XunL
9KjsTbe4SI+CMXas1BWWstl9l491G4nYSuMhF5HtjRlbsDynxWTOKirKVucAaraR
iHugz8bzck/GYMb8ELZ5huUxiJBnqDeQg3z2Dcfk3gLYZlHFxka5IBgiKwFUlBtG
a9FxbZ5+0U0F0VMnKFh3+r+EJ2Pv988j2hOmu5juvXVYxMQboP+DFqi1mY07E7f8
VJDdwy20Us641gjjoKQQVpt9FRy6b+D+ebW10t7c1Mk5VlQcYwId98RyFFeLQE8m
h4UZeyG3R7wViaZDALIQTiCXF2A5GqeZAE1wpEGudxDwN2YpWUxvmU34j/NDWo2k
7AlOQNxdQPYPnYtqncEH+WuQEiEnaheQHZ95UzaKNn4UbYwFCGTq0bRF6NividiW
FqLKyKiTMhGBhI4otcRO5QT0BLHH6ePv0FvOO2lmYgte0EtPhJb2jmAe4tTT3LhS
LGkkkFN09Omb4mqx3v1FyScR3IlKGSxje90D3fw8zDmc+UxXMc9K1sccbyepdYUd
0yRFjFCsXlVJPyE/RT6U5jzA2uPHDKgT6vJ3aFKl/BGDl6o5yXhcR9Zr/JxUdDVH
CwmHevQMc99sTXLRTWQNoaN7iKksM1xiiewEmadW1txQ1vikLvggpdnXMaWpVgy8
3gPjPXExt+rG3J7sg9f2ErZEYew5n7nReXJHASFSYjuAiiGigzWYysbj12tQtZqj
lJFRKMad/eH8VpAAbhMu6pz3L/HypryMl3t//y0UU09RrsgNAhYw/nongPLEb7Be
Au2xDWbNs7yIBGLNfX1beUf4JB9M4mHW8ahOy7fNYST92f0htd+5THB28JDljwDi
dDpgLkIYJYU1k44mxnFqBDF8c6JrkXrH4Z4ti2c5ER/OsGm3tlEZWpU5ED1IjnCA
ZjCgPehyGoSmaJppP0qIh9hMH/p3c8SiVJWXuEhW9FhiyKPSweyK8msZQMAiILF9
1o7Mse5V63h3hTQXPEssse3eaS/i4guGqyZc1PEaSjV6CYK/OM7jbnsTLCqhKgmJ
MjhOLBSOQJukajUqNrU86QJs/P2RDxzFIa5B2pqMH7hXZf7oVh0zwtnqaW2NodZh
SKPQaoEE3h2SbX/Ogm7LYPmTCwryak3uuRFU/VDouFFem4d8k6PAswp9H2XZ6HSS
3B3wK045dwG810VjIPjxL2lMEje08AXHwR+PzcstEv0+XhF9IE+9zdZ64g/prXsm
1G4PXblWaRFz4FKnd3t8xZazJn4WNtuYF7/4FId2TZZb8Xb63yjk8z1UCBtJrhQ/
eRm/vFpz3BwK93c8S4oX6cTzvb2Cpi8bsIb5llv03ZsLA1e8YqmYH2KmRyG12LW4
NecxwY5iXG2EwdsUtOJ+oFa5q91U0PZCN8W3zLBREPoe0HdSfyoySq2403EbwcOt
uewOOw0fEAvkQVjxL/nIfbEILgC17DHjjaLsCsvF7tlm+4TbZypSeZdWJHyXSvoP
onW13ezMcK5e1c6Sv1a/owZHPpikMeI2vzmopvkCq3jBjgkR1xWZsgKS8Ok9h9ka
vnh8eALwSZBt7D8JC3VX1PTb23EKb5roD9GJpt4Pq6c5eRIZse1/h/iPaVIAIrch
x+KOIUdmrPPB1CcGnBGRkhWPGc01rA6PinAS0qg3UKXsoZZLIh+Fe8YMrCqqvshW
PwH6O28lT6cxO+SXR/pfWWkyyBeVZYvVybfPWMMYbQ3iqVDrohOOJiLKCYdqMoLp
QvJgsNh1sZvAXeh4i0OOhtRO+O1MtyZXSdpn6KD7XMFTTOLv+y6gXkGlOgQfNW1z
I5ODwfrKppoZP1iGn+bW68O56qxd3S3PzB9+T4hZ42PEe6rZNe42vP2ziiFygxta
wavl9hJNm4J8LfpWPhUduZP94FOdfWdSIUFHcrPP0kHGnIOD/ovfoEMZuNmY4LYU
/UD07PA2jm66ca4FgYw5eUrXgoAOr1iBiFVwpawT2ER3qOmy/LR3dzglMAl8j2I+
W9qvfa+6e7yeAKwXp388o4N6YR2VcQRQ5rmP9n2v21TPoh0iQJJBe3AnII+s3gIu
RPRDGNMolHXQc11o1lYKeF38V3+jP+IW7Jf9TbyNiPCXaRF4/rSZIVialgxeQPpm
D2cuebD8y/tiLgpkwv2jU17lzpw2eejKTHs9XIaee7+AuJEsNHDjujGYxYsGAl1h
rVKYOWw+zNBJOpRpwL6T71Zb7tWx1iLe9siif4Z3jGxYIdz1SekN8oYm+2WKELRG
6VC1Bweh4kPBxzCbqzS4mpIHixsSeE+YJH71EUrEyELacKOodPua5by70SWu4sm5
TazRrg8Ix78lMtwkv7Lo6X3kWwqcIfugA7zcCEfSbF9kYXuKtB2znkPP4kpXZ0pg
COuQirn57tHWuGwjrz5xjHvMDyeLRHnxhSK47pVKb6kAWyzHAxi758gylqROqBca
5Gkcz1Rfv2be4QJ6ZAK4W6IlYa2iIDmHIxTXhFzZE4uqZwH6mevG93QbZt9guiFn
K/6DY9qkSi0UWnK1m0gWMs9dzIzHJqJUzgcGYucp5hClZ9D62qeMr1+GBOrSYfJs
0V2on25u0KusrBKmVp/xBR+i6y56Lk53mh7EqXmKE6a2ieFvYAIhyLZy07GrkIfK
1PfeHCKs/lQTvbx29sYNqQ9PKYtS+eHtRbCZ0yTG7Ho2xoAGVYVa4NlSJRok0oBb
MRdBG8qeW+9bnYvm63xPqTuawLJub0Bp2Xw8rCtNMRVZN5jCQuE/aDX4A7ACmg5z
KbPOUKK5OMjnEl0HyTTaa8xCpTNABj3HiaR7RHQQ5TBZ7L/F27/OEBH3cg4pf5ha
VBW7jL+SHniilnH69iKKQNtjqa6OPM7zYHsx2ZgHinCU+L7HR6evsBJjYL/xA6pd
6imuJL1czYpb4zP6eb1+w/tkDAIvR3VYu/B+SsbHq9F5LWLYhW7YAJAoxvLlSyT+
SmeqTNjVQsZvZoueq70Uc6lNXSwevLHsFjks5dMz0qpknB3wtXQbzQeFyWT71Vn8
1ggyMKx2EjkFZuJ1LCnVpKVZZml7pIwsS8jJUdjlObnp++ilA8FQZN+qw6qn4dqc
0rldwycwXE4RJL+k2CnlKcnAOj5tm+yY1ZPbXZM+qen6PDGOf5NrwZMRZWDx+9Zl
wbgALK3OMhCoKVATuTTrirWrg+QtLaz2OG7eoceKNPHg1HaDMqerI3+zSmzfD+AJ
eJ7y+zx5asb1qHjCes3yY/HrV3o5/vCQENJhaEAD105jKo09b8XPdkf/mM6G5dpZ
QGiq2sh5Pv+RRo0XPWwnPskTnEZzkysPnXV0eQWPAuaOobKarboLC6uyqp8iCsr1
pj/KWlIZ1jSu5bqZPB7Lg3c/UDBY6dQ/4INd7iI66rtyxmXdq9gHgukTv4cS5j45
0W4kCkht8CHo5uoI6giHHOisfETIFtfRG1h6UH4zDA4/jbkWiyqBPBMAn6WyP929
1bYIHaUkA9y743TC40R+0qosXo8q2NYlKoQQWBJiBD0JA8qjGY0H6Dmrm3rs3G6f
/L/Keu4Gh6yYa8LKnaemnodcTutZSO0JFVYnpF+iG+kk9gyJU++xh47StKwNi/Eh
4xX9Yipam9dSCWvZZVWTWwsdy8Wy+QVKo9cCfVDqM8e9J/grFg9v828arQQntH/t
79+0REjSgUb4g9wnbv0DAwDHAUQ+ZMsumjKVpaixRtjafulNTR3ithA/ku8OgCkP
w8H3URv19cNo7rFylJCDA7S15OCH4xyZQ21Z+OjgwVljouRfWt62LfVHfUcWgVlE
NtCIv0JmPYcY5uzC9IoWzctZWmxv8d8BLmd+1EictC05OudcpOcd3v9av1roFh1z
10+dL1LhT/42z2hJm5Ry5ttNuRdRfrKiAA5kYGEaBS6yFi0+Zh0l5KsOhgarNOCj
daG9jM55wX6jbsX0QVnoz23F8Br20hfW1Ng2r/Z3p67qijyvVAQfxrpd3ueL8IVa
GmDqC9nfx0PfnLvJTiAyurT826MCTnTy+GSOCx+wQan0ZlUaks/Q6X6th2VAIEXk
7NAS3NOKetr80F9SUlYc9W32phD9wBKDO+7XjaE9I6NPjhdlAZdpiXMI0wciPWDP
6ZtMoRwkjlDD2mG4AIDjYHr0hJk9yTjn6F91uZOrZVXaTJ87z4+CBosazQj+BLrh
IobkexNWIFSbm+FCH+gk9FNVJWoo1JN6P/ll2oSJLpK5qF7wCcz5Adf5UuC9VzPe
o6smUkAzgCx7bTCy8KZPMKXxrIpZCjyDv5B3wBpid9QmtqA2HWchSizQ5LL5OZol
+hfnk74tmNT+B9w6Nl9JNjlfeOPrfxLflHDCS8MOSNQuDuxwlBEhyrHthg6+0tlK
xw/7alOEksK0YYyqaB/re3IDNUWbjYAztUWAdIQFhCrb+WovqBWcUkzL/Uy8bA+k
rhEsrxLuyc/yzpQWViyM9K03bi+2dKBDRUEjellyQGx6Li6e9EYc8OGW2fjqvraj
fl3SejQpn/nE6PRCpypaFTV8nNYzZQC558jjymQ5LlCBg8SC8Ti+Cc7o1jPJdZ9z
aBvzs9Q07KQBW5ynrV2nszOeFzCD+1CVEdlsYHVrNvRQ78dQmdIQPugTfEbHvHES
ONLU9Sw2ywbCrUARP61DhtkYpUCBMCSVoZldTOF39/EPdAbAQov8NUSEG6FK+nsy
gA2lbdQpmwTUZkUAjmo+VzApE2dZMloWBYkv95kYDkvjhDAMMUvo90JedZvDOBzf
7LZai69M7TfwVISR6EfKdPNbKJDMqVBj+TUU3t4OdL6H4yyUjNgd72I7OLMynVHH
oMNFXXppsmgZVVO2izTwRc5NEO+JEoOw5LqUrk5ro1GuynJHpJfmKPUTZ5DdH+Gg
PgGxHDYw6ABdRSaBw8o3e6XQOgDqrAtWBAfqSfPb7Vuk9JXGE2+UYB5ApyOkxJ7j
eog+wHe5kJToR/mJFFsvOp9RFx3QcdUTXvLAm6JTehcH4UBJmCdE6AV53LaeT+3x
KIfw5uwPdqnlKL01zhqFYsrScl8nsb4VaEc4HoH2f0UUtXJOdAj+7TTmaGjakoOC
UcAbGcrYsEaIV+CO9D5eUo1IU2SugzEab0liam0HIe4QSsVSt4LfNC6MF2s1DWVK
qq12+Zb2tTK3aC/YsGo6W3p/nWiHsi0UCOVvucGav6DCT24B3HHmuqlG9P65w4Hy
TxWjPs2UaedL1CbpII+5Kvf/Rq6i2yNdefXncUpL6+MtFeiLKXWkX4RqWwfKi+rM
5fpKoyk5PT7iDTc2YqgWwvSBYmMGMSVv/dCq7MM9IZLVvEemYsOKpBRE2QibbApf
5+vmg0A4YRrtHlMO3Ri+SxKPxZ7vhwQcQTUezl4zwGiiQVZ+ppfLBmg/d3WWSZrN
IX5GEkh89o/LimS31ZAY8oCRZoPJIWctO7vAZGEQPZVRRKJ8uJFPIKQi8m7Mexaq
iaHUfj6ctlFn9tp+T5q3VWwbj56qOfZIZmC3Cb5mxNrsBPHWGKk9972WDJqFbWnB
afFouRfh5h/oGTQmRPOp1CfYRutJhdbxyXcZ1to522RZdIoIuPoouCxhJd0EYZZV
C75iYkVYDxmEQUNO4MGcDQr4LCMI5yYCCU5TITcuBYrKCK1VlihosiG7W0xfoMI4
fRbFzlVMDFwD7AcD+or9ifPfPi9IhumqGVh77Kb/Ns6Xj4MtMYL7xpEyK0IRI8nk
LlBkRj+ZjGtkHw29vmT7P1udn84WzvVIwhARx7kXaoS/M5ReBHUhhpoz/NFv5HPh
5YO1kDP13otT3WagQFy3rj3nBaVYCR0XM0D9sxsm9WYRRlrSsd8bCLm3biL8SrkW
38LV9pBp/OJs0S9KixpDdYEbPTLPOzB0HHEoUajQqzrSSSlA0a9THqlJFWOqj9vF
zMVe8Ol7FImyc11AHTAzkfkU0ONcBgq+f0cadQn36CZ49bZqxYd6V7Rn2q9JOB1p
1xfYUYUEVbira8bDQnET3iVtq1N+pOJSUzpHFChwl3jjGOMo1zbnVPINcYLw4K6N
jvr5lSafRYEnJULNxXWnW8aYcCX9QWPOHQpdIPyxbWPgNB/cZyFdGftpNzeXDi2u
wdEfxGXhY5B3RoQjdjHUn9HHFlll5TKu8kFLrq+/s+K/3B1tLvLLNHWOUUhFvr6c
/zv/B+Lk1MgkXdWp9UfQVEqoK8s9culCR8pGOmVSnDl2aBZ1yzLVDhhhNuLdq2fK
uS5kMDACK9g3Z8AyFUwC4az+coUfk4UFF8SUA2LU4QRqNfNZFa9YY7gUlGIckZrD
sk1CngO09jlVebDFZn4UkRbWaKKN53bHGgybbQ9plkCGwAaMsGJTfWn+7K7Fnyde
r9hMu/QTTFZFTZBHIPJnMtushL3KX8lYZrQExqhPcf9Xd3ssKZe6U6ThFWff/Mc0
JSdvQhvitUdRTWVkG5SusQDXiEeX8iYH/8P0bOweHL6cn/2COuyiV9jaUzxAdG/U
nPyJEjhiMQEDV+rwCQfdFb4mPEW+Mp601XXfik0nM1Ky3oE7DZRTe/jj3ipxJrBb
AbixiM3k/K0DQjVDKrj6cGxtMPOE/UflaIcR9NnMN31krmykLUWCGC1UU+eXfJU1
mEtqGAuOf9A72VnOZEcZQEB5vJ4mxWIXBQ+Y5cjdjxSJS79Vk13CNrr/ALjyTDFX
5cb33qDy3z4BEVzC604fnphq2QZaMAA6BB4LLvfFZ1LI5eVeb4PPvNCKA0E5P04i
VCEAnwn8k5Av2Vqw6j/JMyR8KEnnCJqqc7ompBTgeQkX8afg4YTf4lti2oH3/L09
fznk00B+xefYf+JepkjwB90WjVUaEeKtNFx9Tjqt/26VsvDvljyOpIkHNHzJtm80
qTl2pNr39hHnIdP0kXZIHe4EK9CC8PegEzp0DbyP5J60tKPSgTgYAkDwM7yw1Nys
6uCCgzOCdQ4l9BFjKhhkg8rG5TUD5kcx/KtA19RmUDzuuAwTMH3ziAYNyuc3xccI
uiuEzyXy+oEjXJxy3con5FHfyIw6E3s3UAWQSr4eeEyW5vfaW5hw55uclp3i4RYX
ZmyCulOmGSDhlAPwrsRfp9He6lDmffWtM16cEf5+0Ri1c/UKHyzE2H+CpKKmLnFv
1K81S/CsY4LXKk63vsawRhTkLKCuqLWHYse6bhUxI9VuGNggDukSrg8+tlKQmRFD
3mU2l19RBQZCFN0/8W64hOESvqsvHga68hSQv8jMJK6IZ9QsOLUzba8pTyQMK9wH
9+nuAx8lYVjGJCc1CRFY5p73l2Huxijr0/t+KZcC8WlWGTAQV5fZLt0QDXZApu7Y
p+MkO2h7CSNDGGtQ2tyS/hIufn5oiBdOiiGoi877tNxRBRZtCUiwxmRuQy15H+Cl
POWpbS1i6tRv5XsZxX82cHsqc85d/KOzH/t7foxlRxTU9FUVP4egJ+W6xzJv55Ao
9izGDWnxH3URF4rNeCEt7Gle6uEDeeIH8/FoNud6aQToddnbaggLvAv+Mjj3Kdh8
3Job+vnBCFl/HS3dZGkU0q2Q8GBTK47NrE9B2uWl2hokusvsWXmRR6NLrNHDvwmj
R3yxcd5rsZYqn66476bLMfkesY/7QraICVMAaSolPaEZP1/jSJ+tL2NJV0p/QWpb
GUL7tzIvbFbykQp2uJoH3Gc+vzx0Q+QcySP2fb5Z/0MrBxiEZ0WI3n03ZOgzcbbu
/9+kMu4wPEXJlRXV41K2rHBna+nG+PQUX0plLel2sTCehlhBfqoMOlJvm/SpXuRn
2VdWd+aApGtfFB0Bp3wXEwxcZULRiKuvCkSbiTh0pNPxwoS0eDhL58bPcK9/3PFB
PteQ98G1NoR4w3o4hwlmj0C/Is1PxJ9sbxWsFnpLuOdBv4t4FEONnjPNraGIkhmP
ORLOAkLeAO5+7IJ/UWu+y54QTzrXtS/mXd2cFRSVe4qKGNHqQOVJNxoqCWH7quIy
crbKJJ5wWEIwTsQxevOZGBSggj0+rhrD2k29mDVv6z2HfGVtcnHJFVu6iz4Bwsnm
MIec/HLUgCBg4HkRa5R2cXdR0Dra3ANxoxJxseFqxScRcO8wQYfpWUB7SYL1YuiP
syaiRkEfF0LzBMEy6gmmKDv1WJnMJ0VsAssJJ4pVrwvh4YKNItulwt9OzC9M7geZ
f9s7QSTErhF4E6ScnkWExXkyj7TOwQgRpfNP6TxiX0CkYNpeOyRvSBLne9ejLBeD
WabN4las1QddL38o/F/oGVnvOIjztVWkgYCUXNb79/bZAMiOzG6uWaoNMJUHi5BB
eTBOJYt443I806erBIwgg7Cf8ddsoHiGORAJ12k6SBBMtBGBqYohB/4mIqTrIe9a
HNOGoRYGPU7AJFjiawz2fgkphOI6JP+Rx2WHqL8fx7gIg7emdFDrJuk+ZXqc5nob
qiQefixZpcvQ5kWOwyEXjmnykAECW90JXZtPBV8doUVQVVtkqrWYpM0crj1Zz/Jg
A8evGo+ZpGtepV8217/Pbls30+9AFTtdEvs+WbjUT9fZtZOZ3SD1XN3/cqdYjH7S
csMCjYAX2NMsi+ptcoCrfGDm879DaTMoKg0uoz9wrCSYslKtAWnMMv8EFwz+Zbwi
OyXyDI2faTqJMX30mia4B6SgrDxIKDNguZUPpN3hMmQ093VFPURT86GaZXNwO9ES
v7EyzFRmnLAL5qpeF5dubQ/kGlK0TjI3AKyaEz1L6EJ+Plc7OYfRU5Mm2U0pcNcW
YQ36zB9a7e5xTUGNwa2/1Szc7D9mu5MP0/4l14GCAdUhi4J8xMlXs9ZFbmhd0os8
IqmGxUbGBnCF4dIQ4F4iLJ9/CDTyuZ9HcEndyIqdZvoy+ygAlmTFbA9KzixIw7a1
2qJKRZdEplzY1YbRPy4pg6bfxqVJQK3gVArSjfxjCtbLryhh3APVyRuqx02qmtOo
2Tnx+UDDXruMGro6HZ55Uq+ZkdY0ZDBIvjlz6x8LFzWZdwTD/U6O3W9l9QpBLNal
D8/Ukr3ltDzkqnRCE660pkYhw0bP3rBo1X65Xgi9e9xHkMJwkkP0FPUEtYJT8Q9r
WjTqBmOGDqESwoQ/Kl7XHjAUEzi8JUMhLxWy/YyP+6oSDsJi1mbsWlUvQQljAQGT
BzjXBLR39rpxk7wWEIfnXXzEZkhjcnhPOkV3pGcjd7RG8xRLCk5Z60uZzvxldIg1
qB006tKc3CizABWr/E1CFg+wgLBcxVsFt1S3Xgiijxb57wn6Pojz9OwPoz3PNWnR
Ads2m5CWeRgmoZqwsNpvN/L0DSt4VmexiDeaYDrobxZ2kL/Y63wiBeIyULbuODke
r2vuMzUPOpfYKme1ZJhX1jRuXzwQFU+W26MkXshdkIAS+gmu35Cr2PHBl5L4LOro
/16pN9zBA2mToOwk/cBxGiGLfYPsah7hBQWLwTxZYLDrQvdAaETWGUIZ0KJ/lp4r
85rj6ywE4j1YoFFtZ6V3XkSYa7xTNwWehzEKh83Se+BOK0qiFl+io7iOduSz/rwX
rtC4VbmHWljiWCYyeMVYZk1BiX1X9Yc4MDMwIwOMj7jSRs6u2z67DJjrLftDAs88
avjaByexWdquLlclmh9j8yYEocz8Hd8RvwfARAhEe1YqacvvVZJESZAwtmqj2cBj
Mr83Pk6srAqMr5Ln3gWs3VhBtVLaCSqy0+1lCweaRChACOM8zJ6+/h0jCJEPewbk
sjxlIHjyeFvBZvJEnfqA0KdaEMVyFQOfyMWuoN8+GspGl+rUhz3JcqR8mreq8jXB
NrGpieXMouR54iQ+VLI9IisioN3Hwrh63S6LMcdJ7klFZp6bimd6teEUXqkkwt8N
ti0EuWRrGw1RizH8Q3MEWmzUQ9GHZzO6RNaKrHMvieXKtx+LfA/mW7nsFrQQsJ0J
G9GR97HolZXHQG99dtm7VazoGoEfPYoNf1cIbO7aV53icO8TW65qSpbDmkpi0wq4
2um3kXuF9gDvuSZTAFxVg6p0t/SjS7R495xZKxxZfbA0/zG/yAJWJCG3y55HpbFu
VrGcAd4UI2/GGhrI8fhU2AgZk0vEAdPuWRJhE5/Fvx7A4TEmVt2apGK5RhjocmeB
Yoj9/GaR586qkCB8sBngBAiAO+hQMrdPJZlOX69yFzk9+W3Dg7+Omtb1hibVAg2D
TBuNfuEWyBf9K2krw3cBwAmHCEyWK+xZaA4pcaOV7vJnNkOtlBI/WLhDYbEVgCaz
37v9uG9dsxLGmKLVMajiRtS8lN7f+3VFD6tE917gozrYg9H93vYUyLu13X8eDaE5
dApqKYcIaF8q3lzvEQCzXzVnbJ90mcUZDFI2p78JbXtmXXQtJZswpiwRNMbjZEAr
ROHlZ63X34PCTrVhwXeNpQN+n6RT3q7ccWSyhaeZnF4ZP+9YAo7wkdaSGHdpx9Cw
yWXuA5QcdwkIfNwZJeizv5nUV/8JTi5hpZ3QNd5kN6iK9FU9zgBzSk4txM+5xDVw
RjMciHYnjyEzrfGfmnAqnA763VXK0Udrf0NoSY4nrLRue/KRnW1EbhRneYajK7TR
gwCBeGPQes6TF+Vp1L1jnIwN5c7Mb7b2fBK24wuF3zFIeWe+ZLmU4lrp3vipRoUw
H6QA2n5vERmd9dc4Pp8tuNQBGnq7TtqhQEW6GWMFks50XUkwP5x9FGr84mE2L7eJ
hyqz+VPgAsVSvYJqagM8T2z5gPW37IopcYYEH+M3PDQMcBPf0702u32utIlYA0Nu
rxG8Fo6Hv8wZOXQUvv9I4Y6u5Xr2c62wmtg4FQLBQkpQwLcNwxR5Z28Nbr1Q4ish
hC4VROdt/uD2CBCqzfN2bzZtenqdR/WKQoBy36MLTUagVD7qqMG8eCpJgrHdeM6Q
QPyFuphl0MiMEz+NwRA3U78bWy7lf5xq/gDHM5uUFKVNc5csq7UuG+auPB//8f4i
C41btxABp87tswUl4XycET56GTN7cb+2dDInmyUbGVnawZ2zEu3kNWyjaxCizR+l
0QjAZMCRGoSq42irdXDYB/wJrM2IDcsqV6r03FqRQr49pSexfH+U8TOjWm5JM5Zu
HeB4Y3DrCThWxd/ZlO4TbkMaOBwmsHnJW1UKSc3bbfqy40paMkienfsYsiQRbewj
ru+B9K4kyhmqp8JS28G0tObNnothOSkh0Q0cP9QYNtrpCVZcpiXhZ6Wr1GOGMi5r
TcTz6e3DD617UWF6wS/sQ6EZ+/32X9UY6BFxCYEdegofUzYUpEbCUs5jwzq8nteC
qQfkMGD5feIorNxn+mRIo4YGSshmop+D++hTqPQ8A8BBVH1LUGcNfrkxyv+8Dxuq
er0GbpJb0N97LAge2hzQtIsisCN7xSxvW4+BvRt+T+VeD6dEI2wQ65B2OTLcllPA
SU7LSeURIAkJuqmQwnth93p3D9rG/sc/7fREuUzM/NJfUS8KhMIm6FpIoFHgiTQI
c3Eyi/4qaZC8Ih2XcbwMtg8aiRYv2cfOuvPq5h0E8k/AUCdYelzs9Mv3BsbSenJu
fkfzeVOZSaFQKwN2jocfQGvlIi4u26O1OXCeNtPSwGZIdZ9ro5oIn7MAAekrYzic
KowpRlbcw7vCHuDpkgEIEN6ibXQoaTem9HvybMTlkWl8m8jiamrFRgCo3GwUrOfP
qJUwT5bmJWIUtf/zZpEuMiiG1NQMKPd8LBreihDtt6H8LDv0rnibGflbv9CIifgj
vZVdaypj5hGpglrZEL/4Q5DDA0oCIydScvn1MwFUs8Q8kPeuiLPJvvwWkTVVCpe7
5KkD/vTFOUVNlIKfJ6BEEIGmnRqfwemxi5gIKJ2I+xdNf0aGwQe4QEo3LUHsmUd7
E0JZGhF9BsTMGaBFFjsBG331aq8Fj9lfuAbSSWnuPTUDLgLwqxAMbmsqum80F26U
7vT0s4PxWqtiUbBzCmyq0oO5wdQjJb7tV6ffV3tNYldZvuipmI7W0OGNMol5Kc03
F19S3dDE5B/57Mmg9GvM6KaYFY9c+D3UTvpqxEk51vN4dbRiV+j5c/Syc7mVxZKW
9JOHIrpNSenNGsNzDPjCcX8coQvQh3gTHdC9cMeAHeb6uJs1JElxgGCBgrw+GJNS
LOGOyF9NHx3G2XpViNwwFb+kICnCqdfY0+9bhLoHQGRSV1jQQgEOVt1ldqPzdfJX
nM7sAIXZXmR+u6R3rsj6LG6K5SO+n4mKITvPIevKw663Bd90BkCZdcKas/reScwB
XpkPBOUy+Of/jYVp3w3YaD+X3VR+PBltZMOFdpUnluA2L/GuVaM6a1kfRLs+S2E1
THcUvEp+HXHEXYftYdRXn4sRb0hp0LMuEygZO7VmGlsg1CwgYaSbcSDDSFisCeKX
VhrpWG+LjUlQswSpBWA+ZjMhXTO8/+eg2naqGmzF/hi5pPdWjpRVEs96ce957Cit
au891wWQshl1zA5NxPS6jQVCyuH3fPw32OFN06cCQeHs2U3eXMMgzY7iMCaw6bJA
jEwbtncJxd0JY9V5gEVWFV5doNd5puXpe0yLpS5hEeZGB0M/yAaReNYvAu3a3Yuw
GbEV+JrZvfwOL6YsR43D24cRLI1c9/j37516HKIzf3owUjppUQhscjAmzJZEDi+Z
3w57w9rK6WdciR86Ca/6VNN59XqHyXCF0pShRWqljCnNYNyS1LMh6WbWXt3LPAcB
N7tEV81gMG5j3i9iRY+0ReD07kWh4omuN9SJgWlRFZ/NGzXGW6VgxKtAqxoAfrWk
X09kumtg/q9abJ6f6cGxvCu2NsvJZV6SlgBFRtNFOfakFeL1qILag+tmDTwuXHT9
wd0alVDxCntFu1APAODD76X0wK0bc6E3OlhRgUBX7NSJ7Tv/W7KyUYXKAgLjkMhY
zCZqpFf2g9P2bcUBIkDUPmPdAhku8Y7bRqF/aWjrydRHdgH1JB+xv/3hoQ4D58AI
Fm5eXzjDkelw+vBC2PCNzI/7PbbXs75dxWcnAUEJ/0SDNGaSvrU6va1OBwxqLTbH
AJxKpjXBoj2REOdri3hScl2sPbFS5ER6Q5aNzSsnUg+n26Zi2EBKVS0SB9IVaDWV
1ZUZkMIBX7S83FDFK72DNUR1Bl2Bo4N0OdtWO4Wd0PlhHJS6vwaD5udAvtvL0qqF
ZCUfuBWtogUJ7WA76EfhcTxQmpeLU/VNZQcLxJcYQ6h0JkoLQtkAbT3SoZ7wB8NT
Grq3KUglBzd5s0hd+uNL4pQSKdbvZo5s0QkwJXollup6KJ8F4kEMxKjXlVkGkvvV
abbGT0Z+2WAZFbYtYy2rSnj//nGLI+lO719RL1LNR4oTG3onZVI621wdAmnkSbA3
risgbEja3jPz+du9SCFmZ33SvFTiTgsA1SaIMV5VdfcAm9hnLj1YF5rAgrVsWf5i
p/ZqcPmhe0r1YCaSa/H/LPYYgo9RzPh/u7GJnOIWRUy3BaSfWhrrHR4xOt6id0+6
Lt0n6mb8/a1zDomp6VwwnKG8WiireKGivqZx7y7kCXe5/llDYro0OLvae8pMmLsB
gH+o7BNwRu5cYlnv2U6Puldzde6T2VotCDzB2d0m0Wc1qN6ZF8FeCsfeEKOVwETK
ni8uD1XYWBCdOJ5T4vPkxbauXxdebFHCBv89VECPqyrL28nx2DJnpqg4v4enuzOl
7EWIwwU/SEYzeZs55eGe/arAA0ThpJSIP+m8gE5mX5eeVAJ/LQxplKQxPnODPwRn
SZ/3S1WJWWAEvS2DF0YwpYSf5J7OPANyz3yUeWzwiwiCE7WpI/i1kwR01TbhbQ7b
qvtxup/9+fO84XOjgOV1ywQ9xHPcUVVqehuCbxZMo6LUpu5ag1Hj8ORgvSGURxSU
mkTVqacqURsdUTbBWENT9kK1q+ohb6BkDWE5li1eS7egnKQmbkY4ULnE1RJ7YRSN
IoxLGsWloqziP6r+6VSmU/D0sM8uAxmbtSFGOHSbKQPtRTsML/z0QCQT+iviJaWb
n+fumDL0xVNinRSZNTj7GCUeX6iG1cEG6vmzPb/qbrifN7d0OOw2g8oj6Vu2ndB2
pc38t+yNDW8dDVsbE+aicJB/uLhJwt2qrkkC2NZS38Hdh+5hdFMY+h8z0DlIMfaR
oP1odQW0WEYM4ObN09VQOfWuD/NgW2y1x+veu2N0gUY8MA5B6JH98H0yjJOi5KmS
xDbb0KAguJH2KiVaxhLVQQUrGHq4c7sK5SzV4TsHASkv5vfyJ3wWCLDF5PS3cwhd
rTvoSh3tgP5ECDu4Op4yFm7kf21t1j8wUl7zmcc6ehR1+1HupzOMgJ4LcnVjGJOU
U6hxd0mHd468OAjcA5skMOFSVndWvVOVfFMqQkSQAsA7VXFnwP+NTp3ZwH+wGBXU
eiW4gpyhtzWidFcL7LwHNcENs4nJPAgflUZDPRsXC9aVyhQUNXJFSRIfeDTCLFNN
ZZg3m7vhYpPpIl0NzY5SWYvKtF4odFyOaRP6rV0aKPcboOjCzt9+wSPMSFVrK0gB
gi5+tl2ERtIvaXZgruNxozp+fYNcjYTfOt9sWqwA44JJPjHA/7uKiRcpjHgozO2C
tMmAJ59OnodaQtUq0FvOP8GIH84xUYSy4KUqwQCh9RP5k2+XPW/+GdVNdIPlopOh
olVdQIPuizazLYJBnXdtMP7zSfbmokunyCajioQtEw7jXezVOSw1bho5CZ2SMHi0
M+FEbvS7OcBG58pLnnYbfwtJLnDjix4BgLr6IWYtBjv0njtW2+Yh/ttZ+8FVzdrJ
dOx74tENNlFYel+Oe7GmDVuh3A5kuaOiXYuQcnhjB385wO1i8SuLka1A4fLJPxtF
cKvxQPDsoWxKw2mGISjPfiTj3/OVSW4obNNimmw36Ve0zZbCMxYgwQRkasat75Xn
6h4vH+dlvTfPTphCM+zszz1c57PahgmhlKy9wYQYrTbnCzLjhrYfMxHWmk5RZOPi
jgLiNnosBK5tjWqCmX/Fh5xrlKz4BLwRuSBUXlmLZqdi9eZmv6keheqSP4ygr+Y8
zhQYMNtyYIvRxa8hSVlMIYI0A2R87VpufAH6DznCGL80BXLiZeKuThO+B/+yYO4A
nxi8h1n4w4l9H82h0xW9ZgO+OnuFFuxR9Pj79WC+hTJETTpwgYPse8Yx9zxMDq6R
b6koTydU4wOBhz0xOFcAs3iNISGz4Q0OE9TcdZ/yhzBma4ModGPmfeHOfLH8j2i5
zzugndArYOMh2PWEJnvPWHRzCb2XCAF9XVR+qmNdM5qVWKeki7CBuV5GULvLyCxR
OgkPmuDRryoTmg8yUn36KSOW7QM9jhzsXYi3yHwKytBO/L9gcOG9EQod3T7fUyPS
3I3WbiV1hqejwuvZQFPDA029l8xFHCFTfIrxlE9EJ60IvBcoo4iyFLU0eRstKOK8
UpxHVLVIr4znuw3LmoKZw1CH5ZzAWNzsv7iGQnhWAWelDAtBX8SavZQxM/Xfqoe6
EJFrSNfR5X3kcd09jwx2v0nqVo8WwbXdDGLM8PD7hbSjiHxpNxf5a745hXa5Rg9+
lA6RvrbhqIZHsx2uc8B4FExmHZ7NKAhjHAZ9RQuW8Xp0PoTa4+jzAvPx6+IjLy5y
AgdJqNlMUKanVmFyc+jOiZ+/YRhYDNyMHZoV3faApvR+e3ysQmL6OZk2Yb1jTMH/
vRuFt5/qFX0LJ0muH/Qy8jnGansQB+8tEkDZM7ZwGVd+mQ68BC81HVNlCSDFBdfw
hkvyQkXWutaTZMgNCDm9iOSI+MAvU1q1Q1YSjdlea/E2Bi9r+4oNFdn8ybdwhsm/
ah/OWLznAXESrBgE2CO6m0mYuXOs4ymbRP+Qodc5HF4Q+l/+cy32MKZNPJxzhYNq
UPzyGm5F82JnBfg0OB7xmWQSb1s5hlf87UGR1hTn9bZQ99Mi3F5XJ9lX4/b/2gcC
zMO3cuuK0rBn2/SHUK2txdNDN0h334U6JS2O5bIzQUYcB0fDrr1qfiHZ1Lu4Ei74
ifTL7aAMz4tUzVdFQZO2g1hi3SREPPnMcJXBrv56VpSC8ZlWkHViOJ4iZEQ4+H5N
pTOnkClDqQhLwT/fHYzXzR5UL2DKs1s8YcKOql1ZDu7ZLCV6PA7oPYOYo2I8k9mp
jkeUSBZ1p2aIjVSJbs9xg3rzM+RlE762nMSrPmBydlRDwajsxRwZ8O1evOWhgScF
rO5o2Qa4GT8kQyFeaMZYV7IdHbrgMZ2rd3DhcZnKGfs0SOirYSj1NVfyD7VBNthi
O8N1qrmuEypx8I/l4Af9kLVua+d9BZHO7cMF+wv369qyXqBoriNTKkOGFNga2ZX+
+9l4QpkEobluhRLBB2zRkor7iHY9JEjpRnujbs5yGNQPlifKNoLnaL2uFiND7UYR
tbtXROUky15FFljh9ea/3bC90IMDc5pwD9tUn2wac9/6O1bgVyArlMLQtYblHzXG
Awo8g1feeeZGHvm+Ers4K41zu+r4uMB73wkT2YuiwrCPQaKK94OizMlbgaP/GQyA
3vg+B26Mam0zbcr2CoTneJUE9uRLsJim8/4ELSiLK5rykxPmJMafNDZqjRcUtKeQ
eXeo5IFsLTRZPJT08jkmtpB9MjWWV7Fos1cii4cfyv4Xty3yYr+Mkno1TWC9Uz1M
06fBP5DLZz82Nx+hehH+HyWi00uKHJ0rZmID6sJANsMEWCxzyMryNw0Bucxl11KB
Edb6J0fj2x9IUMrphR0OsE5DNTUIXr/OXKWVVU8CQXE3vvOytY5dnYYxTfN6brhf
cPR2JEbyVi2JN4QH0BtlJa71CdfIxEOueNY8SEpcMDDCU2ik10/T3de7ZhuZIUzQ
QjvXn07Xjbx6lB/5a7euzX4eyAEWy5hZiX/X12LC29Osx6b87Xk6iYWRVhoLBojc
KE0dHMwTZYLQAqoMAWW93PiuaSOFuALZOQeBgScRDFHWB3/FumrkcsQVCAZhPhqE
EUU2q7KNyrqO7R6BzsWaRLF3pMTJ4VOKnZ1vjCGj3CK/B+7IwIgshvMWba3PhoN3
xxcQxkWhdYvh5VzZKBp3rfsrsOwA3cOVgc5foYYOdHnHUgNYqsjHsHAIwmMkiHf4
bFJNHZo5sUFVYGdZ1fiMBYfuAubTzrG21sQyzf1REJFfzg00PjvxpY/sIQLZbfJm
ey97zSo6f0LGT/8v9Z6r/oLfFsPVl9RZytvZfI3xdJ3+5tAk7mEVie/tK+Kn3iKH
fKRf3nx/x09Ag3Pm6PymMJ6JoFjM8XGqwB0bQt5ETHtPinuzK64EIqkL5vfHdKX3
ETy12RO3QGT8kgxlHgmyy91gYN03M4qe21vWZ2plARAoXK3dsiYwpCA63L1p4FlL
3tSCr/Nq74qA9Xq9r9TkTS7mD4Xrb9F5JkHgkfnehwok9r1ibe8kWSh9OwnNFl/3
Gm0pnkdCAVFoZw7Y4mZUU8Or+M/0ePN2ohaj/oMLu5aAtgZN2F/7yL/R91/yL8Yi
Z59wqBoLuM+VO/1ynuAZYSy8w0aPm+/mq2EtM0Tvfrhpvonaf3W5cO/KOr+Zrqmd
aqftSXb5JvKmMlZNbyryCGvSkQKnfYEWatCAfXOsPzFD/jbqaM+NIVlhV9MBbYMP
LsyLpwKInu/MKKwqu9NcUtpHtzeMFQsT9j8dv+q+gbXSSEwmxnWXFjGS5qcrIBw2
LePPm4skIxqs06sp7ZUQ0+Aywb6rt3CkVc0CkKrAaIlYDHKgBsxQda8a6jmt6DY2
OVzAT0dhAOB8IlHjhxFgWP29Wy1uuk7Elp1fzBfvV1lN9vtI5UXmpSskJJalrA6L
iZcGL6qQtueW5gpqz7NIG0jy7qozfdcw+oCiAJFfPZMv3P8smMUmUGjytV0K0CkC
TJF69NX49+5c3t/RTpEpyFh2TSqkBxEiRURJlftOpoPPL6YEguXuNJJq4pQ5S1ye
H1jzQ9wvsXpLK05tUIqWRroqUHLdUIHMc6yX11xv5rDqA+MQh2dEUHGOr2EuNapX
cL/rj2Ty/93mkdK/AnI/bZRdOJqY9+O2nePGdWV0+3sEXl3BlcCnidWN7qhyIZF+
+bLreu1M2A5ka3xMkPbxwmvu3iTfOrmy4lM1suE70qPJA6krCutTYF01Sk9TcD1w
aDbq7LCHAlg2N6YMv1YZyeIZ6OtB3M5pocTkiREL7d3CUA8JED+Z03dGA7F+SyHC
ZibIf3FeJwTMYCVt2YIbuZC5ycivImiS8fNKlkVSTcyrNp7Qz8GMRDqX7NAenYXV
IBG1U1lWMeah7fG9D3lLsROLRG8865isbM1PD1/1reHiC7M0k+PJUxD39rOfiYWv
Pl0JQ5RkZSJe1OPaQEWGOLDV7nZ3bGKaTPUR+xrnStalx7bJZH8xGxYyiooWwpJr
DJlJSOe0V6y2ADCxz9OgY8q9BwUKb3PR92ItxHYXotuXaHHOCJNKfn2A2sYKhvtR
CiL3ioq0lruIIHTf0ghQ6Hi5OapS0gomRNwsT7bcVfQZZMXpqspVEiz4Uu/Y3caA
Ux4iNSwoh1vSc6UmGvSRw0XXq/agm2Qih27Jf0kW2l/5CgVBzuM+Q3O9OXF3TgcY
vJW50UzQKjWCU36I72Qf1k1cKnzny0P8TM2f6mtwNH/OpChW6BsczvQKIAwbuZV0
iTeRd5ksXB34Sx3oGJfWTmId5Xt2om3bZremTIq8Z9W0F5hcbggHuh5dUt0ictSs
bAVbQ3/O0D2uaYozNB4FpXFE3NMdvtap8BFbxrKDx6+ieFt+Y/qUIaZ6MWEbvx4A
rcJ6iz8IH2TJVvJqp5AxG121xHF6RROomR9j1gwPmtQn8KuDwMi0GSO0kEjSDdBU
GU2WpLn4xXqNsjn4jbdv1kCmzO24OdICKaZmvnldyyGhkX9wt/z8k7KzByPbeGBq
ICtQNb5OJyxKEl5hyCr5a3A3g1s/cj7s1D15gxqb7kkIdl3+YvxVIsZ8n2NqjPTH
DIAlSp08r9MymZeRw4vvRoC3vizBX/McKz/F/J37n2C1wEHPgwBTwoI8aoQ/Xfdp
AhgjXC4L1lyTkB+/CPaz4UL0wzQByF6AX2FLNbQ3I3v83FwkqE18V1u5HukkzzdC
+sAz4qG62aVzH34a3C1mMffEvgKl+2Z82a5t+lJoe95L/XLjae2EouP2r5j2kd5B
9KugxLftoZbzZzY/TWkZDFajcYJ/XT+BJ1huFO9HlCCVbniSOguk2+E6JGjkUREI
wyHafrDYrwl8T5nB5moI5hRFfyZMULobKiu3smG6CZ8MC8E71fzyGHEe/itOcsAv
+dhj2pVnFEGf8txmTrttL8EzvhpC74QyIdwcGxCo2dgru6cz3TkKh2AuYH0kpvSs
YoL3wVffF/21AB6+cOOXNf3v9Hz+dGm+MR/dz9uQ0WhUTKMQwJKKNfX8BqYVasaN
B3si0KWd5RBdOYHytNJmutuiJ7ZwbT8s05Y6+RruWBiEXtAsmEE34AyrxWfrk7eW
Chl1GLKYukZrCaR3Xie5VIlw/q7Vn+4j6T7xzuyHxyBtUn9TpyEnqXQdjmWL0Z4k
iN5RunpmFC5kGMzg0S2PbbE4cyVgO15qZ0C56e7fclBd4I9JKSdojUmBkS9BU5N4
jqxghnzKik/1WV9hfVq+pHli+905VvUEuzwKpn5ERh6IKvfhnziX5uz3JBvwnjkV
D2B6uI4b6SyXMgXKsvwQY4MSHrj0f75PWdYciA1C/BTxEW2Gcfe3LkI8q9pUKTV1
FLWIEqHUiJofBUur3djy8tPN3KdhRgXOXraMky583BnwmMul8IjZbgAdlOWYM/RU
ENY8UyLz12W9A64oqsGMQX6cubgTU/AENuoaobdmgo0tH8JP22ox0hgK7jRkR+k6
INuKk29l/gAcl9odlND7FbBv2wgPgPi6GiYgtk+BWacXEAvVxbupmEPHeOBJ34/8
S8/H2XkxtISYR1qimR16dMHW8L376AhQubJse9UmWMY7G/+uQ7HhWiWZCWxvbJeL
iSp3u1j0jQEUKTONLLSwK1aw310S2SLDgvBmklH/dHwTdmSedCTMXlpJ3gOtsjes
LqRVh0wcHZbX1+YnLbieGplMa3BbwhZ3DoIkPZ3Cv9Gwc5sFDk9a05MP+Rs5WKV2
8IquCxGeApKQPWgHuu1ELBh57sd7dZMjXd/hU6SBinLp/zqkjll91a51nz+ye0Z4
21ldSglKrwtZjO4dTzsNjrTX5JA29GHtA2s70mobabIJw3CNsEcJtC/XFhKdGMpL
3RFBUY5M1ESVvCeupe8fgnb/8FanRiH4zukB8sTiMzKSGn9tAaseAV8WdDxoWc+H
HX77+3Tzlfd4lcjGjjyJtj/3hpQSUJ4CDvSqRg6jRFpsUZ0+4QR5743AZmX+FXgA
0Ha4RfYopR07PSUBoD9mbPIw8Sw7rX3G7O+GEI7K9pk9DLASzs2Gn/Nlhq5rwKqT
/Z+fjBw805p/GVHN6IRX/4bc/tFiqzNWS/Hg1+6Sol538Kk5dqRksOdLgVNhv/2V
4jGljxFSr4nt/a2Pfa+H/qtxgpH6F71MuC38BTriTlVb65QIGB8Fute757ezT6AA
nZuXvgHj892JSMpB1XoxnR9K3yxnxMamnRiD6tmXZ3RNsV4Xw1F+qR30RdZW18yl
catExrvNNrpyFqgTGJCIQaCSknc6ZjDoVN6pognNlcjAtgx7v3Zngy4mSggVwBj/
H3L4pzngYMP7xGDf6pOVNpjV65qtegKBJ3pvfmDBSd4rGjhtQXWgYhk5YP2Mhdeh
FSALYFISYpPlt0twTdV5F21LTihvz2IT1Y31p56IGeJDd+euy7OVgc/GRfWpBCod
5CknajwQLom2qW5gYHl1Q9I1AP9k4M23hvGJgDH5dmTXcSliKfVQQPODgRgDIntM
hDOXr4yUQadJJP9V5ZC7kELTyPDZp0qUcqSk6IpYl/7i7GKtbyw3Hy2q7YKZgred
GQ/d4qRSmlEdVKpW7XCHyQYM+zB9FP75gsWFOvgerJJxmthHjzk3+BqaO+TvoYAY
CNZ5cDSkAJMMMrkQQ1tQfPTbzQf49BfWDVcVI7vcRrTuEbj9MjkwQELSxMfEQYvB
zyfSz/9NUX0Ui7nJWvh4rwKRywc9pPlFUfFP8y4MquveuYvUsIVcRm9ceuqEihvH
8JEtjGIGJWZHeIdLx9DGT5kAky4lTvfhbEKtYRg2h7FkTS+0asgJPQtXyCrHGAB0
M5L+gqYc4mVA4qHIVbz8Iq6epLHTKxQMvTz0zkQB9irPAwuQpM6oKkNvgkAZBneb
lO/70B7HZJjca3di0MGXShcvhS6CHNPPgH7yUL3n0QEza/KfE/bZM/qKW/H0onLc
82sctOw5Qhmy92z0UJ+jwKkQfX9G/UlkXce4PMI9fIJoAGX3O8IyKwBVV1mDXzGW
11Qp9rNvcS33Mi6J8fzDCLNT0hccQtoaGoc+UQuKYsT32CcrRYrb1M347IGvSfI5
2PKSNhl9yZYX8SRI71bg5+b3I74idoeXzXjWeaaC0UDDAycCCP1ADaO9fPo0RG6Q
F96DMEhP6hSWagpzyfSe0hA+Dja5miB3WrCq0AM6bc019KeBGblTTPlheF340nMe
RKbKnDFfuM9Smn0KJNEHBIPF7DiVT3Jzj4WWIGSaUoHZQW5OOVJY2A7qz+g9jUkt
HuyP03+f0ZcrAUAPMx5vNJ4am3iAEnDeIBUiZ/n1VVVrQ75rueeTIM6tbLK5lNiM
CJNCCTLShIOuJrVqQNgalFKd33dG57KsaZFN6NmhLRUZr2uQQb5/lUWo39cKLJxN
pwFi6AqEf9oAeV+vtzM8SVS2eIYE8nwaQjr3Ja+h4UpxjO91uqjNwlRcD+hVAvtY
5Mt2pCx763IX9JXh5ZZSKebDIznbA273s3SYfrmQJzi8I7koy2eyzxOqOc1QqqxP
2gXNnXPUKySz1SvaJIEzp3PXLDhuruUMAw7McI0m8cZ58M455K51Qzr8ccXI8Feo
WPJ1N22WeEArMKXO69bM++xFwGyjsxM7NqtIzeAMg+lAi//7ObQtTabvDMCOfbT3
rXV+FSAB4NtjLVTMLj5lHEWJkrmihv6rQLKTbkBTdN0LVXezqw2YNusn99cl1Fhk
kOA27EmarST++H3zM7ttfkJiMT63W0bMfK9fev3rgjpWMOqxI72qAS1mFhoNb0v9
KMMaJfRMuuD6g7TJitIgfxN+T2kvBC6r2Lenb7FQoK5sp2DqS9L6nGWmUdYSlaSq
qRxyqKH7BVqV0VuI4gwGGZx2oaeYnroyI9RwGBCe9hesjw7SlYq651GCLDv5ERck
CYEVw/Ik8wpZ7rKU1gel6HCUhrl/chF+ZxhTdDgdvOnhD3+M3qgdt/+F7k359kry
1u+KezJ4vurArKmCCNS7qMjHiWR5rmTKF6JRUbSOKbviye2SU/cBgPvDr7lzhpNS
QxNqYZB7A5SPyRgj+ie/6YduoLVZK66T2LhonLv3eryuQqFtDOur6g9xF0Ri4x1H
4nCz9CNFJAH/eBbIrsZfn2pFkzyCemE+p9y1dWa4YZG8Vm3w9ukMLfnH9hpdDCSQ
qFDfGHpyYgaElPO7TcZVJnnD+SGIA6s8dwnqjAZBpxOzRTIl7PGd9YbWam6h4NAb
gRs2cM/75fprl9F6DzSl14T9iz7maBg+vtW0NkWaY5KXBoaOs6+b8AjuBoa1hzXh
c4HfUTN1Sq/jqZVeUIA29IEMEsdeO+unTNk7dGTRUcVdyLziEya4rN12dZN4R60l
BPkuj275/A6j/Scn/mHScWTHdqlngJULj7ByUejWOAJy5EloFoLoPN0yiRLvtvRw
dJyfUbn/B1o5njDVJYKVcvR9tKzMJ0aKCWTH49mbFgmZQnZpazhD4AmstK4NdDvo
aIjR2Iw89ciarxdOzy4DPsPWEVvibFOqBoqcGfZMKkhDsJZPnpaFtIEvLUh3hZnT
ataIlmJs5keEoe6VtYbHT8oHpyNC8fS61lEioaeXcTYeZIDi9x8j+EKoiAfp7q3F
nFMO1KwWMhJhNNpPbB7/vXPegjCZxSfRJTyh1Id7WzMJvEYZnmxGgfl0Bszluwl8
HVGpFQ23R7W0y2D//5fgbwsznNgjnKNoq36Ix8ELb2vBMACW1nzniTT6WpxtngtG
ucwZQEbKeO1w3KBxXfVl3zO1IXvppmZ1CABYlNS7OxlFwxZ1xHoEqnU8zO/fUUkP
+HQMT3QHnvlIk4x8VYdSt4+SSljjONsswcg/XRE5PXwiDZjRi9qF4+nAnIK09prp
14/nbJ3da8zyueEKbfFTb+rEwvajgkIK0Zfy9krzeq3V3vai0h+hRpEzugKIuDPO
0M0LF3T2wOEjqfSq7GPfNbUunfMQ2M3QtadSdGAQSXoOYkiq8qzyAkg8mJU042kK
BL/lZctNko7xfWkRb9U94UB8wqNZkDNTeVPhBgFN+l52M/aa4zBvd7M1fYZeeeaJ
wIW2yLhkf++TRFEjteLCaTFF+Ju4SamMWRo4FqML965FYDS1Hxef/f9FHTGZ1r72
sYgEL5riJpt41iLHA+F0OOmhaCdJojwP/FmjmEkKVnQw+iMNexTtLG6HWkaNgUIf
F+shf1Ez4qvNriB/h2O8FAA8k8VSi/afafnZ5G57EQ3BQoTKSw2/PwmuBCFOMSbY
W+Mi/D2BMdZ81PXmffMMCgAYWVscKQLeU+1+/QF7gg1yZMzvwcALDcnsUx5Z0jPy
v5onVvNg8+Oa/mxUBE4EXjrgWgdHykF5POYWNmoFwxQBBTaBp5OMCRVUI4OYDXXa
kqGD0ftYv/y8h8STw8lzIryzGfRlWnP3A2k4y+rugT3pwEc06JGf/PjZnbB6wPIo
gykiEr+q+H7IsluzI2BdpjrYfKZp/g3v8y3OkPXT7GhDZzw1/CZWSafBDeqBclk6
+Ox+3wYRXNuwXmVsz+MU1dKqi+pAfSOgnZq/+lY8CjwlmoZ/AnYgjUXMWo7gaVVQ
VCrIwGxXRLF0Q5SJTCdbQcoLetme6RmukQY54M0NCir22/hmHSTc7DOse1zJrDwp
jLDNbcoJlqYfboVpNn5Dj1VvKU+r558aduwNNLkG9/g5Nw5MMEPgTmfnpp/Fjnn6
5wrfKXgJKMi0h17/vn6ML0CZMZpWUuGsuSdBjIbvLPds/3Fce4ymftka4X14TC9o
qd85xV5oTyDuNsANs9wY+nYh2W0nR6Z+eRILXPnfrfyIKH8K+bAFTm4WCPrvWbmP
s1VwYWN6CgVFlt9DMBRpcqYh0pAJAIab1iGlL+h2VE4dX0l07owNAmbCaQ9krrpS
LR+YPDQVrn/5XxOLNbqIOkcyctyhZSJu6qp6rSuJ8dQSma82d1OaLjt6tkMbW5jH
/e2q4gkCSQ0SviG+F/uPpYljNx6+yCz3jnlQP6d2IpNiYmFHOB13VZwYJkLur2gN
t/jeD7SNrH5Pfns0sSrGQc5lArAtXzFtZDosMa99JI/3qzgPMJqLwyQbtxIoEmOQ
slNFh8cXOUUAHdXU/4Be63S9sK/lUY+IzENRa53yAQvhuZILiNkCh3/4IhXHXQqa
pj7R9ewybYfAserrMgs/oZZnBDtIk0IK/SKaiPd6ZPL4Z5eglqcjXCi8mVYxXbL5
aDYj99ygoxsIz1Fvv1omKKd/EGnj5TtcIJ5dTdfltQuHtQvq8qkjmZMtFOxGrz4e
AhaaEtZLqFn+y47d7PeHpQuweittdU22D07kKhyxZYv/37tbYmKPN1fVUHqd3jie
g1Tla3gY68K5wuXqxlfisI/9QArq2MWDMY4/jvdVYmx2wpx98jnLTGk33bDGRt29
uEmd1DGaEOO7Jh5xO5CvlKfr5FFkQhU1JBRb6mhXcliXQzx08G2zkpRJ49wPaDD7
bqxlzbqOJF+eZDGb26cs4d+88+A5ZpNNiGjYqYURhyKLn3uK4x1S3z9R33y40Tz/
KpOmSoJ4Zc8pVrHQ4bvEeaWDgoGuAGyesQBajzzdJWctowQHQaFalxTM9gX4neoO
qZi1lUtDG4YwSZT7XvsOaF5koV2vSv/7N8v4TAdlqmLxTB0peNBxhxnuDEQ7SzXt
bge6RJu+GSR8rf0zZVo3cOSE8FZG16Ey/USCl7tDyGYbtjKAOpELUJfGdbG4znvV
6Z4xmkdUypnRnfoJSOA4qkGGECSH+oQIdkISy5hKucdtgG/eSZR1e7kNdUc4OKGX
LuomJGuWssTW9o/t14Wba4IUls6ZNibr/EJW9kpkYeT9G1o1rViNmAxwSetsGbyY
0NG9dppHQcOrr0PeFo/xMtT4q5ZPmeKlN9splrQgir4YGf1+IChRlH2X4hn80tyH
Sn8hRn0nZL36Ve5YHl1CWbT1j8g9y3grqGYKF5wCfdokfDQqjHnlD45ZdFL76ISa
5qYtQBQhO/XISbkmEkGaUvH/kHkdnHxSirPust2V6/PohOGquCdY+ijevXgUDZOQ
M572KO+R0dMljWlU7XyyAXwKflL32wY1v/3xOWWC2VES6SaizRv62XO+s5hAi/h4
28hQjI7JkqSj8PaTLM1rGy/g4f1Ue14fIEMLY0KQbjf/EEOzzP9ChIbdef34K7B8
A0A0FaX6bW2GNdx59I9JtlEcPMbkFf1gh16N/SbJhuHG9lDEMBuGO8DGBUuM3YwL
RXyOXnCq5/qMUDcnbak5XUTdDHen8jYEgahiJFx+P6YOrxu/eflOokulZgLtCS5p
K2YW4YC3Pw1xK9X8CmxHp9S8yI4V0rvpf9jX3Ygk73xv0ULlGNA2aRfp5Nl4yVTL
PexFz7oi7nO+0EWNzmud251ecqzLfX5PcG2Y0DQSn7Ls26wREvIGya9K8Tbdd/FX
LeuO9S6k7FvFMAG1bWsXDoIcF3xHv3U4eBF1kc1727v64nukDIQ8YJ8d0TMmVR8M
WatepK2UoPhL5hFkSKejCVtJvJb+i7TMnCAqjyWGy2eW+y2N3f53T0SkhN6E0BRJ
1Hk3DXI9ujB3jhEpX3ncI57mPmCHSjZpVs01coYbCk05GbO8Z73pR3f3jJDB40pO
Z708qG+ggwX3yXa4R+sgmcivkuhwrBmBnlQzFFrwZaoI+t/bihw6hn80WXo3FeCr
NoEtYmX7iOXAFCIUvAKHyshvW0y/vXfNfYMI5t6pJ71YMzDfyN4+sSddmWoN6qoZ
SCk2LOHGvcCqTqVhWHsOyIvHqvQjMe6r+eOUPuGJkLQuOhPfopvX54JJR5h2wgkI
/mUGdIwoi2aV93PNguHJB+JEdwE4xB6QOD/qNFrEqIFLGkQ/58mIat0XbFPYSXyk
YyFE/+AExgQ/FTkglTnFnHjaTofPRkH/+9C8w6QKnBqbvpD5/i0Bc3p0yDzTcbIx
gZXOrgo78IYmbcl8ItD9IEdLfR7r+UbYy6IMccyfXzsRMzqyWSZrmO1C3UGsv9Bk
WZd2XzNLFIVfMDSY9sp4wsa54rm/nW5v/0KYNB3YrncwRsPvJCXNW1Dgjl0o4dFs
y4kSqDupb5F2MckP4t5lJ5LV4GbbB4Alh6HRiHRS9nZJjvOFsmy9hRVpu5uwv2HC
he5NbJ2bT08VmtTl6+hJDkwvCH6G03Fs4Wxq10JteOq1h5T8EB+vam4dEKT9Gkxk
UE7K/fQarK4D3aowNXmY5+2aZrXsUDYI+xuBGdEe0wOst+oH/H+yuasc+HxVElKx
IcGij19GPjXF1iR6DDvKKj4xYLNR9qcKKJ+YeG7VqMqH4mucmx7IjcaAsLsyJLi+
BilSllTzoNOCrvdDj4Q9yMLPEJNdxJ8Xf40CIzUqqr5X/qkKaF/6QjAL8oKEJ9Wu
qMrMD7Ncv/TaYida57sqfA==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BPtkWfzQGbh6s6fZXO1ozzYOWbToo9bfVIBFjpDujwojbna0gRzZMCFAocjq468Z
+eKyVK8df2acXDtnSDlYTEyvt8hFE+qctGv70isLsZ0zF/uW19rEPy+sU0U+93GO
X1TvEUgnXtKUmwy4bYqDpWjAfIdbFZ2dvVlReyBuApE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2240)
FhWvMhCIsayjikEFnSpu6I/PkBy1js3kN/opt0jnmR0irDbhWTEb3Yf9Wh6JSRoA
gDw3d6blk+n47dF1QmW2PYM3M4wSLJQXOIKFhxHTWyB3I9g6/hBNxKSgFNOr8Lvl
gFuyyacTQGsZBN3T4K8LCBA9p7sR2+IApF4fzI6MtPwg7l7FaIOWuknI61ynDKdC
RI9clQ0OecsipAWpVLpzTav49oiSAaptx+oNK5xbGTR6fiR1PE8FdPkHbSlG+/jJ
ZzEpVT3vwkdh/Bt7osJUFtBzmg0Ft1brHHKBEr7dOl+Q71qAuu0I7o+2tIyikla1
mXDwG6VSfL2n1V95lSwGGND47OAdzVGVyMECB28MWucP6AUeB3d5qJdclodYvV0E
E4IyuOcl7hPKtCD7VKc9HJLDxVzj1wcgK5PCvCVv7nUrtDTjIkj51tKG/jfkkbxv
y8iyJgZgu+hmwiTADXlM5aEYK5ky2Qni4hN/OWrMMZ6oSPFs3VQAMcwNbrRjETz1
gIyPg5Tt2r1/hCEcPkzIE8vd2QYd/FX7GFZnaC/IkyDB+/8+f3Ucq6W0MoSFr4HW
qCeFDEng8i6jAOtNT3Mv/XYeMctIrpKX0p+i26pko3zrYK7KmTOKplzxHUBe3dVE
zPTzWHFTNmxyi+rT+8S69YYrsgiZ7pN+I1Rkj3yjcflseRn7ZWvwKDFzrwASwhnB
1TErTv7G3uCYuQzXMbZdVJg3b+8T2mSWyR3KQ3kA6u4IS86NyJhyeLE2/nUb5YnD
bg30GiZY7S/4XvO5cm8+z9bcBkWUnVMUQQw2W8coNwdlMyHja/sd7m6em0kZ/0yC
YbdSRC4LrRLRpicDYrOiRLckSFzw9Ow7UzDX2jbuYeLyd/hYEAZ5vxt0lnz3p8sK
eg/3OFpndzDqqv2jQvm3Jdk9InXBXfTQK3uneIFCfTJtlhtDzoT8/cBeuL5eybgI
slaKzb216BEktoL5WiPoUvBtD4Dhh2cVpQaPQYT4pthIdu06vPrZMxt16KvB4a5Q
hVaXznwT1YWNIrym1eCnZtSSZLSgJLLT9zGrZyl+4Jddp/dUhQ68vnvSkm5YcxRr
J2lkjJPzcPSDi67VvSqANbp00pzXqGiQQbUkOMQsI5hw8/uYRR+UW4r4VopxV88R
O0M07ldjsm54xmeunhsUW/r05PAPISq0huJr2djlFWnNVBAwMJfQjBRQegGTNULN
WlHG6xsxDY/Dr+f2i+ULy4P1mjVdYIkak9Dl76ySdaAbyOaMgDp874bEl8QFf4KJ
c5kNdvmJepBcRyXUbrrRZJ8TFAAjNffzuBQmB5oZvtfUmvsMD4nU4JWdFW5wA+jC
EBT52HrggkRmz4gvgNGWxqn6tjMF4LJmcfIApHDk04BYmMQH+v/al+lcAqRrw9OU
YWBegZmAdJPKaan89Lya+7jucsx7sbbkcG4oQjytUX++IoChfayDFykHE62V67qq
99y6gvrM7kpiNiYTW4TD+LigPJPa7UIc1FLMxZOSLc58foYZwo2HnubUyVvrX9FJ
Vf8tLJe6clfNEpKhQd6wLYoTbGUkJ+2p+RNp3dsx/VQa2QiHaKU706ANQ6K16fxX
PPzwKxrEbr8NOGKhtEVDeTjih/ze1KMzg4SLNrucD5oNuBuewqHMAxMjsFaTFqo+
YgOot7w2/U/N3MOR80sfIjxghd3umsBIvFT3a/gJc1X8iReuYpL6p0h78NR4l4rS
l5UKcaXwSdYP0qVMrYRC2Zw58i7ogINMZ2FXdrna4OcNMrpTWk7NhiV4D6sxcQ0J
84y5Vv3bMxlAUEU2wdmdqdGqfxcIuyMFy1Gjv8sc0K/x710di5H9xevs8THKVYd5
/1xVr/JrHVkDITK8ilBLJrfQYaw9iIl24H2mVHhsU8FaNaGP1m2cAlZRTj7PoQPW
00BCZGzqeTkUuoeNrTVrjW/6z5KbgoYyhRQpc25AvbQ4AgPoyxU6xHwxRfz8Vggm
VFd4QYHtbPXi6rlSqs7Coezx1WPEtz5VMzQI7ANACf6yO5o4VX8Ik1VNwyfT02HQ
zDVbx1MnVFKiwhxV3qtKdjVrKZ6DGYbl9/uIUtywx0mXyp0KknM6MgUKWq4lX1hU
/pE1khM1TycoHt9UYUEyoS4xwmdFgZ/Ijm9uJePvZ+bd1qTH2kP0MxnKx9hEaGy1
iuokkBzrqfTflrQTSwNsVJTwPhZk7a9Upbg+FE4kippBnU5SiaqHKiVAtCiIOAPw
haYnV83xcJHC+85IfA8hWjxYh+Uio5iKzaLU5IgVBmQMXSfU6ZOhgMoEGJLAxnnE
Lm+Ws9qT/P5mdgBJk10tb/oiK+0+qxhYktAUa3rbMmrHyKZvYzuJdP7qmk70GH17
LPv2hcsP2HD800EbIV5LaqNNsjzbTbeuVOxreof00KS9IVJklZx2NBvymjToXvht
fj79MiITdcU4t+3drvpytLXEJf7pF7HwSG72Jg0BgfFXWLcCn1IzVevGOfGZMj6g
F6+x81J6c7PQBUpiJ/TgfD4NpLY45qjhFgA59Ykyfiw+QyjdDL9AulL4kzTbvVJ4
grmjPMAkBhyiyryTTYPQo+K2Ptcbtdfz5VV3XGIVMYLnE6ND7Fny7g/sfDv6wH0t
5c6zltFBueIDiNTCAwCtcofuJdhfwInD0RHVPyvlJNW0wCB7r1CY5DuGZOqwqKhQ
thXkOOZLmEfkuo5IjwKjYDCRTuajGqFaeKeqA85L3OCLZzC9a5OdkjOaAj4l/u1i
Sma5Uy7CEBoi+EdU1HXNvIpv1O0c7B4ZQzwZeAImlE4dj2q1fJ+c1IGeppM1A8Kb
nbftjMSnzH+xJ0qmpo2+ucdEGO5XiwDEFGWGdM7NAL39olk0R7is2CC1pgRThez3
KraaE5WwuvZ6qwcPGmMJwDIIHMFaNKy4QxvULYASrSAYc0njDjo2hTkdndugIYaj
jrVoQEVqsD71cZ0D5Fvxp4ieD7HgMM/8CF9KQsgb0jg=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DqmE4ccxkbY9HcSDCB9bquOovmZ54zruzJvckiFua5WE7pmJYGb0rKLlkOSK0WXq
vaUdzHtyERZcl5Thj79vGjeCShppTBOreOiEjah5mxqSPwJJY+28sAX7+Rweafkp
UuaK9pBljhtHvk4KOLN4NyZr1YoR54NwgRokUKalnVI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 32976)
L5dqwEBrXIFHWbzeh26TEvX6Ys0y8FTT8X8c+8+BeZD1cDjp2MGvVm/Pw7dDeU6V
zmOGV9WugHm897NI7pEB84YQDiTEJuKi0iuCno8f+euB2SIz1xUkbuZh00rj/rzs
JAh2gV/HQHkNcprlLoGJYxucqpMYJLbn57xPZYNsD3eKE0gWTuR0N2QkhKu13MIQ
u4fGhS5I0XRdnPq8OibaHvLeLKGoWhg3I+Vx7i6NiZLQLeo+6LAxk7fgpj4sGI6o
KXGVG6hGVvJnQABEiH/V50RyocIoSTMIi9F+jyXmpeGaFvxHnnJZgfDur0+71E4z
sen1wLx5VXCutSI0IvMecxHj9WOF8ozk+tCCHd12AVAQcPlRfidfTonE6q5GFz8M
D3FDcaeKKeyDvXjTXI+Pe5bnA6CvP9OHi6mX1PNDkD1vcQLBPeYMHXX5gtPTC8GO
HLIuZCHDiBuJpsu4dAFt1+2h4YOtZSyoSMr8Dp7mSZ45625jPVQXh+JM3X7kGvnJ
4DrUnpTVqo0dZ4ueilqNZ5kte+IzKoZ1FhghIKKWs+r6jO43Pm9mJ5vfAJ/SodcE
vTYI1SFWzcHiWZKfIXvv8vdu5++Y/zJriemAgqAeUSrqTCtdb3ag4kVfuoNMV6Km
PNV2p+mosrRbwSiaEBnQiX7XnkUqL0gyIqVWq+t6xCOaDyJSWQrFiAHWrwwcO8fh
iOZV9jlgBs80PVxL2x4uFSNgIdSrne48UyN3hrjK4g6Tna8xnJbJaVfWMtxG6EJx
SFyl+Ib0JgyIPWHyFjMl+vpvdds39J0hk30S39/Uea6VM/nvaWLlaxXiJpTCo3C1
OAxCBuVk4pafNYINGMEeCfIsAZIZAB4ZgVigBDpHCeAToH9CobyP15vqe9b80FN9
mZF2qPZcZ9lkc4QR3qWL1HbU4D2cbAHCodXQbj5Zb0k7iMN60V+NlbMTSxsiSKym
ex78RB0K8NnPh4cAayS3XwWBM7ZyzD0FQ0eWcT6b2IGHdhKg69RqqbTcg7hELZ8O
aD2BJSFBcG7VOXQC/RAcrV9KPyoWG29C4rkSLZ04gt+xeDT06KqJlTsuG4aUQge3
h3ooNCWSRiOVITZcLd1zMLRAR6OWNPjB00IS1Lo5a4dyLURk3Huxez2gvixTwLNf
vxz2DVmOYqZx3zA6Rgs8uF/bC3RxlD+EBqayVLMojEaSH72zbYfUW9DVi3oYJ3BZ
Ft3Dbudwbjjc0wFhAms6uIKOMQs8nyLEwDbdHJgEqsVNY/SHk9SCqOUKiGAcmsmW
vkMUPUXQSlKbJHa4ZGtBoTNn83m/ikvZPQf1OjBlJqWR6ZALpyfWcurQ+U6iVa6h
4L/MUKP5efxh2eD/0he8LVWDW2+620Y2yzs62QAsEaM5yjLbIZMTUSR/hpaqvrqB
wC/jtGWhV2v3DnOcpBzC2FwK7MIM6GA8C/J7RkjCAAHlp8EwM2LI7bIwbBBGiglC
rhogiPIshHTJFlefDPrUGC43UrDF3uej8ad6xM3H7FMeemCcvPkUVTHUaftZV9U8
KxLRlmXDWWRDnGPHYfnB0wRuGuimbji+dEjACqTP+fjlPWcqNa0BMhR0hnhBPFBN
t5xdRU7PrNrRtp0j4RfaDf40gmMuyJgVAryyyZzS8x6FjASt0TWYmMsl1JxwO8GC
PlgaefYfzo4oBkvirPB8QszWnVlERsGCje04BOO1w5an/0RRIEum31ILZZK+CmgR
1Tu2jNm6NFkMUwrRZvJyiMSzjD7v211VjVzoOfb/5qKzKjNzlE/B4rc6+/gpVR7O
sdeFjWkL3RrYOpc9ofjJ6Yjdw3Eh9ma5fZn0TMhu7a2J9usxzgW2RvWuq8aULXzj
9P+/KO6VW/qVh2wsAy0w9TGP2U7YNaTDjaZEaccu74wan7AWBlapaGYjLnzgKlVq
Htjy/ujoMrarolM0RP+xnvvrkCHDWZB5oGtbvHOO1sb0nlWk5FIuns3VuClkeNPM
MsTxikaaYalY2hVBUhdETz/CpseZiu3XzsUMR2OOrwLEMC5XZlSgeLqIBVH7PW70
/RYYnxkg7vnoB3Qw0O5krEDOmrS+9KWg227x0B62a4M143mfpf89LSrq3BxbNrKV
1HC8+DMf8hSupNb/bNTGcVob9ewD9S/haZ2Kq5EFCwl3TS7//2DQMh95m0MA8O28
1q+Vg1kPxN2ABKQ+EE9PLE91sgYm6wNiVgm//gd2PhIcIoEw9vGYpHfafkRI1gkQ
pnC3kO99OV6QXZLkCFWp4swNbm0S0RrWi9f0KoBAIxD4vkv4wvx+K9CXf0lhdrgf
3XuPZhwUwK9PLq3NiJgl+EGQBkEYYYoZaIoQErkqz4KmZ+KeBbobP1dyVD8ty2JC
PHkENjGVGCjUQudbnMrFZcTWA72KFgO/H/8msqAhKghqUdBlE3Jj5lPkvpAIILHC
sicqY/rtlHxP3sCgpvHXCpGdbavQXovS8OM0gCazAna6+v9oQSwX42FoiE6qMH62
zD/zdAOf7Uxa7F67Gh5Ry/zEwcQccjdWxsLiFDge4Mdh1JXV7rS26cWJc8AR90Ed
5sodHvEA75kCdxdqvyYXhAP1h+TlkKzXub7n0UlbtIlvex70i/unkHDiOCKTVu/t
/ApN4OYBcb2wieXf2091cCvIZiKcTu7WmKa4M6vm8zs0WzndTr7Q4kcCD4XdKjR4
0ITWIP1R69mSUF6DoD9KcTbDzP2ZtRQYctTT9wt/aY5Bjiu4kzH0C0QlblUdT+i3
+0U6V+yJkFgFwkMDgPo6VFw39352jsxbelxdE604QfpTYh7sRSc3Ipbt2dKwjn8W
NDTUXEoFo/nshXz2P49uL3iphBO2i6Kc71olLJDkbqEfkTNC/l9rfDMHHgwo7wQS
PIwW7vq99MbquM8cx3O2M7Mz4Hcwm/d7ATkYe3C/cZlCAdvnyMFAofXi6mteYfU+
Sn95KXXIOkL5+gajVFIX6foJBh2yB5ItTrKZabCnbWCltBe+85u/UyKvEJOTZIiC
wwMZBWOboN3rEWFaL07xU4wOw0j5/q+G++7cx4jp7lDc4t3lMmMQIV5m+XSe7hQ9
YailwbAJkH3pge+5ZzickYHbJ76mxzm/O7uw4jw5MDDMU0cLJsYW0ZPB/fRs1Zff
IOE7/WQ2Y6lBf2aNJaWrY69ROS/zqr6onRi9w0rk1iOJI5xUxGp+bKjzyH4YUxJ1
9gc05tgOJJ+dhbFhu+vxtYovkWRnqL/UbaeBEJgSrmTbrftLxVRGgdxjso4HJSRj
3IkEgIX5VAlfIOkWozfTxlpXQRHQfekUBlEurqzPknkB4Ji7nL+aOD0xfNLWJEGN
JaWib2WRq47Lnw5HTsENRo1FuiaukGNRhuU3ZOAw7bUIHW9mMBtOYYPPXAACaqTG
zBd+a2+xiILTOsljIoOcad9ssRShRgTES+1CIllNsxTtvKHflAsAesqj1ydgJB77
tsQtpvD4zTDuTT/pRvrfe8lh4gZqIlrMKc/4Qttp43G/caeAgpNOstLeG0YzQMu9
lsY2e5gDBrkdw++Ck/0ef210QkrTsEY2LgNfRY71pPL4Ir4jxJmeGKzH2TMKBA0W
j2z9pNKM+/CyglmcL8BC5J4Z6OW5KURMJCoWm2xtzRVuy2+LBW0sPjWZorWMD3Av
Rzjmz7tgPyqi4q7MSCcv1i+wYq8wQGsmOh7dHEKrpSj4o+aZ1VuZQrOKnfrX3gHV
5k8ChGY2l+7BwdKUmwiRzgPKrro2mbwyOeaUlD8FKKX8oVP8YwDNElPVbLhwA3pj
AiIlkzRiQBgm2AWY6CQUwKuKVwr6CkILD3NlRjUY5tjhGji7a8GmZSCCTdx5terL
f8mrz6hNIQAqIPiXo3NnC7jgGeGpolRPF0CcJNuDgOkhkttP+KnYBe5HuBE02RRS
6VF1mLvNg+JD8NWqJ7rUrMBEWMv+wJ4F640OYTANE489FvhfV2mFV9IgZUMSgryI
WnBCfYSfheYjMKsKwW250jkUcBx4yQ7xK4Ye4Yih7VCOoxn1ODjdbVwHLcLZiEgm
mDtGkp+h68qF6RuEKJB+SRyhCaQMP1AerxTxtRZkgdpDTJfZkMxKFVSOkBWrTq8L
+wR7Bk6wlFWrdC2vaMAYJ7uZihr+idc1PFTf0VehHMdV+ETKxf+zRTYvf91ISPia
eT+OyU7jqFt/KY6tIUwl4EWJKOhR1H2gcFcrODr4rIAG9hP2dPfDvBgOtVg7S6XR
JaVJSA3X92EM85EUbnzzBVeIBdCZV3ver9pU3m97mkbtvBtHnh/e2HYlwVyzoOHA
b/0J4nYVUcMY+VySg9zXkHhXYOgKeb8dm895NixK105VBPiooO5hGfc07jZcKxzZ
KDSToeoXw9PZYewHn8pPkb12J+4uNr5o5OaPdGHlbOWmoJzOSqWpyPVMe6RQ5aDH
/xNzl7wuYp4gCrHaRy0e+d1XtTPqCbFAbeACYtgf1E0LtJ1v5nmlVgC/uuL4qqKU
b/LRDPzD461CqskLRs/eLkmHDj/n/34e+jxNwDAi75Kll5HFLUdRM7B4y/oMcOJE
3VTIK75V/SZIVYam+pNsW0uBELTPsy2HftcaP9f19mtebswUygcPinDlD3xEBGHZ
20V7bV1PkpBcJHJ1Ea+pu8LINcLaALk63Uy6nBcab+TmvzQlzf6vJi7XgXId+I+e
K7H8PVpr6tvKTK1chN5XquPrDH10zVIp0PslRhu6annlhyxpURZt7C2wuQn85TWT
HSuIzGO5mI4P+V6j9cmncm3Nv9uC6VPDI8eRADTTSHwlhYjcyfklIYGRa8Q77NF6
yUdPSUZwnySCrGRCEMxFoKO3YWM1/iqFUMmD09BVbKrfQ1lNqxqbgyFdpuQXyv1T
CCsp1YB82M8Blsy9dG6gpJrJR0tfpQTWcwb/v+ItL3sC6JEfnE4xa+Ay6UBKXPLv
iq0Af+t/NCeVF94TtCCAT1uaMyEVfXB68XcpPzpUNnWxmobUDYZCI3CwFzowohj3
THPY3Y4X5PPkRWDiDP6xj1E/O2pZyj3ACr1HQkk3ieGmygwKyvARTTmGUdYWBBaQ
cYxFzgSUzZptDyFtmBjLpwbtZ1pC38XKdMJ+zWQvF6bs2UXBQNCblNzhqqTOMzcV
bCB1UQN/wcNM4h6GMHWTjaKJRqQ6WTapOFi6i54o/2rC6gnf1X+XI6ipxWwlC/So
y3JB9axaJDHWECQsDg+x/R9TneZIudneyVWGStpIU4b0aaSYXS4/I8qNyCBhTtM3
HPx9sAiAGrBHY4dWVdXdlHhZETocTjZdaLNUVlp0AjBjKCOzvv38yfpX9DyMGhQe
ZZ+v48h4ECXNmyy5J+6Y0FDJROVicmGfE4HMgEVZNahj3NA10qrgG4lPT8gLhEXz
Wlv1WbtA2KEzZd5yK0fPgCeOEJ8ApKyrr2LbdwBWOX2JxXaWCZ0/81kOIl7iEecA
6AYOlJVPaTjc2H6r8WKCm6TFoKUdNPmxN3NrBczp5vzux80WIFrGumJsLDFPkDSQ
0eF4+41YX86CRj5c8GB5f31dOqekcvHOsguhRg85aJpUeDvMHvsK+8u0BKlUuX9w
6KILxiC+Ubqr5Vhah8XXM8gzDxtvgnkY9XgFFID1mOPTXMC3xv72B2ZeWvL3HUYG
aDtjo1zOQq6a7B6uJa/a/11xVESS9lYc7o66PT5zwOWfPeEP1GGfNJnGgpxBpMHr
rL+u+U/5CGiGtIzBYEMAiOcvYefp5YtCwdtPg7+Y/KXsx34pMZEnaKtR0mMQER2v
Cmm2O7L0mTpvHiKoz0PubXZUAaBKxogB5PomBBqyQVAFamEzL/tsm5eDMqZrq4If
V6duhNivlmYNZkCXhy4ayUS9/uLZu2xLEg3+QQ8i5BUZGDzh2k5SQht76SAqt6WJ
+/weJ9up5fgwEYNi0R6aOMpwbPeA9Dd/htd0bap+mauyJBOA5l8tmrYo659C0t2c
pa83fGktEys0xOV/2G0tFt+XKpsg9k91IMSjUmUqvBw3q2UqnnPAAut9+vUnfQYO
nbsD2jgoGfpbRwTBtRD1bUVdv2PTjnjLZfNiZfEfYVAY1M5NyMcSmJDgWZFaSIKM
ke9OWFWKDaFS1NupEh+FISRcdqOZ3pIoCCrXSx/Kn5MG4WQFA6so2XTUQwGBxUna
ITXcc3P8KJ86AQlwDB3ToZG+UykLy/0PaIfIz30SZ/IJr3jQjXc9iBMPpaSlTTCn
N50Y2d2lm7Rl7ufsDSO2qvq0ve88YN4BmMvKLvfS9D4LU+bzCBBnUq5dY9sgwivO
sRapCg0fp0EuUTVtKYDAvckTnA7W6Rjb6nfvFQGZWwNWjSZigvrYyHA6BPfT7Pb6
m3G9Ry/J9Trzzq99l1xgFrGbFLyPqMVDJ8hrJm+F5VcNAgDX18tVgl+G1X/3tJc7
Xi4GFmzYm8QblBqUpybGho7cj5S8VIzKPCCSu05JJTExv7/xB4TeNjSsW7MpeU6h
nqOviwLC80uWyYqDeJaw8BXzIZMEmWVhxN002CIS9HL2eVx0EdRgcXu9oeYMaSG6
Mrqs2Ieth3PJNAhTtjPSBCNMVqIwOkJGmhiIC9FNkjo3T1rh9846UGokvYvNOcgl
lpv85w0V2eybNRYDa++wl1WvkkuIkz3PoqBQUxFVZMEEdya11HjZaJwAMnz2Ycvl
PE3oUExI4B4V5Y3jlY6xJPhF94xGjwhiOigmQBEI4LdXl4gKSnjKPlLyo7sZbeeo
92n8wW7aMSQOENe5Do9ah0YMdezQ7kRFwZF0qB8kBKKvT0V3cZ4Alf4NmXis4Klv
gZrE8d3p8yxbbevavUaNt41nNLlM2PELgjSqhcYSgYMvdLoBf5MG/EWQtosFvVdw
DdBUeiUp+UxgdY1zLduIYWqC5iOC2LjHO/Qlqi1aXqpi4B10Ru48gXOC83c5W60w
MmMif3yN/nODBI0q/85bIlssLmu6kaUHs1dj7Yv2A0fvHKp3bexpkVcRlvJ5jdJu
3WGHiodBJn4avZtKrM0YzfYxGFCuS5ORjXxMu4ACxxn/OIJeJRdBq2DABSSS1ilB
VxRQPvzfOEVijsEkfh4HamquAnEWl47j1/CdwLBlq00NNwhv7z/vNKgnLKyCDM3D
7fqqaZqta1RqUCO0TFrwbB7O1HVUCHaqDyJG5bHFgkFZJqOjrO6MBeWrYat65mvM
tVIrBZV93zf+GeyRlzt/02Du+6Uns7zfNbi2odir2rIYqy/XRPnhINabypI9uzvt
2iGyD1sATIvw6vmybpJkL91VV/CaAu14FMiDxU+fhK8COg/fRQQGR2h/0AJ4n9hi
IctIJMkHoczptfAGkQeQmp7ElyFuFpvdvw/JjNfwllupg7/Iqnyepf+sq7CACP21
U5eXp3BrzakaBM29p+IQoRiY3lH2HkuX32YCoepxJi7wlZdBxaEcTY4Yevf65v/p
7QBz9iyDFrqle1wHrnxZMIbRWAXgOkIuBk1XzrZnRWD/KcBca+E2VWJcBg3HCw+T
g/z8dbPyu4FgwYJr0DqOUpPkqriWkwBMZN5nu5nikAAaUoQFw+ewOuwoRU6z4v8S
rd6/y3li9iCbjOyV537xpfWw1d40HOWMlfdViAZ2E2lCgjT7oiLRO16Z7q9z3JZU
OAV/vGrHziWKqgSPodgQEGcnEGsC4BXy/IMlmPTOXh72dxz4rknyHqAWZC3QXzPT
Evj5EPYFMIqJKL3zLiM7lzeRWmBoSLq5lSgfGP5hr4a9xaMgBecyfxHWQR2uZF5E
P/c+x28a5jYOT1EgkxDCJeCHBgVVqllYpn/bWkiB7fx50MuZgGLfxvAhIBPYI4Vr
LrOesS12YE8x7qsNJpCcUeGrF3ZgfLDcGLupgFW9j1YqW/mZVjPEA1WsL0IRklSY
xevCpETYQij95QDIriyM3JaufQ2Es781kaaRBPeiTxesjwp1huRGcmEcGKYbgBHq
V5dS90f/MZITHTUfnWyisJHY6rTZ28uO+tqdDuYlVrZt44UcGF9iI98K2/p5kj2u
oLlH5WrbSBnky3Djl2OY5q1dqrjffnqRlBErjgiVuB8T2VfAIiibUsqYHgwu1a1X
1Qk+ryzZSjCx1sCra+qEXoIJzUDXZuPrs1f4m8fQ1FwWURQJrQAbY/NYy/CZGw9j
T6icXuzDhTSN3th3lgUAsQ/gdRfKWQbDUu4EK1tuW37a5F0PQ2wgcHh9BdZgub/p
PKT98p2yNkkFG7eBJcrkrCkApWPdCrFmjIXPya8rBaRvrsddnEM1rK890j9Q8qhe
d3a9B94r9OglZLGkuIvAx1E68UbbUA86ar08T9OHW0hadvBdSSJGO79wipUGb+y2
6s1qnzo0eW5OKnUAUperA2RQQBycYjeMxfJ2nmhciwH88qAjEfSRVGr7Y0IevpJT
U59xmywpdBVhoFEDTad3l4+Ehcco2yf64H5hCm3gnC36G7LZdST0xweujTEg/wbQ
PyiNEsXHs3gezXlwrVNl1oT36mEGu3O7XwqYgK1PBoBKaPiwGdllO6wnQWMeDCEo
ZtTGv9i8Rs9yZ/UaMVYwKkcZkoW6+xI9YSQstOnklrQzThoGnCp0CEEgPre8NCPE
tbyuBxfM7VRZAhocDXVUJKLl2a66kFK64CKg03wK/kOXYmnyBuHvM7Ye+agr6NRf
xmjeh8BxAM3oclbam+vdLe5DN70Cf2p3OkuervrZsYxvpLI+gsBw0FinJMsfbF3F
JLMmUaIPX1lQJ5RAGZLwXiv5JkRWqiQu1dGLrU6VvdgpjcLQ13n6CffODTHvqgdP
FJuFMkX2yCLV4qL+d+x6GxLdgm21uQrjqIMyKC80Nns2/0RRmhSIJbuTi951hP22
gV05sBxiOZMl2HlJhYwA6J0wtruxZFrnp3ySpj7rVgIIOcMqeiyp1lN9c2fFSiBJ
jDZ/0eqXisbBE4bhGfQ0Z+gI3ZuJBkGbu9Udc3dR6T9AHMqSi3A03fNqMtTY2xk3
0fF/JXXCanKPm9CAvPjSIvzapHYVsPdwxelC7mqLDwZXFGDu339o/5qrfYbYaHAB
qf7cBt98SCxlOvLjKzgxdQ4BCDpdr1Kj3qrY3KlwSUQH8LuYPEYth1pgxjMxgjTk
cfc8mr+hMZQUcMB/m7bRnmsI9xFtANRMcs3OOMtHrEqv99oMLwFkuHAFbxeEMKl6
Wqnzm+sIl6y+I5wFa6U5vVfIGZwUGcgA78ycRGjZvXquloin/MU3OqB/qnbwDp7i
eBcFtefeN3mohaKQJh1aVIfchOQLugGwXJtsF1JGm0muwAHveTdI5jgsdGfWTJT3
CNfl3aFLhrGY+8MHtGA9/ibOuAm1Y8mLedkk8p+VIl3uV0U4rIrYICrnIQk+EmPT
OLIa+Bv3/bpeLd4O8jL65eHEMTIuCoJMFEAPktgJA2IohEFwb8sdHF5/CtpAfBJS
LWL/f9nOpWDeTh3Y6pepAQnnQMACg0jha5vYlQIwG/AIQ0P2VkwIHszgybwTJ8bm
JNuU+ccFbsgaSq9KOs7DCa0U/RCgCwK/lKcZMucR/FZltjSH8KGwpb1AVZp9znDu
SLyB63zMla1mw/ch/c48MkhmOpOO9ANRcDkYTcUEAbzBpikh0XioubQ5QBe6Gn4f
+eXJKNrtkOmtA1M83YNuWyxHxXn1pAYiVPcTgKD8hFSvRdPuAdUh/i+uqb+g41FT
KI9fj+6pcmvE9McLV6vBH1zX+pLjN+bz8sTZui4ipn2SrDnVoC5Mwlvoj/saWkhc
R6pKzpROi/dxzU4UvNpl6jlq5YJ1LoI6syQGeOOEJLDmeQCh4SYFBEx9PJiwPDVX
VavWf84nGkvmC8FBqUTZK5YN0eBf9eNgVFAJ7qgzjXCrFST3LZxVCoAOM/c2DyCq
VSbtWkGQi2KcqF3/zKA1/kF5Jn6Igy6JEMDNmzP8Wtt7Ko4vCp0lxCABB5Z0Xrkk
KHNku2onIopuC91WK3phCDNuFD9WQoxRewb/0qUSi7dwt7+6AZFP29wOzj5GOG7T
o4LMtXugekUgtsLZene/GLAP7FHQZFOhEQxEHCGXg+/Gi2MfBZden1MwYII501RQ
N3GWOVtQcD2eUKmoImh/dbS9hZrA6of3ej4TNzPSQt0pMby4jdfQPqMAfaT/OXjJ
gKcQuA13Za60y2YfVEnf3qAukWCFzrgZ1Q5FwZivzdR7AkTTnZX8Y2WvXTn88UpJ
KQ+4kc7mu61J1iRUlzulYajcTdAtBpr04jFHvJxFJVHniw4TRbTRYEnbHGY8FatF
bJgv9CkmrCSKVf/mS98N0iLUkXp43Ncmd5b3I1hSNjL/2uOUB9SdnkqFuC7i9OcA
36Wqv/CwwKU7BdGhHrc1137WwWE7ZzH9ci5h0L2p2A/ei3mkT08b+6JSiNa3tXxj
V7Sy8B1IIZ8YlFJb/BYj2gmBiwXX3Q3ZJHXnQpMqJFglXta4esxWEhXQuSX7XZG/
Xa5BgMfe6sMiZ+II858BVHGtMcQEzmcIG+iDkTfMyurPwhNhmZPePAG9bHvFuYSo
u58J1nHPYoo0By/hx01UxBelCgZ62euu72ypQnKNG1Jniw2rI8IRzgLTd8hXtx3D
a/oIgEUC8jtCLYC6oPC0/GW2J4ZkawSU28ElHZe15yQIq7ZWY1Fvazjbd54Sh4PB
bORXDoZcSA0W2GSsLE5lZezQRsg1E7MaBNbVie+yy9x+CrAFjR2oBu2qDPs8HebU
+PAFv09HO+jupEnJ+lz9HK+1xD/ZCdoH//toFYnzrmaBFRGtz6FQT82OuA5yAfAY
fQubQdgQrpPEf5fttIsSl3u1GijqtFFZ5+Tz9OP5wgbXNJPDKS0f10vHVHqPqQl1
F4T7xut8xvVI/V5YHXgSyfIOlXMJRmlCpGih5cfe84heRYgCj0n2JacanpSERVzE
cteA/u8KcqJJzcKkpvQ72lRq+bi9S48n3BeFIjYFEq7+FpVFMjFI9CZCMJwBCR59
LppEycKhsLVmzfhMRqwzIEWUy92Hcyg9wM7NEqD/Sshh6LGMmKRS5oVUs1l+I9CP
XDs7QbsosW48LTyc4vmGoL1WAnzznUlv06jxvoYv0C17j4MkqbBKc5LTzGN27S4z
TNH4YG1wyRr0ci2Af2eGKl2xzhDaF+Uf4aCc/iVkjOYYRAaukYSR/K74vMsTMPKc
ETKWxEGaIPa3XvzuGnvUV5c5lElGgUcE+tDYwdAP1YB8Kg0e81A5MZCA+gxpaMXx
PBzPH9+y3MCuFyeMrhMUDcEUkoFbizsKvZ+DJz+LAlAV/EEEHe3MSKbBffAAUaB3
qpP6/MnTb9xekeaOSPttpFFL+SVMdDh/tpzS18OLU1mXi4dmeg0Bi0mOEL1elAd7
Eh5NT8/pyjzz0wvTidKC3fzscz8rio6WJDoR+jd0SY6VlaawPO2QI5/HFYhJ+Ie2
qF+NBoNATp3dIZ1dGoeluti46el4haWXtvrASwoifdgaKR6W4aMePs9KbpNwUK1D
l+WBFgBYPpVjoPicAUoKe+/j3ma4dZgvJ79Jjb+VFUvAMFx07M/SkRgwesMtLMiR
YGxZktwbvujsCULaJSZFFMLNxtShVLvjdx5aIhENFLUM1IS5eptKlpBmfemaxZVT
kkvqOudBXp9ictpSQmkw4W6ks297KzO+2DBDWjUK5enTbUVOkmkkt9lpFAivGgFB
C+F5d3/MV0QsL58GlEu9I7PDB+Z/tPybTJw1WaMeQcpdjKOJtdiEG5Br2viuyhCd
yUup0fppMPi7IXrx6xuLdS5fZ0lN0AMYRB6JEmGkJUqWyxlDuX8hMnZ9pnvSHcN4
rey/TPFgMX4hqVXBXiVGTR+xz+ApmfnEM7qL6W4xXZs+vET7SpHugC+/dFk18r2P
ervoQNkNFywn8gKLbhV0qY4qhJ29JODS6ZgL8IXApfPylRNl15wNei891Bs1n8Fi
LUbJxfQynfAXEn6/Zd0QXZ1q7fK/XpmRD5cowteP6tm5q0rS8FGUdbwpVLXMXNN2
PKyBPqKhJr8/yVT6JhTvxTlrux5h65MEZimEm6uK4FLCN9OfpFKmUwQ7zZmVHGbk
GI04KvtJ62gH+Mmdg+vnV+JZLdWSv1f0DXDMewUD9NVQirtL7KADDk2LQ0m2Qy62
B4nGRh6RH0aE9M5rUeNO7gep2r3QPiP2CjYxNpgF+NHmJ/uFItkU9mD8OYzpMm4r
+dpGDrJclay8cxkublAcYuYOW0CB/LsXV1MBfvEJSJhgqD+yw6DGMqFDQGx4XQuW
UUVWPINCLk9OGdSzJ1LSvMs/mxLYxqq2P6QXEkBvLe5GxMQbhdS5JpLO4fJ8ZZW3
7ZtbpSJob9/lug6X6nS8q+rZHKe2hIbQBmxL84vDFUg2nVlQTrXevDqiMr2rJSo1
XEViPCMXkARgGrysBa3YP+mp1C4ixGMrq8rRL2d4oPxU5cupOkyX/DSkqgL+NKBf
wn58B6mrEBMq6tde2bCTweIjQE4539VbJtss2qFgCbbReZWcrxvgQsR4pp8nACM+
90aUY7Cji7GeKmey15SWgxHRaAvfG0FVjrxlpGQMYVgpwjc/vBE4/T9e4qVJKDcW
cfsEBNpeUO6/OL/F7cbKHOU4ylVEHhuUSn/X/Zu5ZW1ugUBIU+Kg0BS24YQ/bDau
vOSfM9oziFssslH9GSdcvs0FQJoTpvEJD9hkaAneHYdWeCihGerJ4jowEBpBSwvX
UPAmqV4SOtldhJQpEKm721Yaq/ykipAek8coZ4ktWw7XuU9/OB9KtzE0BQ+eSRBM
uCuk0gR4g/MQ53ePp1XLpkm7Mt/gIW35rjlO2AQJ50OCzm9d/th9VsjNMpKfYaNc
xkxlv/EQvKwGc60JpN6mgYbuiIo65xkU5MAChxUVDAwUb9A18x2Ox7g4lE9Px9Co
x3tCza7u1SWIi3gE0f61RHhAS0d+pfEKlEbLj6gbnotq36CxXipddNd/e9jOB8WJ
rrrbswIIcDCW/v9+zUrDY92dlP+pwUUgzlS3nfUH/Sv6ru6pTKb1gOmsSVlYCl9e
Z8+cpmzlC1ZptqIE2KnfeOLa/3cel/haMaJi/vt3maQ6sWiM50cdJWsOqXfA9zJp
ggH1o3+yWfsxuSQCt/Eul17Bjde5H+2S1OAAizv2tspiV8pM9p/Pwe2v7mWwqXUj
Rt1Ln/GBzJa/0s7Jdvfp/DRK3eq2JmB0HKzHp2jQYc3vqnZwnPnNvYRMzDam9Xl/
/VUexkZhRZDJtYdfOBQ4cWk4eCj+wIKZlliLmGtfZf+AD4Sg/KR//AJm1wtCCdWe
rsFIFoF6TfLpCwQ2qbqdrnhww9mCurUjxI6nlrfPs8Pc6bD6VWOmtySW6N769wnh
B2RXNMpLUm7qVWZd+8g3ZTrZEkaDV3VgjlfuvyjqyrSw/20jK06FvyPC6DN0178s
WjykWACr5Iz7pdLBjAfmL6Ho0n9qmxdqofslKSpAJa/Z5renb0gyJqjxCUxhK/P4
V6gihYTfrfHIxdTV8I5h01MiCCGSZRRaUSoAsVgmuTCmFJzsBvJO4AiBdeBxtd7s
WSCyeDYMsn6cEH7CZeQ3aPNH1WNquuSL75UeB3aBtjoHLTysWERuVQoeabcZNIXL
nOmFKDs+h4Z6AFnCQi22oKfyQ0eJe2jXCdCtYxQQl4A1cas5NjANo1FtFg7FkFbs
68swsMQPVw9gV0AyIEEHn/eJwGAqGqTYORTEGwqhkhXp0ZpnM+D3WI7HqSNhDMSL
1Jtybr55jCnC3HHazu208VWtXwdFeQNbyCWybzhMsQblACqPlSscCbRTRcl2CLdD
oi96L4NFDl8pygU+bNExl3VQiZbqtVhid+HA3aVbDl8P2RQ/gmzsYmhNMGdLaH1w
SHqXb4D+VyYqm6NhDJghl18tv/HGr2q+OscNCPhQu1ZPAvyTNh0fbBdPUA/gaLck
f9xsYwQGVw5Ir3kutIf6NQGQ6Ji4Z48Tzvis9AzGnEDqP6nUTw2ruYp65PxOo+Xg
3SRQu4+7BtkFGbo/qbJlZSPesLBhdy/AmjpoC1FnZ6cu06cguyytaWSPyF3KQ/7Q
PvLNd9jCxZjJtLysJmBfmG+AvyXlEd/l548sRjaRPFxjkzxF7XiAgOb//8gIki4i
wGCave01M/c79WBNkjcG+04u8fBTyS1L1n4rO51p2Af7caTp35aho7Tg2+rgeLev
+Xb+lJQvPpdHEK3rNWf7lR8Fmmeo20ttngxI1LiO5X5vaUzPDVqD09klW+YKX9f4
vDawK+u02v7AKmDb4YaA1I5Aymj14S6PpIHYRl9pBBok8xCxBDnrpZtF6uTL+ZF0
27ZGlRJnEfU92RwpQ+f89HJGWILv5L4mDpLi3ByXR3qTTtlbFZlGCTkCLAPGc4Hb
BeHj9I2PPMpbNdGQyY73cZQafejDm/34TGg0cH5f2xlAA4SEjQ8VauxMqzv9tPOt
rvBKMeFz3wZ1aqtUglaXrRe7HPeRGdtTxc83wcI1TF86gsOESH6DQwWSCTozweC2
MyeBW5oeq9hZm0CdnZWeshUJmgxBlt4CVgL1xflat9MZIHR4QxXXTG/8FgjMQHbd
1W3SnWICiaPEnNr7XJj6vkaDTNIZtgEII3V2IqEuuStbaGKrJZPgoRD60U7N5uB5
eVgbh/sHalHaLzM2j9ruSGPxHwdVp8tAogFI8iBhmOKXBwzEJAHNEOKlWXu0QkY+
RrgPGwdKGuvjyra2qJKcq8Dp/SZcaclGsfXVTg9Li5hYYV51pQfe5b7P3nhCCC1f
eP0jWDYJgXpR1xG43Np3cKUbj0kq66bkoUUC+Xxc/cY2a9t33CFdIk4aV7FScNe0
Z5+789ImoxhtGJyVGeTVJHIpboxs+QKs8m84oS/KNqzRI8pAvcPq0oaJrpUxVlkQ
htInOleIFAiMkV78ReuvHk64mBRT0guXHYL1wygY8qizuO9SR0Fc9isDwC2cgtUz
74ea2o4UmikfzimE4YaHVznL6sMnYD365olmauZe9X205ED2XVjCkEhMpivtCKDD
i53f+fBlPJ8Cwk8Mr2Z9sw/Yn3+EBvUgzM8lqi1GzydbMbRrcnLD/fZRdMQ49iO9
tgrgqJaKOrOaaDVfP3+p79xPOGzQsLC+q70U95+2nZh9Qcs2g3zyJ6/qh/n8OPzd
Uqtwl+k7WS8eZaAunXBMpEYpHNT3adftxY6TUtqrE/Oo01Pzy/icmu+WpaG1acA4
4LCNvI0g7v4PbxjbLZp2lDen1uEiv0p8MuRFmuxPmswX0YQ0nNmJJYEOGYpaYwDk
G3pt59WP56OSzRbNyTMcqOzx1qMYKm33ImAVvzgwx3i7FC7y2c7f7K361C6ouV/Q
rYjEOh9nygIwgSGEUQDRB/DTRPou87DwcuEVOa443AmXciq2GJAqDPWuWbQo40u4
Agxp92o13k5KjbaE4Ln46Vv5Wl6L/iuA+HBi7Ta5sF5Vw4YNrRVSIXwGa6uoJoUa
4DjVoFcHtwNjOJ+In1hUfZRy6v8CA2dqecgTZLIsMyGZUkqjyS6MMzfsYcusg+95
ERxaxE5lPXEbwLcRn41nw03Iq1GqlMj4qveYVLTpavRPA6B0HjwgYsAE/2ss5jlX
GgayRduhCSJMg2EDNIhILo+ym7V+4LMClRRHzr52cSa9ktpZCAvkBXCFq5tH7hjJ
IHgnISsCDwxicJdzCnbIMyfZ/TDzpYL0JEJVxjEi+cIEWrLXmeMlfpzp10Ud/of9
jSJUtj+xAPun+KbehKbMvpa7ZimCSmnl5aLAl/Y6ipvUys1IAius9Z8/bszFmWcf
TGQVzOOfkTblY2wYJw+j+u9HxjPRLCWvqoHfeNUJr1RUvbuiIaE6BeVVKHeqt9BI
EX1cHyS9/A/0hWkgjg+cIXz5eZtWUFsoIlMOatzNPuumM7IYV3XE8yyCqS1loigk
c0WamWDYz5vHYZq5uGHoZMQTUNTjpTDc5OgCCwHoCnJeyFtcbMqsHS7S6W4eeQ/J
CtdCFhmROTolJjXtPKVX2ThItgncgn1n+rjYZ5pOJviJDUTcOW6mj5vNoNaAvmYN
QWW9AeNOQVWAbinAhPO60kapkBNqhgbXjkmkJv5OMN1oe3g2UYO9W07fE80/+uQh
oNINjWxRL8ng0+mhRyhUryBK51QytHO27MazgcJME7d1ATr6DNduJZPnHoIptXFY
6qIulH7GfvrAGOF/OtCQcX7bYVrPcbNGbVJv5HeHTotNb0PevhLIux6FzcfWvZ8l
M2j+sNu8csVaLMq/O8koQyjt4HL2kTPqcM1OPxCzoTNBzVz1By1ctokFRd2s8zPL
mgemd23+fc24sDyOT/OnARF8EUXaBVQIAnmShuiLmxhuUy2WQzItCSk0L2LMeo5Q
dwNcb22JPwD1sxQesL6xtfc+KrJHGy8QVWRWGN1DTaKXUruhollrjYMKSSnwg+UO
EFtn/Y/T1suGs7NqGJV2Lx4BjvwPZuY73Lai86sFBPIO7BHtcJPs/jWv+mRKAdxb
QBn3TBeMjSLMg7piTvmdT7svoUOAFHw+javdwknEVwJBZCkHaSjeOF+Vlwed1ao0
YssttQYx3mQ/f8ubVvE3mzDBMEOi6EOGVvKbAfs7dLE0RVtsBL82kFpMO6fWkH8B
ygL6+/N6WUFBNcP5ZKMu8fskK1buL/TqByYjdR3bx0ci3BAr9LyRwKtfZF/fjzOQ
LZ8h9ioE+XaYovgOqbVdrVAWCwnDtGcS5tOUj7sXwQyKH1aK2v2GRX2r4vglp7rT
+Olpk4OFvJLalJHMPavfn32wUlrIEOn090+DW0krd1dBkTFc0kJgLcWvICa+AXrW
5lWsHRy3dAWDJmun+nRGCqtFMvd7/j4iMA8Nrxw7m+8pkZhK5erjtjfNTGRLX8QZ
1OdFloHgWDRiN3KzJ3/RA1nCBododrY3lvUxN7alD525yHtdCvY+7bUCjsCRQd8T
wsQgTPpNn8bd48NIzCldT7s6uJyRkNAwOIh1RU0atFwKWL/8H9vcVbAB77e8PZvO
njFNX3zNbqcBAyuU2VXoLT9cRBFK+Klwn2rZfm2OY+mhNrvRkqWQEp4sbqRH7tnH
RFxWQaWgU1dz4abr/4JqxF59pm25AUWHdoIkdblpFPshqRmXoj9RpLjsBTcfmM9c
GViZwUTNlNFvBUpvpBOpYOahmkS6HnXzXF0TI5mLn1dGcpzB9P8UPogI8Wk+uNyZ
JRWVNo4YPlunhUapFtm8McD8IH75/jcrvL3YeG4YakZXc7UkBN/Lbkr7dSz2OpWU
4VzT6fPEENqdMMjKeP8/FmACkap0cSI/rrpmoO3dyoxyYjXb2TuJ2gJ6vMZklLY0
5pBUHvIDNb5Gab8vHBCvgFMg8fWP4azJV0q4IZ9dQvt5jrWuERN99UNZA15RE4mU
/KrF+f/rd2rQZzTxHSC8c6ttf/5q7LbJCMoxA+Znyi/eurc9LRo2SD8FM/sDlsl0
AKnYCW4Gs0jlNi9TGOVeA1zY8YmU+FKfbJK5C//Pbe77mMqrztxcAYFx+gUAYcO+
t8noQ2K05DGJSBxZpHeoz+NA/KQPmoVxFJCs8ImKgAJ7qTCkHF72QBM7c5tD0z1R
akoR3fZpf74nGfLYEuEXo5vnpkf75SvnFDxXyvvqdrFYer9up7HNWHEa3p/LxENC
5IYo7832rAmDfK4/kV8iJcQ/JrC7UnwTDoAb7aS1/3xutXiO+nim7W5pEH1vfnDO
JEYLO6W/BygpOwSVR31aueicj1vhT4BgkZub7B9xWqdItsyWSJojxK7jatSArke2
g51wtinlW5F4Ac1cbpwKl9HUoQQTNeBqfvhD2is815ZSrFjJRUlRDUm71qQaMXNs
35lKdN8AyS6wfID8Ubym5rREcR+R3t2NsRV3FWnhm8HBOA6VD/C4EUytyTiFEyCD
pZmaTebiFQen+GgpIkuFWZAbQztXh8LDUs7c1TwpbOvo6AlZQr8R7/7VJGJi1msp
5i5PNntQkYEFigkd+Y1dqwbkpzXug5XFMXh9zsZfRud0luf2N5HH12l0nS6XKzdR
iOP0YOSnM4XHl7e6/9vg2VPPcqo+NQ45KVJzk4+hyS2AqxCaInf8Zowr1D+bQ3sV
6UiF/sGlpPo4gNEp1qBBcAIALMvXjl1uo3va0qXtpIbmwXCG9ISDS2RWoaZ5KZiG
0CVM92SuSicMIZZJXBjYJ1RGIXC9NY/abmtCo9Gq1xaa+B9JRXH8w4XtmA5addU8
tjUpsEDYuUuDdHExxOXrwl3AZYd2If88C0rskOCJRDCwv4M9t+DJRICJ7090GRQA
aTf7sy5UDYkwcDO4k36vQ3y1YyyoAoKX09xcThemUNGfi+5qgOjkrHTEKG5G4L9T
rVBc732Luldxy7++OuHoI4d4PKoodffxzsde7qM0hAEXkdWAPfkv7jH25ojGCrLJ
9UJvwos2yJwmd5arU4Et3TfIWN6U8hI1HL2ApsxxfygUgACey90kCKjiNLShYsZe
MrPDeXWuwNPpu9xvxb2k3liQXf+v5W385n9ck6aaAXy2Ofl53LOR+9Y3okB6lQBS
Ffb/6N0x0wD9HUbHXiV1vwZhkQxuCcjwDvfsYfeyInJNQgLNGqTrzcFc3iF8LNQY
m+roLvEXpy6FNhaD9uU2SKPBcakehr5hcZNJ2aLdAKduNStrDYLWl25HnE7AHEBU
zBRvXwu6CJJjOmM96Pnp3RYINyVVSbXoTxdWyCf02Hk8MmDZz50aGrlgepADK9ca
jXQQy50T9p3MkynyjbWP+6g2eNR9Mh0ZTIvi5tlf9caKxzoMc1nKwSU/iqTW3jy0
ubMSDXE7zALtQ5lsPcB9t41tZc+VQDSzERJvuCFRsR0jFySwt3R88GX2Ndne8XNQ
1tgSGY8yxyFhfC9v0VOEar0xB4ZWKj/IPz4ahrtBTE9op4CpV2T0vFn18ohgUo05
pp7GXNU88qCDyWsML8fLdSEWgT4l3YMUCiD0fWZeaFw6tEaEEe4I3d2lds6CmSqw
hXc8PS8Kmbh+dO+h1890y5IhfwURoFckRt3ZcU4znCOo0h9kZw1s+JnUjvbZcb2G
IN/rQ1sNSz6vODv7RFOMgrq7WCeUcBgmxDfTWOMTtxAKQ7fP+wWV0+MtwQXR+wXt
7HVRAHWQdqKhgOB/8n1fcOdh7hs8VzGRNjRp8rMhrJb/zmyu3bmJShyL0XBGW595
dpJSv58adKi9bstGiwnM9y+i1giNtejjgtOUxcQszuMXW0zm/cd7sRu/E7UDNnKA
J1H3rn5+4JOgYXk7nHY2JK6rc2VM7PqIREd6dcTP5neDIJBWvpjVxDNDD/fILHeL
fwFN+NUppvrE1wLiPj2KrAtYgKb1479iTa1KyEBcje9ic5FtwXH6PPNfYuS6IzNl
WhQnaSW2Nnqb6q0T1qpDnkuWMGXFKM8kNEBv9SHudevgPsh3YCC07hJ8Orvu2sjV
+L4Ke+53Q4gJRiv/2v3BrHb5qdfrvU09L3QvNKsWejigijt9zvyDazgrdP0zCXKZ
UrS3wHTCn6Dl3tEb5h85y7tWd0NBZjX0RbIETbzjgE8YeUgCImXl4OIVJ3YObvYo
dbM0M0Mt1YM+FLVamhs1Ju/JiXZmE6R21psAtPyjwLFPq/EibC2sPpTiBoXnRVjj
a6ypS58ean5kPVo11ydBtwERgfNJAV5T/00/ZH0bUmDLKp5ce6iddq/Q5rsyevP7
zu3F9Qg//LzZ9SiS8UXbZfZBiLm5zwHoJg0RZjLVQZBI28gsUFe9BJzNpAdtCcKK
bzxp4CFFvDEeS6X9Vgn5oVKRpGL5N+2SSfJOkA+Srk8I3M0dtk1yDn99JrKNWssf
NuTLZb/jYj7jqzzo0pfbm0TbYIUPfaPCtZvZ98Z+1RrR78NyoqLu0PtcczX2Zf6D
veEOZ1uV5GGXxON+945jgONupWOaTsFO3yQjc50O2/fYUQDGOTOVRHf7M2CDevKl
QlV8jHU/Ffdn7eubGPNYjGUGpaHn+pMZDypn0lvCvO/glgFgQEaBx1L/gPr7WErx
ylPDRm04kKYmpb0J9gjx8Ct1XYjdjAIX4uEv9CPiNyzEMLHSGUtPIfQlBCahIwHG
AMpEt+Ai7JCBk2VTDe0ybbo2Re0HW10D3vlfxJkODgs05R5lSYMAhNDwNa1OwugB
WfDw2xtFpB77Fl6g8kWRarJyT1YFPxj8yveweYIltJ/nCf/RnqM6rRQZN3KYW0lE
PTmVnWZJ5/Rb5uqw6GXItjc8riKAf+phcTPTXmhc12SxgBWvycpO8mt2cUHziTqM
OCHcFQ+fYt868bmvKIxiFRNy4XqO/WNZqTFgEL6HohdZKPMaFYeZsjDJEYclKomo
rI78x7CJAtY0D5NySjVGn/6x9rtGw10EjqYtOWbY2c1LQXX/W0m5QhxhoFL1tYqe
zOyWG87vaQJ2x3joVyNpm8JcX1t84yKWtgKyuB0fCyQEyDyA/1TGYf9RIq6P91nF
VRXjmqE4X5mhbQxRLjeH/XzgI4Czz8pjgvMzZ3hNLpmfuya9nxKonmTz/MJe7RIf
Drxo81mZG20VodupN9ess2Ig3qyjWDvqKVMTjZ0y5KEBBdbDEFd6LtVoV4ltw1dq
150C1tOdVaSkPUIs9JrugvIiTTVHqblLKrdPDJrNsGlUjVnPP7VANP0DzKoI5nec
7yUKuN7oB4u8bDq9NTv1CwwRdIethiBhW6uTZKbnbWbg11A5f0scLZkicCWVmULD
4ucckVIEudP9gVLitw7EuAVyhPimj2i1dNAUzpJXYKIOaGkItQOHHZfHp/mL6ro9
9AG1eu00yVKwkvrYuyuODMRSYNDpylCmVQO52bp3xAT0fMnhy9g6d00T1KbBMhoG
0Uq0B+ICO85KvNQj3jUNDDI1FSkh5y2wOplZONIZBH3FmNV16se+9k+Ir7UdZdeh
hC6cmzt+p2S0fRJuwE5QAz2dxRjrxeCxntWT3XE/qdTujmanZksE7UJlvI0iEsnH
0SmZGTopabqZFlLEEA1cF/P1qrm2a9V1FY3m1s4ka9B811kztz9YGne1NX/SUDob
NCJAHCcbVBX+Tw5O7iB7ZDG73BrAxuI5fxwnOflWwj04g/kQjgd7yo4mTJS45YXx
u9ESKpgFXEQkcugQPIE5aacnphP2qdSGrzBQ+BfvYULHf+LDYdVqy0NQW0OWkGMl
CRS+/qsh6B9SXyw5Xhbm+Fkm8aWXDLA27bT66+RLMjdy7/B0mhMSTgkOWbZk9oXk
ne+GDSWEAH9Z2GLtiRrIBnYvbJ6osKm3gYfLiNHClu6e3FblptH7CjRtXV7xIY/l
UNOfZMA+HugGMWtT+0AxEfID7sqepOUwy5g4/hlw5EK6aBVP0GtJXUbzM+1Kmo6t
6D4yfMJvn343BoBrOgIRGN4jfou9Px+KseO9HhHByfHkijyx8jncuLi1f86Oimne
90FGS6DbkiTr2fN1FbViZ5smRxfxwnpLDDT0U9iUsXFwqkA/8uyobfW/mztv3scZ
vP30BqY6SJ0dMEolkAnj225fwC8QbQCj+4gVbpeB41i/iJg3kp8GFjFIg6Sy2Rsu
eb702gKc/2BS2ROLdOzDzwghrxgqv51Jl6Di20/TPPEGzQMHWo8q449cjXkjSI4S
QjVUh5rpB7iQqZK2GkJaW7NNLcn6CqHHWiXVgt/ueGev6QJqMdFC+ujH3PmqGYfY
6ErfSske0NaK6bQT6XhdWh9KnNYZskgYzZOLnDbEH3pSzTiy67GnGZPxjYGgMRmD
NBDtcypE6c4uAuYfBijmNIohJPNu6lryMchPWNMStwVW6jjcT2raqkfX3AAjcSbv
99AvKcsmObZ7/x1czs16XNsIRokbIAPMig8vjgUpXV1zzuL5LP4qc6UwUFmBk1fr
xANaKS65Hunj+VJwLJDoKpkXLW7L3XUHFLNxzWelcA7JWQTTGFAPr0ZkB+ns4FDP
vW+8RTcoVpXSuuwgrca/yKVaBOP0r/PSnzBLFRGlg4hZQwM2+V90Dr/mvoDALnob
S1Hj1tdj9S3KH2MgMOCMXfYvNJlCB+EuKx3ELGujaM+q3RmzCURocbLIAEUYIKka
K4UcqIwqw5gaDxbUEh6UEdsupnf6VU6TiOVOs6/ojClvXY7+zo+pVlyGsPI9gW0W
IJrAFG07vf24CaIwldy0snJ34ImP1xPk2vXAHfFx2iwTG8wiGNXFTphWJKpTtq8E
heeKjO8CHilX0oncOc5wdEXtheL9gYAi89EVETCs2j8/ChzKIK0kiEG2ey7mR9IJ
0EuTr9nWwTZr6Ir+q9IAz7SZwjdszj4ZKrbfatguZa01jSWsq6lRovPfqMYcN9Zs
qkTqeVv9S9CHDW5VYayOLdmVaEyqpT1G9ehAf6wPb9FHvN6ad042zrY4KFYMgacw
sV/aCzgxiyXjr4zcmMyU8mHiCp087Ew0fVydNENPCJPiaH375UNMWhmUe++Uec8s
KVumH/jpCVUy6GsP+Rkp5V5YCfTSUh6zAdBt3KWVEClwMHUTITeISD4qhZqDa4JQ
SwN0alrHok5PbCLShDOjzcmlhts6MBs1nQPApI6QqPWUSbuBxd2k5BQrEkCWaEwN
ovsNvvFqpdld/ObqbDg0PrQIjHHvEzgpHqNje3Rf5oS/RTdy8vJ2YKOZqJ+bzS2j
r9KM2iqX/D3pajPaFeE4jUPkfquoBmuLhCPxcQrflo8S+e04IxnWf+AgmNUdCjUq
TplSBtFIB3Xr1Z62qHfKvWlT1jVxgF1QO0D9jfwvwL6z2ogYk6M8jzx2O8bmGhGk
0lYuEpsPCrjxgMWNOzOqNWoJLF/iw5cezSy10Ct7RcKlC2vadDbZmgMbrKu5SjHN
x3mkbP8G2K94vBs7DKEk0NUORlHAt7Gsw0Q9S6KN5epaqlFOVGAmScJrEozkJKVd
KsUX1dlpWKu/56L2Uzg4DE5khIsTYObh658mDlEELY4e6hQsQmX6vazCLpf3NGf8
17eLWHqCbw3BhNqHiuTAucWS5D4Qgt3ldBOZA4dkNdMZrmjB8mgUeWZRvZx/N1sf
IRB767izfydNWz8M2zcKgSaBJ7lfVMgfcBkwTz/qu4Lq58D66xC/cChsBWLSouhr
+V2FnUzr3IQ0v6a1qP30I0v2c8cnwUwKoViA251z04bK491/f01j+pCG2Xhwbglv
FgNRX8oKHCpm2HHhCgO+pRi2VLocTlKaDNmQpWonNUew9cRoefQPxzOYPKPKizgF
is5DUXlIbktikJXHpobIy7OkorOf4CBlTWArJPUNMzerAFps10ckVMjhnZi5TlgV
keLeWJZYeYUB7bd3Mz2Y9Q1G9dyXr/gGBdjHMHcGczPzCRNuroVrxiIaWZ4b6avG
W0pn/qe/DLsyyoPWVM3Jp845YCFyBPLXnAScY5YBtjXs8WZIqmS/W/g/0DF2rdtB
q5azja8eyH0ehHDkgCJ2YSldBrC9ZBMMbHvBeIJoFD0MGyXyEP0+clbkViUWk/6z
44wKCtE1BJLkH/zp82nWlu6Yv1Was9/C0HfiQ41LgFsYEBcaI/fyMR7W27MFcqRJ
zZYVUzSJdR1Ri2zdHh7NQCRv4XJ49gsm1cqYl0Sv+hhT5hKBLONBq4ow2GgBycRz
6RZtGYVYC6ntNk1ajTmsUR8/41PAHMVci7uQsKmJdOgZVkzQUQGVTRj6kWSVrofW
KJOtlNbzVA4WNPbdJvXZaeqkVsC4DH2J2mmMRXgLQA8Uc/jHnLOzSbF4YCeWqVxm
oMYC9mkwzITvK7fkGDE9Z0xcVp7hH5Kgxzfrz0nr1M9puUTD7CgsQV59RLi5avvy
cXVWOC4JHJX7N6tm8+YMakUAdUPDcCyyOmq5MPfi9ubFJrG3M0EGdkZQMn/F+mnn
ci93muYfFzpREGSJ6VvIN3CZdbTYb99sxl+Tdlqa+YWi4NRUIpqV04PIexVmxGzd
7pxDjJUPGgdNWd6vZZ1A8GTeYHx7RZ+9ZYBa3fetGTC0DNPkVaKyoN8MP9Up2XgZ
gBybDsSr4pInW6zuIS9OcQQzv7PhN6u6AINO/5MDUa4dWqZUC8eHj5Un8syuuWf4
MrC0ngBXa/iZSmoruX5eaWfC1pfJH1kyFPUnpE2j/0DwnjbruV1hFbFEpyvnSyQE
/G3n6Zrl8XbkSBm83YK87jknL2OkGGwGxJuZBg4qj04RO+ga1wE8oHXAEyqC8Bdn
gOZU/f/YTh6PsBs6pMadk14uzDTm9omcIoXo0a1coNkisAKj7cjJQfz3ZP0ehWC4
eWPV3cdoC/NI6qhlvZDMgDrkAwOPdWEJx773btSA9FqqnsaJfFQgMQS2FMryO/PI
cGTeewuIbZmqY4IF4DU1fwUJsGsQGbVjXf0xzOUeRMD0It3mj+tSKuz99yrqMoHb
BXPoYb37c8d1LnK6+ITznIvp7K0Pzqi2InmYjvwlX6CIyaCS4v7sAdfn/KdTRa8U
L7teEkWXo1ewzoHKl4JyHnwm1B6ZQv659CYlQ8k2tgyywd8PI4sc00ieMhwFzWDn
tBb34VFZU+P6Cb0Dl/S33QRv/V8rOEioh3x9dJ/8fTV+aXAuB+bgzL10M52bqWcI
kRHubUjJN/sJgWlFMsti3sgN1Vh9Mcf8K1WMDEZU3jYhEJpJ109YuxPrAa/fIIJx
5ejqvUd/lrGWWdls1PmJxFiuACxy+VhnLm6dzy1BC9NPVogVnp0K9GPpjes7kPui
A3E8ZosGZ0dMvpCaZDWKHq+ApLegsNVQD1DdSqGK0CP+OPh2ZGOORPmFQN5VGQwH
v/Ee+jDUVxbCcQHalP1fevchvwHRue65xQYao/JUP/UiYu/ly/C+BV/HbXVICOd/
6MBjHVbD93UqF32qN1X1yITVGs3aQJDmqM+9PwlQxPXdXl1lqPcKH5/3gWvHtYjH
YdC0QcabHiCiBHU3I4aWRLWFKH5PWt3pZUYR5sEPz1XOZ6H310eIRukVwWVZHoC4
8z46b/3mz2FrBfJyResODK61AxB0S4SQNnZK5PaZDPPmykjsyJ9gxSRLNAn8xNWy
PDcvpfyKjBkCjgRdH/JBmvEHIvU/CS0cwGPCY/2lnurT9u0MCmRLgsiyr/wFNgnD
xj5HmQhGTjwTSQ0XSjvlYV3y0gk6Okgp3HMdQpHBdXRzszW3oa2bXb1qeyeZ5UpI
c5YJZzUBt/a9W/fjlmjYzYP7grnkfIN+egJe6FF8DtwrlpoHOFS2hbXO7Dn6nWfi
RtQdGIYk7D48qxgV7LSVPV7BUal6jHfoOWpQd2+q92T8vw103NV1UZbCPSY085rL
CZKIzWi1Ea9l38rX0F4XYYMwhY7757y3Klb6hKozN/GpFdgIB/mAtm6gqHm7sKfb
E5cAHO006J+v8c//msbSj5qFNpGAZ3i6i1oBrD1MzNsrZlJy5aQF3kmQ/ATEUiVQ
DnO7DuExEtF75pA+6Fkmo02FVnMFogxDf3LDmZ2peENoamUiTaq4oPE1s/3C55HI
eZAwtDmaSF1RDReYbhuwjBfJYVhj60qnLMOiO6KSMSJFhCF61d4Mpi89Bl8gEvV0
tclTvI31Relju4Yu3GpJqS8W9xVdjP3hhHpNlHyyQCSRba5H/Avb7k4BiXqu1Oh3
EeuMXO5hb8ELUpZfP/U5gjhF0agFX2bh+5ot6iQJxrqCnlgIodEMnaA5HA8NpZVr
wPNKukFfi1QLCc6RrVkfDC/oREulUIshBosGjwsD7Qpwn+/+Uy9Itn5IBIgu+4yw
CwB4Q/TRh8fclYQ1nfnJdBh8XI5v23mXXwlBtVwo2M0wuDWjigTaUjZ1fKDi2oP7
aAawTSi40ilVWbAvP5ibB0rPXnkirAet/uLrLWq2EPuKK5HcjKOF7k4pCjlgVFdc
LamkSLoymvZDWlgkM/jDCgBb/eoNkRjC192DXqaZcctwX5q98n8cHV6pZV1MOFv1
m7n+FeEje2zCBMFYxQzDQ0hdJSvfkXtbNplUl294y4L6F59M0e9bmPGYnWy+FyIc
hQftsWOS72f5LLAP7e4kqLoH0p1GS50fN4Xur0A2IxbJ4ps2eXwhD1BUU5YMRHaJ
MLv/Bk1Eo5HAUQFdUJM0H4p+QEIXEbJLRENF7lq2+jSe0nCL6oLqtH8BYqxrXfxv
xcz9IozKaMWY/LsdU0j7bCW1KKy70umlsx4sQklLk0z4M1XeKoIWerPNn4TJIdO1
bCC1yOQEA2aWxO1u5xP2vYjCyEk9v3kPR+MChWgqa8PS3AngTpRABkttKvjQr11U
atGvopinlfSERWSxAdu7tds7IoKqRKdt7DdPvQzZT36YF0XJyD9wNWTdcR0CBsDw
kl5+vqPy9J9zdSu3u3tJFQcF11GXz8Q748W8nCjMFx68pKvw0qIJPXTMm4I3dd2S
XCWK2ETP8wLEHAU6SAY5Q8EU4fgP9zqP6e5iub0Cb8k7wjf+3V0nG8R2kSUk9JAc
PeBrd6IlTK8/ABPxAX79t8nQDZ8YBhZMcR1MbTXGQ0PA5tqFgYybnZuvxlBAL1w8
ItfUUt/sEhQqi+Sbb0z3F5imFS3+Q8N72hCyKec8OawgsnpNjUkvICPLvm4ISeBf
Ki3nXrYagEdpX/TGfzDcphcmY/wrsOfgk2RmD0ZolNhs/RGf8r30V1SzhjOreNMa
IxCkgfjHiBkm5qpFPoMxRE1F2BElo5tmZC4I50MV/RFMWQLaQfZjX8isiO7d2mJf
IUu6G2lht1VhEWi6b4+v5ZD+1ZGZPn6VQq0BY+9a2qxSMKYOCuv74yU7slAAv18c
BEBOhoCP5cTi7MTdHYi0k3MneEoG8Bv6NpUsb9WREci4omTu2JtKKNJMCly5Ny8S
7UeHMDTRX49XkRjaQMZ5QKf0yhI18Il5E76tL7y6bmnZVnVW2AzIPhudMnGRgjaj
ctnuh/0OrU18hhihsbkr423cRVkMJ6Jxx2m5+g2Yva4T6FkY4snFR/nP9rIuV0qG
obFC4/r+ANKBnxBniq0qsbiEHvr/h9SXDeb5/h4InSMImShMMfYmETF51okrM3g3
jrQE3GSrJ1SaJB52RI+NZjV4OeXt7WoE7elkeGX8kJ/Cm442t8mpSfF+F4aRsOSV
gtqNFoED2ZYzSwfs/5IK7plVOu5VnEfLzzfPsXp6hwzwS/Lbp/aBehqlLQQ+6IXM
uD0VgBMErAVmo+nhkwbIEM6ODXhkZUlEJNp9xucEGhdudBcfrmZrP3TStx1xRB2a
/TaIlzJew9iRfRS333DIDea+Pd5L12v6+EYniI3umczwEnH4nubeAafPb167DNLS
jJkfKRZ3LL5ycVfTBtXLjH/99tH0ywjyaDYo4P3XBeXSniTKa8CMcoT0ozRyErDE
5vypz39tvkE8ABWNT9fY4UxNtbh8IuZeq4ppECjDjYbdssMievzfa3x5/DNXdx6F
zrMoRrcdd9swzXwVn0q0pSzrOfstReTwkZmc29ovl5Fy2NcEcRMsMWooSbGb+/3T
vihh/a8z761852Byang1a+XG9Zf1sVnsUKwTkRj8sNKoAuq3p3WJgrfY+d0hkJEL
KoV7sFmXMXJc2CU1bmSvT6qHJkwcWzpK2Lj7U3q7MJozc5JOAe8Oeeru/aigeyHy
VfWLAD+xF23y9/XoWA2C49qYE2Yk96d4on6zyJ4ZP4uFPtWkmxOJeEcf8lS2hxoH
JsvcQfg4Xa4+LJJQZNyDfiuFQTtD86IVg0USfyPSxgNokZ55OtSN68uVb/hVhV2D
3+sHs21Q/zDITxgAYjwaQ99T6TFoRooj+FR9FAs5A+sK1wE11+DuKR1Nzg4G8yNG
THyDE4si1w8aepHklV+xSQvEf0qeodHh33OiqUT+NwWuqyMIEwezDO8lTwL6I6Ye
irgpngvQX7K8MO93Zp5YsHkpTfg9J01WIpYFz/fue5qf2zdOuoxFFBY6Dk7BdSCL
Eik8yFgs8ngXsKqiE2ORKeyMuTK51SaPP0Q2SlQA5IOenzmtIseYlb9u5uKVDen7
lbPRr7CcJSx31tj/BPw/6tw6W7b8Lj+FclKqDIRZPDrxpLyANICCVJDd5nYZc/h8
MOLTYgDo3S3rYaI6YEsICqWjTi2wlhxoSCAiZAibGHLOFQwmTnNPNyBz9iQppwAm
70EN9SPsyqViv7wJxe5NyIxKplAiM2jcW/2AEzebGxQZLPCwsmnxarFEWemI1pEs
Ak14zMeaP0Nt6XW7dKcXV4iQpUiSU6lkzP3sv77Wkhw4c6hCmU5ETwLcpmVnT8So
tV3H4e/N+Ca47gAMfPc6TDSlWbc4vqI1luc9FUEkHHDcb8rz8nbRf5TO99C532gu
e8aEsLlPnSJmPJwEsl2dhHUYCA1SrSQlofU/j4QSZDauop4DFla7VYjK0cURWsBT
F7Sv5YL9cnW5Iy55KqAEC3LhAd+8/MStUzGjg3E9hCas6jblTpaGDQNdpvI3vqrw
mH3Bfft/mlH11l3WPgT5yJ/k1j4cflj2tI1s7pcJoYS3qUFBzfNeVsfUoTklp1bj
yt0oPqu6M6CRAxmqNNyanuTYFM+ATmuFcjpfyyXMXwVt3QIzctKZV69JIPJscRYN
whkNPc7Hx1mQyyS+HYpkbBEdWeDrbANA59vxayv1/uH+eNkWJmr5EGLsXZT7zZAc
P15CmTUqdOzuiWHlOZFpm8tiZfC6LWwdwB5lhaMuJuX4O99L2IqhTvHXsABabdS9
nakb41qwtEBukMn/Dwvl9uUsEpt3I+NbFFMs5Va6UH7AxHnLoHix3TGrj4TGX+OK
iqZsVvN6NuxXWdpgEuf+O9nOopnn9Gme0nj8r401Ue1YEmm5HTFbhpjoARaXwhcA
/MBReXX3Jfe499HnaD9/iRvSKfh/SW2J2tJHcRRAYTU3Rw3eanlr7zoQkJuY1/mR
Txw9oXgd+LDmtH8CRWPN7G6vSQQerkQRAogwc+Wesl+jJ/LEx+VgfgE3DoeRvRAj
mE9WAYCd9/zfm1BKZbTGUchgPjhu/RRWZSsxTGVV6li2jOaCbTVee83ef/n8v6Xr
Ee3MwCcmT3mhvdxGAhSU3KSaB/ZeweIF3vL5SAqCY79Mu4AXFoGURx3lDsgUewgz
6WEjnYiFAWL81HXcjGZkcrD/cP0dxf9rfUklbd6yFOAmzgl9APwFrL5ZI7BIwu+k
ZT2uLpVgR9W5HH//0vsRKAIHmyQgAmueEKBp+N4zueK8jkvuhWHlxzODOLlyRkMK
mY5lDI+LtuSgGpxJQlSQIWFDTuIreUrd4vDNccqlqwKlxSrlui42rNJfvfmArx1V
4kvhCx6EOAn2Vwe2KHjsh9E7nEI6rt6rszAoWbR3kuDXZaTfh7HXwoz9kadvrTw7
VqLaSSpgbvupL6AeV8v8n02oy3HkihH27O4ZmqVJGztmxUvVL6JgHAFUmhc1fgqG
W1cXuqkI0bWM8Gh+mGN7Rvt0q7ILrptMt0h43Wz0hYsA/ztIORLP4fh3HEEkD4uc
OzRdzwTpS+WRVZL7XafvTXkjyUE741dwUyds6+dlC+cDCyuzcxD58uXjRyaG3cgL
3kE9+fombS8euSsMsJzSpI4kHIV7l5Y0Xhgy7wY0qnKyEmhLildTyqkC6YyvLk2m
wnmMsa6ASnlO/cMLmpxoIf327lxoazAKM6TAD6WCJ+r++hxr/VoApsrtldXWxyOj
hkHGRN6PSqwxe5RK0Wfe8otOUQl9wss1qkN6Ug+/d6a7xCzd9q6O2kVqiLf/CXTU
9gqBeSIN3Sbdput/79Kce5R6zABcM1YruWuEgrx7gO+nV+VfT5b20VG51i4f1Akg
I5zTCpcJUN/Qy58gcpRkxJgRJW03k7cPxlHV+aw0uNapFnrT0UR9NL0CFuJIw6v9
hZKJJlMNQxqroGGziY9FKY88zjNvIb53+W/aEa+2QKJAqPFIXZYV9effnrGc1AOk
4mgXoDjoYVRrmYzPsJ+ZlO070noCfILorR4lqTcigOmcv7+91cW2+IvWTmXjdSHL
aTTdzkoPqsvrK43vqpEQ+ZKKDwa1Jz+hENwqZ0m01SbQv4SbMA8+m7SdLP9zNVrZ
FxFf2BDIAWcMMIROWy6RIhz+w2dZamOqsOFf4fdc/7ot0g+CGpqXq5JdOIK30zrQ
MWLc/gklfH2CVufMgk+1lpjdJ+GnXtjCpM7nB4sucVioeVtYcSXb41+RcfKEx9Ku
R2PuikMmDggbNG30ttUugxyzxfHsbVOCvM1ny61Ys0/OcO8Dyw3fD3cadVLzcjxt
mbMxn5CZL/LupZ2dXZseaR7ou5dDpE1PfI1rHeJRdNIHG4Z+9HkkSHrP+etXnpaw
3u1y2w8gr63A72xjgQpEXzDeQuLTkAa9n27o0LEaB1qcin7hySH8pHdGx8p1hyAZ
dx8GZhoTO0TpJ60L8qNAzbE/uKC2AuJGvwwxEhVyp55QirL2iJzrE66F+aDaTOZ5
ZAglOhURAPVF2G/qBpyXsXCscG/lwVL7yKwfnI6jQgTJbq0pesiZDXJDMr32SbPE
8+8OpNfru0GhQw0Ln1IHdcs8TPhRPvhv4bQSuDXMhnEj3+lBuYz0Sv+TdKE+uKRF
7+zMofGk5MnINOH8ZwYCa1YSGGm0LxHlt1rn7iCZ40/ra0GZ9u/LGqjGlpu/6cfF
Iqtoo6mpkHV1jz9o2cfIYcTUyuoL+n/UtrlGD4Kyw/6GNm6AIMlGJedZoYsYlfy1
dQVuZ20AuNOu9nw+1WSFQslaQiU5m9VbS15dOpm/0zZKuXCCtRRmRdrv3gFhBuEc
5BMYaa4qSSTeSiGl6kSW7HI6Y3tezC9PNUix+ON2S95CzPw4fRu5CW+ozOnXdZrF
jCR2ysG3yGyNRTlyxw1CakxT15qKhO8lpWirvekELPSUZALNHf9bb+1qnQ4Ra707
0YysrLA51xZMm9wIocyLCVzZZ087TqmULAU8FS3reIkCIt+LAZHwXjGeJWz9hxgD
FAfV9UyWgF9rJgUNC/ohVlxqzJr5M5DEcaDVUWaj0fxAm1GoNO1Q2b6JiM383Egy
4sXv4aUag4FQ7PmygmgrO7EMFSznOygK4szS53g7Y3jQn9WuaJfOw8rq1IE7rxsG
l4Zcbu7QYR5p9PzAbwU/zhV2uSZQnB7EstjPnPSJh+JHVKBek1KN5YwU2wDUzmNT
x100AJ2q3bT+gFk3VKM11/XErM6yudEAJskldzKtv0eFLjP1yQ3dPGRZ3RY/s62/
HySzZXcWiTIwNtRGzCwUSENAoaNcM6fCAWpfjyCq31DaSAoBchELbL1bRXohySTi
wUEAvSTaDlwA4nPyAqTeMN7iWHG3SBWchsEHo2hnTnxLxCYbIP6qBbtV8EvCWaYz
Sy9WOBR3DDytxnto5b80V0IcxGlVz0Pt6U+SZyQhta9thz8G+MwbCRo9hMXA1egc
ud4njw99ue5LugIvWg78MyhZxxoY+SWQsoukwSptUZDaznzmHuFs6tGTkJXQkeO3
730v5evzDXfBUtrGvHzJcxKw0YcfpyUhrJCkwLqn3SerQb4GqphdY8TB7MkCn7Ga
VFZtALe866kE8LAmCOj8XopdgUXGsF4yDqKjjWJdEFRmWEZ0YZUOCRaUXGlReUAw
FXjxwkGNWaTVL1SGLwP8M+QNFAlMDXBhLNMijB0pVZ/mHiXMa2o+/c9lmpgycxCG
nqZmd43r2QB0NWDlfQlZrCob63WUrME0JLft1n57xdfvPAORRB8lP7HzQM5UHF8r
Y5xeRfB4rfwxiJ1CmWJofQH+0/REm/XnqLqhOvmnRgin+CO+ueQUVlr+roYHb5hH
6nYAEvGFgG7v9Pc4x7qEhzmxds/urOgKpoS6WfES0pd9+y4BcejYSKktizXS6VBE
B35R0GwRa5uhuoF+xBqyBGxEBSJm1DA1omHeU9opXRPCXhnK8haSiwXCCVBucafy
OCJTCDAWtXJGca7vExedATz9nYY6pUn0UE0SXdKTcEbskz1GEMYu5xvb5n1X8/jq
4wt4yqY7ZO/BoimPyh2CWxYMJ1d40iBA6Z05Wpz4D6LCJ4/12TP+mIqEdlUuRLF7
L4fdCz0GCxYGkqwPgIqyRmt5tDOAKeAwmFUdJ/YfZy92HzAtMBjYBiZwA5PMHlWX
wj1hT9kiBaXz9NrnlU92BUfC+jb8QONT31mCnPj2Rm4mXJTPN9OLtzN8zRkn1VHh
wUXa0EmOduQIVDuW2f1ac2yBWb/r14tKcJoeeIL69AP474XTd1sC5PWPCs+kivCF
ASDorGPHNLVhreveFmxR/FFYhNIIfsbk55QufJ99dgEVoym1WF+aWkpNBYnXaRkh
5lEoiWiYBchQfXhZMSzsTTdqprwsbGyNK2hauu0wpmPHsMZJ64UulfXHYMOoVpzt
D60z7QDJmbpVoFrNV+jZwEeAIAz55TUXuwTZ+sDFssmbL2KBCSBOCq/FrkAjtx/O
SNzA4kkR3EQcl9B0sjm9lgtMn36Q+r8UfgSuZyA+tG+fHpaeCGrkyEtPIakygv3T
eD3K5mZEktxG7bonpFBshrd5simsXbAiy4xnzmVJKLqCt1J7q3YeZN8kPGKy/qqr
7b1tzabOJTlJhE5jcy7owpNbFsOeyqJZajACYHPl0Pn33dIkkemV2GZnraCDoh5r
G/kG7b2SYMb6dVRTNFmYDH1pNSme9fTCKycrrJrXJzjbTDcuAAIXGtlOq0taJiOr
pstOm/Uiivf2Of9e1pRHG/RS9HaM5VHYPyq4y24QxIL15cM97YHV1XdRTilo8y2U
ZaG2hLHFUchBAXXNrbAGYDKM13qGnz+HWLlpmiInRRt7oiU2pWrwGOAfDyF5a/jh
xh4iUDTOSfycxbILAIfnU6/jhrUVIza45836X3vhFbDh7hK8dErdQJHIS7Z59Jeq
aIZauv38tATXBUfSeT9eBvwxs7TzrcVnu+0b/1OGZRytCwcBLOsejlQ4UWQc7d8b
sVzcY+b3KxihNSqP3tTJ/K4eYVqj1ZTU94wZFr9TeHaofctggjs2Ms73secQB7KO
bufgKKgHau3RvIWzshqGgN5PIOpkwWER+FPq25hwDfinAS5b+7BC03+jLvxJ7R2c
6CK1Iukzk63s2Bvmlrlvz74cre6RpJAvnD9hcy3jZOIGZ3PuKmdpWj3Sf7C0dNvz
sO/Yx8tIcXzB31cEuKtAwaTySZqBSfCcaAPH4V4Hkk2JLaw8xBtamL5VBjX/xaQ1
GjPZepNprfmZZcK9uXYHJVj0ptkww84CC3YyQ7f5wWf6771992YY7JkzeAK4TAUt
OQtoTUfy+xY2Gqlgcrm0G2rMDwWjHoCma0/5oejh8pJVLp9YhQw1H1R1a28DfvSf
Zy8rqydmXJbVS8KFM5ca5CE+vjVpRDj8E5CWxC3herPWxIEB+nWufgcMAhn7bURQ
cza8hDBG5u1zB1wUIzshNPecmeOWJbDxps1AhviUZPyK0IzvjvvSyaue7lPGzoG7
WcO4EKnFvn1H+1YtiATaLHfRC9g6tWnmxE9JH/K+f7ISNkI5a/1sAZWwWFlPQf7n
NojAJnWOzUVpIbk+RvreE5wkGZ5mMJU6rvHcn0sNsomeCaqx6wJ8fV8K3FhIiI75
uM9I7LleSmSRl67CHYJ6sKZA2QlkhJUnnW7/Lq5MoWKyeyEirVdnNhnXaMI4n8LR
TFsjpXk0YvibioyeJ8ipKlmILmValC418bNceMlylWxCgyDs1BDTysumysQjgGwI
dM36GCT6VhuTQAVn29gQhESV6UReucFUJKQyE5G/LasX/n3fvU6tWFvM36gnFLRJ
/wt2+tQWH9BlYbqIFl+XEdfmSsFWI3a63Q7iowfHHHl8bw/0DVDucoxdOWkCp66u
1/wjRIqg7Eq+IAjT7pdwHjrUMnyrisT1GtJ6t2EIY2aamTQjTae9X/nLUAnj/1ba
oROu9BikA7VCuYfdeaUOagqeFABKTCFNOjYhop27H8fYcUtEq1j8/OAz4hN9CgZB
r5aQ0Gf+jU71FbxWPA0n4gmC5CjEYir5Ijc29Rx3xnPQUYka9Ymr3s0v7O4Ek3F8
7Y2dGxfE4uyRyV9s092o/iZgUXgJP7PEPRxdGI1KcICGlMvblC/aehR0IYoOP1ai
C7mG8kJ4MyOrdzrNIphmR8pDLW6ZvUNkkbvnWpC9/rsuw75XG+KGW9Na6XQD+C4k
0qAdDhiLq8VcmDoCXS0K2KmOUKTTv99Dvg2G2GMdehkLMiDJHpz9mWBvJHNe6zcX
YKiLGmLGrrOexWzQT0wRd2Dx3eTi5bghF1+xSWoZTlJOFcfgmqXJaMU0Box5l9Ix
5twmgYyvaDf+7rwZ9LENwIwrGT+Bb5BpQ+vna5O7d7S424SkH6MaVCWZIZAjhmZF
0FC0A20p9DFwLqk6qB6jYC2vXvn8aoEtvfSW4DSuxWP7Wj8rq4wxgH+YjoRsp5ME
UHQ+Wb+aXv26lZZFv03p4Fs15iBGmr0/Q37LF9BNPRoRdfOLl7owX2qL4BD5p4yu
umLBMjwWGSjOgGRGVu80G2VzxnQ5n1UaYXyIi5GMeSAKNPFvhJy5OMhcn115D9pT
hGE8tIwoTlR//MtUZsul61MylCi1NYGM+NDcoZj3IJmCwjBp9Vsp/9bnrN+5ZhJf
+X2QySRhcMKsvFMdfpC8wm5zj6fiAJMrVlAxmbQPH0IGOJOTPoByPNJ7m9PHt1im
9d1G68zBBvGUKOy8Dyq/trha9osaNQPs+Pg5q7+tXefGn6ScliIHULhyD1VJ9QKp
gYtNztZsW/eiwNccQVXXZhKSlR11AzIThfx0mFB7tIBo5R29Wkm8rUyXYKrnB+JJ
H1vOvu3KTJNXI2LYckZIvGsnVLNlihIEWXA0ZTxpvT9PIFE24voB/NhGxLEdOHVP
MfJVZr1javfnIwiLpuso6CE1A8FMo8oIx4RyHlcBLMdBxKIgaouRlAzPD+sMzEcX
FHBHTfKKqtCtBYW7W9gcV7+RdzJuQu58vtQHn5zPm5iAFJvXJ9H4KulcDplgzY9A
3eGk0NFGfAxv1IShRnxyhfAbdGPd+BLvBXSfDRHqAsKXHXeMigfp3GEbOsJAxq4z
lNu+sng4dZ56T2KPMAc632ODsVBvXDgmYTWokaF7KOqlv/qyT4sG4jiv2XNI86Xc
JpUYWgUQiIZQl1ngJ6fNp8P89aGzGILSjGRT2MewXAKZmTc3zAi536sbElYpFdo4
r4rTbYCT6zJI7zd0+qRevGnPGA/uDeQW7YWOyQu7AwYdgOTE64DAbRApA94KImL4
xpFX6TLwaXcOV3HBCGnH5wAQU0rNB6GU7KyqAPY6TPuqBAr9fMf0ujGMd/G8HwPS
YVwKrfkLEimU91nDXSfdcpxuRdYbqJj2yqIGGS3z8lFxxOgxVjZpN43d7yqqG3+J
4Pezkw9AqHogGTcfGNh8hqs+L6nG7jWkM3HrMqZY6DnX6hbvHWIOaebZoPjE+YdE
CZ78VCW7VADp7ogaSESrPA+CCGSPv9+2Cda9EbHX08R7bZUjVzt3palWrgFZ6qX2
QRYcv3cLsfdsOL8nyH/hFvnodpwFv+GBMdWuIoErHKkO2NQmNOjsDCCQMajXfSF8
b1OjlK8mC9QUN22NCwBXyPLUN3AxPSNDwl/QNgDlTy85Futz8BI0cteFMpZS0WZE
DqXqYykEa/4STWfJ70JTYj0I0iaYOnkXkovEM2eD2FpYvPXnNsFehilCsBIO54v7
LbBkKyPsstIFKl7Sg9kQM3tIenhMdTkvY/ZbO5+NlxJSXjDfBKjGFjUSfA6/DfuD
HC92BRrC2K/W5ppaxz4DrweXSKwLuEDUmK5znOpawv10DzjpAHTF8h5wdVetdGA9
zPho+bKXBq02QZHjTcEonPcQ7xxMb9fFfIF5xVnMAxkuOBi5wrgIoNTSRs/qs666
ZsBl97iqQM3WNg/wwbizkwlRdAr1odOvtwetmGNJuDd14bbwb105XNoMbZYzOtKd
I/AFSJIjfn9TziwKHtXx9plII6N+DiDCQaax2dNbiXsYszxUuu7LDpEO06NWyA2a
r+hui0ODxbaFwdMYid9dNqGQktbcxYIEMICcKZyL8VIguuUchG/pX2XD8p3q/oPU
LfNPse9H8om9aRamrNQuv0X5nZF8M8X2JKbFTTlkH+NKQQvt8xO5lq//VXMIoCsL
FoMRMqGgp4+SFo3jU1Zci3BgbK1VwloBBTOFqTcnKc+oANYJsBf6h7+T1+ChO1N4
g/0BSrZyMOb6MlfMPXRgKQktJapoPPqpAOUWwp1jHWUiIK+RGrIbrjAs5+SStYa8
SGx1wIzPEgqKHMjI3q1s0BxILO7qNA7Y9xrneUoFfJVpLvXBUXsXJIXG9VGwG0tC
i7QgoxsbeYw7b0jcKytak3zZzOW6UY3B13N38IgC4VrpbFZgG3judHw60RRtUnFR
rp5ijuOVE9PEXmSqaWXS1oBzsMhFaklsHQEUMGufJ4QcKcbbe3/WhboOcH78y/1O
f/BZAnaFVKh4U2ME9p9wkfwkfR+GmMNAergd0ngmhG8W2uA99QmPKMkh/uQt/ui5
BahueyX7M7eLcbptOsuBnlopxIS6I3o2FK6gI3oGTRDSElq7ZMBY/scx190aA7mV
h+ejFjLCDxpLEdx/A9ayNp8Qlmf/d8XHrV+MHQYYqLoiWzUmZPkCopqstPI/UB2d
4b2ctA9Up1gokvgwhlOtzMY3Rzpv5Q+L1z9sKAb4I+OBu3bImH6eLPVvk1PmSzd9
l20sjt7rBmSR4cZ3xF4FoK3X4HYyq94NgJ8rYe4ImwtzjK7HBEGFt0DlS8iiUqkW
sa0m+xxVNbqurf26NraPURvmQcNn51vd/RNYbYeJkC8wTqNtcNoYcUCVCwherhFt
UzF3DznAdz0ynhr7dTIPgQWk4H5mYmkHYmNyiafpcvybPpHd25K02cJSidDaIKvi
chLl3Y/31d5O/UNZj+KLCVu2ryAKGB5DZuAKocASxgxqzZ+OpKlnSyWpE3Yozny6
VPQnI6tIy40Kqeefo5i6j+TuXEvE7ZyDkOGj31Frb2tpDkr9TuqTNhjzRbOYuKjI
DcSevkoFtnmZBgeWMVZV0WiAN4Fkr+OitbeyzRNFALdJgMbTr9oxL6C9J592yBIN
vTYDitV2hnUqtyFr4RFVHzoKBHFOhhYeV0QcH3QBECRWI/0sMrjsjuGbitJ7pPWy
Vt/V5Lgq3yymG60bS5ThGf5GFowBSz9+kwIguKno45rCKKhIjaXtUj5atmnqnonv
/w4rhznPrp1Vaf6F6SUeWNo8vuzo6ubFAiLJLMQz0sPyYc1X7tl5yX0F7x/8RsGx
32HDiASjK3K/jthLv8TH1GYmzUrOHK9xKR1Tvz+R0WlxpxId+e2+BSss7bK+u+i9
0/ZDoUf9U/r+uWc6/yZCg4hKJmdFLNN7qAmE0+Iw6k7oJw1RiD9YuiCD2NTNkE63
gB3OETefsFWxMYo75yS7vts1zax2pBiMx49AvjdLUsHSUsm67maR1bNLYjIZTKJe
B/lhnT9SCToU0tEIvv2JqtBzQr0/Y/Or5BuE3wGb55DdGgM18P7nNGV9/ubwa6ai
OcG8Ny6FdLnnpqXsh18RtDB1yIEUWbo9US+NT54LT1dQRPF94ncVX2dGj42jslqX
MP1kyn27GR7z/qVSAsMSEZbboUMknxEOKq3JXI+2+gahxC/WWG1J870kGv9XVAmU
R59y6/JkzoRtlPmZoY/1W4+/L/HCt9OB+dix3Nbp0+wK1Hgy6q9eRX2+dNFpmcOX
FFjpY8bLzZ4NGsgFChcRfhzXIq+DYdjA/MBUriNhOvSq81Fe7U9VevFpVF/gInSk
DvXvNeKjij60Xu8GX06ORN4iE25iC+0OFba7Ux1l5yqhGU+L4HAwRvkKtxFrajUT
PORfni3CIQvwqWGelLYqbC0hMgfBzUe3gw1td1sQyDQnW//VIdl34tmPwleV6SSE
00S1OoGGFUR/sVIjkZsh9VAZBOJ2KGcy54FWONuc7y/ynLodfR0Fur8pym2me5j8
xsIy4p5Fr4zsdqYXTAMoM0Q5bvKs8z96ZuRoNgGdLKxx5Xw35CW5vCFhRXiDj2SO
QfXZSoNn0OjlqOkgxsDudyLIhxGaJ4Ilkgu5Bxt39ZGcLODHzPRxMSKwItTWOQH/
TAQW54Ri9gJHBRWWxJP/28lFy9bOS0YGfPiycdaoyObc0hxrfzaANEZBrE5va8w7
lHT61yN54B3gc77Bvbcx82Y0hAjQ9pzJRKKNW1iUASEQ0tC4v6AI8ATMGaDTmgXi
yrhTem3S9FLBOi2Fnhyx3BsTOejW8lUdDBT/Ys26WFDUmEYaJ5mexTlBbTxr+dV2
1Esy5dXt+woqRbxmqoIo1i85IDAHhWQMCdtjPL4oP96jfAaVS9viGoTIT7sGtS3V
Yg7rjULj0uu48f3PQqJY9Uu9ycCSxCJ1tCMMt4Co1FmBM9XwCSvQlonoLtmjhJ6/
+q9yLtLX5LGM37LxY9y5iQhm0Ii8HSRQJE7gFHfcgxTSIMi4Hr+bpxWTMOVNugTj
/jJaWZX7VtCyaB3gEBUD93vCF+CrXpn6+cD4bFA1JPkhCQZH/XQJ090dqH2zWWju
y3SeI8bQB886/S5k8/buIkUeb1GEH2waav0LZP9ij6UPvAfSBGC46UUraRWdvxoY
qsf1Xj1Pi+z1rxcsNXZBgVe1o2GDHGcP5b5RxMx4cIbG1oE8jtvSCYaEDdtwlst4
3Hi27URar/za5hDVWzJscopwF71LgoZFcP0tLf7R7YFUctRug03ghpYWa7edC7rA
Grl1QEii3kzIlL78TClFDjgmjCLgc4yrlL8C0r0BOqNe46rJQkzxCwCdosqQBCt8
W8kV28C2gEKUFTgJik+OKfDcpuCaaJazrYJWIr5SFbYZy3bOGG6QaRbO/V3Yl9Ty
yEH3o/3D1fqF/16M+PCbGQBJUHYtGfqNj6/L0YPemwJOzuMa2yoWnH8pbIPwegKt
9KPhVYVTr8mFyL1jSYQkf13U6LrtvGDeCBTxxyu0kDPlhgSrbvgj/LCFovqSSzic
HMKQBWnZiN7OnV54F+DByuMQvBLl2uRV6s9jKWaW4whxYTWhefTBi5+ERGkckUgt
NS8rehEb6tfHXNTRl4oucBmT0zQsuF/7RINaGv/h6P9HyeaElTku/+kDcBsvu5yD
38mutxy2Z37HhUJq7JHABDLRDwz1tUu9pxvzNv25XKe8jcFi2Y65drWGUijEtXTL
OhHEdIbs8SMGNmOd7+EL1ctNgqpnWNyzJRd/M5Rq2zX8LSQhiMGJKbG6PRvmcveI
8N+uvGmkCGdNtyp6IXsF9epTvC1GQ5P7KnqvOFBfvHwfCnzCQlQxacJK2PSWQhd7
XJC4J699+82gx4XObpbeEx8cB7feBh73ZwhYhm+4coOqoyHRnPGarXN1vqZP/Jcr
LPIvGIQfH0nlmrO5W61VvDp6VYp3KOPVM34hzV94tz2eqqFZInRuFiBu8wIsKMjE
TnyQKAMBgbcsj9JUjYyVnT+Wjao0nkx0hIiMkxJnKbS+mdKY5cbVzIr7wDig7Fr4
byitF9PGaCT0ZsNLE/C8h/2ReVhclzC9W+VS2j2uBs3QrRblgwbbZdrrEPI+u3bZ
m4UBXkgdXmiSF/aGuy4jblaXSCZcNX9lZp7XFVr6gKhRL/BQVrBnw3e1mxf5R2Cv
daOzbYkauCfOQ0yE9IdPf/lWzILpaLGj61xmKZsJV/KSRHBXSX8PlDv6BLbp8eJb
RFgY2sJZiD3eSB87LfdhBkikEiiMWQb6qqGzHxle9jRlhYxxfNkoYohWEuBzAre6
QZkPyMnN/Vjwim7zjCwHvS1NOKcRqqQXj5yeXHotQH7CvdGjZyPsbhnbc1SMCbqa
YCMbp9W+cwx+LzRqzblgZxokPPC6Oh6eHEPvuukOuUO5mrEJy/SW6wsCGJSSB0PC
sRXlVN5f9AjzXNL03HcfpJarqhAOYBRKelz8hGsAvThE6oNS7b6ewp88whFPTFez
99oqHUNNGHXCRfqhGq/eJONHSmfg8ALOKhGwqRlGlxx5sB7C/lw4V0Thc+So8Fph
oLzK1PUX7Dl7oDanh6LIU2CMoCgWsh7za5WWUhCopwmCIRM2dganmacvw8JBlmi9
AfbUscN6FbF7T4rmM29ATdaiIeJpx3Hj1n6wWW5szLKUfaoqhe4pXp1hL/csBWix
tzUKhs/fhLFd1GKzXBj8Z6c0RLgMXmVuVt3PIPLUgOqVYvHT8+r+wpPkJiPKqXR/
yt3NGLc4LvFhR6cAkzxRIXMiXP9Nk9LXFGUZhIWStklleM20bFv+rVx/tjj4qPog
Am/i1Bt7CMqm+IOHUQcV9+KvMr5e4bDp2IXKTD74HBWaBsLDVSZkPBxBfgpdhH/S
V+VFNSe6vwuITEzzYeekBb5uIGGYx3XgVHYe7HrjEJ4ZMcSr6dJGLnrmUUBIMFM+
uAyOeJ25/Ph6N/ODDlOzEA23MtiIOcbaTMvdVGSNwlOwMEJnfZcdGOQ6PpJCpOYu
JoVLFMao0F5fdy8F/fGnFHYViNfZFs8f1IID5ZyIKRROymOZMfLdc/EUSO+p5wzt
aSs2T/M4gcJIxhHhIPWM3xIu3yInAs6Fm9cb8RWxWd+xSvEVAjeXQgNvdhtKEVwV
Wf5E4KarBjHwdDy8wu4sR+4Onfpu5DVX7wzTz481cP8o0Ko8iQNI2TF6Sx4PKrcY
3xPufZgXhkAMr9uwlG4tenZIw+aSK2uVD+SOulP+UYNWcygl1QjAfNlVsJU+Ti/J
N3wkKEOsbdkE3wKjXyLGwWl9s1gl5IsKisnfgOC6+iX4iuh29LjQWagkaPjfv/f7
o0VYP7lo/Xm/2CcJbMVu0ExoVbqgieqYLWk4WjxaA1w146Hf1SVnUgYo/Xrvq8Jj
4Vr6ohUjxWkvfYXrl96nYnJ9a19BB7BpJYDZyvvWyG+o7ZR6bxP8F0kovF/TPzeo
Z96+pOyxKWpdpcSaXGj7qxfZ106KykS83poKdS6PPGriksfS9GkWeE8hN7adR8x+
ToLh3zF4IZIdQ64GASH1KO+QMW00/eBrTMVHEA2OVvboO+j1TuG6bVth3efMDfip
nVVStMtpHz1KhXjmFbPOGQCCCQziAa+Z0WXNsD1w7e7BpOrPY9A6GTL8keNh0mlG
5ZK2FYCdQzZZTna8nA3G8wrvxBe5qXrozriHJKWP+ZHVUxlIjxStcZOD1WPREpYC
AvXGofBgWyFQ7tLctN0Igu2sGZKVLaAnUiWJel/mHSH0OhC3saxl2BB+9wR6G2xd
e9+RSDckyk2/+LrrPRCDDRQ8CAxLLRob7koOVoFCR0L3ZCDv7lFu3pfSMpU8Zh56
PmDMq9/JI59qdZDvJCdj708pbm0b2tKKnYvMaP7WhN5MA9cVLBaKQbq7DDq9LkeF
BnomX7dkcWSKM7MxRK+z8FLUghBdrg9WbkLG1K0RGCcWuaRoGQ+iowmpwn9EigcB
UvKGpAhmQzpLf4IDSd80KWeLq7K2kueu+MH2mEeZSonSXntqSWysHYybN6qH+a57
zcirWAoob+AzhzijEv6PVvRaHHc6u3F6ncwsXgN722SyYhPR11nbrob7AwSEtRx5
y1zOY6267N+183tLuifxWous4/REfnhySbNM1Y8kL75UzJwYulMRf8biTRuTLQNW
ahNMxdyvyUZI0Z02WQVpSHuPmT2j1fvYr0ht+unl+1JO+x51zRGjgl6fYdEHs8PP
gl3/EzUiyellOHvKMV3hWf93VSKzuz/HIrkQcsuLANS455hAAaR375+vQYGq1rmE
BoPYRo4eYIlZxZKZYqyBs4mVdkSYC723ARumYBI2BpUlgYc3EM32C2vJaqpa6n5X
06j0M92zuKbkSGG24PnIU7z10TX5wxmhY3eUDTAAJpRLvL1AsnYGDIe4fnZaYbFH
O4R0fb0B8WvAtIdA7tZTqOTTCtHrgQbw9bEOql0l79Q5ZaqSUzMTeSNS5fWvXdPn
+P/JI3UhD30ojmhp7gzq/yKkZGG85hQZEYnNLPh+fh7KrFUG+x1CTLmFxplrykxD
rFHpcK4ovwK+q5gR7RU8lYGrmIVFZ9TFSkAWmwmdUqvl3eINlu9SWTfaJni7KnVf
R5gFOMwnQH2dbFsX/mP09ptvUfwhp338LtzSGfbs3Fx1PpKNCmFbh+IpKWRm4+av
+zHei13Dq2o9jkHMBE0mCb6vfdKuYZDEffJsC19hllhjQi29IOqSUr96IxSOQ+zS
I5Xdiq9es64C7TNjG4OHwWMe+x3nM2y7z0UNsP0ptlA4LuSYeL+wQayyYUlUOttW
0Y7kMGqLfuqD1+RYbvDeU8cZomhLbSd+1F2cp10S67lIdwoiboQeDPUDRv7lNJk5
ducBSz66XalcuyDQxr2iQf2PGrEov6DwsoTcgqLIg6XcjdIK+LCqdkzdo1JOBPG+
EE6LHu/rs27im8zDBFptGYYr3pqG1NsA/r2pWc7bsixXHcB/gkL6hNFgFNRpOe1w
IFFq0VBaT1kAmt2eRjvN9wF8/5Vmr6jKGb/8LKpQFIBYx2qy3tJdwIKdmk4I4i8B
PCmYu9hWZGp80puk0eP9PMMVceNMzt020cLYfg3AjkZiGDK27H5RB6eJbgRZQVN4
vESaVn/37cOL7YXTWtBpsKhkcgP0TRbg1W0eJkgXswHyOG7nKqXzNNmQzNCoif6i
5TUiOaib0MGiILIT2U8UfK4mpWCm5UhagwmXLlsE5hkwrmTX9bOJLGu7R2LaGLZr
NoE6l623GOSncbe/efgj411+T1S/4stKqXTnNmc8XX3fWEJWc8pqaxuXzmLcJNzM
vE+RiO4wv6qVl9FDEM1nlOYENKuUD/17n0nClmXoLq+naQWrI2hsGfHl0clXpH/y
A/IcDvfns5UdcXXGjfqLwTmzH5iKI9Y+A+lWLZDHEvYuhUL5JRxT6JYG7y+be7Ef
vg8ESxLm90OHuqDIEJLHvJR0b/zo3JcL2S0/Q9w1EsIF9YihXkW+MKROZYX2/Muz
tZRbo8pC8yPty/dcDM2KGKYuJS2Dj8kzSIPTLjakJCelxKxZJb3KPwZDfSF9QWa6
LXRn3JbkADEnaBc3Sk+uwPmTO2WMU59O/Tftb1hM4wWOcqWNLbLaEGOa4i81lAUr
rG4Pfvru2iDOG4lNcmm70F3KifCCPQ2rhIh2ZCEGmImQ+kEg+ZnR11PkDRJsdj0t
WmzraYdOkpNMFgqHvpsRD55Og7+Qu6BVkprB1aPvoqMg9+X0Cr0R4TgWaqW4N5uy
Mnyar9iRwD3dllLGTKzHp5WSfxTYlA3cQ/+vz2+9RTGY7Btbjhgfzs7FtGQ8gpEz
z3gjaLnSzhduKk9Ram3muSC/9oSenXyctD7/kNx5qUW+u0k5FIkqWCr1tmz8Rec8
kzlNMNzlCdcBBukLUZoL1oSPOAja+6oEKC92PDFFmUps3RO66nUP3p+8nrTU1DLi
kWflaIdz7Bq215mDQoqZNMJfiFNg5mO90yR/kt7jeh4imGf4Ne1eN1GHvrOh3w3J
r3U81tCEZ4/i0OLcd1pPC85LLTJNpm8YRpxrI2RAf5B0qbmAEfpV3tYX1IWJ6S+u
g0MJAxuK6MG7FwgDFcRZR6iRZyShc05LAqEm7m0MQK2PW9ZMQu3sbZnfoi6iqvUL
l+Y9OEilstTXN6/DNXci0+45GvkvZEJhSWQzxcB8zy33sZGGZYMI8gmGy56HlX/Z
eXr64rG5EO6Y7dKdNEdHdKMV35hCtPZkH4vnrIxVbEHbkEa68kgEKhRcUpKLJwQk
jY9qHoPVO/vIkS41uQnyqW9+DxXBBwxQfgbQ3CkmVLjtrn5mrZDdAQVA0C4rkxNW
E0YJj5SBYtdw8IN1sHFzsMz8D76Et+dfhCDnlXtYKSNcSLR0Lbu4AR4EKsJiIGo3
gEaBz6TsrCVLnf5ejIKDqnlkLNqg0VvPMvKRTva81pgSAF6Xno+/zbejAdnloAaY
6OzloxZro9Je9XzHmOkL07UM+uP4pfzVi/AaAINcQiXgP2vhcEDRTNR/JnCKVU5E
fBKvgo+QGClv1x+Pf/iUTblSim2NyAmugN12QxaEk7UmyBNK4eqWCo1Ok8xvA55C
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WA+Q/F2r4OfxWXjAE7bNm7CbLjQ5DMoJA0AHmTHVlCvuCnh/oc2dcIwEKEyDGGdU
vBOspG/SoiSX0r9JiDIev0JgvgKoY42xpZicC+oS0XmdSNt9SmlMI1hz6OqtvgbB
H4HgkSepGEpQOy/sS8Eyv62KTr1uz6pEbiqTDUpQs9Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
Q0MCWLuojl8yJX+Z2G/AAMvmsJ+rotBW0IghtcCDflknXFw3C3d3Pwd9Guxm4h/0
oya08sR3hk1Y4xXUG0lzB6SfGCj4H2+DtxaZl6KqySPn4ZjTOnThA40+yndfxmyV
DTBMQv9TmnT2n3xm/AfoYz2DzrwGG7M4qbBe2AfYOHTpw6eZQ+hPu7eZ8TmJtl7R
nqEo52/n0Xu47kQxGIrWnLrTXK8Y0OfzUo95tZJjEThfdhDy4qnZe+yO5c055Ge3
cIlrWA9fZTfGPJhP2q0pDcOj/dIhwYjgIXV8uJGiJYGvpI2EHLAkyCD22DEOZaRu
08mXqxm0PkMA2CvmBkY9cctdTcCvPYTd1Q0wWNSOz1IQ0V8xF0Ci5focy5BsC95/
8O3NtrMLg1d++3aEotkhjVqAyJPL32OtA1Wdnh0BILSUqpC96hFtkk41hPJLemJT
slexY33J/7XUewTjRMX9Bj7ODx/b9XTUfxZSUHoy7ih8muAG569KUFFPBGJQ9xf1
s1UJD3mR/LzFqBd8LJl3ds3uP6TdgFgRXp7g3mKwZ4ck35qVvMIaTM+nIbHsred3
ZVcwNfh76oIRtgCpRar6pWngkbpwLqjQjBtdZmRP9iJ+xxZ8uzGHSUdtABINL/zv
6sjCKXJt5Qk/JimWevsInkYkaIsSD3PcCV49FKNjC86gJjrZ172ywHW+6y4Pam7s
1w1nGZphRqn9Xjl9YdcSyC2UqWRkIJBtb90z2q+nXTUlyu8lQetN/Xaa8m10StE6
zX6sKZ40s5hoyMch2ow9uf4vLp7rD3sbWFsHXSzpYzUvG9Yz4+icwQOw85qv5umj
AwPV48aribCo27AiSyG+SIafwvAi/ErW/2ul2PCbOms9aPlNaucxPJzdFfX7o13i
D+AwVYTRQMOM/2KnLHQ9JoqKAoFg/bviiKAAKbBbZ12HomXGConPhtYyOg9llk0c
edf6AFfaEY3JPQZv1cTgKzNoti/qJSNBWJA4mN6K0etW/226vL/zOv6qo+c9h4l2
2ofzR61qVJ+eSvx33t82TopPl2XbVgHpYaiAvY/mWaybhuFqeq0jWdgNynMUJ1rc
wSEeJ+dcm3e7RGu9JEjAuxpPhcw1nJZuuVL3tioRrOACa2HULa1611wthEHc9mbg
Iwiux/4K0LFTi8NChzNGihES54wELTf39zoHtbKIHNtMwe3foKsyn3Z8hPdLJfhb
eLNOfyyoJvsZ8n76cQ3E7PL0p7OW/0DQo4I93rHuN2Fi1qwL1bE9hUX9MuhUlaaU
GtvA8HGcS4er3a6mafogM9wVhxyqqfz6IctCd3qzYSZV7BlU3dQpTy2Cm2wUvBDf
6y1R4IoZiKl8VVXbfyKMAyS/q5Id060zBtA4kVPsz98bj/nXv/HbTejIQjETnk8g
HrZ3ig9ddnlLVEadB3XiMm46LWh9qnmHIq29wSgTLd5Mi2G7r61FzfPPrlLfF22q
RNsZTcQ769xlUXkmOVgZPZIgeqy0WvFZQdV04lYQ1ojZmTnAnq8sTZeJuB6E7VFz
iBW1w4nGfGOPahE83MGPFYHJpTqr904C/kDCW+uQWvMGFe8RNRokrrsNTxlqj9Ou
25CSKlTwMZmHmjy3XvSYAoG9af9mm2vm0QtaR3mFkbPxTR+4BDKuF0M7jPD1EJTX
tD3r7skqOTK5YsNqkBBz+u3unvjmpt7DoPQwcnPQq8OyCj6KNzSnYhxVuEK1pIhH
zv/cirHkQeu7nEFR8kgFY1JIU+wNxa2zi06pd910nCYKclWjmWIESCbqT1A1qnE4
/132fIzwKWHUfc211Mt09pcT58nQQ6kZLl+FwkujEF/xLGtDQRhaqd8J9kLNzpdd
ohrftiKRuoev50xQeROpH37BBcn08/3UJVSdJ2c4wP2zI/H6oc5mBmzJswDxHrFX
IlUCvt8LJvrpMgNntz3THoK6Zdg7jZ4ESgGd8v4WZH47wAJOqutABhdJ4wHdd1NQ
4zHYqFzu0z5NDwmdDb2pG2EFakMMT5Cbhk2UCpvdwxVLDDf87MwCecG2E5oQWG9u
bNXAIhHssaTLhieDN6nZtz/1f0uXDSwEesXKvnw4nWuzehFdtMgwKW5NqPGRKAPR
hTcfpI3XlxgrkyOGzRVIyFMfG0ByR7XP5XlthnsREQm0IvtZl5wmu7gN+PfRpHVZ
CInbtGNlz7YJRayEQAlrT0BZfh8fio2Zd+Rs2/vo6vxGzW0jQ7zbClAjAg2DF+7D
gNcVcTtF6dj//lY5poGdta51nnJKsePkWQO5imRtPQD9mE4ggp5VM3AJhbWS3Pjv
xz8b2U4X6c92nB8ZOy9WGKr9ETbJiscHi4fDx9Db0GvDk46YzOTqYU2/m9IiZ170
bCEDALZilbNi0ms/47c8ygichjbyFFpl3ire1gGcpl/woxihzBmKd1FEOFYTFJ2V
z6ywcx6frL5qq/R25kHfbNq8yYSPNBQ/MRG00JiEtgFSDtCiNWdvKx4amPYkiVUG
rUDJr1gDs208nF2CHsT+vSJfv7JKM1wC//CVPiDV/bH3hzPpfqe1xU+AjS7xtP/C
nmOgkzpVhMnendOqAT5tQJDTLf05Ya3mRDpTGjph+rluDZlVDOGfkZHR//Vu5+86
+Tf9WmI/taSqAChYrGU0VvR/sbKx8eHSzK1isJFgt+aC7scUFIV05zzGO97EDyLw
nuGrrj+g8R89jfZANcXBg78nmHnTIVdjYgMqXLPLRYdpnGuWM0BMYh6qUg8O52DO
aI/F8LKUE81FQn7akcJeVhztdf48/xffdjEah2JMqWbP0zirpL7kTKDugnVsNGy0
l7lDFS1r0IdSFt+5LApg0bCcxoNLY2NyATGuAELtZAznjfz3Z1/M6ukox2KY5vQN
ijA+m/LsezLJIGPbwzPhnWCo76KxrX5jd9wCNhSYgphf7G5j6hqwKzZIZQFgn17l
II+iCNou9tObXOvuTSKr713zOBEjmdoAnk7j9zC5alcVo9o4Q0jA9RjYyIIh3XJ+
Ur+oEyii5t0LXo0JR0K//Vwoqkwbnaw5ZP7DzrfXLpfcrd7Jmei2yuw0DAW8w/S2
TIejFL8wYIT1MEYmKzvbfACS1XMJah0S2OALZ0AAaa/KPGkU1OBvM8hwD+3gpVz1
BKm8rYEt8v3DwY8SRUFgjecjat+2DkHzWlmS3Do3iMZkEg2zk+MlM9UzQ6TnfJsI
idTgid2zviNOBEaYBzdzie0oxgWMhT2KXb/0mdBsJPdiHkv7XtDjUa5o/nEmiCm5
hdsfIYDypeh0PDVyqRZEWP7pde2CImteFY/afF4vYdvHqgEwHmDV7DoV7HXXPIw/
e67+YG/mQHctojAPjTs1hT15jPDihUrpd5r9gfuwNSROb1JaJ3CYiAtUJotv60ow
M5/S41IDYP55jqrCbl+aO1j5m+uALJcUpc0h5+zfG7+K7EuXpUTCxEpQZG8BDxWy
ABVXHLc3A+qi0AddyLWOJbApvQaMbU7WWQS1xozWBV87UgWddGzNwPhdslmiBsnG
ZVVI4/9mOVdT/tXEnoCas1dhUsqPc4Of2ME8ZUj0e0h/R5qrOxOaqyoyglkh3zlw
83RpDvHRO+/5LfHk5mPcMakB7J96wkb2ZjuenfMaMHMNnduOUlrw06D0I4tZdDye
m5QsMLQ/Nq9tSII2tjW1sSBtZpZP3lz/Cedv9q7dJiKKdBccqO0lkbSE3TwQs1ds
m39eHMB5OEfkeDVyau5LJbH/9pk3CXdHrOx9Bzwn4J70KBe1NNchTFilbN4oxCgx
M4/uTbyBSB+FFopnvWx3HyNq9nTll15lNqZ7jI5kExU5QvHAbZHuAIa9kCdfbTF8
MKHgWbQ8WbaLxys0Sh8UuXUx4kdvu8gsjpHeA8u99qtwOMl4gr/B88i3rPRyDRyW
C6JLo/IFtZRae8Z0gisAub0GHcxZzjuP3xRDNSvJOoWJGSRSO0KURrs0ji7pJHj2
l0PmP9dQTnK2b+YrhgjbkJnfbxmdKZ5u4m3JzQ2Rd/ZV+wWktV5sW1RV2FpNYogv
3Pq5tUzNOapGZnVfKMUccKkkTJdzoQdpHCWOWuL36q9YuSfJO9evzsmbCZ8MJGUG
4MezfrhP6qbOczTXywkKFSTaIWSjZY8Yx+oIZmU+wK0VToAi3hu6QRPwa0TIrJkq
Fgt594BE/N8nLTK2D6S1ZdTApqvCJ0zXCAmoz0thW/dTZ8Kvlj9VIRcRTteLgHZ1
ud8MC2JVdEs8bVXWYTSnc0zNp+2iFiAowIAfP59GB+lSI3A9OjwuPMnbdmhpRRrI
1Bcj73mM4XQ7fGEB41kmnQp+Sy1tw96OgVrprScT9iesmxkzk/rPDtrs3vpKnshk
A5EGxiSmtHtXlsbEU7XTr5lgweP8y/rVzWceig9Lw8mY1gYhpz2ymw91K3RlyCXB
c5ZQsP+Qru+H7Gj1wBOzRQNvMUbfISuvg7NdOb3viJ8kJSGAzI6pXKk9Vyfq0HBI
y+LqU9yp4oNHPdkMm8shR3ipJGzmJNjJ3No+uqG4jLcBPNmDG1Dtn+tVyxglqhoB
3JRXHPKLjG5yCK+vjYC03iSxdO26vqn4GN6q7NFP5wxb/d+uz0KYnV/P1/2xiSpN
o7QspOqPT8ThOchQ2k9m/0eGgTSOlc4EvFuJ1dhJMk4Vokhq5Wbeekh6Mz3rIRxE
HX+yFUjHS1dx7lhf36S/e8lQeYoHkZrb2kPZ/PpPv7wyd0+5ZxRYfh7tDCsVhuHh
usAK/oJ5ocL3DO4qyK+io0nUUvTKO1mLfbxp6W+cN6HQxB8wDFgWKwulTbtRJKKk
QDlWBdKti6Wue2dBoZaRrnsCUehOv6wrmcoajU2dJxjeDv8Tsf1uLCTpJPx+XJBz
rvJ3tjSkJBgCVxxW4k0SRMKoEyomYxKBjDUa+Bx7OoD53d7LNHJZBr4ZyP13JN46
caY9mf0dnXsfm3Y7SnjbJTdzCgRu/MZFyH/8/94PvqVCQZst/qlJZht+p0Hptwyu
BV1+nOyeevovflSGGFqrffkehJz0zBlvrTfC1P/PIMpBaWCmnRLwXm0mqtvKzX6r
jM/mSgFjaK9AJGeOnLBHtYE2+JA+ajEM7MTT6uyT5ZAYn0DSEf5RFzgEdWu/TN1p
OdTqm9N/rZwtvrWay3CG7BAdvQsZ33tXPk1LaXiQMqNaYMLfaCdWn3vhK6zIewtO
qx2iYy7UBsOSBoMjIjPCzmhdkmiNG/hmvsFmyK6fyaLmgh9eQOJUCNeL8WPi2Obo
7bAsX8tf0Gca8aWakIYpVjTEE7IG9F8tkLapqBUtPl5WnPtsa6yfnG2YhLNXVyBz
d9ggXhHmxoDfWdVoFk2wI5hfb35jyFhONoi7mnGcHHKlGqxsmT+p3WRfGgLUWmW1
DC4sk2RM9cxU1fs2omfQBD0tSELz1Ng4B0vnYlyma0SqfjbMXp6BbF0xlaCvUS0S
kQMc0ryPQU8SEn15ztsyntuSVvdYyMSV9c2JKSD976J5KHtQ6clA4TWiXO0/Q+/c
uCaZEtftNp6fYCq2oowjt5jMLyYlZsVphW4gys82Naseey1SlTK7do38yWZyUKJy
3S8FjrV0mOE7EM7D8PNokPTYEU9Weemh6SwLexgCiYCYgkIPwlVcCYxiKzTCnkKt
3nXCm3DQDgi54KlafW2z7LX8b3l09k7QzHD40Z2JdG1d+4YnKJndRNHkHJgV/F4x
1Mg0y8CJFXTjQkuYiLwoMYMkDWeE5dxdIAQM+vLiQF2Vs8ZvHFq6QlABYUHBKqhR
lDAKY0oepjLqeXUIQkGMt31lyQW3RHqWpy4lQHO/zJ99I2uJRArYhHMtO24CbZDx
c67/PqXsJ6o8Oie6J3/3czuz6UGgrwhq/iKIg4an5i3gkevRo09t8vUAv2MWyh4i
XQqrrss0iKelIG1WWKvwTVS9JqCfNGyLX4tEWJX0UROcv6rpf+i6ANA4Zi0Eryo/
8MJT1qCXtQUxEhmJW3QrwG7dXV97/B3zstn8Nw5QQpf9s/JAlOQ1mIqiKDFoTFUe
0qeB2p9HSr1DQLf33NbS3LLYL+uZPhUF0VKSZlhge/5xKcpt5Vba6MxBshqhKZ1z
Yj1ryp0B7vBLk/cytZMG9SBEO9xTyH5pFl1MNj/7h5tLaUkUKExYTrL3rTP10hAV
ZGzt6a1LKU5dE6EG0wRLd4c6cCi226qiFJ5zgpO/p6U8Fm5vfHJRWlW3bTIbqgFo
tXn2MboeIhCsjILXoF+m7GdOBXIk6yeT1DjpwMdOMDpFNBZ+XIlfiiNOECHGQWCZ
C+y2OAH+82lXlicq6FNZBzERbN/xteM5N9gfYYs5gUirMSvCKmO1GVQEZAAwj6Iy
8Wezgj+TmtYYqhCNOtN7VE/tsK1Pl3fOLGV+WRpjZN7kXRHWSqgYET1tJ82TFqnq
zWMRKOsqrjJoVGY5KDzGrt+K2iIwIeKYDP4Jfb+8kixlBT0DBIEOBWKFJ0qhAQHl
77GkxlZQ2JqKOxdxe01QNXD9tFEZK3Xsw89r13LzlQHp9s5Jtf3SiEwSsDwhSwLi
Iweu/l3vXWpQZLPk6H7U9QCj0Dw4/enJFQ4Oo4CpEDb4tuT3qqdmOPgFdG6ne8gn
7z2Gwzo1uTHLhjhOZV5787cyGdU5Cf+PO7MEhU4BYXu8RN7pOdtYy4uSsdWi3VA6
7BB3GvRQuJIlUKRnMXwoPZ02gHu6NlBI3nIc2SvMqAdphSfiMjJ4tmDH1FO+LeOC
npAS3xcuN2ExB6w91rpOGXu1lIQbaeyZUvMI4BMGi5XwBlWFIYDTPPAnpRRiYrER
s893vFkmgLTIVXM/uNZhUQZVm/Nc1qLuJyrnS2ecDmTv826TO4lV3wpv9ml34Uxk
FCihPK9hvfv5LDopxuaDd/oASYeQQ82pJ1ANWSQOMxYeIxyvwsxaSL9OkCnri5Jp
6NxwW8o8k/vjm3flBg5ER7rjr/doXpqLdMLLpbD0ouhUX1PtSauvi9cw5CiqDpba
CnMLt1BciYqSfBMSpYkLzkRfYSIPkDzSRy1GmrFEdiVp4SA+zIQ2R2bxHpRRTYxN
6r1v0F9m6pI5WQbbpJcWuLs79/3uvsb4rdjw8BOcpUR5OF2NbwX2UqKXROQq396W
K0IRVP7RIEstdVPSKqsdGSYVhganuWEUanZSmdsMUG4IvCRyeLEb1iWmCGC7mayU
LNAA5aRjdQCDEVrSJvoLzDUX2f+a2W4XmRssHNLkkygGf/z9MNb57L3xGF6/Pn+w
sdlj26xDmNun40o5UBoo6Xnbtd64d0JomWAmeZZiBQHVQMf9AtQWHRIgNw6QR0hp
oTrul6y/NFDGKhQH/LuwIgGnWeI1zITLknqDuW1GI7mi6W1wJvjgWyNcm3DSjjPw
+8384NGDWzyyYC5mRRXZg+lzIfrnwq1zOtnuEhzW+JTmZXNZBktVi+rxmrOMsAAM
EBc/Wys7wG/1JfIkLLJBeT0+Lo1wWc0biaOH+0u4OvZ74Nbry9VcHfEJczeCfkb0
d5VgzeHVOQLs/6CQ72yDstEELwYuP6YRlMv7FHIk5d7/EZLhAWK+0HCLUnVoe/13
`pragma protect end_protected

-- megafunction wizard: %Deterministic Latency PHY v16.0%
-- GENERATION: XML
-- arria5_phy16.vhd

-- Generated using ACDS version 16.0 218

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity arria5_phy16 is
	port (
		phy_mgmt_clk                : in  std_logic                      := '0';             --                phy_mgmt_clk.clk
		phy_mgmt_clk_reset          : in  std_logic                      := '0';             --          phy_mgmt_clk_reset.reset
		phy_mgmt_address            : in  std_logic_vector(8 downto 0)   := (others => '0'); --                    phy_mgmt.address
		phy_mgmt_read               : in  std_logic                      := '0';             --                            .read
		phy_mgmt_readdata           : out std_logic_vector(31 downto 0);                     --                            .readdata
		phy_mgmt_waitrequest        : out std_logic;                                         --                            .waitrequest
		phy_mgmt_write              : in  std_logic                      := '0';             --                            .write
		phy_mgmt_writedata          : in  std_logic_vector(31 downto 0)  := (others => '0'); --                            .writedata
		tx_ready                    : out std_logic;                                         --                    tx_ready.export
		rx_ready                    : out std_logic;                                         --                    rx_ready.export
		pll_ref_clk                 : in  std_logic_vector(0 downto 0)   := (others => '0'); --                 pll_ref_clk.clk
		tx_serial_data              : out std_logic_vector(0 downto 0);                      --              tx_serial_data.export
		tx_bitslipboundaryselect    : in  std_logic_vector(4 downto 0)   := (others => '0'); --    tx_bitslipboundaryselect.export
		pll_locked                  : out std_logic_vector(0 downto 0);                      --                  pll_locked.export
		rx_serial_data              : in  std_logic_vector(0 downto 0)   := (others => '0'); --              rx_serial_data.export
		rx_runningdisp              : out std_logic_vector(1 downto 0);                      --              rx_runningdisp.export
		rx_disperr                  : out std_logic_vector(1 downto 0);                      --                  rx_disperr.export
		rx_errdetect                : out std_logic_vector(1 downto 0);                      --                rx_errdetect.export
		rx_bitslipboundaryselectout : out std_logic_vector(4 downto 0);                      -- rx_bitslipboundaryselectout.export
		tx_clkout                   : out std_logic_vector(0 downto 0);                      --                   tx_clkout.export
		rx_clkout                   : out std_logic_vector(0 downto 0);                      --                   rx_clkout.export
		tx_parallel_data            : in  std_logic_vector(15 downto 0)  := (others => '0'); --            tx_parallel_data.export
		tx_datak                    : in  std_logic_vector(1 downto 0)   := (others => '0'); --                    tx_datak.export
		rx_parallel_data            : out std_logic_vector(15 downto 0);                     --            rx_parallel_data.export
		rx_datak                    : out std_logic_vector(1 downto 0);                      --                    rx_datak.export
		reconfig_from_xcvr          : out std_logic_vector(91 downto 0);                     --          reconfig_from_xcvr.reconfig_from_xcvr
		reconfig_to_xcvr            : in  std_logic_vector(139 downto 0) := (others => '0')  --            reconfig_to_xcvr.reconfig_to_xcvr
	);
end entity arria5_phy16;

architecture rtl of arria5_phy16 is
	component altera_xcvr_det_latency is
		generic (
			device_family                 : string  := "";
			operation_mode                : string  := "Duplex";
			lanes                         : integer := 1;
			ser_base_factor               : integer := 8;
			ser_words                     : integer := 1;
			pcs_pma_width                 : integer := 8;
			data_rate                     : string  := "614.4 Mbps";
			base_data_rate                : string  := "1228.8 Mbps";
			en_cdrref_support             : integer := 0;
			pll_feedback_path             : string  := "no_compensation";
			word_aligner_mode             : string  := "deterministic_latency";
			tx_bitslip_enable             : string  := "false";
			run_length_violation_checking : integer := 40;
			pll_refclk_cnt                : integer := 1;
			pll_refclk_freq               : string  := "62.5 MHz";
			pll_refclk_select             : string  := "0";
			cdr_refclk_select             : integer := 0;
			plls                          : integer := 1;
			pll_type                      : string  := "AUTO";
			pll_select                    : integer := 0;
			pll_reconfig                  : integer := 0;
			mgmt_clk_in_mhz               : integer := 250;
			embedded_reset                : integer := 1;
			channel_interface             : integer := 0
		);
		port (
			phy_mgmt_clk                : in  std_logic                      := 'X';             -- clk
			phy_mgmt_clk_reset          : in  std_logic                      := 'X';             -- reset
			phy_mgmt_address            : in  std_logic_vector(8 downto 0)   := (others => 'X'); -- address
			phy_mgmt_read               : in  std_logic                      := 'X';             -- read
			phy_mgmt_readdata           : out std_logic_vector(31 downto 0);                     -- readdata
			phy_mgmt_waitrequest        : out std_logic;                                         -- waitrequest
			phy_mgmt_write              : in  std_logic                      := 'X';             -- write
			phy_mgmt_writedata          : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			tx_ready                    : out std_logic;                                         -- export
			rx_ready                    : out std_logic;                                         -- export
			pll_ref_clk                 : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- clk
			tx_serial_data              : out std_logic_vector(0 downto 0);                      -- export
			tx_bitslipboundaryselect    : in  std_logic_vector(4 downto 0)   := (others => 'X'); -- export
			pll_locked                  : out std_logic_vector(0 downto 0);                      -- export
			rx_serial_data              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			rx_runningdisp              : out std_logic_vector(1 downto 0);                      -- export
			rx_disperr                  : out std_logic_vector(1 downto 0);                      -- export
			rx_errdetect                : out std_logic_vector(1 downto 0);                      -- export
			rx_bitslipboundaryselectout : out std_logic_vector(4 downto 0);                      -- export
			tx_clkout                   : out std_logic_vector(0 downto 0);                      -- export
			rx_clkout                   : out std_logic_vector(0 downto 0);                      -- export
			tx_parallel_data            : in  std_logic_vector(15 downto 0)  := (others => 'X'); -- export
			tx_datak                    : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- export
			rx_parallel_data            : out std_logic_vector(15 downto 0);                     -- export
			rx_datak                    : out std_logic_vector(1 downto 0);                      -- export
			reconfig_from_xcvr          : out std_logic_vector(91 downto 0);                     -- reconfig_from_xcvr
			reconfig_to_xcvr            : in  std_logic_vector(139 downto 0) := (others => 'X'); -- reconfig_to_xcvr
			rx_is_lockedtoref           : out std_logic_vector(0 downto 0);                      -- export
			rx_is_lockedtodata          : out std_logic_vector(0 downto 0);                      -- export
			rx_signaldetect             : out std_logic_vector(0 downto 0);                      -- export
			rx_patterndetect            : out std_logic_vector(1 downto 0);                      -- export
			rx_syncstatus               : out std_logic_vector(1 downto 0);                      -- export
			rx_rlv                      : out std_logic_vector(0 downto 0);                      -- export
			cdr_ref_clk                 : in  std_logic                      := 'X';             -- clk
			pll_powerdown               : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			tx_digitalreset             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			tx_analogreset              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			tx_cal_busy                 : out std_logic_vector(0 downto 0);                      -- export
			rx_digitalreset             : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			rx_analogreset              : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- export
			rx_cal_busy                 : out std_logic_vector(0 downto 0)                       -- export
		);
	end component altera_xcvr_det_latency;

begin

	arria5_phy16_inst : component altera_xcvr_det_latency
		generic map (
			device_family                 => "Arria V",
			operation_mode                => "Duplex",
			lanes                         => 1,
			ser_base_factor               => 8,
			ser_words                     => 2,
			pcs_pma_width                 => 10,
			data_rate                     => "1.25 Gbps",
			base_data_rate                => "1250 Mbps",
			en_cdrref_support             => 0,
			pll_feedback_path             => "tx_clkout",
			word_aligner_mode             => "manual",
			tx_bitslip_enable             => "true",
			run_length_violation_checking => 40,
			pll_refclk_cnt                => 1,
			pll_refclk_freq               => "62.5 MHz",
			pll_refclk_select             => "0",
			cdr_refclk_select             => 0,
			plls                          => 1,
			pll_type                      => "CMU",
			pll_select                    => 0,
			pll_reconfig                  => 0,
			mgmt_clk_in_mhz               => 250,
			embedded_reset                => 1,
			channel_interface             => 0
		)
		port map (
			phy_mgmt_clk                => phy_mgmt_clk,                --                phy_mgmt_clk.clk
			phy_mgmt_clk_reset          => phy_mgmt_clk_reset,          --          phy_mgmt_clk_reset.reset
			phy_mgmt_address            => phy_mgmt_address,            --                    phy_mgmt.address
			phy_mgmt_read               => phy_mgmt_read,               --                            .read
			phy_mgmt_readdata           => phy_mgmt_readdata,           --                            .readdata
			phy_mgmt_waitrequest        => phy_mgmt_waitrequest,        --                            .waitrequest
			phy_mgmt_write              => phy_mgmt_write,              --                            .write
			phy_mgmt_writedata          => phy_mgmt_writedata,          --                            .writedata
			tx_ready                    => tx_ready,                    --                    tx_ready.export
			rx_ready                    => rx_ready,                    --                    rx_ready.export
			pll_ref_clk                 => pll_ref_clk,                 --                 pll_ref_clk.clk
			tx_serial_data              => tx_serial_data,              --              tx_serial_data.export
			tx_bitslipboundaryselect    => tx_bitslipboundaryselect,    --    tx_bitslipboundaryselect.export
			pll_locked                  => pll_locked,                  --                  pll_locked.export
			rx_serial_data              => rx_serial_data,              --              rx_serial_data.export
			rx_runningdisp              => rx_runningdisp,              --              rx_runningdisp.export
			rx_disperr                  => rx_disperr,                  --                  rx_disperr.export
			rx_errdetect                => rx_errdetect,                --                rx_errdetect.export
			rx_bitslipboundaryselectout => rx_bitslipboundaryselectout, -- rx_bitslipboundaryselectout.export
			tx_clkout                   => tx_clkout,                   --                   tx_clkout.export
			rx_clkout                   => rx_clkout,                   --                   rx_clkout.export
			tx_parallel_data            => tx_parallel_data,            --            tx_parallel_data.export
			tx_datak                    => tx_datak,                    --                    tx_datak.export
			rx_parallel_data            => rx_parallel_data,            --            rx_parallel_data.export
			rx_datak                    => rx_datak,                    --                    rx_datak.export
			reconfig_from_xcvr          => reconfig_from_xcvr,          --          reconfig_from_xcvr.reconfig_from_xcvr
			reconfig_to_xcvr            => reconfig_to_xcvr,            --            reconfig_to_xcvr.reconfig_to_xcvr
			rx_is_lockedtoref           => open,                        --                 (terminated)
			rx_is_lockedtodata          => open,                        --                 (terminated)
			rx_signaldetect             => open,                        --                 (terminated)
			rx_patterndetect            => open,                        --                 (terminated)
			rx_syncstatus               => open,                        --                 (terminated)
			rx_rlv                      => open,                        --                 (terminated)
			cdr_ref_clk                 => '0',                         --                 (terminated)
			pll_powerdown               => "0",                         --                 (terminated)
			tx_digitalreset             => "0",                         --                 (terminated)
			tx_analogreset              => "0",                         --                 (terminated)
			tx_cal_busy                 => open,                        --                 (terminated)
			rx_digitalreset             => "0",                         --                 (terminated)
			rx_analogreset              => "0",                         --                 (terminated)
			rx_cal_busy                 => open                         --                 (terminated)
		);

end architecture rtl; -- of arria5_phy16
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2016 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_xcvr_det_latency" version="16.0" >
-- Retrieval info: 	<generic name="device_family" value="Arria V" />
-- Retrieval info: 	<generic name="operation_mode" value="Duplex" />
-- Retrieval info: 	<generic name="lanes" value="1" />
-- Retrieval info: 	<generic name="gui_deser_factor" value="16" />
-- Retrieval info: 	<generic name="gui_pcs_pma_width" value="PARAM_DEFAULT" />
-- Retrieval info: 	<generic name="gui_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="data_rate" value="1.25 Gbps" />
-- Retrieval info: 	<generic name="gui_base_data_rate" value="1228.8 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_refclk_freq" value="62.5 MHz" />
-- Retrieval info: 	<generic name="en_cdrref_support" value="0" />
-- Retrieval info: 	<generic name="gui_pll_feedback_path" value="true" />
-- Retrieval info: 	<generic name="use_double_data_mode" value="DEPRECATED" />
-- Retrieval info: 	<generic name="word_aligner_mode" value="manual" />
-- Retrieval info: 	<generic name="gui_tx_bitslip_enable" value="true" />
-- Retrieval info: 	<generic name="gui_enable_run_length" value="false" />
-- Retrieval info: 	<generic name="run_length_violation_checking" value="40" />
-- Retrieval info: 	<generic name="gui_use_wa_status" value="false" />
-- Retrieval info: 	<generic name="gui_use_8b10b_status" value="true" />
-- Retrieval info: 	<generic name="gui_use_status" value="false" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_enable_pll_reconfig" value="false" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll_count" value="1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_refclk_count" value="1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_main_pll_index" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_cdr_pll_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_data_rate" value="0 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_freq" value="0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll0_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_data_rate" value="0 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_freq" value="0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll1_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_data_rate" value="0 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_freq" value="0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll2_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_data_rate" value="0 Mbps" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_freq" value="0 MHz" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_refclk_sel" value="0" />
-- Retrieval info: 	<generic name="gui_pll_reconfig_pll3_clk_network" value="x1" />
-- Retrieval info: 	<generic name="gui_mgmt_clk_in_hz" value="250000000" />
-- Retrieval info: 	<generic name="gui_split_interfaces" value="0" />
-- Retrieval info: 	<generic name="gui_embedded_reset" value="1" />
-- Retrieval info: 	<generic name="channel_interface" value="0" />
-- Retrieval info: </instance>
-- IPFS_FILES : arria5_phy16.vho
-- RELATED_FILES: arria5_phy16.vhd, altera_xcvr_functions.sv, altera_xcvr_det_latency.sv, av_xcvr_custom_nr.sv, av_xcvr_custom_native.sv, alt_xcvr_resync.sv, alt_xcvr_csr_common_h.sv, alt_xcvr_csr_common.sv, alt_xcvr_csr_pcs8g_h.sv, alt_xcvr_csr_pcs8g.sv, alt_xcvr_csr_selector.sv, alt_xcvr_mgmt2dec.sv, altera_wait_generate.v, sv_reconfig_bundle_to_xcvr.sv, sv_reconfig_bundle_to_ip.sv, sv_reconfig_bundle_merger.sv, av_xcvr_h.sv, av_xcvr_avmm_csr.sv, av_tx_pma_ch.sv, av_tx_pma.sv, av_rx_pma.sv, av_pma.sv, av_pcs_ch.sv, av_pcs.sv, av_xcvr_avmm.sv, av_xcvr_native.sv, av_xcvr_plls.sv, av_xcvr_data_adapter.sv, av_reconfig_bundle_to_basic.sv, av_reconfig_bundle_to_xcvr.sv, av_hssi_8g_rx_pcs_rbc.sv, av_hssi_8g_tx_pcs_rbc.sv, av_hssi_common_pcs_pma_interface_rbc.sv, av_hssi_common_pld_pcs_interface_rbc.sv, av_hssi_pipe_gen1_2_rbc.sv, av_hssi_rx_pcs_pma_interface_rbc.sv, av_hssi_rx_pld_pcs_interface_rbc.sv, av_hssi_tx_pcs_pma_interface_rbc.sv, av_hssi_tx_pld_pcs_interface_rbc.sv, altera_xcvr_reset_control.sv, alt_xcvr_reset_counter.sv, alt_xcvr_arbiter.sv, alt_xcvr_m2s.sv

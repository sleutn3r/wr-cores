// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UubtP/uNkjqpwrcyWEz+C8zTX2NedZE/erBX4A6AL/1wos3Hv3Z6lmqIjy1WLZvE
80XCacGtQTseCupaG96RzbJP/TcKJPGfMit6EZW94TdW6FccFhn1aH1gZxBuS9Vx
NIlTctiAVOYyZW2ZDHAMVkODoNuBu/3HIJaFC8Yi+vw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27680)
Kw90xhaKBOzZzOnaSOji1nmSC+zZHSylW71BdgV89TAChsyV5UD56LhoNo9o9CiL
aT4NHlV1kEzVtW9+uSoprttdEl8pQqAVhjQdVsx31WvGao+3w4iWtPy6b+ScYHUi
BdheKxEmCafsdP4XcuWkBakHClaw5rNDaNP69aexeHp+PQD5fpEPGasPyRJzpuEk
a3s4DunMxZSc41LELHxv9m5awDPjx+9kHe1Od5Wq1yug8ouaMfMclsOO4lvRYR9q
yfNQRWLoeRslb8K21ycj5LQ+EnhTDkZJRWF77OIuk0pyoUBKenPMc2L1CxRzbQ5v
i8eUbL1HRyHPYdgqZ6ha2d/1ufxBDoq5z2g1iw0pM+NpAuPwe8ML1a3mdshx+feF
X62sxURx9DGh/iKhlWFKyfnKgxyO4Q+Ijv/VBhV6qkg3bAEhteK6Et333P1AA1Eg
1TCdxaFOUslBQ792xNSjEmxzOuRe3IGT3tg+oNmtKx9cgtflHl+fZRHnVdgp8LwL
GGkpBVZZaQwf3J/dINsw+FDhy4Fcb9pDHcvHE67lWHZ3iBfJNF8KHi+OjlZE+WZO
WsXs30tUfTQi2P4SKQP1k/L6p8I3vqE/yUp2wYbtlKqXhgHUL7NJEQrHBzDH/RB1
lfNvweVT1euRejFrbgks7nbBlJnX7KdCTFWgML7MHUD8UFRA8is6jJOjSvK0VnLr
eYaDs70tsnXA2puZ8thEbOinFWaoQfx1/qh8V6t2ndDeiEIYEtPlosxnu1UeDrfy
MspkR506nVCf2Zmj9cfa1p2aV3TNGJ6i1sBoEutOp2iGyrSpwQ9+1TqaKQir3CLy
cpaHSCtg54LFGEYmHF6oGPyhChyZEY+OruO9493LLrIPowmqGL2xILLioD6bL3aL
FFByB7fMmmH4Mn1/tPPxFwAlbBvBFB+HnQC00FIc9B0kzFQTjfL4GQH0D1PDAb9S
GtszpTeynHfScQmhDo3tNgQrUNkSsuHHVtYoWO4DZxjLHu4lJ4HGn/72yS0TW/yr
PVn6cT+La5fbcjJHIDI88r9MyYfH3qYjcKUmeyyngQKsKDO9DpslS6eVNmqVaMsk
ZSO8vIn3OPRNwE+nQMNdWDtpJ/753R3fpAErcv6PPMHmtmAZjJkLNwUQDUU9cE/I
LRfL/XmmHJQ6TB0yl8u0XJWD5zR4HfkaY/Wlad0x8XcWUrBx8JvrghFyh/JDlnSB
FQ0NgRNoyzZ51tqJvFbWhqPtnGDbBtP6Q31yKcXtWfMufHHZ0gU0whfyWZjKgPgo
EGaVEp1LJA4e0wb/ZoeBHxILmN/pEFTX8mjyZe+VhuhLNxh4n8vtyIysX+VoPfDV
jF2Ir7BSFAVRu1CBIpVhnfNa3nugDvQ/gDusbRW1u5sK5fRHwMR2lLcZBZvDlAHB
zo95F7XisgEjm+ifVYxE2Zxi/cWJSmG+lU3oOCrikG+Okdd+vjTbMs8T/nVYL+iC
mnb9A/agD2xA3q0Ky1jtpdiFATyV+jif8nGmYH8HlyrN4zGsLbgeKRCtD2XvyNpo
/R5C/OF6UkxCe+OSsin2Wdqlw5of2rf+oBzeA2wDoUYeqp+QR1VNPWXumS+xzT9+
SdjxJxSHOsQUxxtWpYal9cDTn0MnUkNPq6h/j8PZFSvBSyGw0JLpFg6xKYSnAZfH
YiS73aqCAvua9uufvgkVv6pAYXs+tudqMR9HqZG75jvhwKpZw9nLm1j5pWr9wAaA
soI36J95DIEDJ8E7YybehG0nEIsVCh8LyXMCf2fslC2ymOFQ2KnnI4JY24wZZo6L
Ni1JgYHm/K+vgkGKyW3xWqHfTxhw8bOhuBPrdpp/cjQ5rh4IR95AF/h1aVBde4BK
qdR3UjHqx63WqcPiwI4nYBo2bKite6Fo/EMm1WCYDeoYH+OiX9GQyzPGsnmNtd3b
J6+D2m9+E5sg/7axBN7Gt4EgwNueEY0QSx08/ForRL+85HLJ7Rnvb6lCP4mzKOgm
rJSuVb6pOTj0u9IJ7/oCqmvmG+Igs2vDXIBJkqWNIFU7eVvOTLlpuRxbpDP+xzdU
TLWT7vArLQjCwSQKei0REiAwCVb3BYrBfWg8vFzT8+3ZmiN5i/gxExyjtYsW/lDS
V0q6wnZuwrlGH4WyPjH5b5y9iifW0fC5jCFylPf5UeZXNYSaI7Dgn7th/it4fsVK
27a4vQZ6iqBpG9ShYs0H/g5K/hozevGMXOIVK/McGvd8FoNO7MbjXqOehXsmAKX0
dL9xX8GbturlYNP4X4xuacgovkVCLMqzouwAJJIVhzA+hmCcmJ7UokJrh1WEomNY
BClFw9N875JCZ5lS/WBwAP8Yu7DgTB3MSsJz3ynepc+t8pSrtCllxvrmqpBxlP3P
LcyRqROMaNF/GZrsvoX/fo0u+w2WvbTPOD6pizfW/dQzVqPyoqL3XaDaFweYiCdF
y/MStk3TYOeK2pyQgpQGUPzh/tC19rCxAcarjvH+1H/SGsB6Dn/qwyzZ9iLxQlzf
fz5DfWrlA2gDFFatb3hqbKePVT7iXT+mrdcRl6aoDYLyd838UONd6x0SHmjfeSsg
BD6OVAMUwAVLekbsJKjh9mHFh71a/49goepe55ruPKJ+s9ewLnzcLPOWQ3FQwjLL
gavSd/Z0JiuDTdind4XFxaf+RNA3E2qRBT5MLHCBxiy/A2h/Sf3PCocd9A8Ae7xG
xZnB07fMtrkxIMQy4KszkVmvRFGK+QWaOHP8JBcx6kb7ZQ63TvWxizm4NUTV4Goy
Xfd7pH71EP1sFaKIi77iLTFFLNxnn08u23izzKCpw5xmFDg0IcvYTC5SAFDbGFUq
V7wRn6pVhagqY4Kr2GK8RbOVKW9/xlgdp7loL7iwpoZrw0QAdrqhxWuPEcVTNQkz
1MzjakvD/rrrzxEBabIHD/2wsVSouQwoJq/NLo1VMm15uyVJLZJ7AWWdjOjvabcc
Npk0MuinM/U4rfQjXuLARv9KGtFF4+IL9rysjL4ZAXHbzhQAoIfYNKoFcx1l4Dpz
bOCrm97ELOdfiGVWoHI+9ETQXoIGk70jV7ZrTIHDebBh10y/sZxyNcb24MWgQbRj
uZP8gTswvpSZHaCOFsw86h+l28OA8L0iR+SkmjxBuzvbu2M9ABwVAJCjZJIBu8KW
Zh5l8nCekbtXAAhDidt+pcCCYadxRlKkbXiONyhO2utmAbLoN4mwqEiT7BUAOhlT
MvYNzblKU+L0LejNaxCLgIlwiEE3xE2Xr7WGEZfpZ8ynqJmSzU6IqETIlLqQ0f4w
YzQHWZ7Lg7wUQYrLeBl++w9tJOqjWKBVH9A6ZcDuNFBj1bxPQpkDIpN3b/pGwE3m
XZYwfI2VHSLbrNso2+cKf3lzB2vKmY4BlhwF9rLn1ScVyVRLlbnbWeYJJeHjXWcj
6A/xUSBcJxiG2uJJpT492OmV2jUgr6qdjzI8EBiuSEEnjTZGF3aJZ50N43mjLIIt
Xaxzj78HUTqU3auPTHGWrlKa1QxvRdHAH2tBplWQlInjpyc5UkAtCCuB0O0azJvd
ksM+Det2Gc4DMvzsvh5fKUWf3ujgI5hbMsJFX1bLfsct3ZxqeeD9V4QHSXoU7GZ7
e69+dyT0maNIvuRezhDA1UW8dJ+hyPH5npAxzeSABJzZERiDhrR5WyQDIHFChL1y
K2xPNRgWS9fHLJknHx4iw7CvOVQSjgmPswlE0VISiRwrbRpiopQqQkuTOkmpK6/X
+Dc7Nqhcz1Z6ZEUFAORE61IqIBQWGOhBQsgmBVpfZCKc66CRTguiOhWEMdaSfBsU
7GnrE+5tXHeOV7O09goKMP9llSOciru6YZom5jQ6uXr+XLc3eyHBKu3gNmY+D1Sk
AxGjBHbOKEWE4TWBzM/ywnTZ/Gx/i6h+BEcqBaHRwbTOioWa/Ofxx+CKe7o178j/
vcoAen66MauoKsnuiephP3zlfFWV1fo/xcfeZt4ndV+PkUqRBZwuisIXXwL074rc
LT/6rkR37j+aHAs2IJXk/vXqbSg6nU/3nDOH1nRyTE8K3ia7I0eJPqnglEnSkpIq
V0YI/g61Sa2wE4SOy62gRdnw5vhlSRDcKVvEpvlVtx7OyuDi9m/qd9CRmTOHg1BW
fg42WlNxOtykmJOxfRaHIhKA/rIibW35WmhaqHq53xeUsCQt+tycilYituVZ7vAu
BfGd49KfpcSAEXbu7Ajkg39UYz7u2wkdyJovItA7BjE1ZtaDo/jCgSSbGpsXxTYJ
TxgC9y4sf+S5pDEUHBfQdRK0eKQkwtNDBmZgQgD5eUBQ7R+UDIdmCb+RDj8onDDz
rbc7tOQM34GnDyVqgDdJRKDRfhFWjch0O0z1ejEwCf+swWo+7xZNURvyFur2T4VO
njQa9D9aPDJnr4yrt03kx6JU8yFhv/kPIw314zAMI1NNEmFBF8NS1LbVjgqfx5/I
RY6NXylGHJ4tHOkuWxoIXmMrdtEWtR+STSNOUINYWpb8IAwpXoSI0CxRgiUnO9Nv
TclW/ajRhNTZtptpt5Bw8bBuVXVYVe3qEC8Mjqu37hBWmoNKC83qBotx37001agh
+rwT3RBa0vz6vxsH37/CyzF43i/WgvdYNa0gG4r3wJCHYCF6kQ6l+cHQnR6hBKIM
R/RtThH/s/IP5raALU/wWDwRFW2HrdHs/qcOMEPKOMovsW6TSA/ZlPuCWU2Dvewj
uxdDw9uDHp8L24Z5N/d0yMAZWxWmfxtdpr9nJIeUHLJKnmqjNwYmEWatX4TTEjFX
bxr9vVBe2ZXErsWsE4obLKOBT80Fbaky6x65shShL9kOBI/gXrNdqRLTadZead9C
WzvLS++7fpk8N8xNI94OWRg+2VjJZwjv++mNyVhkyJr0MDiv7YbjcrWanmxwCvWa
kNjLvTaI5ljZVdEpBw+vOJz9GZIzt7tJCMeoZHPLxsImeHqwYkHZHVfo2Gf8H9c7
ZXjmacmIihZKpcuWtAKIuPanAU8BawuKvsez+NvlRbdfTNfnYpFTLZhuFB2/SZVV
IQ6F5WG1wgpMxwiK7iUNvBpgrgWwdHlaqfAScLTofhyUAlPYDs+p82cza1q+nxAj
JYG6fAXKYHmGTugVpqv6THl4B9fRyeWyMj5Bruo4k/qU8sLEQCVZUqkPyKTY1V5z
raqnn06yycqYoOXFOlbWHcxl2xPE1v5eLmv0RSwuUu9DCyqrn3kwccDZ1lGsJXoE
s15FyDG6iY5KufzqYnX/x74/xoolG5PaoyIUdFpy0KjH6I9i1eRN+6/+GKtGGOb1
q0OhIHp/AzUl9GiP075bFL7XwrMch6oSpIqdmvJWdzBc5BV1qNeb5iic4oUH9zgl
vh88t7fvGWHY4Uhm3wCpNTlzcyZS0Gm+6ctW+Tj/RyMfNy1fSi41lQbgp3xxL9i5
6RCRYmZohfoL2LhR9NRMYof1QwbgJcr5pNxUbPJuyN0kA5aNmFWvf9QPZSeVsVG9
OnWPTylUA4Sg6Lk9fg2JqX9p/xpu3qRWusPi0c1M/yD44k08D1LSX7QYT5iAOzmz
5bbOZp01rnmGPGTNTrXqNnLmxYU/TDrPvEWJCZZ569kw/Emdle1weTyF+hx3KOgQ
RLuccPkEqj0Wwf2M5ZgVQHWiCPXLMtIJez4TcSTscIr7pwCglXhuPUhXp+5Ynx+l
EKxDq/HeXVnl0vIhbhVu09rKoWtkLalkWurMmi0O0JLt7QePYgcMb38WzLgL6rsB
l0ut1hmI8FZB5idvd/o9ixXUaTGU3lmV/veS2+FlKYVgZMnpYTHnDUcc82IF1odb
IkIl+bs2xDstfz2mESO60ef2zzPOHZCkMatmd2IQaKNzrm0JMVw17buFkO1RjX1d
GjcnaeG5kOZltWC6T1z87bReLp1fF9L3J7yLa4iCtzTjZ5jYEYoef78eDtHLzNzq
hvwwngmsHBwxWGjVsJK80+6+PZoLegrgogs0tWrgnFjMZ+gEcv2gZVL7A6jAcAx/
/S5++5dV8lme1fXzUvUiLVSIxyCk+lD0w+I37sDpMXrFGUH4HBAVpu2p/3QDotxu
0wE8a99ld9uXuKu0W9LAAzo77XKoiezJkQRcq7IilWvsCsip+IqyyNIAEgu1BqEU
O1SuLzt8nEBcX0FC6qkHhN7tMh3FVLQlc20CumR45HjWMEVlRGk4trVycvYDxDYw
ieb497gORVfEl7zNVIs5KCR9y113xRozGJ5fYMad2kzmhI1aByV62vjMf5u0il9C
UvG/0ExxnGN4qYyAI5LiMOhLEAbmoKUrIVopTg64sh3M/Rvn1Xb6A5b2wzMMQciB
yUdAPmK80UOqNRR+rXCqwl8jba4Ff0sXIbqZsnEAwpIDxfTKzmDw3gq5yIegLEQW
iftbK46Xpu3+AmzuNR8ClXEad1NPwBWf+XD5NHl6co33kgkl8V3SzFRxerXykjyS
3udWO9LrlgWVbg/tN+2k2nJjG5ODp/X+YKfNmk/Uqxl+rhxEETAT4CTUdWdKn5Ef
Hj5/AojtWCdPDzpCyuPbVhFDammt9BKdKWclqBbM7dZ3ahZ5o8I9VDUIw8hhUtOC
Lhi7XEFtS1hW1SOqqX3vUKeq+AXwL2Ihl0Xu6lgyg0UizHqZ9W/21ue9c8/g6EFK
skRm20HlKfUc8wtVinTbRfmqH/gDxPQVJ98ymttpubRetPGWyAoO9voMnSz49B5s
YkmreQAVMWKiZq54g8CjgK8DwMi+SZQNbNf+cdp4pExX4LZPt1s1oDHT6aEMqSIQ
e0ZSaWyhE5Bvd07MzVrFmdNEuh2KEtx0jd/JoLYA+vJX/ZfCtBUv/jqUOaEq8LQp
NX3yeKnz3ltZnxatJw//+7NzqSehlIsAa6JguokvLKkdhat6kh5dVrBqcJ9U7CHl
Ns/twM8jX3Lte9qhOLL0DGTObJBISsLru22YgQm0fIVTxRJ97s6PNEpqn5Sz/wCh
aMC+InAv+t39vEWRqZ6gWqpVd/vuzyExT//hw22V/8X7ut3mVptR66kVC4E1Y7RS
PRBu3PpRyOa87rRu6ifw5lah3yKNbQYmAPfU4+mQvNbHZrRxb/p9EiOXmJkawJkb
7hLyrXdEYOLZEDUVVILe9430f8a/XahXaL5YRZhxlPW4fvQ+JnUfg+SERNats7ex
8niPQkvoUj3r3O+NCaym6Zr2mlGzjqbj52cHLUIskzZpJoQH0yyOm3CaHjjf9pSb
YL6HuweNp2wjfuoeMUrW6dzM2das0gxUQMo7jfn+C5UjJgDBoVgdMEArH1OHglH3
mROxS+B75gmXoboYPKjoxk/1LRk4KuunSZV6seRGtppl9d0wl7VP58UWqk04yHiD
AADbgNqo0ex6ivMBzEadZxdr46KV/nn2lQVZ2weAIR/yE+I9IVCLXxU/y3yRmZHr
Dt0N8gEI+ZRNc9pMdcbXVoubMDG3T5XhaYOegFXwTysUw2YgKZFEmjXH/WalvjEb
0F6WJtYs0j8rnC5sjE/5TpFU9k6h5Sh4GHQqv9g0NUykxT+4474n8g4zGEoSIrvM
wkqdE1vAtib4a2Xiq4agrU5XN2ySpckRfXa3l/Dyp4Sj/fCBAMxq+Ll27d7XLYk1
6QVXvAld1X98TkznYXaWf9P8nUCe/R1xwtNMMkRgV0fhEHb7cIwGK0DJm+hgmK2d
PMjgt954GhyPlSzuX0sTrM9hzR3o8tTvLcq8Ek5HFYV1JK0FUSLxqsXKaKDik6W0
9FI9zs+qPGeGyW8pp/AiVXheUpNRXH+4aNDt/6BLpZFHOUxEc3gd8c97Ulnz7zG8
TXOvqmsewdTczkfy5CivO9HJ5Fg/z2sIgwpXU355MIEVSSid4R3GITHYCFbSDR0X
zHz5YYuQbJdNKkaoHeFAO3/KWznG3essll+V/diqVczanfE7Fq2SiC6QK81ZHtjU
UzVkBTIgCaJpooXojF0TKuPfejcEekSKBYp53y9ldu/Kfs1IB55rANpXHBHGk4a3
oZmcI/XieJl3suB0IjOsgKQcLMOW5h/JVBRfCuexQtalqv1RGaMC0XiWQeQfwCbz
B4wKhNnocDvxVF/+Yu6BPOx4QkStjMXwH6zlO1DDEUD9ybyrbpHp/pSr2TTEmY0Z
AFiaWGwCbGxOnxdO8C0ipAaYVwkRgpLRmotU+QRVzXbwxmCFvAAqPwjIJW6HCIZa
uSRgF3AwJw4GfK60gBOzSP3HEBwRAdsBCVuMkU1ZCW/0glsa/nfL1IJb1xyOUZSe
e28SCGJozBMo8I5IGAI/05JeHU1cxTVk4qhKapw7Neu3HfzRD+0ik2G8LVb6wz2x
5S9FZt8ErivK4If4wLiOYICi1aW+KIHi0vbSOsiI97Kpur6G3JsjZnKcyw3t/jzO
fg1OG87fNUrnty+wJc9KiL/RV9O5TRBRDqNFQeDJAk4o2U/e/tHNKr/Fq0kIQZEY
1FyXtKI3jivy3D6zquGeaoePLr5fdbal3cr4UV1tXXjcISIFKsu0mlGOwQPHZHpw
ku6YGb3H8ttyTYkoLaU8t5QDmDWMKTfM1A1CMFoAnzvawf8nrERbj2loKo7aN9ts
b2FZdDuo44xYfZBmllny2K2forum/c1LnlOFkcBUJLFD0g1MSWHrkOmn2p+No/kw
UnbnRBsWBAGaefbk/YKZSAMaa9+6Rzv2hqU+4zxSFvN9jPtRXVuFDseLBnPajfKh
R5oe3/fne2pRZv9DlbpxXM5K/uZrtPX6T1PYBo18PYHRYWHL2Al1ZMz2bJDwJ6/G
vQ/mm8wxYHSJuro/EO/lHXQlNFvZY3J0NAuAJTVKOn2+athZbYBQ2l02YnkHXgBG
3VCTEHg4gywG1JEsp8D0YRyhuamkBGGZ4jb2zGjfHJDqCB5o14+Q1WAhDaNewygO
L4GFMNLF7wllvr/BDYdNsE59QYuNWWTSV4zezdIV27T8z/2qEpo0SZGEMqBkP1f0
k8pypjLt3y/JEiIjcWwt77SXBEljUAr7af3QKmFmRnO7TUAPoDLdwazzKlB2LpQf
7c8rOQmBGxs7OnSRBmpm8ueSxWsag7XE2Yz1mtNGGYMD/D/axOjZWUXso7xzF4RS
ZOIrL9h8SsGG3z80/oQQzBFkRWfWXxyCVWYoOMe+ULV+0vKHc1QIbs+oXpG+PBYf
LHJ/0eQ0zBXlwyJSCiqpe3J6x6/SEBsEGfMR1QGiWDsYsX6mji4/7HuCRlDGBDkf
fxTZVEtVjcSy1RyNDohOZEhCeK98+a7mx7bZ2QXCvv/ixNtlVdCbk+YveFw4if98
y0Fbba1LkEARHShLJCGsN+lljZPwr0VcgHzGG1OceFXPxFQbnBDrsTylx5V6XLjM
Ie1t7uwkkr8z7J6cHA8xqFXrGVqqvUmbhiEMSSi+dwTLzFMQzC8+JwSNcYrCBnzT
Bm62kVbITnRM2lzjZy3rRr2gegrV2dQ+6bAWsF7upll2P3XFMwWrNINwjVBs+IrF
HXpz9ioCzPdaZg4zPJlATAENim7qsO1dSk6apZKMbt3U008+qVEr0s2wlIbyLXEY
HkatLmkMURHZDAwnHRXkuke/fpwOjPYdBiiS9M8yo/C0Gsm+25A0R2KfqqWEP3LG
PLxK3GA5SKfnbCJuxma1lutqOk4nDLWqcvSyF9bZenWATdlaEGOwFYgT5cQKd8h2
wOqhKcp4ms/ov9F3zRrH/4WnPA6kQVqof12NPbkB+pqmYElN2rIqGjv8Y85myBed
OJiiQR/YrzYgSZJfDL6FSDydXpGmlbmWD5MmzA8djB/vGKXWvCrMdnc82Nii2axz
2gm+VdEbotWbHQhJpj+srTvkUMsfgJdWxeh5ajGij4sXDn/Ev3pap/U1sbM17f3Z
gHhJlpJrEFrg87pZH3pPzOyAZfiRdmj3YKsBml7hLeROxh2sDwUU0OOIcwJLQHfO
RINrmyIoeQv9s1lo4eLgnQj9+W9nlzO6LUO6zlnAeKA9z3Xm3OluTo76EQlOytpc
SZo3reTRCFaXOroThvR8rP9cZua1VViYfXVnQ+GMjBeNSjnN4plWq8q3gzPyzmc9
CR379m2ZCcZ4ZDOfVDokUwT+sbdG26u9eRu8/ALSLWnSEAMzIi/rBLM90PrpH1mi
ygxrSUPML0+MQdKAh8IuQbY9e6nl4moV7iykkgnQeVOzikZeLHXsknshDlEat2pI
BpghikyApJunIn73qgf4BL2bUyvRvBWOhLQydSWT/Q80UfIxVGM7ogJt1Jr79FQa
6Mc06AkKpK5PuAEr4q275O2rndk4xSgSEF2F9eGJpaJKQqrh4VgiHNyq/2QSSK6a
Iq8CF+btvLziDROThI8BDjXi0dLdhvm8hEJtSXVwXth0cdlC7d/EMJgZGAMtdl7k
CgAR9SIkoI4Fn2MJ52WVjuKXQDTDYBboqvAvHeVauOxpJCF/w5Hr1p2TB5PoteoQ
Vpgwe76WPC2oQtb0jzuyZSDGgmk192aOXq8AWNkMX6m1PBxbnaYUTt5wFabDCXPD
DYiN0ggZQFibxOoCby1vBKajpZp9AcfRQht8NLjk6f9f6tqau6p6v2Od7CYcb7FT
cOK8A/0qIhluuQSlpoLpkcCcJ8RX539m8aGf95G/z7Lxh/UmmKgl7HRf8kCgooqw
2TqbhTDT/g5aXkGISu06pLi0QUPGKR0BMpGNR18dK5RwFgmxCK652YNxZjPlnF2R
apYVt7EnjwsfUA481/r6fK+dwm78DvKuUAPr9g1OAf6q0eudU4lcBjt1MC7PWgHo
luzIlttzKSNbf8MwCAWxq5GJBUI6ghSs37dSDRyHu6nlHbHpu0mOyhvXtJ00d/Ae
Wzjuycv36DA0bKrdIl8AkEtXoPqY7tefcdurnguq0H2JH1UdzwbQ6fl0hhFUujgy
G3AjN/3d9eYF0a0wutpQCkb20mrWeWKL2/zenmq5ULSEIsX9KQG3WG6Ea9Xk76Tb
Az1PbNi+LGo3V4n/+kP3xHv2AJMJIBjIqttprJ09YyDvNiuRA7HZzZVdxlk9+Blp
CEJPQO82XP4/4BrZ/gtwbNgkyKX0Ooxzke85kVnu/SWy0dDtsnzz6B2uCZKRzS2G
IqVcHjojDBTl6MwH0fRu0B6n+PQVKjw1hxtZfPgNjbDVQ9HrnoMNU9Fi/0xWNCJJ
dk4kD9LNBFA8VsNedv+O20RlPALQzPl/4BT5HyBzwLOUm3VtmwilXCjysJAYIAJM
NO4YbJ08LD7whSWrzG74st0ykL6gPKkZJJrPEYU1scIK55zJvJnW7Pvsl1on8bFc
nEOGJEenpRm0ZTIPJKmoSvHbhAegoyaajduqcxGkggMl5/YIMOhfzjpRZOa68QCD
eIBh6H+Xlwketnfh2dkNKP/0rxXEmcKevxAhibLXBugLZUhrPai2xulw/0LsuHLh
g8K7LaM93LWU8bS0zJq/DibvARCj7oBB+D8CZwk/2+QHAACtIwP44p25H94x1oPy
FBBuajjZBFCt5Br7FoTQvp+Jfx+UgdGTx61LnvzIoyejCoAuaj0+tgSpx0ltvMHk
vroT8/M/T5EZ2Z4CdAf5nBtyhaniltCXsgcZMwKe6KBuzyOstHZNwI4OQe1FB3It
YGWrxMisC8cgq3+vGVcR0cjzccZwY6pcnR2GOBnImu9Um/nJ0TdK4PolDEaRcS6y
yBErJ5DByePyjLQ6+mNA4byr7+/jcPnJ62vuYa+SYIdrasA6cdJNlv6GEfoxXYLr
N96/ZA5yUcDvTZkv83EdLhuB22rnRSIDXjdhN7C7Oxf0RwhDUwssLygaprBVe9hg
KSKsyQsklPoXbkqhdXBmG3oIw5C9iZ5H5ISJAU0Wxya3TK8Q65qKqnvpx//nllw1
tD9aZ89BKg6LR2ranbQkagQ4s241/Pjsi5bh7t0m3woZohxMZjjdZP5uqy1C2BP3
CEmuwenu9YjMhugWf9vybojtNAtddAPoGdseyD7T5q3BXvo9Gz5M1CcGf2HulE7x
ENfVSscyako0m0p/ServhXKq7r4xL1dTgvqPqMRGkIXg5Og9zc7XUk43kd+obywD
4JDUbhsbsst0MAGr5UUuRH/euXAmQNsrCU2jjOG87PXpfw9ZKIoX52y46vtZWxtD
vw711u/AKqtMYwGv+BGkve1pr9Jg3W16hUupQ2ZaCkgP5r2Wf+81EzQGHSNbo93z
B9uvldziy58WYyH6x7Oiyt4vd8qwOUE1f3JbBad326CPa+wTXN0NXkC6XqEjHsdb
PPa1eb6KId9pTqp/U3mdgJc/V3RcRcp4J8K94Q3ZSUP28MG/tBm902yCqoDDiuq3
sndVbAIeL0WYDM6Ldt+542weI5GG6ubCwBeF1P0ZTKIzwAQOSPnmBPKyU1+d7A9m
hvTt9Qkh1or2A2YmZ/0wBBYil298jcIlgwUaIV0Ch6GB3X56+DOGTvYqYxW11WtI
HUU1lAPoJk5n3dBBjdhBaE736AaOWsQy93vHuFoc58Bduenaqszvdd4VBACX9m/h
bFXFIGkZifky2bqcjLProP+e83Rfq2OiOQZicBRNMGu9dM+z3I/mXQHaPVCYLIgv
UXCb2sDQwlDZAKJ90OmYAgWOvrLrO85RwPVgpKZ+c9vIV80FLnjM/RnMt7bJVXJb
yGiO8/4XE+XvxnxXRvtqQ0neMo63gohw022aL9ZoTcCatioLXCx2RBAv3fwaFSP0
6Ny6A+2i+ZDLzUr7hfM1HbvwsAVUv6LAV3lm0Xc1/s4o3EIXtfttijpDjEKmf2qr
mayBHnVo02LWoZJmhjIiqV5HgsJgDkmibBNl8XC5XWPSzGTIcI4GxE3SKC+BwTkc
6xc9ec+KhlC8QQQDzfcM/UzeENPB8olpy0Z4w20+8cbo8Uf0qtk2EhEy6Fdcvef2
LO+e69jWwYE/SSwQrw3V7JX/KjlXrRJFe4Putdlvd5ZZYQH0zn7SPfmHjxGoazRx
AcYI9XFmLDpbz3Mxb4tHbbjyWfePohudbYr8QQ5INTmjMTUbtM5LHlKPH3gvrOG5
NmeophxcO6to4mfgDQbeU0GFPspkyrJ2SGgDCAFGFh5kPP3O2IjjcqBilRfW1faY
gJ4vHOKXHfiQojYARfhWeLQAkR+FUAdbz3zrGivZabElKAMNo/BVNw9zyQJBhriu
UU3MEjSkjh+XSwsd3ywKn23EzZFIJThnpNCQcedFSsun9blLp/b7J1qhjjvHZr4k
CZP2iz1sdP/nF2ETLVojCd2LDfQ1jUSlsgFZprc+GnXSG7Q7KfX2Xb+7SjqibgLy
WPksHrhknGJfYycEoWiJm9Pf9XoxzlYTqn9FFogA+nXKYc5w3YHjREWCit6tq/zJ
5uhvU7ATcc1EUll7mR4UOfY1z0eCZw6F45Qpm8KbLVf5oCnq15S6XVuvtO/d2iLW
a761g+36pnzr+OQlqE0x+GIrDgshxx8YMheWDxiqGdrTgVmT0xahaP5wpuGYPQ5F
BO/m+ajV4hN2eeDozZGv32xiLIr6cxD8qt7oRrlU2MDynNCSDSWxHaTVu3eP2Wio
4IiGwocljz/8IpNBUPsLg1RyZQ80Eia1PNhyZwwaWBh0Q+JHWmcm01Rvw+KaNWO+
6ksy2rLbHxU/E1MKJ3x1xQNrc/w+wZU3acYZrcacQVnSAXDLm1z5MQJlXnKjyRjk
kSu5hQGMdijvqQQYfLeRrrISGgZYE84Kxgg9cT/cSzR9hdGwAuyXz43uu3WZfQjs
o9dqZ6Z2rWNdLCpuAoV+gO6eqli6/TlrNkxIwj7GS8yBOQ3ohiKX1uSuqOfrEqg2
5te0p0Iwk+JjwALeH8UWuzFxo9C0abfCbMfVa0s6YqEjbRMtg3zqhRML6omemSgr
Nw7dROFnHkMHrCc/X0H3wKd1fAelNwQuf9Pz+ghLjg6PKC69L36XVXU/GMhsA7Zy
jHF2wbSuCOQwgcNtom8kNxYz1SVxBi2FaoX3Vbi/04u7Y0zlFv0YHwDJynTqhBRd
cyXGJGkOCL+u9fzS/xNINr7dr4fTevs77sNezWxc7QAhMsc55LOhv+uWcw+PzxBu
8Gq4t4ouKS2qr+FMfTQjTvH/cF4WmVxC9afeJ8gUEAcW8dVwPYnh23dF4RyWjUbz
jd7Oz/9N4f1hLLU2WaY9syqCcWC8bs/HfMSAieWxH2UqBfA5dA3V9dV+WEnm5SU2
jiryEmGLrvPQpj0iYWik22eydrzAlzXsY9hJ5ziyAI61FihIULljDFPKS8PBwAr9
qQ0xj4BtdGzGQqSBsvrtnuzNLcuOh2QS7bTksILV73iHnx0C+z+tZh54dooiUBjF
CpAFtEeY/e2kzA/Exys3BHyJsKiomRqVpxP+5zZ6zwN+wPC6edKTtNlHqSMiLTin
1t1gDx+DzilU5a0nTd2rXFLlbMpfXnCIOPaVbtLsCQKFmBkErj4QAqPL48sPM3wz
qZ4Kv3EwEzPsnkSGVp/HLi1FgzE7Ne0CqpazRmOibmCdHPcrZSzLcwsGMjdSq1Fq
noizVSniifyWdIqgEniPeRenmE3DJ8GcgOAGuaSIgapoGuGtluvPlo6owv9VC6Z1
I2IERsrxD8LDJJSkNqPcclcTaTWkO8tOZXFcGlnul2UuPE1mhA7v/nSZP9F2X682
Tpmgosq6arDVWApbGcNduq87IdbB9OF3uDsa484a6wk87ynxlzS9tSf21B4qMknf
calsc/9192Wtg5YTcn7MwGtPfrDq7YaemZR3qJqxSYBOnCykWgtt2g9SsE5Cvhar
0md6ky+C3RkXlwQZsQu3Y0HkCkrua54EI/mWsqwzV+JXXU4j3/Gef5XB3cJZ1z2o
DiA1JBQVUnLJluy1lI0EPFtlDgUEOAEY1+ZSRk9hyKKqrEvczjeDf5yS9/3IxMDv
37A3YdVzR4p3Jb+X9ygIL+YFQqNXqeW77DQJJlx8fa7QLEbxE8qPiaobv47qdpnS
kLNVroV7h4OiL0r+vyw06Q2qu++uUyiE3ydFOcfWJObwfe8upUTYz6+R1/GFyWvR
FbMEROvc4aAkQxjP9Fpj7g+y0yB+GR9lE3MuDBtcMHisrfBZ8O4p0m07jNyMtdSn
aKCOq5bv3kJOvgdmQ1zyCXZO0FwhquLoEJtfKhx1aPPLSuGyPPSpVONwtjfUkdxU
UOPJTYNGwnfJGfL5fQkUfa6ufXEERk2BoEdbbuNAvX9IbVUuCvN349Q0BP2IFRmJ
CTo5aZ4zuVDqpviMEqMGBLbzeJp18Gg4QccjQ4c+mXhKorE98db2spXcdNfvCQhQ
Lk1IAK5U86MWFXGKV766bqRlVK+u6ebJbF63A12tgkAq8e37leemMbtIvd2t+cqG
IouIGCbhHZMtUB2dS75PoJmcy3EfAtt7S9QtCO1reXSh1L9H4cIRWn/6YDOZtZhv
oStvscYVrJzIfuVcuoOee+nptYv9kdc9tKl4IRdRot5LCsXmJ1txBTCjQTZS5pP6
Se1YBnKZwrex0R62My6iMmAZdeoEPU6YDI9G37Au3S3d5OZCYqQkOvnXftiggQo9
P639/BNggG/9hJR3M90gUs3/NfGOwfS+3tTLKjue6GivHtcM8vi9E50ue2rLaLGg
tfOcBpaCEmBK9NgCl7xKoeYLWcjWa3vfCM7G6bIe7wmXnw3CWQLPQX2J3K6mwLzZ
vas6SQS/W/xcxTSIBwoNBN9OZUgnyIaKBmS60/8kFu/nBekm6dO0XE/YfK+PWq+d
Opdz2daIku9e/SDlcDCSmFGfzZIv/xXnBP9ZLRcL1Zdbpt2NDJRcOxIaz0o62HI5
wQaFqljb8pgWatYIPbKaUOlBE1y2sZvgxtDxNdRvS1/rzFMLImw297ubpRYF2hsI
AOQVK6r/Ae5xGbmq+huKjOQfbOkduUcFgFNBQGGHwsQUI2kS+AZafnJYq9dkfDl5
sX/6cQ0nCNlgf3q75Infqk96lac8qUjZxed/zFtySd81OXy2fx/SlHfjwnQra2H3
jxBm6Ckr+BV4qFj8fNjiutGAfjFVfhHI1twYDGyAh3yzDAqKBr6itOG3GFXKkCDy
DmenQM2F9DivdEtdmokj02zunwPFMjOR9cuHj0KHrgqVRNMdA9t+ifuUFt6UlcvK
xbpHXnZmoDhnbDLB0WAkxae0r2kWDx9mP+iINgblKrm1bkbHotPbIZztfaVBGS+T
7DxipnRp/e8YnmVEhGRF8NbcDXKDwvlTV1BC6fb6SCwaFPD0JWueEWSis0TO/Gdc
TUcIArfukVZ914jT13KxufEl0p6p5QQyN6y5WEbPg9nACTQ9tCAmHHA1ymsjGe7n
W3bomQ0ItbdiO9VfzS7EQdC8jb7dfLkYhSI2qZJIXHn0fvYy3HBHa6ml7k+KSfxL
XRYyEriHYRD/FgXx3A7PERmEIKedBMOGErhvpfOPmUysnCsopm9LcmsKeWqd3+r7
QYOfvTq2RKLEha5gWs9Zs+HAnVLCvBdO4OamfynLnI9off4/onTQUvqvB4320XaV
vyCbLEZ66ISBwI1pmEqbHUQYV99gVhgBUB1L9t8PhXSavcwA0s6cXtrznChFhc7R
INY8A8xRVEDY6oN1DMKaNN48RJGJxpGtusQNPz3ikoJRr1ZsHLK6vSYDNaAy+FNa
OmQKIA4mHkB1IUkPObmwX+IxPjF1Q9AsrvZldmWyMlrCrlXv2g7g61MYSw/WsHcT
QXsd9xKN9pIRUXQKVU86pbNWNwiisggrFTjvDwq/NRsaxhlB8PMoSS3h8HtCvd/s
Xx6QOzGhjQFKoT0bgl9jN0NCNxDPPxdIRVV0HcDeYjyrIQAwwxjtapAUxS/l263+
MDO7LHTKmMXZ9prHmIqhs40/J5ea44sCNCaWfghowQppZLOb4/AoBTkfOT8NBwg9
JaPNBgE4bfUjpqRss+5Llgi8IbvPb6zeLw+2qr3dwgnZ+infBCd7xhGJPBlET+SK
2txdoUzVdpicmQD+vOU5mzwqjqs+zdYNw8+KabPI2eZCdWnyD2qh0BPu26QQO27X
oG+ir2WxP8PVmeQEAgui6npwTFV2gDUB6MYrwIHsarwmew0toGGKosrAPwkQK6A3
aOXR8l7Qi6FR3WWrLf83oCFBKyQiJTer1vtMVTwiwIhzGEf02NJqVPn2NYLtZ4N9
NgNP+6SDKrSlxSv1Gnc3b1lQ72Q0hn0uTKLaS6FI1fKcvdzSUfIxC9F08jqspeLi
iGs5GGoBqQd5g3C1WJabSl5451S5vFlaXRGh8rIx5xeIMt5LVGUbdSejHLRJjRQ2
XmqMsnAFh6FEc+jxDLQRc9g9rqVOiPpFZfPrhLGmSa/hBlRF9iHgSqhX+iC3aeYh
5k674Ir/wOI99EAUwKjx+B/Ij5eIwjj7T5lbpbV25I7DwNNMnUD80I/vC94pMUql
Ls3X5Kwp3qw++LcE9L6A72evc0WU45I3qdFH2mPv2+L8S4I0KquEm4vdg1nQvRGj
GAHQ/E3X82zh1xqMBvQN9GvjfatJjjb0DyK48yfgXjtimchw+pTYhUDoRLr3txL9
glg+QtBjpg2UeC9UE5iDmw4wth4mspwuWu+EajV3wYoddy4hIQt2n2WP+Jqv88PV
acPEVx8jlf1oG7gA7SoHoA3UKpXqxv20zBwoC5W90edsjqR1ErLnkSVgpgzxr/yM
IyEXgx6QqqD4KmGjagF1gJOhpi+W4d0int+mrF/kGwLz3KX5t3sDV+TBeTNsCcpp
XsGub7u/j1sMCQQoXGG+R6QRiPLDug3dbq5wmP9146JFPzFTmfLOv3E3Fer8YPj5
Uo0vNKfEYhqe88Ah751Xn1ElL3OdXYruxl/JRvxYOnkiCBxuilcgZJgDowzxt5dV
ZB9eaaOUayylWXhRsOCS1ctbpBKS0o5NSwQ+2wXIupP+mLOqfBUwPpVA5mquvL5L
rbFDjDEpefbJdPeSavihlldF0FNGmaegzhhNYMD8c8Bicc/PKu4RbWnwaU0EuSHo
gOZwOR37ZYjq+XbLLF8dGwWatcxa5MhDhEoFEJp8VIiw3WJPqLEdNCI5NDFBP2vV
QawWKXYM9yp1/FLpIpviWTZJ/hmsffhCtT1LZSReUqs9H5Gl42glAT722VvvLxpK
556Rkx2fcLUBF1ejBuBzEMDhjqg8FVaX4WcG9RRyBW8YLtVTLh4/W/lsTCN2LOPW
ZlBIJNIkzrsbf04rdGegwkFVFc/Am+mxV5tPbhhdCfhz+1ZR5kNOcuw4D6IGY993
AJSFijdG+ha587t6oRppmVrSZdpcQSddsvAuzr6Hyge47Hgk8ATtSnV/WujHGck/
PZlYciaLXREuwR7XtRy3YSqWwYCVJ2uteNl2DZ14rusrMxaFqpSXqClUKATLUUVF
iQZPStk77MIFWl3DEOgKSu7zDE2jBfFHB9kBc6bTDwBeC3SdFhYtVslJVsmy2Mx5
UIH1hRQhqOwE7qDH+yh0LKeLsqasZvYILSr9iYjuoImHrPnOc8taNpdZ4TaYjFir
VEbMGzXr3giVwLQSSiUCcaYmFhtL8Ny/D8ufnk1iumdT8AwYBnJIwaI5tOzEkxsS
/OXOB/sBOfrCLdjsdGUHMlZF977Jny3cYbWIzcqM4/K/WqBlFi/qEmfh/5T0UEHV
Ha06RpEq2A6mlhsL9UYGt08XG8Rh3MtQs4uBH6eWfS59jEy5XHdlez+ByrgQCG5+
SSnOPBJjfux1H8ez0fJEHVQv5eyjLNaZwFbjQBJqF26PDJo84+dZfy6bQiM08j7t
VgHTUxE5u49gOYx3F0Fp1oXAQHM1mX94LCHXeCzGZh2aXui3JYNC4EjY/SZvE8FY
zpPXjMoBLhsndGE/nYaBrVyUBQJNSuEfCU24O5ocHh6Zf/2PRBHtYTkjYoTogmNl
g8aOEw8c6wc4VIompyHHliywfyy3tPOuFHKt5r6XP4YgOcAq4oWFJNDTwJHq1oRA
tw2AioquE10erCzPmHL3jOA0tz/dPZ35lAAiE86XsfaZkeoGHPZ5C1yEGs48VSyF
ba5EYPa7bcR+exBWUVJSGzhfikdyaWWmE9TsZOr44A9mcfSW5f0FYBT0B35jBG/i
p8SeCoXXTGecArXWeKGoRfwdI9WfsSWcLktxknLc20wV2jeWsYLT0sthZbG0K/Fg
sCGBBuPAw7iGQAtpnX3e80sOkwsWkLnrhny9X0FDU8AIqpwPEB0ZLehUEHhGYxRx
8eqhWj9ILYg+RrrkXbbNr0wPx3WfJsW+oDbjEjwxeQ+5sVGDa84rnoamsuY0BhjX
7pG8BIXXFOP/LuZ5GircDARJfYXAXhzd/jr5RU5X9RLyWFXvhX/czneicOFvddfA
rZFDjbtG2zyL1F4POGKXSLRAutGUnGCYiRatJYX+rmuma0jC+sp7Ypldqjr5oAtL
iOiK6PwFRer9wugNCxWS+BqQp0fimHwy55WhJGI9aMt7Nd0pIBiNeYE5i/QeDGq1
S1VH7bzbGQ8TGIUYe4hLHeC5Uaz7YQyOFcMD8qaqAT1LXEQnkY7IuJLs9/LjufFE
Zz71SihSHS/7HoJX7UWdGkvlAaQwLum89Lhhm2zJ8XvlXj694+fOEOQIaAuoKiin
NXAlQcbuYniZ0HLI8cwyY7HuBrOyLYFzMhg5QJQhVkHEvusxZUJeQE/peR946wRd
g+C097tx8d50gcUbn4J8GmJdv/A0ugXYpNwkfOXV8jgl9EVDYcqslpBEgkDaSlXg
5anhXPnqC/x/xS93UTZFD7FiRLZ9s1LAdn1Z6/xVqZ1bovO8GYV/vN8YIj2E5+8O
Tigbs19rzoxcglBXRJ8KrpotYqY3Npmuhrsg0fyRbYm2j0MWi3N23zsQxzVBnqYS
hZn/mkxt7MzGLBz5/5lrgWnp5VcvEjlcCN7AvfNne9ygxmZ8m/YHV4dfJTOzaV7p
5zog9UQHYbUOQ7Udl4yqYxT6ZdzEi3VKTGjb04PUYdHv2yQav4Z+GE20X2uTw3mD
yFiiXaCPBC0CvxLUbNZYjw9BW+01HgKZZevByRI5wVRqmJTRLmLdaSBZha8nzuY5
mpvqO7gNKHXizPbr7c6Wsw/duwnBfL+2znSK3gJyrWLYciGZa8JxvtMy9bd5NCMu
FneMnflUX7jdUAyHO4RJ5KaModXXKCVMghuZ7J48d/PV5b/t3WioXsjfkUl7pedd
vKW9GdTM0In3ceMozDwhamX+IOM60hjjip6RXDJwULL/U3/5Y0fe4eNvhPsvSCHF
3H55KBxR3zp2JT0l+IlfcGwVlJxBWKl+m+V6tQfR4uJ6jhPqxUXSybkF+Qw+h2zy
gfvZybvTYYp9drUxgCU4I5y+8rdyvK5CjnHoW6AIvERauI3jn/bvNG59OmgYV4+Z
9OrGAn3a8ucfAGCW0PoI0LzWMlCv8mYhSUm7JWaZG8yXk9M6GN7yYrQJFe8L5U7V
Y2HA/ymDWjBLnF/8ZzN01nHvzuNKWLOtnzOymKOmczbl6V8IH1k9p56ZvHbhI7KW
N0Lskily1cD0OrA0GXLsPUYW3xdpY9XX0FIa5E9jCLU96bhINFDc6W5I5miUZSPu
i847Q3MKtcB9G7dBYF4Q84n7hy77p0ln/78i4WHAOpL6hG2UXJgJdG4/3dCjLH4A
zE1PWM5ApCc46Xb5tzzazZ11S5pFcf1pGYJK+yTIn6bkcuwO8Irlh7zPRxAkcPRw
G2NUwNc+CdWqoHtlBEKvLArozNQq4jHGekk1NwpMVbqjCtZaww+9o4DJB9lE80GG
hj3yAV9QZGqEfVUTeT+HGjhr5A7pltrciiMhUCdp+XTlTPvaYi6J5iDZuvp5O0ba
F6l6p37PGSgywV048Y5ZUDyLTMr3MHku+2YNyI2gtHyKbqiYtgzzlyxmBREu6n6e
t1bxxj2prMQQNOnVUrSpJfELovdzAxkUYbeonnqigzUrMcf63C+NO3zR4XunSxMR
3gaxjBGMXsFIZPNXhTcUkeRfWZLnHGCD4FR326nqjpzNwXK/c9o4u5wEv/RK0Lva
6nWuRfJkV8Wfp4/ouErKMzxsjmyHbQ3aRXU5PfT2axoTi1UlxpNqJb8MVvuhwX16
O5/LTxF3lfho4gYyWGv3mzuBILijOeqISbBEPG0L9EEYr4K7U7vAS1QzuX2026eL
e8wGuYFcQtiQsfrxiO+vMS+vMwz8+kim1jlYR1StohyqD41VvS3k8QnELVCFMnOf
2+xQf2jLykHC7yYeew5NGXoMPwovdAsMAzq29SRwjlEuSUB9a4yjC7XyFZOg1Dye
hbk67IW+6wxJNr6Y3u/u02vX48PKxfT6pOLlS8K/DUZ4XA+GaqSR5jnwyJVnURHV
y+Ylf/0BX2cJXN0e05N9JTZuZz5tltE1+hvFA/WVSKSiBtEPQzMxMnPcYkFrwGZc
0VOd1SqLXGlbzcNmIH1OciI38sjoCmFrXZOptGPu6jTgnCotTpN0AotZRKLRFkFm
kYxyeB03L0k5KRjwnV4Xq/asrbhngKIbrRMg0Ax9ygXGOS3U06nlX2yd0vKroRZu
SHOb2AWGw4QPDt2PZadJZTHH33nz2MysCGO8FqYot+9OFniwsOtZ/BRLUdbKcCGH
7Zlqe68hNjAAABitOac14gjargAa5hBlbi0l27G5Vznnvs5Ulz2OAuwnDO2nR8hv
sAqZCRqiWj7LjKUq2kbATSBWfDE4n5Wr/4ivvDtQBsRXlCrcREkXLK2Bfqp0HrIC
pRBfNzdybM5o5QoFEX/67ZlMqSswxnMF9xSOgc6WmUe/LhZEBirUEMZbfEZW/rXf
CCdu2yFlIgQFKmG152WKAnI5L/kYiXCeqZymUhlKytAZPd0am9nWjekQNy1AQKBe
OscVNUYO+G/R71ZZsVyoqunf/aYamTa1rrPG4rRWs+4f5Un6jd/UKc/EVo6XLZmO
uDcYS9e38IDPPOTucWh5c0vq4oCNlety2EWXpjAWMpeBygKQ6Z89h7DY08XSkSbb
OYePlJFkEhpt9h2x8mG1oB2LgY0+7PPSJYQHdSlybZVJcQf3SGTbeM65SaDTUHo4
5RxpsA1pxIAySVAkU38ol74UGyERZdEfYaiNPI6IiW5RbA9T9LYYKrd9lBD+xUJc
0BnmD6SFOswp9seFND41OOXneHkzls+3zMTs8VMIx+ZICB3l+mEoQtQ2ROINvmUB
HcJqNL23v2SALBKUtgNp4qX9cxHrtq9nqyFPuB47q/d6xm2yIMjWb3iSdbbk4t1G
ZuFYP46EljiW20wtRkhzPiIFNjBEjFNpuxGeIZFiJ3d/rjskX+/QU9y2svmda7I1
mLpkMwNF6RaGwb/4H4hs3dnx0PsqIbUMDWWZpixpadpyObtIVJ5ofQFtvkkuqPPj
d9r0VzrRK8RswVk3xOwClhtiJsqMbgqTnzYRmse4aqr8J58/1gh3TOBYB0/fbZPD
4N2HDY5mZqRdEWSg0nTNd+DIXJVgyCGQIl25J/yzb6cp5CMOiGvUVP55P1k27TQP
vfoA/SOJ8UtqqtUGUiJMDamU/ZbU2MYR6PDwtzLtzoXQDSoc/G5S+XnzLrZzeMPG
eQEzyyLYy3NH/UovPcB+cD6c2lWDRhIjIYsW7e1pvm3jrSalgmvLF2xoz6vL2wLg
jMDfBdpR4L9csnE7fAnIse59ajlfVK1TkTx1KiE0KWzvUqDQhpFw/h8t5+bQt09q
N1hJkwqctXzyKFHslvcxtq0Qk3mlTl9iwQx+tUSxcJ4fkbT/MQFDELuO2WDQ3cNe
Fvm7mMSv0oOzoSUEvhS99Etl7IYqkRWKs3XNEPE6nxJYo/nnOpCOJJOdq5zb0r33
/QRMlfwkpwDK+/YfD0bqApMNZG7Pp7ljMDZoWr2pPXHzwGN7ZO4h+8VbRt/cEHBa
YxaW5VoWOIn1+3N7O1sMPnLq9X0/gZxpk6gzCCF0v5aCUGHn474sgYpJOUEx4dqn
tpz42auTy2scDQapj6YyrF2clcFO+Y55zBRcezBfb0xbNwTOG4P1Ro4BN884Y5iD
CWBaxvc3xqIvw4Yeb5IDJJrzap/yj9iP6Y6N+r6bz3L38z4lFGIyLoZHCv3NZKnJ
ZMCBhBAsWBp/Wxf0AOXIIUPZu23w2qDQT9JBR5nNYOXF3p8AukW4xxqlf2DwRdsf
SOibJFYH/p+SVeyumZBShmD51nBgLsYBg3lNcfzdN2s4WDss0K9a4iue/VjQ5eyN
bgYB4ysxxJR06RHIuSB2A9UIY12cxEVYcOPPj1v9+e3FS/1hE2O4ZCAQxPXgCSBE
xeabFRCwYOVEl38Tc6eumAKg6WnkSYPUmj7CxfSsAo4xl11EbjlXI8wwow+ynQz8
7nP/92gHixYtq0VS8o4SXRL2iaqV8hY+wOTpbSeJRmiC6Eip99KTUQB2AWmqjO3a
2YnsbKWO4XKQP2BFeJKJWgbqHGPhjg3L+GdnsHFTY/QGGWIHtGukizdsLEQq3rLe
W8iys8TUdhWPhpLpTpm92lxoEKqOSgaPJA+wTu/ChWyy3GAYgO/qCPaZPV99m6k8
yFsVGjOZ402k6SfKKLFZ5Gu932T5zdfE3ZrfcHkiB53fjCHFePOVwGsBsSF0hFqI
YYKY+nYJMwZG/rGIjUAiHzuM+op6kGGrLz0UUMbI+P+tqDlaiclQuE67vw0FoT5u
Fpp0KfzBpWSwbBGAoBZoL8wjVug2+9B1ioQargHzR+qgJuOr/jru18qgjUGUZAOS
qJofsLoEfEbre9PVOIkzExnNd3s7AHpi1LM3Pjg3aaHldZNtmV1Px5d6AdRee0bQ
Jo6eiwB5z4v+I+O1a3vnz000MjGynp62EpyO86MPdREB+gZmy1905Hekvrxkf1Dy
gsrljvmDdvtzGAKzAPdMMFe4aCeKeFbTQl7I6QNl3I2+Y4V/Vb8WHjvGqf1pVZie
3bMFkMuFqjCN8bhsjfiocDbOPnuOeg47n+caiyGSzx7JPBHapIOl7NmivVLcEDeR
jTk/U4f7jgBv3o2qEs0TotSFJR8DWMpjYbCwHyclTvPXRMfbNgyMFLvC04sveVlB
EXXx6ARibonVmW9CNv8cqlo1TZGJvgYxc90ApCLNUz4QO2D/E+P25Js27YCO27uv
chr019Fro3Fozz/WZznJq6J0LzaponohWAUwfEr8JUBOaqk7ip66FhBG4KF0j/nB
gKDUpV85dfPkHKZfnsfN7zoblWxRD7tQg9Nl7/UlZuJrlXQ0qjhFcjbGxgvm87OY
vN/QCqcCITGP9HDQ2/ARzIrgSsdx+zlS46NGjsAMsb+e0JUeXIwBBs/awnK/4p2J
JL8krfBQPbr0zGxvEfoX6FBtHk4pBiOscJAjKCM5Mp6OVoVLansRdOZpvpFEESAO
BssJ/FHc6/bIJY/7tcTNboxvgdx8xrHOfFwWf0nqT9paSzq2hd/kS/7NQft20Q/T
emYkFYJFvSxWAXJgj6cpaqi9miQyPHETLMiwn7iMWvnyMoJMne9ob5mxttWAU26V
ShqYAbQK/TczVga6ls9IyItzW7BhDqk4AvYKn/dvjqw1gVw+Ta3DVwKfaadT8Fii
z2f0zKWNnUqH0l7ak7m5MUChduccXAvR4vJPwxq5GceNP48y+qygk1ngg1zhdsVX
M57usJJBw69Zd+6cOaC8+EAJLr90YSWaYtQLUE0CmTzeFxmm2SzjxtXk+c+akfqc
zscBkUgeQ+/FzXlZjGVF/DHulG8aiexkg1wnzdm/XzItXfJJvkn8DpzWCghMCzFV
tTfVE5AFAIREftK4bGl4Kpao5DWrqslyB2CXv/ynQFfK6BL1plS7oXNTP0ORoKFR
kg+lJRpKETkEWoX4jmvpMXOLG18xHHtw4KFgs456fuNo4htH98Y4RZVWP9Q9/HT+
l4RsBSJrKFMeADXk3RZaRkUaVCk7gSF+rmWV7nw+ADguY3KppfivbIYabzPc6w1C
VNLZEXltNfp4R64JPaFHBuoIXuH2g5b2+dYyWccQdYwSWnAlh+B45WH6LqX+wmlD
1fNiBojlJw8CIifOJHH7RS1EwJROyvjI0/GVDxo6uavoaRBwK4bsSOXNrsUIABrJ
ChBKfBhSIZWgHwN7Mm9PqEx5PAw0qub8I/OT/dRgnfPfDbNyk5Ue2a50aBX1EO7f
kHnVasyZNIKl7QhTST34GsGUKFngqNT2rnFAwIW+TKZ6kWxt7iWeD3nbCd31a5c1
hZl5HeZNd9m8Tu1QGbsTHJO0Yozl5U7JkZ84lHWxbkMhal3dyKEGMnr0qqs6szhK
kL9Z6hzOJLWU27cF7BbMFcUaNi4Z02hzJ62tYj11ghMED9dvxi9gSpTfP97/tBWC
7QRuj1WLtDmHPGQJVhI8NfQDOu27sZsnLGw9wVhFALHD5dkgbJS7P5lFszTr6vTl
3nvILCLg123ltYJEYsPv0eYi/p/WbQa1mp83Mdz7hRZvlnLEcQANrZLd4TOPXJTu
VVXoqvIJEI46+FLM//qgvLrVTmUlpzGmjPzHInW3HOmPZOebNKi3/ujTG858gx/U
KPvSI8p7Ocf65rOQXQh2xbnlg3J/C8tViYHueKdmUau7kC8a5lwdjMqKK/azLQDx
OGMegG9oTjts0r3QpdOAJiX+DdiLFH/0Rm0A01krrJwT7iPREWoXkmj95qplnUDZ
nIS7+2iD2cFaNpDVlJZoi9z6FaaE6o0N9NjdUKGeRTDMNqvKaWJFYHVQHIHVhUuj
2Libqe2XIGUo5bi26Yhe8X/XEHh4eCHmng+HPSNA4DSM/+mnCCr+V0RP4QerL+Bi
DY/VLPb5/DYwfIONrpT+8TrJznH/uIOyWNfRZdZQfehHUzXDH0NfR0tQ3HKBjopW
bhPHAesCXxVoKOwiyDbMvhvWUdoOYx9Tjq1N17HdQN0mD8py4g9joeXYUFVdynlP
DfB9Ti0OrHZWqx87FiMCZK41PtKl4QZdUV5B8GqcjfeLChLxpG/yhJJLQY5F2pvy
oLA+an5SPJzFk2YAGc/klVSzb+INA6Ywg6nRmb5WVPyascaXQJoxQxpIQ4DB8hLo
a5JoPCipKVwNa1hgFm9iiNU6XiOJeF99WsJ/xL0ZjRony+ZaJn3+zFXUtf2RuCrz
AFY/OfvPb36nGevCPz5Ddya536sNpjh+mFpqX9EdTDZZuUILONuPfCjOCk6FN6sW
ghaTtMs0LU1yho3tjPo5NY1knen2pKYpoq3c5foe22AGfbM08bnGIx0nzZxEm4cY
Np0OlbOenwhulbKQ4BO02H+5MdOwt/wNQpo5ZRQSwJ+Pt7me0S+gi22KEdmABck6
G+9fE536nB8315dUtZfGIwNzVzTYEQppvoJc6VrbEw2mucGNWviMOZOGKPEUvrG1
5erDKC7fDO16wB+I0zw40xilKAgPWfQ/apEMTX9VxS+ac06oW1Q+mgCOolEJn0vs
3F3spCNcJkYHiZONJJlJ1MGbRHxoVZp6qom5pUgFcTQ8K6VF8V9ZnpZy7Y8E+KG+
BCMH5OeunINzSB3FkYCghzYsQsYrqYNbc86PnNyjx4VYWmzxmCfs7ArW8ygfoNLc
VghMaoZfoj/PCR3Sdo8uu7uzfFE5BbgPiJsF7uII+lsmYqAqymJHUL0drS2QzIXW
BgMZoemw5m343Z/ZD7a1upkiV2/e9sS68Uu8A0X2/LmAkVhaPdcCnylXyJnCow4K
eCx/ytJa6Nhl7+40Gd/pxj1/rJMHSUkBwWurDRL2wVyzpg3Nq5skQ22zRKG+jlWJ
RhoLfkia/OoAWh3UXPzzG9inJvebcjgYbS07djG6g/Kc5Wq7RjnYA5yfqL2Qv7PN
vgo/VjYPjbpdM/gDdYa2c2DlrmmXchsIAiY00/OaDvcUydNZ3HuYRmjf10n3Is+9
M/3F5cvKby/6/MJ+9sgyQf19rO19P5rIGrYmYbZTJm1cXnJ3yQMr2oJ3r623BzWP
CdyQ6KCfnU9hfq0WpiJllJorf5E1Nv6/wt3Pc9LHpq3tuGgmJszH5VKf6/mdcMrD
LjcUuVRJ7CbKt83re/SBZlU7V5wLrXrXT0k/Dh5A1nJrWwSHnBHDB/1U6ROPUiHk
KJSCbYJIqUKbGuex/sNscEJUC7pWJLao5bNY6pDdQrnz4ee5a10ir7XNyMsc399X
mcoZ2JPDiaQptgEXfMw5rrI4//7NeILNRnCJH54x8OY2v962uRfh7cng4jOIc3/v
+nFKU5S8QEmIIKI9GOQ757zovtWrRh3xboEo1jOcL2Ot7L7xhp1OHK/h+6N5FxTI
Xz+CcBbOOZSBTd94S0KrvQVLDEHl89/YJk1VmHXTIJSu1nffemj+WyY79x37b3Q2
RxKxamSFG1YbFeoOPy0aUQH+pRq+P9rO/vQ2+hhdYIHQ7r+B2CkjgIAr7mi87xSr
udLHDppNGhEe77b13UgF/3Gl5Yub1UpR/FaGvrZFBRYglICNPUDdQl5CB9jI5h8T
hja52YQbgIXVheowwWBwJO3wq+NwCJQvgkJI1ei49olfAifufOdgnLVs7W0HS6xU
XZK0vX0DiyzzUjx9U1xnZ6BBLPOpDxzvE+J/zXCxet3rkjqU/jXhQijxIG2FyMAK
ynFo3sYe6Q5CRvRZS+n1hkPGaik2yZMg1T2y/o28Y/GEQFDWrXfhhwvXDorv3D6L
SjWho6P1JoLwS+1hwO4e5+H2lGwN2RmNPsbxHKxlU/xmkQglD6eC+XjAL0qeVAXZ
CcjSdU7ZKuqdkEbpo4W0GyJS9VicdgXezd48ygpHKMyIE7003+ywtjKGIsGkodyg
Oe5tNH3vsVa+JNhitlIAQVEtytGUhV4HI8DKMVFMGO27rzvEYnl8Y3WX+s56zdxg
PkLbesUBnCQDwYlDPrQz+lWY5KA+X4DI8DSlEEVQm8mTN0DyEYnp3YbZjNQtvSQw
JJOOdezXg5VlScPmv3ZSxcN6/++RfQwoM4nCRAax4jsFPqo7yqOZKQN3Yj4UVv4R
s+VlRyhq5glgfcT0S7rHp7tgMecGf0HZiElrl0u+rkHUkoIAdBicXpde8JzIelmi
swH+5BTxNC2c978tq0TQUAWR2zUjC2PKVtcPsv2mSvyB/7Kiyvvt7Idu2z/fa5Wv
MdM0NuZbAJrIQ/n+kOac0uBep008tVidQQFXWLWeDb/jxtu6ElslgHx1HcfGrU26
D/NyuInDynX7ougWwUkj2XcG/Y/x6S1tXm9SCV171dddrj5o6tYXKYQlihNII17G
zSHBixrBaO8FwqNytqmMgCszGc1s4zk44/DgZMYMrhTx85IcMAR6OWWpMKdCe4N4
KsC4iNebAG2FXHgPgItWASGy+u1rPiaeR/psruBK2rM/lVrut7bbi9oXcoZ2gM2Y
pe/vXqimqIiXNTJJUxBPXUwuWuGns42WwefaDcyrkQIEzuilLltb37+qkd/hmPG2
8233yA8TLtkHIjbhKgrEGesIpNHrLHnfO7bPK0XwqB4Qt8C35CzofPF4u+2QKaZI
4NCJE9HfpVOHwRtAbBwvpDu+OPHF4VcftpyViZRjSknJpyVVVtymGwId/CJGyKDs
jL2OLIQWizyFnELC2XbaQgMSZl07coJysj5DFscwfkZN9muNPvsxGntBvJNrpLMl
tOmPOLbeuRVQgd8psVoMdeLyso+qgrHMe6tB3uaYTzdLvsVlTKiTVSKJFWKzJFWV
yYOb/KuHHCn+9NqtEF/c4m3f98DO0Kl+a/tZ/n3H/RuTsy8fhlKa04hSMgRUDiJc
5aFTFKRwZD2qEr61QCkSSawP+1DeMa+gq/7yrC3cp+rt8Jmq9qbJoTx5iFs8nAL2
GkKzwHsTYEgjLKCSjiqoUdyIP6gcpGmWw0KI5Tc5zzh1U9hp2EtbR9tLI9fXTT/Y
vvEZLSornlH0m0RsCPHaYDoVnzqvQYw0DwRyZt4UiCU3zaxH6djjC7CVWtW9+cNX
QsgvFyUnQOXY3bZv+i1CxBT1hWM/bX7QPjegDG7TzSerKgf5VRf/zYVgF/fX1kXJ
7I9IwJbchBgQQOZraX7pa2bJdd8caKBRj3UDWYd+QR+81iQNILOcFdk7gl/vlwyY
dh0oRrMsu6rsW9d/kstwQI/BZ69LOTN7Ro5nef0KbAPfMYvroJERNucmwJ1zZl6C
SixSq/NL6K7Jw9u7jiis/6/SkBNTIdIbXnXzVymFzAyRVjv6qpnJgu+7g8eaXtV7
RuZeYEJWHO+eJfJkEUgo8V9UpefPeV+fI6G+3QXclPxaxhjcSh8qQHQ/KqcLl/5g
4NchkFBX9WiGUop4SP+v6k9MKiWFhIpZoFan07TJ7XcMZgWPhl3TPgBlusxbwzax
sAeOmUAlseneL0cBsyLRYirNabI+4gTi+duSFhmS51uiDU34gL6sRUSESPBvTZlE
cpt4+Oy+63ZYuNUH8r70YTpbcNPU9WkmCtw94AkBxNn106dUKi4+JdkloQuIDKPj
kYwqNpd8H2ctxxO+m28fJ47wEDrE6UrcnHXaPtV/pKXQLD7M/cBqf55NEg+4fmpp
yMDG+QAhqgHBwwMqkxAq30QeBwrhSzrkvptbHdDzGSxNkKd8VH3ZK/YGRtZCJwLE
mEoGzl4wNaicNEpI2UQxZFvL6zyMzVmVdox6LMFxWJ9o7wRIpqJilxwu5RQ6jock
Dmw2iG9rUlVZWkTI4Tn64bOdo1WSFqcRIkQD48vDsyZkOuVTNZWaUCU1JbefmH1i
s9gJdslCU21CYYXn9AOdbTUzeY0dymoxQrCF2VG02vk1bT0KylLk8rGQYIAOoloK
T1MaKkMYmbYWmLfrcL4wu1MuOykq7a6MSQ66X4tJW+Jkf9FGKK8JCw+anBotzVWU
EsVAjdAyrpLT1ulQhYlqalGY/aW9M3GldGQfWmMciwZUUhcy5DyBZ10Z1j72g/+P
8W57u1MznLQZ3CjPgOg/s5NeTWsC8HIuuKZL7l5Wm6VyxtpFSsL9rDq2HDLHBSQl
YD7uyRoMABaFRMkqwopMy3X0t5zG+nzimAr4aqiP2+qlR4l9IiH8BRv5fx8rzP2V
GasZ8Ety0SbRhj9ewHnSQDNKtxCrNhuB41ouUdkgLvmPjfkbnrOxJY4J3IrtQpYF
3EPMLSCARCVFHLfH+S41VAAMdz7esXycjzpGpSu1LfjsPWrZDKj/5HKWX2aGY0do
KiOB4IyBLfkz1BGWvxbNNkEQzGwGK8xqvrAwX38z64EEZccee+h9Ccr+8pIVDa5R
Y0mRMcuxpDddjzmJLa3Z6yfGxgrqfnHreCphL8AQhV7waivpAdGZcAYvh9CeCibP
yat58pxdile3BRldgFMHRZktz3ZgLLHtmYJpXkE85Uu+e93fACF0ZtV5izepwRqx
VjcxyZkl+LAYWDYiGCQiVtpPtDhZdxXEgv9dCvF/pvnHnzOVs1AGRAsXWLKL0VWm
77phBVMV2gL4jA/86CTlfIhXBZfmpowHAqqcUdbrG6YndBldmFGty4RSDgKEJM+D
amV3HLL0gCKqL8xseDQQv1q8a1DsxvGd1jrJ8qsuwnvKJxE+UZZ1bfqiM7Cx59Wc
7XZOJUSCcoQ/tPUvuVEzC8mGeOuPDZCKMH5S4pfZNI1dwUvyqlomkuXhn7EMYQjO
BFQoM+wNJNDFuSwO+5qgVu/YooFkCP2vPN22F0uXXr2B20ib+wSlKY2eZjCROXEp
kmKuNRkHfWStmOSiU3GtU8bjfbsyS5hFhA1oNKww+mFweMsRWkSsb0kV/ZWQIRK3
TBIg7Edig7qXLTsMSJRMXnLh0R9Auj9DpA2tkMZ7vKbffZuR2CildhMaQ4Pw8VsV
8t1vLjcDZ/0uqSGhF+OdJw2CtvuSiIaNZ5IEr36lTfXGtrRNqAjV8mo/eslc+gxj
MW/szKOLNUsUwCnOr3bTutJYI4n3Cg0CaZcJvnStkBXXlyKYm6feRImW9UXEKePA
xx2dRjooFPDQ4OkIKdwhneRX6MNKUTBCCSVD07sHHXIlj+mLdL3nxG0KwtoQZTIb
8uUbOhRpQB9E5q15WzfN4xudulRGK7YmKsf698nKItVBsW6WqQTWLL4FD9T5K7wt
fwhLqyhkSQk4Q/jIhETNEKUvj6wgBPDJx0cn7HrcV946KvBultLJM4nQmAfwyM+b
6avwxx/lHik4prUiaXIIK6vjkvp0MgfQbnQ6Ibl+LF8uYhCxSDNDwlw8C6RkJtp4
sTYaXVdwSDBGsBQLzzRupcIQrhuEr19IbKJfB5KkwaCODBuFm+C4JVd3d4bHdD7W
YhUSJ4sBmXB4A3EGXUekRsdw5vCfOv7aY2O9dXA9ht6foSihNsvc8m4/pXZc4nse
vz3BZ4TpkdD/l4IhBqNkMElKCCIwfKAXTTEzsmJcU/2G8AzkMzJCNWUxyCnkpWVw
3uVGqOXki5l0bp7yTKE8zD5oJaD/4FivLs4FUGucaV0RQxbxueB275NdO3tWYi2V
pU67pKI2ehQHDdqKDcVtD+X/x6Z6UnWyBVA8+/IeKRT7EV9zA+3tEt/dNs6cBQVN
fBBvCKGXdkMJhRS+weewDI3sNFNUdaBGvswE+qoEHjqlzFdN01TQ2xKpDDnyOzIZ
g7MHexcAFqvIsD2ZikSLhOJK6NgdvA+Nw2nFsQrMkpm9+8j6B0GDkECK1DjyWIFU
A9nkfWN0kLfM9kZ5yua0uyolRM+M65eHA37xEKe6mNQH7HFLAX9zVigvEqX3zXgl
0wj7az+BjxZpJRxhcSA7FnOqHkKhVzP0VtVVhBhFsmdyQ6qHkGojx8wR8PNTD8gu
t8qpTkX+K3WKK924Amne2pSkPIHDsm/TLnOlDt7sPMMVBwmPz4ZQZ7CRCDll8onU
ZqwwB3Bey67EC2uiMydmEaDGeNx5rbN2Se7gVzqk1XqSV0Exzf12Bo7ovQ5u2XAH
V/bgDeh1JRD8TmDjbpQmAaXtlc9WnS1xAbE+1+9mFpUubdpHUi5KgBPHfge9rCx5
C3UmrYChK9I35YEDMl6BIMHvvF37JukEVFWjR2agSgy+coxSF+FD/VwYt320i91w
Inyvy5lxUfY29Iv+pQfK7/VA4enpGpAxkNZSDXlfbl1wFvwDcqSxKGCriG6NByDe
IXywdoBXHQ1MhpdSGO76wUszfzGJyucKWcYBtR/cj3Wp3FdFcN3Le7cnfljGZjkE
5KFuEW45PXXUqTvWvBuLiHWKzBVi4XjNlhzFx53jVg3+7thPBG9jxJNLJBan8r3t
ieb6N1betAP0MlJD0bfuRkJXHj6q9LRL8MwfKbWJIBFrOlS2dwgD9tdesf259ZRq
YgKfjzJVUlZsWC7UEw9W8MHYqYPvzbrhKRBzxvqtjyznj8ysQvQ5C7EX/i1CUYux
dGP3CwK5Os497fUKwrpV9RF0jCVo4fu6P4ZENSQR+5r0sQDCkF2U4G1Eh0jy7woU
p3FCj38/+DsWDVy00p/2nn83+QexfLHLXGyUxiU+zf8PPKAfl8p3GV6IpKhrqFIM
8dZD5PC82zfy2/irAAbv2jB637/O5TZSEK95faS1pR5weJ7OzXtMYtEmocKc1Q6d
F6nIXhCQgiRM13N4LKU/9ce/ewCGhwfa4uNfdcXL76GBSoUCJAPU29UAmtEd8cLa
DdDBX4XP0JKh2kcZIIGwelUeLw3h7GhVzjRs/5/QG9KrAB41NSyFjDjmngaDk6CP
pYvmf/XTPzxe9I9adA3bqHDfsXxNNZR0/EJ0+LnLd/rZbbQCkYuYoRjXFLz8YGNk
1J6KEewE/C/GGIxoOQoBS+j6p4ORuN1MW1/pvp9HaqLJVaPaPIAdqpL+oLfrFZIZ
ia++WNopRAy0+7JUnYbrOawBnu2I9Ql4d+B5NMIx7FJY+OiNAtg+LmhGfb6jbmCJ
G7NSXaC0hlrQWcbfHcqHONEdJP5iDbzKVgZrOVzlSStor/rBXepV/TB+DiLNy/FF
7Ao8m1VLy6z8yatbzCC+2YGEK0NrGPJ7W0wqv//+fjfRcRgEJGZqLqDPBQPIqf1C
AaYCOFMajV6499C19ZppfOtTAIoJ058EFh8d0vFmuGsMbKsx4zWmQfDGB+aYp6wP
H8K8AmFUR+F/+/sdnSRiJNwgCLHUnySrrGx/MmYgEipz3H9+tYak2Kz2Dy/x7vAo
gJT+NzK8sE4yfXxgeFBhbGPSx4Tw+SmuvlntDQwt20h6lQrK+8EwsinWVV0FwYp9
79sTi40HUSx/S+Row1awd0Gw3qvNuVeXrFTQ+uBopMdR21S6eqIb4+/epKepdNcs
Uh2ItiFGMM0M96Q0d38qo4ZOEZ6T6JoD72Nc2F2dYBUgfXMJV6Addi5Wp+FF0nn/
wDKgvty8nDiB99QzMk9UJY1rAdYfIIyZuHgds6DN9lc7YhQRRK2b0zoaEAZdgJ/F
eBHen207NaBfeRwzhg3tF68qu6jQUSUdaiUzIEuHzmdWR/gf2Roln1FqxxKPLADH
oq5SMLy3Pf5iM6QMKTSgZ6/IUK6rjeK09oXbrGqw7UOYIP3Cxl9ES7QAmPL1dE3g
+V0zS0MP5b7JG/Fv3lPQUwfCtOLJ/PZf9g9JP6gTwTKmTM4AedbbGeDTBrwqvB4J
CU05igIQ/DglAMQi6qDhuUVU3EmOBja9N4uy+XElSDbRHHMPtprKyZ3EjF/UeOAQ
l1p3wn/n3ZUVdbK+hrsXGbd5R0Dnv1vy4OvPcG2KeEh43NCK/hjEbAWSpdQidI1Y
yyEo0I+nUdo2cY6SjvyWGneOKEoCZEVR5v9X25wdQtE6715d/x85IC/ovco/1bpi
srl93/gyrjnbCZo2jP/AU+TOhitXJVgolvBg08z9F0W5iDz2h35euFpMx8xFS2K2
s7P/Z+gzjoidf/fIjiFcNQsOMG08MgpZjBNaCeRUUyTSXtU2jBN1mcMZNXUAWW3I
D9/rAOZMNecq9d5PY9isv226Ky9mYs73wtiO50i/DB6MzvxCz5qLLLtUKaDzuoFT
sdfWcVCcmHZfPXuLLcsm16zp2+IBQOho+r6hRSL8fMm8rj0fvawz4miFUU2zttYS
eaXf3Vl3YJYUrw0Pe9L72UV9qzNb6mPbyjnA2lFpkIQxcL7byd3qxKevV8xS0LSC
7cRNAKfelRlvgWzSBF6aJON/6du2HttvxUJv8rlWJbM89I9McBsefypA0d2EfQ2C
k8MUWe4Ilh13X+e05RlvkxTi5Cu/YOaZ+e0G3DUHLzSmiHHdStNLIOTWGh40pJG+
4jdF51UN0odFNfoGVDXn9S1dMr0EB+VIlY/T3xP77I57c1u/pljM0SW4mNituSDV
nDghagpH7Cs20o55ifS0KhBWIw9zl9MmsoIToHbDAGH8ZRK2sPm0kdUGAFmsRkAP
KD+IoSZp7NbwnznqBo1FFLhfk02P7YkaOGf2oWSSHv/iWPuvPjFBdEcPV8Wl7Hrv
tfPGS4Wk3HzD729+HgPHlczUZJ6vDFI+MORkQDcBLxJvsQZ/MDH/d+eRWg3zCZ23
DH2rbEuJ614L7zb5gws5BVjBlWDwOshW/G0LRUghsGdOXSvaiybHwv9uSA9pCkh2
wmVzNHrGMgx1Xjoqjte1WP+jPiJk0EIt78fGiH4vM9z8i1tZqTzH0nk2z1gtJEK/
dyleQ48SodEn5npg3uf2Aazh6E9d8Sm9xjE+48F4y53UAbSJbKEiy/m/876KsMS5
Nr6yV+0Kx0yMI/De51Xrq6wKvRvCYyysAlOdxYTjx5U7MhAi0AedQD3tlV0DoecD
FKhoILQDGF50o+Wa/w5DvWbEZbsm4PvLRWx6z4vPlOhUAvMyOTGLrCknPdKBQeoY
+CtbWRKrLdsEww1WK3/pLtKgwVYBkBExKPyzjSZ9EvjFj/ktXIJL7WZCd6bHMkNk
uFT0e553u7uh5iZe4QP4XSW1dXx9dT3PbzoGvRcWDtlUaz5FKRAVJ07tskM6P7sg
muXy9Yy/7S6QtdutW3IIAp/QmONCTSFLfGBbfyc5eHOFfp0BEw74eMe0e49J/Vpt
M0T+ddNMzNNHk0P2Hyx2+/2VC5TevVjmxnXjE2yk4vJpyvlXG6jtv/IYYbHuLpIQ
xVj0pTsK3ccRoq7lT12d+mCD4Vv6CDpsHuBqVMKioJ+KFyImtIIsnm9DamVV6TAX
ueThHT9Fkl9YQ7JgXX+ZEyOYL4ibV6b5/aIM1PkVTvGauJIrjrVzFJ1kcPaPervA
pI9vBOAQLIP9mqApQuPNtlGuczdydWURb5+N4fHUOrX/greLz5aitvKqJAXON81o
3Jtvd2/70NwxaJuNBX+wRboGuBG2qUoKhEtj+5wnBiPbATh5Hku9jTPjBfyvP3nV
u0vzJLGVBot1XY/XvacdqNHv8uDwnHM/PYE0ZIkq2xfw8g1Vuhb0Gk0mioK/M+8i
kf0TeaylgsGCUVPgbCHsC6UyVOP0fTi96UVJ8NTkbN/zUsX90HeKSbx8sTtP1mvi
HffTkbtNvQyW/Ds5V2086gJ+J5ZG3x447zSMoMQ0vGfksYZywHr6VYiRJu5uho9a
vH1TKqne04OEZGlq8+ORIWcO/A+tNnD9BILzGPkSficCRKclTBy1Oo/NRhJ/tvPA
JD4qU6sydcxiz7vvY83g6TAlq9w7a9t+4RoVzYzu13LQdWGOan/hjL6cctKhe25y
WgD+dEGnP6/hCX1pzbB/tdWID28ozpeTLNxWAWBL04PHRO94tT6u7ef/KNunKQnL
3K819f7uOUNE6d93YT5sLBeppwDGPra86gbwBSV2TATcqn7zt6cfDkn5MChqP2LG
066O8NbCyK3/nAtCrQPhnVKl2Zr/WU3HJgWjydhge+2ZTJJlbD1IRDNbJwk1s3Wm
eNceRDTGqJ7vOFpSllrGbBk5SW0qVdeGI6SkjzBOkJzksHfzxuVlscebuVoBcyq7
W6jKfyVMc6pbgOXV1qh0uwE16WpdCfFJzM3Hd4mkcssK/Z7kzKcpU1aE2e3BSChG
/q2knQflgb8M9O3o5U9ODx21q1yeY1ol7pI7Mqp2FwBS2rqRtrmAqe1gZRt5giPa
9v6qNl7z1azQekIP221cDr/UhQY+Y7l5Jw7l02BsZ79SgARn34Z3obOlMWQmcM/t
q8IA15AK76I1OZmUj8sSdMxoPve6fgrTUZA9JegN2lFYAJ9LmXQ129DRnJm8mRSM
U0urcQmXTNRx7nLY/SmRz/DUMJKvtPb1eJlWZlxIf/+PL2N8FUyu+JWmFzR0FFjg
jcZSw6TDi4JpuFknG2pTQyIHUJv1u4eVdR5bdF5mXj7qXZQOcwpJJzayAYJl4Xwf
ypJ6q9shPAsNLEdCygsgX/w9xBC9FHe6hCN+0Tl25rJPXeC4HcI5FCSgSfD0lrIo
ImFzMjJW0LOzEZjwHF4aS1H1I54jeMJlqZMgB5DdVDkFkhnUKj4sI3+pgcEfg/YA
XecjdkgK5xkwn5UzFUFDxOjSgzLHQYkn2p1Vj/p7dsTCNXPw/eHKwAGhxnMSXb8U
OnhhDTowiXkVxuRcbiZRi7EbSN63/Dd178BivZbPBFsDSdN0dZPCSZlbskuoFrhS
KDXdcG7bK0T9zCjI0z16oTm9NkEIw2icKsLpLp6FW/48xrgVVuDrQrs/J+/am9nw
yYSeRQMUBfkJmxuxVOQT9v4y7zvQ1CrWlHOZpUAl8NCoktZfenswyksre2PfDFps
5QZ0YtOWZlhMJs31g8N/sQ0t5kmfx23rJA4AvPb20rY0V2e7e7+Ye7kjsxldUWVl
BBLJ2yUoK7vXV2VSmrVxfcREmwAMs4GXuXeHh83HrRy/TMYHP4zpjTxKmqMk8Rmz
+rl6R9cjqjX7JttJEmg5W9nUw9aPy77gtpQcSRlDV7xRWvE1yPQeLLevlBW8MTVd
kaORFNQlcOta6HpiHaPPMEc/fHdp0173WKgrVFQqt26CsNVI7Te3dQsaVN6jFMIk
2qt8SJ63VLLbC0UcscqVAwd4uDJ85pNPCuB03pqp46RzWTrCpwMqMVKA1YgnkE0M
+yUky382+R2YBjH3fR3+45geFL/gDkJy+ZQp5k2FfQdHanLurtGx/kOkdHP4VtVG
3wD2dB+h58IMoH6vf1n/pBHHOGfZYHrFslf8K0sJyhrx4s+C6caa1vyA8oG6DTsm
BAGvILn03m3lKn3B9kFW4//Qcn+RXweWEJmJtY3IFhg=
`pragma protect end_protected

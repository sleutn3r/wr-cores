// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
CLjVutoUmaFIgakyUzIwKph37oKoYRHbFgQNJ7am2rx2qm1xjp8GNdQiHG1pqvzR
UAiv4gtJZPNhs9qgPRixnoFxD8DNtumESeGqjbnL0VoBTfED6o9Q72d/nQG7O1ez
2DwacFwRMFVNtmlLvI7hnTCTjumsh8yf+zYv+dhz7F4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7728)
Uj+Q1esGP/ylWjJyLgeN6dR7rLY2lQIi24Tbgirr98eZB6ifWg61uW14ayzEAZaB
cwPHB9V4bd5X0C8ZwliOnzdXaOkxFZlEa9VIOIF4KAzXShcv9uNLt9lILM+wlJJW
urNTIhFUlvcyxYD6Xt6oQGd/WJY9GecCWuF5BYkd0y+Y/sV5UyZvSQVtSxMZhcmd
XTg+mIOnEyjPxbQcWwTAIMdHKqblopYcSmbPn2SlzZmjpXW0bideMv+MbWWGh0p8
/r1lV4qHw57+J0vrWwl3v2lJ5U6IUEsUuKLN6GNXglz7D9ZEpPvQcNrK83Ff75Aw
WoeySXEhVIQ38CI+oqrMJj36I5OoGn9Yoepd3HyigA6XRGBpB52mhm5AWKn82jvM
3ZLmcPLsMbw5zuQT8JSZJ22DTdKxWD5FLm/Wop9hHAHRIuTTmHh1fj8DsWj8mNyF
C6DIll3LrI8kGIqOqjVmy7VK56iU9u8bHAlX2ZfCCqsoSu81zyGd5+WPZfTrQ6Sk
Uc4ialW92OQZJddP4fJsRdc8rMYJvK5Ny43dNHUtcpndkhOZlJ6Ouh5iG3JSGFD2
UVANofH4hy/X2tQygG/y9TN3nbjn2NPQda/p4eJ+SVTmXv+X41OXtwjYcY9fKYqd
hUsnxC+LeiaF+VyIebjUnLHLyVMHDVdwy8DhUig7zhJVQVfkZJS+fLj5d1U1KNd3
8DhTh6Y5OMr09tGv0igqTFIcvEplzyIlu+NBQsBFV5iKQKbx0MxUxNYnuUmlxlSf
cMarsdnCKyFeakXQqA3mvCROEMvJRBgZXAhnj2RnM2mTud5ye7nzEQvzKTWgpn0f
PE8Buq46OOYfvtElLvewSHoy9JkrqRLD8ibxfDyK1DfUxLB7UnoKa2fz79b//QM6
Zr5Rpcp576D7HD0MLnNNdJoZ6LE3Xt7LangPyx6d8yWj6cLcjYTYrcaur/dQXeij
4y7nnC2Z9Vb6tsJymglwqFcrFas9YfGQjdFG8WU4yIwXJotVYHlLvLiFaX94cVE6
pm8dDURpxh/S3BTSUZQ1aOiPuoJV3+pZRcfGkGh09CCXn76naht+3U+ICXhHK9P7
yHoGEU9ZGZTpjuxl2Fj7n0aIqr8C+aLZWF/n+CbJzSgmAz+4XkfFXvtoC+wOBSSu
TAGYXwXXiFvU6s7ZQzYoENVmHL1lpUpN6GRNie0aNN4qiYJNwi/EIytuUR2MR0WA
bKSSRZb+5vGg9L2S4DC9VD7keIOvpUGitCBlvJYEfgScuUWR78pY9PYTFKBKvH7E
oLftMUe4a4xWJ8Wt5wkTSwAI+a2mpWS5Ijvy7GA19Fu06OsTLHxo9misTgOlJxsf
kpFKRdyDXTLCw7EKwrYx+95TRNrqEX0X8jhxNUFMlukGScFoVzrkbChM8UROvA6G
t/Wy0/WMoqo2cyYekjlbbR4VyqtD2FC/f8ZEmlQByz5oqEMJs6Cn0BfwVf6WXwEy
Ok5ojSA1sWpxW/adiaUhsclg8b3zTJeWEHcC68FUgC2iGBeBuHwGgMgcVn2UnKy4
rVV3dBPmD4SSGDo1PjgjcvPX3Dm7ID7B5LQPGe5jvyYNQwZivMoKVtTbn5C25BAP
YKMzzZ3U2MBsH9s8oWQOB9CDDh/OH+WHlA9lBZbBSs1hCx/QbuiHPA4okdU4ccc6
5iGecQF538d2IarQxXsm1x6uDgbAttAUr/jlQOE6rWi083QPqtoLMYy0WSLnh2Es
Bfxyidu4peNUNa1AmrGmAl32GZfBK9CU27Ybyc2RfavdnhJ7TQGBCWwrSAf3f/0x
rZ7EG10Uhi7A5eQ+FHkFFWzTtUkw9poeQO71fXW3P9Xv5AnWW042vKvzGtf9DyJy
qR2KRSrNLydFPOscmFdm2hFWDBNaXW/4ByswZAW7W4zitZoxpeS0/nzcOEIYrMUI
D49M7vCV6m5hvQNeDXYipix4AELuav/EGfzaf8Q4cpW5TnbfofLphzw2Eq2PegyT
2iQY4fS55wFUDrX8J+C/sufG0dpXfPq+A5cjE56JrxuLpIAcKSO0vvbsJVTMJWkB
Q3ssZQVyliOwUIiV4v0Dy2xRJL/AdAngEgfZRaFt60/suGmAK4STKEiDteSjFgfi
Z4YwTqs2ZyJ15CRiHtOmpXy5XTi7jS5gDLM1469jdj4ibDpCohqK6CEwAaskn41q
blr8NanEUupBwD9Dr/AtGaSWPKuIGzot9ClCoD68fw/YYkE3oRnqFUZOlgLPn2xU
v8zRxmXJnq3C/Bwx/hZAyG+y65y0my0ERp/gu3jmGsmuJKTHRArKJigZSDa/SeKa
z3E2gEG9iu2Dk764D57g7jQy6d4WZh60PPTgmQ71J4h3mLq5l5kCpIJRmfWJhfWv
Q+vKFHGA4wKJd97PIoDh5wcdy7n8rWio46GZvNDAWdLwKB4azp4rHLZJu0HwYMtp
+9rAQMCcLuCZuvMXIPhDLrrTGg8zxOLBQOlX5C7K2rCsn9ePJNcUPKXEXb4UopHL
heNmsMaAV5+VWrl285insg9IpQ4Gb7B4LzoPIIFRvSQr+5dV/msOBbwdVEl3lZSZ
VumOmX9t5QLtqr9gCpWkrIBCpUZHex2fFP21/yNVT828oVcYirHIznGM2zOx3rTH
WGS5CWXnaxSEyYk6Sg/FWZhpkYwjw9FVSzDWT127Q1XI3JGFdOII6UgR9UigrQn1
9ib0qr2gaJVicdJ+h+iauyPWsdjIo/OueZL4hQnLFsvNJS6eLrEd0dYElSR7QeCI
FI+HeIlqm2so3XCy7vdb5X9l9lvchTO5ndX+e8rYZpMEU0+kr83JQ/F8yr0qVkO5
4xLsc5BwriDE7+yH1TK+mAcV6sebvALvTn+O5nIykEgZbYt5GVnizj+OK4WHRO5n
tMFemhz1PKEyIK7bO/75xnE5y5+xkh4cTYoglgAVUojljXV6ifSnaWNVf53CPRPK
ObgZO2VIMqxgYtjf7HVfcwtC59SVdwaSsMydXnsT6acchX/xIbMBYSOVb+HiexNS
XvbkYHwSSCzS38YT4bIMWTTQNHCvHFZNJVerqy3m6y8dCzkT3/dJ9CwP1CVJMueK
lAvk06H40zSIxgI+tZHooFErPcjHx7Q6cT2PsOOjolWMp3vYHmi854+ZJgMc1lDJ
6CjyvrL7F/k47KQOOX1HAiCJWhN6oR6JNAO+3/2UtiNOhC7nt6YDoDyfrOiNBqHo
1oFbRdZJDUpVrEteagMvPFBE4tZUA+OS3XkEExnZ7vtLhcQ8A2KqCn26EiKwjWw6
TNPbCMdwtPe3gus69rdBOAvxTlVNo610hkpH1RM650trnrNYQQ960wozIwh/tE2S
CtiSXdnrnZaR+COqO3oPcHtEmLgelcfkPvp5sZ8Ntd3gS15DjmheHO2TKTm94jNi
9Pmq5Ckoy5c97aOTFjzcgVBobVMf2uoge8eNC+CLsLDJejGXCkEnzIOqXP5UNnzm
J4xqS5YDVvCUseGXjEfRniuCkF6eKW1DH3ZpdoGkGF8bYDSMrSTkRpqhQcCin3tU
JH9oPiiyll54KBOntDIAgkjgTc1CK7hxMGc1T94jRHcblBmeyFrn+1HeqefK5PS3
Y11txI8OugvWuqb5ZtEgsUNkkVNjFKqhox8eESSeOFEv8EiXBrhfiYG0qMwwzPxg
5jfLx2Fyyy6AKHvW9MiMv2YPbvnwRnucENiznXnjbEPwR+wPG05fjqZXOIfzMAMo
dofAWY1PEeRejR/gDXbUzHkr3Iw0/1KZqMHYCaD0OsupQszvktzETYv3jQvK4U5f
uFs0AsqZDe2Z2B26jorfgNAxRF0qDlUQmgPYvxeZOUTo/Xg7xc+vsoRplHU3lks9
f+5CZHBub2GBmjLc4s7K9+JIgBJ5Vozz2UZf0YxsJfIdjVLhDMyjke2u2/R6Da+c
Q1+uvBCVlRqPbL5/fy3Xw/aeyTBNRPTN37/vlOrWJBMdXWrykeHeGyoEQz07Ajtw
++eae7EOLbGad3g+XT4D0CYp1icMyGBRZdjuz4fUx0meGukZQXk7k/tN3UaOICSW
hEMvC4qe3bB7MVp7B5Fpzm2Ejms8BpFpY79Ixl0mqhWSxT9C3QjOOuxFGHe+a12S
KG0+OEa9Pmjq7xpwRW6bkaqZ+airo9jfkm3xdIDojOxdCiI9Ucv2B/1dw4mfByAc
e9RoBQ+BOBcvFyDmi7HyJlSpE43Rhe6nS7AbZ2ehwp3jzmV8tx12BLLKe4DRrCpV
TUOqW1J4Y0haNqBBbnLDfa5Xc1Twr0MsdrplZKFgLbJnL0OKd8Yb/0jL2MYlTXL7
3i9A3AxXVWt9Z38+J5woBwfywK5dwsECJyg67cRecv7uW96qsEMt9bvUCFkp4nrR
6I/llp0rHU3kLo7mdbemkKqUMlfl4taxtSysR/I34jZImhUs+mN7Y73h1DUFFJXy
2fpsv5zqNRQ3bVvAwj7pNrvflrQ9cwKQvc5SL1JjM0IrNQvkh71NN1dKPmRQCNwz
FebPAd2fqKnOUfD3EcsZGi+He29jo7wv1+0rmRlRutS1/RkZdULgxckw4karfNv/
DgE5u+RAM9RLXmHJEUS0UpsvAVtEnzb9IaoAuny2UHJc5OLC/tqZnO7a5/6S+SIp
cT4f5PwFFD+DmxMHST0Rtkng8Lr3v9zNomDfqM2Jt6mEEp/5o/nairkiBQ5LGgnS
PpoOuthviQfIxgYE+hxWMnv5hJb7eWwuspzWKQge5apPwkukcW/RE30MYzFrMIIb
AxMLlyIrhHrqv8JKdwTGk5nPQC+f6ZZ9LpPJ9mxBgdLy4HzUhYjyo0bSduGMfC8v
IZRqNlKQtrSZ8bxbUEXkh6lh4bQbNfMxrrCq7OP/hhajNwhAEgr5NjKqWkYGkgtO
Uw30iGbiO2hjBu8l8jpam1MjmH0+R88m8CTpFhz04byoY5XBEyAqv6t5XaTX5Rsz
KfSS6lHFH7KKWam8p6zjtFsDLma3H+0EB0NCCv0VEL5ul/EF3FHKonuIcEIkp8CC
mgoRs1JMyXL/63mPh7i0xfet3070WTfeQHaBxNhDPb2yDVaI7jY+GLx2/M2yU116
DZAt9dp6qnlRINzqlrnUdfMgPRRX53+c572AWJ+m+ARlIZNNjnCrjsyDeIO2k3qU
olxAwRm8n0UACp19aLahZMX8AmfGTICw3mNPWX91ttxA3mWTleyCUFlv8lkRIll9
1c9MZuN9g8k5UvLT4v2dndmudnMdQjCjFjd9FU5v/VAzYZQGC7kbXEeWUAys6cK2
swYCdUnM2WxwRpaqd1BaEcebfpgvGSGbuKhMOvqdI6+4XfTgJOHXjINbcImy39So
1Wa0iCRk2Mi7/j7h0BXPlpVUZxfR7UyxhXnyscxvL52SKl2NVQ7DbUq4r9iJGYR0
GND316ynyN1Dq4hThnOP9B6AjiilLqfoDexY5K81xzeOJF7WvfyKZKoxCr1dpb7B
dZSAxyr0RVfu2ggkq20F6ChcjYvJmLPewqtuN5Mg1og32VXObnlFnLcIpGzVUYLG
7nwcu1qZsX6hjXOCpeURBtGt49TauE9RYYU9fqFnFtrQn734ypObeVWcWpoSGXy3
RXqtWxyj9sDfn4lsqoSUgT8ogw8vj2DDQrDChbvenLEXIoIrs+Fz8RKeyvtvtWSp
3vf/OsEWoaw4V9Ito1z3qppL/Vwi7kc3TU/fy4uqCBIv2Vvcz5RzVqZFwKnv39zY
FUZZgkr7l8CvAPFeq6QsdnlrXAWC14aLQZCTwAlmQLDFKhDuR5cNMhKpU68AxF5S
BA+0ombcL2tK/JmNnndx826hL0PhALVwHKiuxy9a8mt6YFBh17guIYnNKrr8F21a
FxU01HJx+NYCR2WNQflU+FwRoswhrXf5vXfEZ0bSg3uZlihBMS3fW79h+EUjgyVh
/m2PRZnDywcZCxu5MXO76h9ZqdwRsyCvndxNk+AxKZH9Lszdr6XWdB31+t7VLkyE
5MiJaX1+OwS0PHft2HoKr3sBh1UJ4Ft9/db4WwNG5HTwhbtDbwSjiVSY88wUw5Cg
1lzvcsX9L3ALdIpf8U6yxUaBHLtKn3bYKPtNCEE1+xWdHqJFtWcm0m3KtbPDoeSs
zIM9e0vJ43L/ROt8NMuVJzVeevvd2jylqjaT7CdPA0Kca78bhPE+VVA/oKtM+2Gm
Bgc8JC3EvRbK8+YEkaB3wKic0XGL5JLh05LoDQPhvoZozSRHQrCk7uHJTm95Y8rM
jfNZ70YQXgygmTfGr9VmCAkt+fpLD/vib+kvGpFLUMWKJNzPlaOY7ftFWf9t49xu
DexxogOLqaEWnTnbTAz1cAF/07V4Ki4YO0kubz5IXy/ctBR8sxYz8zI/5+eZuSmV
2QEgV8JimL1DWlCspZR4UWo5J+hznS/48Nwldoe2iJfxpwk233WxNc6MPDUmJP5Q
3/mzM3kAyP8qdneGrA6eTPSruvTGxWU+ucFuyFDqJztUg6dxK+S9j/YuP2e4JSfU
s94o0cocAPj9k5LiV/aIF//ltYak1z90+MY1tEdMrxioV05V1D1gd6QCJEa3JWBQ
XuGnnj80calcXoARLFYoyY358TjuvpR6HJ9KviOOAi0kMfKIShqMJInp+cqSnWxD
1y5R09/JjkEgOleWIfChLyTuZuJ4W2Lb+zYfjI7HEv8YTRntYX9NFtwHR/bGRU9Z
5BsXsQNSlrH4gnGNUGCsJ3XiZ6kNvcqFyE80OTYHJsuRNFxsVNDK1ZDm+wLKS2df
Mmi/zntV2yBq1f0zux4NvF3UkOMEuRL9Oxph1NuY9nOzqxH65whodnrMMqRjJF2B
korpbb0jjQs/K6JhbnP+vBGo8BnIUX/8eqDaEfwVeZmefA4XtWmI5CSWgO/IqleK
99mfqO1s5dNPABkPYl9AIB0iofNKmq5DGDp4r+PFjgZHHuB93GGNZwO1wZsyKBWk
INm1kf903FIiDLwe7f0vOlpI/ytErQox91VxpQwkGmCmeYDWOKieEOewMjIl0oit
0h0MfEJ7UDb/+wguTBHy7Ewr7rBsezd0oPdlK8yqQnLx6SIPiEzzsmdhPDOa355s
jra7+9iT5J7dyM1bEHHxF7MBXl8bpoHXe3pIMyfT8k/bZQvufI/xMZTMBI3rpobd
ywXCnZSnm13ge7/xfnAnjm2hMwu2w40RbH/rLZNXtZVkfPM4kbZUjUySCnkqcGu5
QbECwnq9X5OOuxrtrcdHR5P7MjM31s2SAFzHlQplPBYi531o3Uly0Qkmd5+FFJqn
lXag7PzeFcSzJqdpM7/GYRMfdv0WLlkXk2O3ZazI8xqt0jIG+qgMrYEf4nvYlear
BwhAQxM8Rfiek+Ze2KxpvzWyiSkLwRck+G6ov6ugSIV1t5H1zOtb1+/esUjlXHvQ
H+8kyYZT231krq4qvOSjoYvX9PvLoJrQxdVeuWXT5ZjrhT+mV13MViN26Y05R8qM
f6ccG+YVLgV9+4zX2kc0HC1JLrS9efw/95zrjXjPbRNt8kyZPiX8+ybb0il13u1u
6ag8nyuaLSOWyQq5iPXEb/MwrvMjc0EZfu9ycsq70rG0TgVZMdZKo8O2bsbgoEap
Pm3Jk+cqSwoAu/HmRFVKZXsAymRFw0hL64AsSj8pv2jPu8JMUDC2weXD37wVQMDv
xIwqrzMzKXEOJD60/ZHh3uIAikYeE87xYWCJDx3UQv4FYWndFqs+MpVjFkBwdd3E
C3aqQRKTX9Bz6JdQAmfOhFBadFfFDJfwsvZr/MIqbKBC1rXpUM/A0LYoR2WyxKcI
1LhyzjZVgtoeK/l5MNyA3X7XkD4Nsvr8iQvVlqRCBa5yxMd9WGLcERuWxNnlOIlW
CW1lT9jFmFUa8OYzBnC0R5Ws5d4jDKQd4/d8d/irtdZUlBA4Y/PL4riMGVFqmRag
q7T9CM+K0QQwkCy+V8YOJhn6kqqnqWS26GfkAvZI22mk0KBexSMXUta4wQX4qcE0
O6PLqu4KxSOMvx4+Uh3uQc/u2rfJ3PKKQRxAvYrxqola8btqiEQ7fKgXfo8NJN0B
AiqP5X/AVNKX37D/cD1iR3Gw0GHwOFpqfUPFFgQ9e9c+c0LaPjvdgkwi5rXt1qVl
f6a3aRrkPR2osdzftYl0LbSCkTFnGa/zCqHZ2PECM+Sz8pY6D7APPeKCqPRTht2C
sucvqBsrBT9tc6IZ27GFiE0iMRzr3fn4sBTd04quFqhrcIkR9SO7joC1QiNIIYop
3olulJ9DRQAiT899ehFvFEGhJ9+6k7lqFIWiQmh8XH7OS9L+YqNYGj03vTLPyD6J
fERcHmhuTBLzf9jm+n5FKjaiUuxR1NLEr6kmr86YbyLBPAy1FuTmsNiVLrIwX6Gh
BB+7H5xZPaQ9ajXCFpc4n0r/pO5TkI6fwUIAl5usGCJdPVY6T+ssNnnQUOW5YFZO
7vTobhHdUeM1REfy2n/gGX00bKQeNCEMIn+ehmnCxs7hRSX3WUJYmG4q/wgJ9nYW
n6Rg0V5Y15zwdlJaTOcEicHGZvvv9C3XgyJWlgAV9XGaw7He1+qWxiKxhb+cLbdf
flkAJrqUCAlYib0Y8qIhvb3CWtLrgxl9CSG3rpiKZaKoIdkk1ymRIcPF8x7M2Rd0
HEWaB++Fgg+OoCa2GnaUwhtfODkbvg3bIUJm7VKlfRCiJkRM/NkJSfKR6kKYW6+E
fAr1NOK3BE1Zgzi/V3A80v0+5AARyxxVDchqEnDcMldL7fVGaIa2fIVkmhTXqnPn
pY2OlaZKOutFdT3+aRaMbVfM7RH+ATmhPaQnoNJxcSryVETj3+UkdY2Y2KrEsVoO
68u5Cd7eu4MAaQ8n4ft+OHXvYILAbrtfCsNmyuwsWDnlq/DFbR07vKMlR5t1PQS3
Q/KHWF+lFSc5K8RLi1fUPgflw6YlHr3x32j40DIngqFf5S9VnE5ZCln6HD4WaKVV
2amsw76uvLPYJoZE2l4EsfMsnwSmlsb3tBfHcHo0jTbYJuef8DRU3pgaCLlGD95k
pdk3rI9gLQq8KCIg1pi0mORbVmFmvszyDi/6mcNxGCxxiFx/ZY1ywwZ9SKPDCQo4
pYPcSfkiKi1MuAdCWyifroZpnMTg30AifltJqGL2lWpzQ169KNqgr9bgeHAEOKTN
CLOZhoUaJ5gUfwIh6b5pEss1ZCCwBK+HqsHPXp25cJknP491vMyDsKvjs2g/Zcny
MFLBdVHUSy4Vno8ySQojgcYIwD/P3emxzJN1UynIBs3rP3ilnggcXMYzpmQ/wKiR
hTjuVm2tBAl+/vSXoQhZ2m43it9+kOYeTzOlCP1X246dn7fQcdptT/CfoauQOlIX
k6+VZWhDLDgGNYzv9PbcGE3eeT0a/3b6YSdxES2wDCbkL+UWQp6Hn0DveH/esT04
cOdSlmVOz7xNPyY47SpnGfjhPtsdBVEOkqTmqepCiT9ynhId8Rg7toXW13taXEFI
Uwidbq+XWZwkawJ5O9Vwhm34tiTUUNajQmsBSA05bMEu1sbNShPOGhaI0B0bWtLa
G5ywNT4/y9b7yEcMwTFHyaiPZKrqshDJbA+1Dkt6H51jCa3ulOQowCE9y3D4Rut3
2/iWKl6PuEj50PqL46laVVH1KaE1xt6rM2/LOKMGNQN8jX5//UP3LIcYO7Cbprt8
DW/abloReshjataZL4+P67Q9WCCbOIVDxI3Suva52VL4tMXjA2uzmzicosWQpv0v
YMXWpb02N9zc+GWNL+g4TT+8g58kKtMOcaCWTy93DE1Y4k1B5l4O9aV4AjUtERJ1
EtMQ5MMEMMynVwSc6VztVxJdP45+0/7YUWhdxix9OLyRtfRNV5x0JmKpnAuvZOMi
EEneLLYl5K1HvGKhcgwe/KUbyOml9voHJubH1srBi7Mk+YMleibblpyAFGFrX4qU
R7MMxSLQgCA1Xv4Q4AuoNYEV6Ev78hDBe6HdqCk0pd4vciwBUshDiZKG8NIxnsdB
KjyLYdK+TiyztoUOsTiOCsY3uplNoyfp3cyl5H2G9IN9EFDhmyKoe06gmd/xuNcW
UKpSe3qGrNP//zF+a3nnA53R99fr3gcIqKqEtPYlVjZ/n7326Us9p7B305NENyf5
BhCuaK+A6tts3YhZElXNmgW+1bG99wVEKcQxMiDk3hIRTX+kQ5jsVBqtiv2sQ51U
AfM/cQ3b9zFinC6vuWzG4NnwCUtB9+kqH5nhENwhZtWIV4Xfxrm6ZwbhDpsYjz/B
Qx8sbZCp/KBiFKGs0IHqZAZWcteXfoQ9Mxy6D/xEti2dwSlDEk0i5qfTwAVYJaVO
wuKrThDvsG+Pk7NgNUp7NrTrkCA7e07WQvERTwCDo7HR2ZYaSxeKm9F4WpXsInSy
`pragma protect end_protected

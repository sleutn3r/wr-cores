// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:45 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
N0WXO1XmQQUSAzddN6oapDbE7RBXUvieQ4v5fq7/Fcyo/K6h/dSnGa0aOC29OrrU
+AFq4W6xLSUA0pEd5EgwCVzyWHyMKfVDm9Y7O5QKqtmFa5NEmr/dErCUg9/cq5VV
3Qa2wxCQN87k92FRJYE37cCTrpiCvVVG8bIvm8Pd6GQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
3BZzUEuIwE/MFHbMuYYbyPqJK/511reCaFbMSHEnHLPNF8DaWu6a6aK1C0RqmkvB
FzFg9XCMdeKZwXjp4W41kBcBC8dYVQKWmWzmAg+1h7VnFzyG2Q7KZaxDcxvntgcN
56R1Xn3s8571RnRRnGLRZb4n2BUacAb363PJ+hZ5/Mb0jGkWYhusO5RR/5Yaa4bs
Y9djru894Keo1n4pDL0MxVmJFXTQ8kErfiPO4+Y8Jv+EkpMPbujnw9HdXPPNW22a
ozup3uEVHxdI0FJy7Qtl4N9DCZE0wFufa3PqrCKFHNrQ1vFzuIYK9d35nHfSt9I/
bha39zDgV1sQwEl1LdPmO1FU9y+uiVVBWVCtA36KYWVUBI9wrb7mxG3UBSnrfZFo
p46cfKDA/iCX2zMxaipPpSE5XT3hZwF9gOp+eMZnJVE6Vyjto7ibgh8kIvGVLJmr
4i8SR6ZoguHSGzhvjoTHz4ouGlcyRIMMAYzq+6rTQl2rECSpkTCb8h2l1dVVweLr
YWdjeOcoFuS8tv/H/oLT88LEbnjLA6PmM2O702ZtpGKs2pq7DRtaO2T8oxnHxLXP
VlE4rnE19qzR3Et9QPQ7cXBhox/w2uvUiCtZer/Xi7mchkGUGhDgqLUDGb2AXp/C
zswuW2qKE4aDMpRvIuMlY6oH/U/07PPY6jksydkA6vYVHFbnSk5ska6gUj8QydLp
ieCmhYGJgwswUycEu1+qDgZKBhtPFx9uj9O8RAYoM15k4gnBp2wRIl5tCahfRLrh
CpwWnGss63JIaSwn4TBc9hhFT79MwiN171nTiAW6QfSwf3OmwJE/wYkwIUbgl8gd
DAQv0n6pgz6DSFhVnWzYwECkgbOyKRoVGOIFmLZsqi8hkE5NonINRiOQubPs3HGq
2FUmFeh9bZw8STcL6bkUGBg0Fv0JFly0f7kJkxlw5pjcpkunGZkpvmKd1pjSdchD
Qq0gdf8f6SiylIN8hG0637ke/zJXey8jtUGizxwjOVXdWxEg8AjOhp+L+qOtGJDi
qKmFvt+LHhp/C8hPEVfcmgu8WD/upGCGNDZEfiad22BMQ0SdHr1PY43h55KnMzkh
Zq6OyoftH7veisPLBe/cANsxKahQLjcTXXQd5sYy2K+RU6vb9nN6Dl5/vDn0qvwk
WkewH6sVzlv0Y04rpM8+Px8PrUo6xtmvjNntfY4UNMIH3TNrwF7H+Y4a/Riv77MT
73eXh1CHKrEKxL7lEO1Fa6eQJTz81Hug+jhs58jg0lKcuKRspVSCf7YzuaWHAIXQ
N1On3T8bkL0/jYH1l4qIO6pER2TDVzLzPZNkOMnGnQKjpsJPODhqp8tZFZh/uzdO
psEJuvblwazR/tR0BOg2Sx+hr0M/D7NqPPKYhfhl6CAE0tmv4/uA7AJrSuv1cGia
7ecdwxtlrJ2rx2YHNqkegzCnudAeSx7IxXl1nEfpJd0cPz+2ZXXb+uhnso0jK7Ls
z3wVn5CuTxuYKsKxMqmSJzYgz1eqH6/HFE2RlQ7SQfblnMtnnYQzanFzhGp0j+6b
elingKdPiVEN4lWHAS1/M/A3CVGnPLN0mh4hanl/AAoCjh6RKuEO9GAekChgi0rz
89sRMURmCmxhYUYUEzpc4KqE1oJHNP7Sqnw43AJLEtBZfUsNvYxrEcZS+GslQG6n
BT2ZQpM4K5249uEHSFN7puBNSeB/MoG2E0oO3lN9FlWlMu6C/QY4SM7M6JfB2qN5
mafPXHaxhfBZB6CspZITZ+DWah74r031fiOZSUQ+47Wjf15eRxA0kNlacLqCmWma
++QVZEsPD+nAO67D4OczrErE1LoalBhV8FZGXUlch8IqidYuRpV3xobOaUUV148T
/HIvUtWbvKNeMVtx7tAhJD4GPnCYw0ang6P20uISIDyLX0hMZEECAGoDjTMz0ORv
7nk3KGHqPxSw5Abry9AQYimQd+8tCeYTLC2zqo/Ch9Cf4sat2kZvNXtWFjjb3KdW
u21I1J7PHB1p6PtUI3SB/K+orDe0KEd7ixRDivgWrsHgk4vVp5G3scpAE3hiUxrl
02AC78bFwXrdCJtwU/S/p0m9G3fJK7Z6LpQ12BKj3jMlFGA/zMQutybLDWK0bpML
ulagLXdP4ajgvGy6FjAGi0uSs2/2l9TkH9xva3Paj7gyqmvXdkwIi/XSx6Zru9Pu
nSiXEN5RBKoCllXP53vbzx3kjUGy2wAW0mDuBH2Efd7WfbdNx4t8Y5qej2eEfTGo
yAsOlTYl3Cbo5GSkxNn7fTvX4rLE6zzR+saD58r05hLSvNhA2HDA3svxYjQOFF3r
FxZ9GZx4WEHxiufGdjK3uQ/dVo+eoLYsSKwKktVVNFvg/u1dsuTMWvVa4fOPUMB/
rjcZIiEZthzXHHcXamkTt/jf5A60oNOEAiR1Fs7TZfz5BXLknjy17rTqjz3v2ECG
pXxFeO+D1a6N99i1R7RROJg8SV2Mds8xpNWvvv+PXqZC1Lo25YGddZaacT8SSBIr
2wpZ0O4UdeSTJqYTRNKmc2nTkLRjw2aq53co4SFX19ULwddqWmwTZlZt15uotyH/
NPE6q9IXUzLT0VL6pJMJa80coLXxbFM4DQdo0wgWI7pj4yNFPswjUXptrBs+PdrO
iigOXBV08OXqk0fG1fsg8+PkYQaT2cr/3xvko3d337t5uG3v9Lph2WY0g6WIb7Qr
eqbGILAE8HeD4dOp7afPQW0YjDeXX5VPcy5LwBekZxerQagsdpQBOFz2AigtnmuH
UXAjluWCrIEc6aEW+anTOpr652ZNI7ocyQCbRXJMSy02q5Vc2DGoVM3qbZ39owAj
RyiCBO3h3oPWucuW6zQldKBDPGrCwr74tmEtwSMDJcNJBkOQ3vyn5m4Kef/z/8UD
Ek1U94F3N6NFDEmgAZ5ThDo3epsD/3YAXhnO8NIfym2+iotR96a6aCpMzAnv2C7a
3ko5yzq9Az+6zK8b9FhHdWeB1W5O4KQZ6FnzWH7hTHg2feYJxj21QQDjiZxwpZSS
28tSJWs5cya8ztRjce/Ml/SlznVFrPoSKOnfQ0LaZx7/GrYHQNl+gvxu/p8JAJxd
XGgZcTzzZnOqmSNhYTSTzvDvR9py22WfQT9YGW1eG1ROsfn1unicUyqoth8IwANj
gFqC4nBK9qPm1wEDJMf06pc7q712UsJ65uwLN0+JFukSLUmBVv/ZcqZIxY7UBeVl
LhOes1muQCn8/kwD0V24yuknLeEUcMfVI04OaXPS1QDnQy3+3QstwLmChSazVAR1
9tFozfQyhRn2Dhnv/8ORTIOgmkC0Vb+JWZ4kAXBz2kxkkPF6q6DDXtVjL/xokKQL
HeMsJ/JMBsmrKWaZiFK7k1/mOkiugOR7yFrdE475qI431H+jXyX6fKJRCsfi2NxC
VHfCDsS4oWk9+eNFhPsNDKrkNA9wqZp3KTCw7uiOYW6a0/RtT3yJ+02ngTpEwQmQ
KODHC7gTvf9dJBV4JwtjguqLLBAyRnK1G87sO21LdN+I2E16pgK20xnJZ1ZpPDBI
xZxM4crhiLjhswQ0jqn3WqaSaMP6bFZ/AERFqr43F53cngik8RJDZwOxmYUm1NkI
MRoc3NU8AArAykEG45Fn5XICehifLJbvdibIWP9FIDy/fF1FyfivnNjTF6alEPtE
JPzDragIPmDYJ7mFDEHO17h6KyFL7yDAdHw7HnCeOThgziYCeMddZ4ShNb1/GaQ5
pftfZ92ycXD3VUM6ZUklmkFVW76ciDWREZSp/37QluI2UcP/YGDm2rUeqU8kVS42
m9SQlAuu9tvVNyCKiWWV8Y4azXqKYqq1zSMlaHEaYFtLOaaQIcai/u2a5nvoqbVw
x+deqslRD9tmwQFEc0eNYLF6No+8z8+3P7Prcrd6+hxGuPVznI4NgE6GQLGOe/Xd
mjnb73QeV1nV0NskSClp4eDKuCpTvMxDLV4oxqrqEVebuwc+apvDst+2o4lArmiJ
BSKSiQF92XbFJGf3XnOVMNsPFAuRzo9PdeZ5CytZ/awLX+ldWTMguuAZo6CLsC44
PLu/fRAVGOrvQXIcMQsIUPDTGZ9Hhlv2Hl+YhfsOqJQcbynWosKdGDKamMC7HLhx
H+Si9s1C1OmQgyy9LUE6ZShw+mL8AC2HADOGOMa1DOtNk0inJZTr+tCTDxt2K/FC
Gp3eSqhlgShz+KSpZFHcDORUs+LaYmhTb8sNu9aJq2v35KDHv71sAAHJcYeUUp3Z
JoRP5G7t/WcccsBCu5pkNiC8atuyDsrrgpzMowPSy1MUaB/bPP95RGUCB47V/ZMY
RsTDD32rFpyvNBhAt7Kq38z3tMC5rEPOE9rrp46VNeba5Hc7mFQDmc4ymmbq6Z4M
qctOJ8NkKEHUfFELbZYMM2RA96IpXl03mWTYLw5CcV9rdvChoEuixCzOQNvKDyKF
WiVduo1jNyCfkB9dFN/4IY0Gpw9qDPSHT8rOHqcFLDs4gH1EpTayR9sbe/aYLbq3
IgbWHgMDgxBxM/ytMoBVUHmNj4j8mOyfDHbmQP17InmgkenTmBIZplcSgVSoxwuP
vEZHprlRy+meovPAJeTq/xX2DbTn5nIlT7UlYVU49+7mXnV4WCiPfbMudgQitf6u
z7Hj5UPjjcFEH39p0prSU5DUHe2VWuipbvLcX0vElfgnkWKbCnSPkxkgOs473FMe
Ns3elIkAu/YX4lErHOXWSqQ0ZPJGx5ceJrUyjT4z+1kaqqrEZl4i/xFdedDWynZW
JIpDjiTyvapa7xJnFItwY23iL2UsyT5yOVfgZtCwMJ82GLET+UMeuEz560AGFN1p
4gqdw1AX3SKVEkcQPebesIw/ueo6Io9C28Q7zVyihCClSt9dyp5b3A5zUn16NjiR
ZwaXIlVvY3aFe4DXNuaIixyDlR2pXuc5DJupTzfTI+ftYSfacG0Bn9CE4hqk/r1c
QwzAKVwLmBiJF9Wn5PU+h+IAI+msMhqEAHn5Jyzg8JgCh4MijvDUTHpYyRhv8Kts
N3PtNDbTXGpAct61bJzwPwpNhfIwIpfJfvo4GI0VioIxTBoIGGKHAJ2oQvc2//XC
CI31veuDtIv7X+GoQbWyvFdorXJ6eCRjUNbufJ1/igc5FJZ1hMlewR2w6qbV9Wj9
MjTBYEjrESg/hhBesWWfRGji7/Gv7VzwG4jgMcGjtzrWeLJWE3+kSDdxoEgtVpOd
+u4XIA62J7poIUBgDOZTrtUfKni7tcUKwenWI1i105Qd4l2sbMwhQ7RIQ/ltcTE0
o4nbJB8O66cP0ZLUzpiKwYEGvKxPnwBevd7oU8P+Liw++eYu+O7l6Y8VFtW6jeHn
bJZBS8cyPUZaSvp92UYEweHoLkATyANKg/VBjgS1FTNS57DFEiqJatlcYrTzHKUA
cyLmo15bQq1mB1swAut3gr1Ypue04Ii/p0IxHMAb88tuJjtWPa8ja99BTdo5otHE
pK1I3igcHnzBcrHnyeKgEwsUHby4ufUcwUxQ15phgLtHr2ElwzP2Y9umtBKAvSaw
NNOG58NzpC9MJw3R6B1DYFRQqZ5JcgvvVekAjXPB8zpmKHG0gNjzZ2XOskHoaNzd
memPOTu6+f+jMSL8qS4WFgy+JgZq6lCyDVHEVcxtzo7REpWaZILURXL5eIUci5VB
VXbs4Qox5byw/ewOmScbBT1tyW0WGlycoBUbdMMtmjn+Hf5oCybsyrCxpbBXkeXr
fA4fbKIhCa9SZJdyZjB0bQbQot3PEvcFPlZo1ui8kAWw3/Gytix8uZwP1re34ldW
2ENnV+gVo/Koq5jyf7D8CNL4DKlJYi0YmPU0BAb/w+m/uSCKw1O7nejo73h804Wd
NzlqnGY4MvaL06MMlgAdaTG7dPpr/i4SuYTn0/a5tIja75UBdXl9br7a0hBYqZiy
GYizzY4Hgirvl5G/jA4qZYZ4lbPUdSHClP2+C04T3piv9molRQonEzYxBipq1thz
h0geWt/ut6PfqOlnLrFQf8+mOncyzbC4ak79sNB91eVagb8TFilIq9FKqKw77fu5
QoinvH1z1Tj5vLVv9/hh8FXYWw1NGHvUEUHY7fPh5Pc2IBKKmAF3qyDWrl42t0cW
GMNkRNVRW9rDGWc+e9uLlRxYF3i66hrFYf+q3w049CsZoW2CckKcjBGFhN9+r6R6
LA5su6raTysnX8/BBGZMDKnPWnUBL2vuwdqPDYouPpIDnYhvsk9q+/v50jwLpEL7
vKnfsnnsM718aBoluUEUVRY5RBBZiN8ZKzbCajrSw807ErdtDEFWUKm9OoBz1hXI
hW7wBipt3RVPocxClIYDRj+FUft2jkr+DHlI8aAQF56mLqHsumJmp3+0mr5Bvr/X
18LnAwpBuhYHCBIwwNVnU+FsDlaeNMQ5jdpjviTKATd7++zOzsGKckmsidEJFPJ+
5GMLZszu7ywFooiiIFjtqwhUEEtnUIlEYshDopIxfJ7EMttDGUziicS7YA+grbVX
GOts13ETSv+YtRc2wYByZ11KsPWORoTjWc/E7N3gOM12EE+lyvqZAWLfscDKtRft
47PwJuW0ndQamAfn4RoCd2zack4pcAXGIFVy/3ElZkl89I4r4oJwk3b205HOPAJg
TgRuCvcWUSHTYkBQ6L8FbCCZx5oKHaYabAUpZ/1CtcDNE83AIYCarMS0xe4MkCye
esJncK+ObR9fd9viOCTulqac+Hj0Aiz0RvZhQe9m8BiPILdu6J2Jqb/UIjvNBHE3
eUzk7Y5il1wuK6yC9oM9rf2C22x1zwZ7b8qoS3w7RwxPYoYTDxdzF4P+0HDeGwS2
r6JI/sZXUQ4plrPMv7VfVNOy0052lf9v6k5svdFhbm4T0VxncyFq1qNxq1iasOEz
AbBx3WHfxnW2aPFjIP7MTcbRCYgEw1tyE5Puf1NxiuOwUXGn3N3NOUdwmEfaBWVT
0ykHB6qhpzU01Rzxo9JzW8yvQeMt3e9RSqMTMkA42ebzOnO1xah8nELBEwbvF/q4
8/nEPYKvHUY55kXyKwmSLgkFufgzk7arOPEBfVfoWsXcYLo30ZsOGLgvIy4MkGGA
h201QBC1RTtOrBrKqsxkgTky779p9GMqffwRBM6HDEuEvVlHwBxqDBnplHMi1K76
ZQ1PSwNK3u9iSwPFpExQWuUo6xzjzm3m8Hhet9DxzUo82GiF7IfagvDNqMkP4CJj
Nt+9hDEZBtQGJo5+NmX6kc/I66ZloLp8GfvHf5sMwWgoiioY8jI+0BMMaHrjs8Wx
Z9291k7H7heEx70nM7iaILHN+XLiLD1EAhaUw7Gmdpy1CGBUyPEEpAiGQR27OXgk
fpu72SuQeT1+G4VF9kXn9tyPoGsmwu9WatURJvWQPxyo8zpg+iUSGLvWIxBHCjLj
RDvN2rzKjLl1IslqsNnMXSV8vpbpx9LuO6s5t7RtXUZ88J/YfWuiIOtQy83XO2qZ
anTBw/6p+c05BvB4kLM/z+eu1XABgBWaA6qJOQesXDMKpziIUdy2kOTQIyW5Qj/u
8Hiwdd7fSICEmiqYhvMLH6kj1cO047X6LQr4GGMyNC2IbliB8Y+m8zPbmxiKpr92
`pragma protect end_protected

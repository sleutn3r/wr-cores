// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
i29jbfpmN78rOwqGYaqV1BeRgyp7F2OuWYMGgpCNh76FBLYSeCLpv43QjZAzWvN8
racoiv1FelkpMwKYQVoqwJC2ClYdU6piXUe+DTTCvbkJxJBIFu/KOPuxbi4qHH7z
gqCkE6UwNVePbYT5tQB+UiwAxJPe8P8zhhAe1zKVtu8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7536)
uM2wSHJMTYY6hYiwv5uROOnG5xNdh93DQx4OC02eLndSVzBtX//PNxVNtpfQYObZ
qGd1sjo39Eox8aDTLbL/3HuK+wlK/U6SK6070QdXnR9W1vC4PWtIsikUmRK/bXE2
zBFRtfSMRv8U1Ed4PVbPqY6YG9onDkwt05IreWKu0ibdIAMUpq1u9k1vZR+g+ouG
QAvv7BD42LCtEfbNjSXZBwFDXkDjZMnI0SzLPv07sa1WchnrQnMxVctBcxitxsZI
TbeJXH1nfJrYFMMav4wu99tQLhOlRw8Gz+WTB8RUTWxocq65D7zWzOkSybZb79jw
tVwLjI2VdP7A5cHadvIa3UJLZQjpkQ4nyfJjX04p/xZL23Ra6T1ruw4nL+qNmarO
Ff5yZ/FeFuOlmz8qWuRpMGYu7Ool9yyWe5CvDgFfHR5IXdMjN0jB/E59OyK5G4cG
emVbUvf4xNfnIwYkJTH30QPrRGYL9BVeBoquzU7cIRznwm+J/85sO+UdiJdBmAx9
0OMdQ+eAu1OMeuXOOvZ8PL4+NkuQ3et96dNyTWtIaC+mTXy0qPI65DipRFbx207Z
pO/zIef1M+EH19LN0QnS6p31zwf9qqcz/PoYQBJ//Ek9AWODojV0JNG3GyxYRolP
sGt97sNI4vpCW+cXwdo+00pf+K4nNrPNsy98YG34dmRULLB+vKRUsoA8YSC0hUQW
dm6Bq2yRGxzBlQQ1gy64Q7uQOG8thltY524qBk1kaOFBE072YDI1psqj2U5gVJCO
VCKscqZ9XCR9RMXPXHM1eXibD0/EDXFcdgN0ncyDkM67R33QG1xMIdd4znAob57Y
fiujFrloVSqf0uglUCMAW1WW/kugbbUxWtuWSI9tA1FYlsvH3cCooXXF7Xb4hU8K
RyubYgTo+r1uOZrve1FUktdJtygaXUXb3gMNamUe+3Fw5SrVRap5E7VYdg0BSpZW
6bW/AmOCyWaZDrqT5cjenE7Dx2H3L5r9h/0e1e+gi++6WlkZM+OmUdfZARu/zS9T
JjobmT2JsV9MiPOg0UKqavizzN21OxAe5LMo5if8k9Eda9eWWyFAn4teDgeSv8bC
jyqTwKUqkwJKEufArl548qstlW1WcKAyeSHB4Pb+PPmYasjyT7IWRiHwKvY68L+1
XHl3PbZxTWqGv1ejFvwH0icrgDhl1Z1/rTQGnWY3MLyWtPcBDKCN1ZcAbokaUrrJ
51P6soJFSrO5PqYaE8m9DOh70lSNC272Cx5AnayqYtllU26lblxEwxlHibSrajZt
A2CuFJ0UYU1rqzzVNs/SzeOF2u7cD7v8nKSLt6b3U6AHhPpCj8kdRgP0Rqw3YPgW
/eak8VPzvIckhc0icC4/l3A3ZC72TKem/OCKcRyZs+bW2zUSkxTREASM8P8KyLsJ
wc6E3omrxpp5ijN32hh21fWfgBDNshI8u08rk7VBJJqToI4w1GJ7B/CKN+8f7sSC
BIVSgAOcTxNU9pU8FZR00C69CfL18OUJ06THwgNAi6iy0D4a3u4bsIZolUfXAa17
Z42c13ap+aVX7chBPVHAaOmqHxQgZV6n0u7AX8OBNfulmK1q8FSyLd2tqPoxMUIk
BaX0S230YoxazpMA45hxRJbmW5ro08yac+vFbNACrwsZ+fToC/TctSGkLcVeg5xF
wFZVA9wyW3W77KLO/7JdM0XpMal/VqZzqlnW0Q57t63OsR6DahNbodErHrkh9zBP
8C8ENnNddGbIV8VJDkvXuIEM8cMUTIFroG54oWPAZxX0EVq+RikSg1vTQYC+LnEQ
1GGP03AYPHV10cfnnyNZKvj3neS/QOGJ1X1YzNBOc/LgjHRpaaAwSh2irhelaUEZ
o5wbXP2mf808lFknSowW4yJf10pUgVobjeWTY1l3mGt0Yxo0udbqHhkZf1C/l3Sj
DmR0DGCf8bFzkpNIQCQ7mWyG+KuFKDi9ozhp2YkrSZxxlNdLvY01ZFvyQl/Aykal
Qd7hYyEostA1Jr+JfbToqcSHRrijXfMLZh5TyE9Ulx2OUSbXWimQLr/Tj1sRVpj/
VdLKS/FfMj1qoV6m0hsnW7LCknPlDWK4IzXF3EbYLNcNChC749CGoi27RhY5WhTe
fkn76dp9FN4CBAsHWhUzClIrb8aT8KDInBSoQsVcxe+R5poSGReSmfVOndIcSU63
b63tBanQC81p6XsfPTbs4zpVz7M+J8nw3+A7lR4iC2eczJwBAhvDpnExpz8iNm5+
57kP4CopdusWz+IX4vmyxyy+gVqZiDaOuRnzd+cSic/tnUfkpEYiQt2FTIw8RIDJ
hbPXXIHe9+2+Fgv3D8nvzC6hwnHiuuztnquH0ZPZDLrzOdA90zsagfbTgV1Fbps8
YhroDH9r3pR4IAuRKuQeIil+HszycRFZDD9PQTdIO03mCpS2yXnmSO68cGLsxzSy
26u410kbJsbE9qAN03wwtqhwP0Xc9vUGx5o5PldFRTvMlWj+yJGjWdu/cA5V+RDG
Yrpw8r/JLu6s0NRESYDAYr254JsecnTKERBAKqr0ZD+cHrDRLpsicvB8iPOAUAEI
NX83nHhNlC+AmmPvdPq09XWlSxKof4YEWpbzr2zketT8sqE8Fom4JRFZL2upffAa
lH+juDkufgrWRGxBn4z9badHQCqIuy2FaOAz2ZMzTBSVs8IXWEq4zqmj4jrpTc73
hwYr7dKmgJyP1Q76/y0abSV16Mx3PMSttbRijIhpxoZFjmMKayzS7Ib1nDMLxMe0
QXqlTJ014FjKVOgkxN4xvGVWB+IuHKsV77l3tbgok7Fg2cTvtsoE1wbX350Zl8Fa
pRSjy5ogDTuf1evfzuPRATp2J940U7MV3vOx+/pLOvQD0p1r5yZPag45ehEOhlaR
JbGkN5RDpbVaY6fFDRN+Wu+FMaDA4qja3p9l5xeBSG1wg/bHHkUBFAucQY3Su52D
8QxDOIDJwMGViOTfC8AVS1tkCsE69d38z6990shuBZpJt8xaZU312bNgrcLE3GS+
gYtmYmNEoheiK/nbyScOoVrtOGffOW1bP2q5DzD2t8V11Zw7uViixcSTMOLQSbdq
6RlmgvvPJ1QkjbMJ0vr6oml7G4QnkkLlNLjG0JzuyrfHSP9UlUalU29mJK+LBLW/
/fOZflQ/vAm83y8qDKuj7zTMhf+5bdLp/y/3FlgHSdWVFzDJZ8Yj0SS1hdBpN2Y/
rlipryS+4MAaEjvPq4EVvyNiWkgqfpzaw+Gv7pRAdHlHb2xXipYEgcOJFGcK1ae/
BuaTH0MeTOqZfu/7G+UqhTA1/7F38AM2DLVzqMt4qgyaDS3opqP3qJ4iW1/6q/e7
8R+XtE73popQ5DKvq46jARPWlal8OXhaN0+gOIb6fX58kRHgXCOflvWqJYGMuHwF
bx2Ty8rv1gzfMbWJVr69gy7dLbBh5Rso86Nt8z5gFmuhR1Cw4J/SXkd/STOT8kCr
KwxlrbD53+BfwohYJvOdlJFgmbF2LL7KI80Lhc7Vh5OPDpHmYP8g4+0PL9ETVf3+
1K3GKziCKmeMOROnsX7aYVI7Kyx3lBg3/KJOt9LXMj3dMnZkoLnHZYoqMyV12Ql1
9VY0a+O9BPF02SBj9ddX6VNtmryirRGvPpO/q/yeSa20taEheZm6Mbvi6spOX5tM
5wr84nuZ9P3gFVf2ypCMwNguOLbsPfgUbdza4KVKBXDsiqcjX2P68AggUvWEyJv8
ZU9qYgAPEey+m7nsXPqhZ0Vb7TzUJAKoRiF72nA7RLh+jgXl9G/aP7BcGSiKpRtc
E0+jkZAutrlZ+BjYOFEIRrOVp4M7/ANzwKLBi7yShOqKyvSCTahGQKGqNazbiukT
zTC9yXdu8l1VpJ/e7ucqWlFGQAcbJdXxkertWk0dEtDTge2GgGuecUTviJA6pcRA
k2V0Gz59YE06UJ05hKjLKKU5clKpZHtjS7c0vd0YL41/4sbR0AhWrizl6+l+h+tw
dmwMArGDGgU3mMQRjCf69p3MYLQtFsULzBXEINo9OS6AjVJtpf0XJMS41RZkrmsX
uXOcbcaP18Rcq8/5jAeDzRCt2nSSUHKWMlYfi/BDBxy8AzZmeAvwbYnQ/ftuVnPf
ygSrCHLYjo2uLgmiew1TdEhnzCXtErDOGwWQiMnUwm/L3QZ4t1/9ghmgh482TUr+
BNa6hQccZYWIWvuBY7T+SsjIn1yTmuS4BM2XFHu3B2VODKBD53dRlKuoe52igVz8
N80BtDMPp42Luz+GDNqRv6xSVvICzwNbe5eEpdzv4rj/NgwBRapEgqdr1fom2MqL
KeiFzzfo0Cwp1ubB76vTg2liEJFT0nx4ctN3rBb9pnK7oDOYQcw5R1QNcVhZ7hD+
F0Aa7gNROai9xn7g9SeAgahOcYiQ4mSdpNDVJseENgWjpAF2KxxRyMTw5kWzElSr
9S/9kpP4bUeTaV7HYXJJCucQJztvmfzUVguqJog8jzapNfhdmHwgP8kGAP37JkoU
F2zvz2h8pDSjfJUppoiVTnNEyApf2gQRu/fbhySt49WY3EKRJZq5Q9c8bi5HomNC
IIOZvOSKH7x6dePsVQFdKUEd9EpYQ56/zzReZRatdnuk3ySRVFWOdIhqjsaBbRYU
4y+0aVGX2sGf/Exu5FJB9OYLuuqwhdCR2785MbOALyDdxcqLkZ7KOMot/cwc4dpb
JBkh6D8babHUgioMFEsVUOKT5BK+rSzkDlvmMi2AkSzdw62+YHU0UcN2Ejip3tpO
fgvbjTAJrhjX+Rsul/DTKCRiV0jHetvMgKiQytVbhn8nbGDBoe+1/xRCQuUhkgQ0
Q7uXggJRoxgHaYEQ+4NKkc+a19P5cge91SAU601shee9rQbQSo+QB2R2ePTaFDCe
VGTaK+DkQgOZOGqda6tdjuCqMQ+iO5xFdD+fW3Fj7e1vKjKG7iJY/U50rqAt4Clg
amKIXL7PviIaicyM1C6XIf82Qzl0jKx/OD9uKzsD699rkBohQyJlg6ENPO/Xcz7b
1pRrhMVEiRMKAETG+UJZ93MUOTdZ8H9V7sbPVl8qcluNpuw6uPvLoBl/wuBE+rnX
g9eLHPDrAmk9p7YlKR0vc62OXr9YDPEo99SAHHfdm3w0PEngjpA1ehot0jG8wRbN
pjEWjslnjN82Ob25ggDUkHNKwHReA8GYQD2h7V1uzRZIIkCgwJB6MbhURZ33E+26
/jEh8XzjmacWaQ0PDM60i/qepGK2ZNdrvpgfac6mAFe11sGmWcgii4RojzQ2PfNE
7ae5Bx7JWCEtWikCbfbMNbb/0VXNbImlqTE6YStJ510QtkNv8G99oZ2YqJqEu6lt
ENHUpnPj/vUBLe4jpYRsAFst3/kmSR63oQa9AFUV7JqbOgvHj2kLOSWibR/DdcQw
ROx2xXDDRUa+x4SaNNbaaHOsOOXtvNxMlrCYILHjjFk0RUT13+8iWwpryyDgPfku
lUq970qD33fHrbfhvRN20SgkKAzdASunTrVD8aJHYn4p/Se+yPUwiAjn4awObBQK
d0mEyHL2jJVRVkkwoW5aS+mnhJ/hNGzoP+DzR41P8uJG/oldb5Gi+LqeuEEDkxVT
PCOyEZdrRHO7r8GV0+CoMHd89w2QpS2REhnV1EFGitT9mOOXxivGUEXjWR1DYapG
F4wOxtvFlYZcwTslzNZOG4LELLcy0cCs83Bzeg9zeAqP/RswW97KGDBtMOfWn2Xm
UyE68751vQH98ES+OwP+Obrg2fFltwYgwELyInGUUlKW843IlNX9/m6DMBXEi82B
YDxNMDNe8pSmaYAZnscssBjYWIMOz881xcw73IvSZVa9DIijbAWuv8/AdHdhOHRQ
6YNtGxC/jeYQNmPj/CaN63+g8seCKA9vApzfyYa9Xlpoe1nb7SaqZwCefR2Elevl
1JJl8tMrYq/mx00teYnbr0rUkqG40EqLOjYmqyOvsPO4Z9/i9tw0hYn4Y5c1vI0Q
9+YYecPnTaw6rBevubsOjYET4H7/8IskRER04DaieHRkPUUrivoZkS/HC+fsmP60
+rm7zfXHbwZu/CUyjMzENPVC845jPIH7CLFJJKj5SXoOSWHBixFhcUBA3MhNDQzp
OcVlY6urLu9uvemT3ito5V5iTNj0bF9JhGUbLNKV7rEQAw8QsG6gdS4S8u61mBKC
0whpRhQLCndfEeTNVoqPS8bcerfiJlFBpQ9nmNTnGvx9jkNfmk0IEptSU1fJDzGd
yHnSx25sVV1nn0p6Dy0qhj8tC06Qd42a1JkYux40R3sm/KtBuZevqeqe2P9YzPCz
kH3TEzQra5QwBVmsLN1hkdTsB3yl3pr/g4GpHaUMhKisymvpvBog657jXZ05tTln
GYYqYV3B71aOHO8f8vwHubwKoMIXonkvON3nf0asUVIKzGLqZ45Cz+eYxWysRlSD
GrQniSfZ8T+/OWVPwtOcwsStgsGMfEcdDlL4bpaHeWidoYhKnA+uuwiW8Luu5huA
BvAyNNOSRILK19xohbBs3i7xk64Xk837qV8mQLIWkqJa/QQOUvZdMjmmI3qaBBcW
uprC0HWtoaSEjl5OKBAqaiwjhdLFCAs8rTUWnPAyqa2YsWtouOWgLA3I7E9BJTOn
OK78Y3Is27Wwc1SNef+vP9VNROVMuSwEXp306P4iwY0VZmR/vk9Kc1UwkwVrPPzW
pO1Q0pVOoKxc4miqhtpTCIDm2lOOYIfLd8+cCTiG6KT1jUt3b7n+vwuLiHWX+F5S
gQCR/+eA9qfO4FWf+7dFJgIwMW3szCMCs+VcCWFd9XZmzoINSOIaAiRPGAX6kvAb
RbL4MDoVNafIVs2sz19HucofhURtgsaqiSgl7J0Yf4khubpauyoZsLdRI5OqIh1c
swnbbvIuvtVUArfPpyB6AJJ+sBqaOW11CwH52Bv5N4mSeZtwHrwO6Ac6+Bk3WSOT
6hunNzanQ77zioTYrCIAdJ/Mwx4ro3zpmS4MKiRI4wy+FURZpjs/G1wsuHW8daaG
hFz0zI99ultg3Q6cy0n3lfMyok/9WUNOFmK43qyUxTcTH/ieWHTZ3BE+jcKrY6JP
lkzkbvspQNRaS52vE+37UVMeLFX2zRskukv/JAEAoUuY8zpxsrjdByjzj4+29CuP
BSAzI3qQFiEr3bfYpr/FhzWtOj/nQxNlsp8PkkJJnjcSTSNfnovzhkah7yhRiBhR
lM6vAqRiTX+MzQnw6CKh5SIgIA9gVUl9bZkNZtTSpXNFnlmzZnzD7VRYKW5BztNN
rjxKhQUQezGNrmJA/+j6ZKBZUqbtAJwvURF3BcQ+dtPfIghCWw2+5UasTI5pSyha
6JkuBZujqZYoO9O8EFVr32MDxUkeUZH2PGerkkKk51qKmkcyoflrVcNzU6LhWcFb
KqfPuK6JLdjlnLWqGy7sEY8Nw5yIhAa/jheEiUSlkvWtAKa+MTuG3MshgkIKnVXT
F7FvF5c9W3EOWHj6Oce4LSGl5+CCDtK2YeFTqZtqZZuH8UGJbSa79ya1+ipmobkD
ZcAwT/RrWNwbx92UdgGfI6jIAhqF+et0p8bJTgSuJIancfdwF8wATHGoxrz3JfCl
F+qhI+MVu2uItviM4nv345FoHQzhgTQ41OfrNsfCAu0TLNFjY3uK7qakVtj6O+hU
HyjH8pxB1ZHuxa6dqVyTlgxdVlB8moceOT1sFVfZJkNyK8ONEx2OXsXuXL1gt2MK
qYgxD0OzC6G82FIZA9grddyT1EB6l1/2l9LO0hLqm0TAwi8B5Ryf2mKTn01sVoqZ
w0WnFhtdHQ3moL8VGUVWt1/bYKuOBoKoWl7SbZIRlPCn7fR3wCEuLZjph3Jl+TUn
peQ8+ja+wBTNl2U742HVVqs1qc4mJd63oWyVDNhA95ycLlEs2lYSwGIjJEAoOvwo
UJ47y3Kc+9kcPBl9UGeEVzRWi7chO+lJ1DSSYf02HMhOiL6fIFj41VSZdKfby7OA
dUZ7Q1CVREiNvtUBuZruZujqWLovY+tPA8mnJuLI+67+0P2Rq2l5rEl0jVXHCzc0
IY09kidzM4sE2Uq9MCGIzJTFWgXs4yA5ASTn1mLMlu2c+HmNtvUE+di4n5QrqRvG
wqBd6P1PcKentHdfX+I1uF6kSmNSdquD1XD3UbMbaXGbcZlEljjTmi2IPLJqHAIT
thJKnRoVeE7MGxzIooovaRhsue8BEJWA115tgMpJIKWY4Clm0HZOC/85Gq4ArhSh
/SIFro4KZ3DhNC5XlVXWqEIBPSWAA8uQf+giLJZW3TtkFZKKlPHfhQnfvoNB5ibG
F4Y76FGZSvWugOgAJ1iJBToQXE31F+LUt7AtpyA6zkZTZRb2kmbHwYn3pYkm5ybP
GzdgmtBmCApndZHvur43L3Mlq9IdNuYnsWiFo6DjJ1HQaoTupYAjfoTcF8QRWaNh
IlI6G/QJtoAju0JqnhnZLq7jHiO9bO9OsewrHbkbiBmsaD9rlhyR7r+94z5drJmp
LW0oNhXdH36xrR715XDVbm10SEW+w85XWjyKqghBl+ndPwMovkQBtWIxBcc0aOZ+
oOEvPCy4NBK9bvyHKY2MPOBtgszr66EvpKMVLH2tJwVsHIICrdmE3oM4slLHQmJl
muq8X7JkhrUc+fUQbvKt+fYyFrZ4HjNrykAJHZujJfEkDDI0XmN0nrm97g0Bvpy0
Asim9cPdTlvVhR7nX/yDsWqnJ/V0FisyAo3yMsNZdd/wxTrAQ1EI8TzBRwRqpFzl
0d+5CMJ3Sb/Ro4v6hEPlVlzqyux5i8hFffSybO/f6rzhlaSnaswBt6BGnDkXRxOi
Vz+fD5Jn+h36AMir0e9qZimYgQ01G+ACPHwARlAfOXXrw5WmfXGxALtdWOJaje2V
DCKmZmyABFLkSyVZtCVSh/gINcp1PEOZVEFuMLwNhfDPEhRXLpliLA2IJt7lDN48
z1Zw4guu3biRcg0Rs0lcBNFnDWaEPIai3vDyl/0+UzDQTHKidncP4thWZnzulqxg
8S4SiJwfGKA2ExIGxWBk2fBQ58cGu/aKMnHGfgT9loObJXN26Ts5h6YFpFg9l/Y8
ZDTdl8Rze1ma4vSyGQENvSqI9hvZqvf91HyoP309zTLmLwPeFWAEUF9mrwyPjVa+
5D5c85pgSSD/zcP3WsRfi3TNVaM7OfiN3F9QquepJVuVEf7vu1OOZQ+9Kha9bPK8
uKuPvSHv6ycnOXorYYIA2tcljWocWZUhwhotVkZR3/YfvQGf/ocoPxND2nCU6WOm
2AVsozApl6KA1Sc17umKZ9PmVsI5UzIq/7dKbo5KLu2tQ/2el8MZrSeU5/pJTHdt
7QqcdszBn6+NmxI2OEV27brgrtc2YJf97IAhlUNQ5Eywq7qdr62Pu5Gz7wjSOUVQ
dVbp65RZyYMlxfGpyX1F5DvPE2Jb3w5w2KnX81vhKFBx36O55Jfkb8RQjtjMqO2T
HSgj33cUKwkxKUdogLOnt71Ca4T29QKCyD3e2JC5292Pa3U/OjyvTJJK2F3eS5MY
yee8O5l4dS/e6+0fQlNmV1OwtUHi1XeHxsZSBmMhNKUOweAxNtvkL8DATTQ065zw
S+e+cayq6rcwAW9YxcfD017W5PfBdoHMg4RgQf23uQEFeIRoLPprk7Bm7WSbmtFC
xUad08ilZKZ3AZJ/k4QRj8Pf55kRSiJShrS9h+9gj8AhwLGYOh5ET/uvoJ3kTv2w
2FwGQxseLe+Jg23aQPcN9BRt6L7DKoYOKUGM4aFyvxIiqXzNvqSKMpTcSg3kJVxh
EHyun/FATuOeOUww/j9+pCarpzbfUNcTW/qy89vNa1hx5QwNfXFCpR2EcK2heyS+
LnIuD4OcHvmm5zc1TnHLSoY2j6SRHn0HXY1WrqttCP+1FJy7M3CRZpPy8OWr+HCR
ovTnqHefHHHwa/JD/hxVQUMUHJ/O3x0tYxyOqB6p/p39weQkWxRGs3p+2oqjqAHY
BK8yhSdeh3edutb5uWEvbWdxYkiGr1vCfJkQOsqmyOyY5tfA7Y/EEJHftZZzrmQB
4bv1m9FLej/vgI1ixh3/UIyrtCGH1a+s1vHvwRVVCsmZ0P7rZFothqTdW7cPSjqM
`pragma protect end_protected

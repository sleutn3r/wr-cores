// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
e+taTlJxXsoD0BHGxc7fc60Z0gl3q4jfzQzhWUzq2s2kHSxhqEgs/R+fyVDpX993
4YD+GMGbCC+by5NNmEzIiObt9y5X5s7aWytVe410GlfIenAWC9hJy+AVIrVmbqQp
0LTR9rtM4KbnCeoLgZbt9T6XMBXYuWPnJDKUKhOKgiI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8960)
tJLZPaz7HE5PfIMHHmnhceNaZ5DxVgRK7wp3XkRg+YcSckMjzTfwH8pidO/A7hAQ
HmP+QCYnVrYDvOEfAw1ou/IuxQAdX3p7YlB7admhIrCXrZLUPek93fVC6dW1XI7A
+UcNjpwnBiuFr0zi3Wg0qqHoiSU7SJR1nTGCs1MsyYon7GzNPzMh5+8AS1jKsO2g
dTYuVOmQkrDt/YDBRC7xup3EaqXVdZk3qlEHxHULBNtEKpJtyWertrm3Xh8Lflbf
HzqS9jvWMaxGlNu7j89zqfMAbaPbRUvo/6CiwSkwy9qfARS8odvrn6biwrNxiaPA
zvXZUoAk4FzOYh9xyVsteGxY4wn0V24ZlX6ep180caGhoaPFctVGpqWW4uIeFvnH
y4eK1iuqk4FaeOfJUDwOf94ewGg0z9Lc1L3CjbpyrjV56xcwPy9z76JfQJhA7hVc
Q//UkyXlNEqMK6f/9zY/esvJEnId00fliORGyVOYzmTQOIn1ro7gRu7/v4Oorlzi
t3RhcGyHWOM0i97HSTB84U3wzUz012TMGzlEq7zAF2GSkI2n2Ln+KlQKSsSoBNyM
+cclB5x97D0Uz38rWz7Hq+LTc1Z7OAxy16b9Fu70WNKL6l/PCEpFZAoNpbHZRg3O
MMhaKGmgB39t/EadXOHez48zXZ9isCbieVmyPRlhr+FyOpTvVI6dIVkpbu5Wqfkg
mxrIvkK32Pc/qFdVCavNpGY8Am0F8lr0mJNoIywj9J3t8uBsnxK7XZ1HNWLxAXvz
NzmHfA35g6B3KjPPnQUhsZPILX/SGZuEcNsw4l72SDvPzTgR3AuPEQzK4GBahkPw
JFUXBh6/k1kGFqNBnWGN2HeX4qp7i2YHgg4E/xfwZpzg93K+/P08S1qaswS8PBDk
cfyWKisF2qfhKX2JDuah1vAXvKgWvyDIty1to5LYNpi9efFRQ76ovihHem3f4WEy
KFXtLP6TmxNc8QJYKJudSdQt8QGckBk4Dv/3JpTt1c244sj1wAXOUcY/8OAn5UXC
IwZ4+GIDTGesEX2x9uAErhT6xUHlUz8xzVlsoYZYmT7q6eJyHUeAfa9J7xxHkTZL
oNhWm0+mmY+AmVxPZGAXDq12yjDME8oxHg5pJFh6OVqfAM16EA80y+m1+Cq95382
E2vKn2JLUt7mM39S10tOd5TJS3yOjWX26RXIkPyte4ZWld/KA3keAX1YXPrKKkya
O5dh2DoUhdZC9wW1gg9BGYCXnbrkCgThHnQk/Kvh4N9L3ZZ5FsO+yw154PB5HhqN
0U31SYrnJY4iAOYk6Sgm6iC1Hp4Say0PV7+Xr+HiYaWvWBxa/istw4Va8r+L97u0
xAgMKtEfTG762TqxzobLsj63jtXkGYDLI7kml88JdTvU6qauWg3z/5qTF0QmSC6k
6KnoXXvipu0j1Douwz9aKvylEb56GFeOXekOjLzPhYoobsJkVioliO3USk2YUS2F
TiapeRZkzme56PS8nhrmlnITk4cgH+wu2G11hGXoz4jKxFWCZwJAvuoK/l1ol2Ci
ejTRcH2Fjz2DH8Ce2tnMQEhFPGZAt++v9L4znEWt1vWJ6owKJcwz/kRrj5BP/Vsn
3LeK+k8HtpV3vTWA0XgN3wx/VQmuuNxUjKY6C+njZcd+Wo6ku3N9jaeVtLRhD0C5
Bvw3eVKqzwPDzX90XReBhr9DJR0hDg3bcbUWSyCudEWvM7EbqSyXUlRj44UjpsFX
3gDeRzPbC6FMlZKm0jpyW58WRuNa4V1etXp/axlX7qPKQhvGGovloCHxvlWTivCs
WTE5AaHypackoRmqWTZMWQYNOngK55h3hlkacw8VGs2o7GZBh6M2/JSIYeAxYpK2
lcxGXevVagLdYHlh8xBjuq7nWGnrql5ETJsvOMolmKfOuQ0xXj5wqUDAWulxl0V6
Xqh6+RPQ9xuUiaFvGgXbFcyiffgEu0C9BQ3jXl6W6HavWbbV10k9MW+hMVin/s5t
N+QcOm96beI6gQ5RIZTob0SydgrgxjvCjhk+x4cyv9aRf+yEOfNwIzUKKWNipmh/
RyR7rd0+zqSfZIDBjhCsIndrrMQ07uHvpwdegzNFOoXThqqcGsqojeG90HZV9JDV
ys+usci+i7c8RzixyLKOOAUGws4XMSSSqs+/0GKNccic6uEwQK6PpSDYbJQjcvQf
aGjC+bzmfIRXdB6n0xR0YCO2KIhDUw5GRTDDqJ5Ax1Z5RokgPmhDzIZTX2OHII6i
Bj66gp1jWH3iT8Jq4gs30j3kzV27sn/PLV4B5Urgfe4VOPFGqvVHrIz2EDVXqHvz
jVIdpV48zCcFvqQ93bDRZJec+UIDA4R3mey0aYP2oEqoYxLfIsvcTyFn/IYV4vW9
s4eobuOItvG6iWXbcUKjgyqeCGECovqW/tybbkguCIHqwxTFgj1AG5SX90UBGSlV
8Hg73V1aS87fw/pbx10NKXKS15Fnq7CG30wnovRiAwEfnwxD9nKrgy2GFATZCqac
QyMyvF/n7AIJUMeYirdVcmvYzJ7c3pJE1QSzVyhY62gbnlYUfUvQ7fAWjLVC8OGy
8gRrpBUt4YuAIsHfFz/EXbXdY9K0OYH96w9wuQp8mvV+LMtyH6tslA3jkCC60CSy
S3DL0IrqXlGV60rdzU60cnJL3VwyOygHQMxINE3yNnzBrCb7ewRFwg9bnStd2+GM
1XrlYkmMxtZlMwHYXfLoM/qFlDm35tpuYOxDYfG6jNBhwGbMc0+481IFqPjL1W/F
Hq98BHPThTibfY1Y8OdDjjY/HqDLqAdnSXo87BO6J096eIVRgzGefb2mpgl5IxGS
tuElBo138wZ0oXvH+Itfitu+W56vrQNHOupnn6hrYkDloj9nRcmvQigMVzh7hz4K
qtFqNAf1jbciRK7lUl7cf01pyBM5cp3ENl7cWY5NQIFvo/gAAk/z+UwX507VHfLQ
8ksAK9AvKR3+S89me8fpvdqKF5D2llnoVToHIXbr4L8F2H1XLcffulG91tISbOVw
pbkhvZjOQgKlrKMGQrPcegQ2gGkJE/HkEYLYR4R6O3GYZq/NeKf4n9h8STCxqT9D
kItQ2ksY6qEIpYwYFYeCr41V5i1z6ic5n0PBQ1TaxdGMahrExchOnqFFMPE9Awzr
ufuk07an2j7FNfhibpjUh9mDtak01P9f3ho93qOv1+TbrBpovjthA9vSHUvzMtEV
ZAOsCKsF/5MoWCF0H00GEeYDI4TCJ6NtyqYsxxRRANreOGyop7/Qr/ax1WM7jOXr
1ckI4xYXHDaQcETV+hjmL79tLyJoXJbeRtYsvELkwrU3xCw1EuIACe+dTNFxFC8a
Zr946UTvF8AI7+zQ6IcQyvp3xfFH46HPUTqHgaFeNb48lig/zoK7ibmmo9vqFslP
8QlNFxjxwwHjlMcpjHJR3l0sH+mhdcQndgI+DUQHAXyel9h9XbkBYp8cl4GoK+no
sY6gsZbZJHH/DcfcD1ko4ViQzx151GxB05cbc+x5xwS94gEM45vLmW/29awJMdbS
IWeyiRpzQhEfEfyPAVxqFVLq0O9w1yop0OG8YfU7LV2sLc9bjG4idk9SPRLq4U9B
4G9fTIAo/bnyLjNfOyH2xyowG7WHwclbRcqv+BjJHONVMBItY5TwvM5x/qwOIIqJ
UToNXUkDT7sMizJ6WRzN0ZR2KNO16iVI/Gz8nTWuXkWucIGgKlyq1AUPo1YQKp3k
Bfo7GhsrVMtGIjdmbSVuSXQh3p1H1hg2Ka/waQ7pK8Uy+RR8/ycEvYAIXE3VjG8K
YIVhh5pa1rIcoOsGbWuhyIcM7apE7ZeKfTSxTBBkudaIyN7uNDh5r/QD3uJAUeRh
QjhfxFcz8DO7mePaeaYcTkgImaL7o68lz34XhJTld5PKlkcUfna3HjYchlWGayhM
7kBSiV/d3IUFJnulNj7MLomtRS1gLrRQyWUTH0smc3wWDnKBXGNVOFkj8goN5RE0
lgTnPH9Oq4kacVGDIKbY+75YM2YvSQNmGzsMhJc9afWNoZyQIAsrZSrSUYikYiuA
9ZmLSU38ysqmRz2gpfZ84y3kgTjkNW0NEymImzwQv5zKeWJuqGxXrKxt44uqE+lS
hB/0XLXQf5H+UYDZg1f7OKgqUs5+Lb5riCMS/6ZaBiLO8/v65DK7ZaoymYxCSe0u
Dk6w1eLgyxynTJi/Y0Ld7IomcLbNq+e3cfCKHFfoyqe0mwnZ7AiW9Q5RoshqsfdC
kLvJgPAh7WmbZXM1OjtdhfolM/JPgIfBTq8oC8bBmbxiYPR4DvEKgQDXTOYoSrR9
9L66oh2kDSs7rBXeV25alii6ueCVupaN7ADW+CLKgrhX4wsQy0C3IKnCogLpr2jy
UGj3a82QuFyJ5zxDGjgXuqie7G9bv6pQqw0gjqDzk2RDnG1jxUruvJuPkzx+tgFb
xf23KI8vBbA0VeUtvOdyJSLrEQtdJ7izMLMkV5oYeUdPovVLOQQtJRqQIIf9Y3Oe
CxwhXkyerVbVjGAj39kiyI/C54xTZJ5Gkl2yMvuxnnd3Kp4DKEM0nUJTJJgglkJu
d0R9jTdT4//vQi1lsHso515us+qs4cmSZ4S+6jCm4OUOb3VNWvqsbhr4d9zqSrIi
X0xsrOprSRCfBXhuVJU0gHyiD0tM+uZQivfwRT+91/P9zqQKog6U59MtpXaeFR1E
t8kCvTR7iyij9XhKGA4MBkIeYk57NItdD2D31p4tAkyEsuFqFJTAkVLRzQa8wbya
zAQaIew8fw50nAWjVzKz8WzHkn28VBKP+6b7pvwqUM0L3+QLlJ7/IGDlA4SwsgsQ
/YSk2hhHMNT45d+jNqcKlTzDTMi1O/3VXOYVbZrdylHykYG3eH9Z6DlFSQ1GoOB4
/o6gQrNPLS4+B5yGYvEAwZBYQzvGYm5G2hpAsyzDNKh3u9e6qR4LOX+kAxQssjAG
MCUIiNoA/Wjxw+jDC7qDr/5r8qoi8dMPEgy2VZbBftBUHZsN8TdKGUzRD1mSMFm7
CsCpM8ntnGAgJjRcEBH7f0arWrIwiMm66C2vUmTMoBl9CL8Ezl1MUaH1Pr442107
ubSs2fUvggZXnhVi7G37dRm1BYnxARvhIx/6zGRwwGUK3BSDl+a1NTK74ExX9glg
HwABMQArJIksobMtby6qzaINYMNfbphFTknKc3lvdfIN7FD5ThE0U87T3vLSfUKA
ttI6ii1uExguKYpgvh692+ztxdEsWyXo68yhpjGUKTzsWDVMEHo2vOQw4ZrGDpqD
vB7lYEZyKLIpy6mEf8IA7YUoFYcU70JKADxauhtRj87mYVFzftzN63nShL4R/70v
m18wGoyuQVO/ya2sE1Pd6sy5ZVgD7WHAAue1GMhKIls6x/yxwMCRP0y64Wqh/Blx
paAMwLz6RpnZN5YUDaxWtgpdAAHQ961lyxjmK6AIT09sGms5PcsrKaZOdDmtvQio
+/Tmk5G9yHgi7x3uDtXupRQqBPOyal1nGLn+DSK7r41PR24Cz5dgKbkzKZwRs/dk
T+XXIEn2jzVaIKI0e/sxY/01N1D3psSO4OzhwVlAn1bL51d7RSF4YjLM9S6xBxbh
I2xmboS2VE9AMZH+ROaD72gpColYueiAuGmqcrmctloyF1x4Ad8JjeU8SrHu4MeE
MnuGs+LFriCRocZVufAe2GfEwV91pv7ia6emVYmlbdTBJPZOAbXbsKf1spV3GDja
HuBG6CVjfM3ZQ+6NLUIbpvc1s/mG4XJGyKnYBBtX6HDw5MeCiAn9/VYdAbJQiFi2
KY7Qmvd4pzkbuOR0MEyFfmdZa3ucwheg0ZsyKyGsErG9RlKiBNS17XBB5Ae9YV3N
mMmOfc9fmqNuuszTASVPeZOEVcrloQs0omY7J5byXJgDkpfSsDOJWc05rCQ6kzV/
wCOCG1V8SN7YhthXAd8AAnDe+n35s0pfmJr7sAnWXQrj5T2bJzu41sueuvAt04DT
QxZAcdr3vbncVl1fFKE5urqP1m9LMJTNA2MPc+wrOOqXIRqrJY3bbNosOoi3jRKs
6AT/m3AX2Qgtp/OsxxOPmTjjEtUdS0g9DqZgykvUd76idE3BIcZWP0cuZVZWbKVJ
nXNWdsz4edCQIkFTk2HhtnRvfX6wFsY1jnrQmKh05HoctsRzi0RVRtC/It9tR6B9
5rOBblMPbV3otyoE+K3aQmTu6GWNktQWINQiOk6J8TBrmeVgk9zaDGoh4bubzTv/
uGiyqaHP+DxVIdo2vYXoRiPyswLAzMTfaS6LRIi79F+4Oa79XoSa/rjd0CQsZOIC
L/99P3MfmoB0DvPIYedKENtr7ddRZR2nX4wyl2BqZtsKsSqt7HRoR871hz2T255p
m98ufRfchd3l51bTkyqvVQP8ZR0su/k/9rVzbtV5HrpDbLADTZJrFKHO/R5ZX3Jt
TcyvYO9+Np457h8r6TXkgSEJ6C/BcG8kv+vMxgEFfPwHgkoi5n/MoDcqX5dK2SOU
gWnQnMyU4Lst6UN1WaU/jIlg8fFYUQCybs42BnBeykTzYbdI09jYKLucbb8OVkIc
2ZY3D+D+8jGlpRrIjhiw9RsiNOUUuLD1dY/YhQf5hsfpt+N8hBU3t0XlhBGFsN1r
UE4b/8E5ZhEoJf8l2u4siS1mn5oI+NWyOeI1uSijn4WFp+VrcTEI8qN2beB1B+Zo
Jj0c+hQEG1bVoAe/+6XYztnxbYNHsuETrRPDx/EASjZ6tgDduVULTrUIICobr8mw
Al+t442flVlIqpO4o/TNTGDck8ym9rURIRaEIygidzblZNC18s/zcvA5R4bp/iPc
ac0Z6+x2ubJFurkXbN6MczAIJkYuCQbcEyCQVYyRyMm+ynFe49s9mRnxX/Wjm5fd
Bh4kUjCdmN1xMtqVRy2lGtjhSEWpAlWE+3vofMynEcH8xDXe5aNoveSEicn/3bXP
H7jR+Tru1IEWVUAUgGAYflYkR2RGuTVzjFSGUa0f9yKghGaF+PkZgVoKNLfeAnzr
QBwJpUASUGIZGezw5D5sup5EO2DTDwZ7kNpj9nflqlVDhmkGUiS4FHGNbZa+kgSI
52w+5AYKdIMqOh6QfZ1IN7Hi/Xkwr5z2dagSZjjR/xgsKwzPW4Kf8zHY5z2C7yFJ
s65lWZvf/L45lxwsz1Uz7r9hC3ZqIcz2FNtWdMyPF8yfUgVQMzHrCiPSwUQ3svHQ
PMsU9RfIN7QWTThgNNECNZ9/TgJVxewhjH0USKLmZVDNLtH2SfzamjXeeG56lNZN
JwgJBoJCbsIzcCB1O5xsKkD1mhVbTYbvgJ7LJxFZxOH0gfB/JO4zFez6BQ+J/O3V
u1ussKudfs1dFlCgFcfIp51U3lbS3fB1WEHmWXlNMLmxd++1+G2zcKurfWmmbVQv
bUSwXw+s5flsHkvTGu7EWfkiQO1ZZ7ibbgQxLHzQH/ynn9FlvYMqPN4Q1qUJHYzr
Lsbq/9aCOGUAJELiqqJ1Kp48j4BZ+AQqdktTg6YULrj1qJa0dhBNCjD+kDGoKL21
vkM1VM0Nm584IbGKspl9iCgCrumdVryNtZ9vN23E6V27mAPc3maUFdKPbQyRu61v
TXlaxqHTKK6OFC4ruLfip7qu22zAobsALOyXdayOhspWh65mhnGLOZTEa/X6kfyT
DGTG9l2vIAuhmJYlCjFwBQL7q5RjN8WnCw0NZKPwdQ9PL0Kz/8ZKWp5zQ6TlfBVN
pnrJoJHV7WlkCfHbA4sCd4K1/Dus2GwVjSTYs+CMpTB0+o7zj3NRDKDeiWLqoN7T
rtfjZbo4cHCy+WVpPR2axAbNGd084oqlFIplLAjymu1mih3kEArZHDls4tO4w4m0
uYcr2OUyVeS/I+GIEDM+F65BRE8T6E24YAfEA4Nr0SaK5j6Kpl5NX3SVMKLe1cZy
NfpsivA8NeZkIszflgnhahWTGuqV0axaKUD/XfbdozQtn/a0djlkVPdNJ31WKyd+
bi/uUrmYvPkDzajZbDWeQWVIoLiDWpSwMFK6Xw3rnqM9AF81I/GWYfWY8idbRXHz
ApghE5pK5NsG03tCya617kCCdUktxqNmkY9uTlu4hvsna5UVhZes57Bf/NAniSbs
Lmv4o1hsRcqC4EW04GtW60wOJsB97Rw2w3DTyALtYRku/vSRpO3SjvM44/fD4Vlm
xagi/SU4UY5S8vmHAGzhA4WbUKySkikdnkvMbjAvykH2eaQSiDCDdjvaP/nhaAZB
Q2q+CHokbmDfdrHxAo3nDso+YnfRHvMdqjMwcg8jSu0O31JjASSmrZqeN2N3a/Ne
hKqXkhErud3jHd0IFrY4uaXylW5pAcgCHY1SrLE7CyofNI8NslZvtH/P9Ee441B6
i9WToYYo1aDkO7wWGCPSmWV8zpSG/M7NVT/YsGF6bp+IaueH7ii4V6CLEO5CLo5A
neFUEh5NhYpVbkKiJGqfAwtskaOrl32hHET/S4Fe9njOj52g8tPk4R8aObB5S/uv
mVmsBrkLUz40+jyq6GQz2/8yX5kj8w5eLHSBMdIt+ORrnyQqZJMn7tlZZJzVPu8I
XzYowgJ0152FlN2ET4/quqYK3pTuam3XQwkai88ZgQ746txMGvwo9AFDN6Fsmcqr
+ezURwoUoKjLBsihSdknhExa8g3nOhjy7QK8SLw0CXQPg+rxZ5SRSg0iD6fhlaxm
NndAJOiSeGhNSK5b0GGOeM8QkSdGzU4XpNoL6ZhSWlrDJhVY44RJTCtU0scqGU3G
2V+DQYRKEqCFGGf2z3xJKB2mfySooO+LC64uzibbiPecPLfPJ4oXyC3dv8uJHMdD
YhKpy7DEHoulJVPTHUCIBY7FVOCoPXgKZRIaseNkUyeI4EMI2AC50Q4UYF31oqvc
8sMjN3MhAwZJsXIyQDmIedtC48gvjfnkDtq8RokotEiCZShLejxsx+E7HmdKTHP4
XaoDzX+GXVjhkUuloA4SSSmorUEuNbsQ7RN27DWv8QXIttyGUDAzZ7A61HMFZC1B
64aX8BDAkgbjMcr07765TgCM0f5hTrIKS7DsO3MP55klxJSvavNO+fejU2Cua+f1
5VfZUXH1qA0pcxX+UJbej0DHmkCnpyxzhBuhK2woOAdCKuPoCt6VTPupFbIWJjra
eGRRztDyE0ucIhE5GFJQGVWEdzEWygLYWscaCnJobBHCxKb/CUq9Q/8vGQcQjAwT
gyEC5cTjidnYwc/oAiH8xBoQSU3EKF/qKx0FRzGznlyMa1efluZh2xqgobuSML8P
Hi2ricXcxElu78nWIok5fqAP1IOa3prCytkj1eEjKJGx5ZHZW3y00j98HNYfbC+w
cRTostsTX1+e/ydq/F81LZV6mchTBCXSecWxcYURFDT3ftmrWS/+xs+4Eg80F5Yr
yUzmlRdGF6/IZumeILYGzvmuIJsXot0mz8Pcr41pefeZ4+U70ZWnkrsQtpGaDIBK
Bui7ZHWe39EzvXA9hdUygWQ2wulST1GAoS23rxafoR/657CQi9JvzS5rGkmuslX4
K3ErSpo/hjpMpQggBWdbL6kEG3bn5xi7Jt7FxnRtTZB4ByZv1PCiHzH5J0CmIZ1z
0TAhYXTxrRxWMjjC3CnEPeeBTRwGyV4+7488aAcDj5xaXAhdOeGsFwOVhK5sp+xZ
76/jY00qbYg30R3h2LiUaCaDewZTCGlvnkCoTkQF0xBaEx1cyap8Cm1yLb1ecgzf
vSsTWRVWIp43rf3q5decTL51sie6w4tmTTBYr9uu0m/ZBP5asUwD3ZcqWbQinrjf
X2yU3jO6BJwLODfJEWFGMMUfa3sOnQ9E/CAMssq7fYYo5j0rGxY2rzgGCX27xPK1
gFEpjqsSjw/NX8ye25o4wu12VG4brG0tUdPmhxK9bO1JoQmxjv6o8vOKcDNZDyPS
1xenwdKoWVJ2JwzB4gEQXZcILfWPVdOPBAej2O8Fp0xzxIklA0oDxUG8IhX6YRGV
CcWpE7Hu4yT+Kc19A7AKgS6tmEdWciFd7/8ZBYQ6riusyxn2hv9OcZXbcHUv8eaL
Ywow1kBuWanQQe+N5urNJPFB0QZuu3uCvcmew9hb5/WMVFIs+PGDalukx3v8VzDg
XOrggehje0HCXCd8m4Ct4/SjkTTyZKYqKMmdYEgm01zFeTyITejihttRkzyDZ5Yj
yDALJwktS3i8AjX7EnINFC4IfrbrO6uWmEEiJcsO836KUyxuksLBFFsiMid9stYm
9zxlGAS/mKm5ZJDxJ1AxZcHx+1qUEd6nxSq/NwUVDKqCrx5b+5ul0h0Qc9Jifle0
yRtvbQizHxCpZ21lL5CYjHBZut3QBr3dr6+AjIKoth8ff+igWWleOT8XciwJ0w32
Q95656LnklOtmlSRrlscRwJaJ9LxkOkRcSN/JI9Tn/GaNmb7ZX3PAEYjTkpB1Mia
yTIhm5d8wWg4iI8d35OPrmZOS9gCftfQzUDjP5cuFjPPj+TeGybP/W3zdgifoTAI
/Hy0L4qa1V98Jcn4rosfJspsVG7icjnD9FFJZjLXKSmXDtGbGOoKiQUIytcX9qW4
HThKB4Vlz6FL7yz94eSIItS0JcvV7pSGFhfi7wC7OchvmXOIGE2sB3mXpOkI9DsE
Tp7KoM/OI80ZN6o2YGX9TyH423ydm6caXH8GHDWBiRbEyW7MJU6Vp3vusb4eWzBq
ED3w+ldcxZqMyhV7nta1RlZJVIVvL+2fwwljfLGfK7gCJ73Xxut3KgH+O2ucLVkA
YzPyqTbna/9bbTs0elv+tA5lN3KIDe9Q5EtWIGoKsgeCAGPQOKW+TXNmiSHA2cNV
//NQ5VGVPno9l6WigTvH151mo4Lxr+z85PEluXs0aeqPpX4V6bTc1rkRt9g6kf62
O75iFUhA+B1rKMjth6M19FIBr4Cs4wS0Ge/EHUzYEBIkHeT36yOMfged7dWUEPnZ
a0KXbUsBjYsfVa7q12H+80tHzfM1hzOQ1kOtLQQTAXvSbqybjfORvqr09n4Z9d+u
/uczdf7vfMAQObNLH6vpswivHtNLHScH32uXnA+U+zusFQKHcQz0gfgL242ZG538
XcqNar5f77VCh8fu4I4Ui+8UznZwzqybBg8nmVHRKumBk4zOMuO2KW3Rxa8GPv71
g3FxJKs5vIE7UOtNedWc7EbLEkPitXXxUVVkapl5fBJWQvjWRvBN5stIS8zJJyVW
fcf1L6XccBiGxVwOy0fu+y/MNEkKIaO9GwFbVRMMzurhE88bt++MJPTIOd+oMgYu
RymIfKRCPPQfHWEViKsMAdtuo4FXhvlOgHPcnVtquM7fUhAH5RxmmjOGCiXRMimo
hRDVN6hwenBEDK9ENq1JpuJqT/ZeJYlquKX2ucGMIgA2HGTX1FH2Fbrr5VgyrgIH
1W3TCJ2eg6EEm4V1KOgy0abVvWpZVXb9DjgBFE8cs3J1Z7NQMTRSpk+a7KkiIHx1
v4I3kS9QWI05JZI+J1dOjsTWR5u7l764ruObKcShZIOgXxfVSLur+gq6q7QyqR1y
SYpv7JuffVu/vXCz1GTP427gQ332fzymb442DtzFrZ9JY4AU+IyNYDIKytb2oqux
c47bmy/2Ld9dm8SmNKuyWA97/uL2w7xGuLaYn6b2EVHvzf1WC2bew71QPJuh0BdE
WEvFU3k9htPKHUDTh40mq4q2bmGozrzD3bT6tdXpkSV/B1x+m5VurNEzsEMIbsPW
bnJfK3gy3y9QBlvArE5Mmsl8pTRkl/7SP1YzDVh16qVoBkv9aLAoiy1E8l7liJJg
p3tdpixwEICQbshLXLkQyqIyVONiXRzZznBFblxF71jhk8k4/mZzaTZu16yGMZ8Y
w5TQw42n/uxoj8NpJOGnOYsTQuz8fTjM6vjzVEZcx2sCz7Q7fFFXytH7RP/AInfj
Gz57iGp5ZYlsvC5Tm95fiHhkgY6XBWeVNM4QbZxzCdi99IEHWRKlpHvzKIGEaSYB
Sreo5Q3TvRCxjhm7mheTIqQr6Is6wGk0onhRr86uZPg=
`pragma protect end_protected

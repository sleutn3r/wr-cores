// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IGKgG6dnYw7WQ69FaeDdxIgOzCft5rRuyACB4EPVRnkfnBVvYNwygJ9pxQAJVTRB
CCydVvT8UcH5KAHqsAFzYCce3+VbVGufGPoKAGvW6OJqi89Ci9KgtPg4nTeBTXz+
rALmJ6V01s0lwIOqVGXOmwXaBebJKQAhHuhqzJZ/3WM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8064)
A16zkvzmsv4S3Ob8CbFHm+tuisGxkI6nldLyqLR9d48CLGEySqQBcQOp5lYqCFqv
dddDYeOb3kJcC98ves8X/QAO44lXtgCLLL2hHVqANmH5QTzU5jbrSRi6LLR0AFDC
zF8mAuvtNAdhVqEmFWAMpv2bA59EosG+eMXv3PP2BjLiDTHR1vnRZ8BMcEVDgWQz
kmhCyvvY+4c3cM8t632aJ43AfUnsGKOqKimUAHa0KYHd2J2gEMo01iiDkhOhqL5k
2khn6IsTmcixf6G0KYD+lng8gRuhZQLS2hGcVBqPI1+sTuU+kJxD0afmg8bzbRk3
6wlqJXsARpixxTPnvm1n3cWmzXjcnunAZtAXxdboL1s1G0b0eO3DTlGrIJNc1IJ0
xu8DoX1WWjwrS8TVEjyFkw5B0beBTVk2hDLnpXA0pI8Rc4fefd80WKUc+I1RM0gH
0YEihYIVNv3u7ki4vyhblS+hyb4RKtP+0JGvLyzCETT9/4lfCNMmI7dXVEr0Bmdc
u+IKHbUws4jjBCRoil4BUTVDRUQ2qVKYu4tbPoDytoHwxaXttktpDhv21i99djpk
a+TBhDSdHO909BwCHSAM6kSCXN6OPXXEnq5Tnl0lrA02FlLKFcsTS1OuxABOmrvh
8lq2PhxXe482wcZkp1ZQ+3uBgsODy9FbpOonVa3VS4KoNkuWfKFi7q0DEvnRefVd
Uzau8u+bvcCWFq1DLMIKNd8JFr/7Ri2M7uM+gVwlU6JaMWT8J9bNagyBqtM+00WC
qmkwtUy0wMSZCGoxmhpYn+z4eEtjMN6jQMNL7K0CZ3vMaJZlJJBkkMov2qkmN5oU
qJuxUeKioqc3RnjLvWrX0mGgPlUvCTuNPVcfyvIwcIlYc0kmHBTbHGLhX7LPLK8z
dMTd5FGq68b5zoTwXRXZg/ucvSVunqwEK/jMpDmnrouWqPNr/ScVOMdiFS66Hd9X
Jca4jGkFMKQfSxQwEauQQ3kpXD3JJwZLIEtrNRnoBAeQyMnDKzQWkuTM1nJQWhci
viWwCPvTLYYohnbfxWendNXXJUhvCgl5b+3Mzrb0Gmvbo0kQmkhlZqng2tRv1MVK
4hI0xGjwWh4+EZsUNikjxApiYKw9i7CDuLjhGhdO3dVe/2I2x6xZHhkLK4FJcZQz
1ZzoXWgZNztJR/jjpTI761RIIbm2/mUhohkPgpoXLHRIfLQ5CW2Ldo2iM/WMk2Bz
KJ4EjEItHJCiK80Wd04KI4BD+PxRia9dvhJMMPd621BK7CwWrk4Ke1rJKwB6+zGn
kC7i1FJyRzGgCBDy9lf7YXLn5Z1TVZb6xauHNzPlMx3XQctoVVC3lodoJ/ZC50ML
nXJ3YSDAOLedC07bs3k2ZqmCr1ztdzKqlYBNyF7REGcyg0Ba8846cJLJLUq5lYyG
+LjbFEo2bFm1ONBZ57vgj5siPumzp8VxbHZE4aNPM0MZIfJYc733M19cJFJpCj0O
CcWHZd44E2troukeDlZKnO1M/+nPCH72oSip9wynCg7IXqQDPuhsHfFfqmx9hPoF
7IEVo6E7OoCvIrXbur9qIuCqbzja0wsShJGmT77ACkB49GplzKj1fsTxYIODQgFv
VXoob3347eKEPoPXLScU83Ip5Ex6h6lxXku0WZp9NLPzUOIKVKDzxfkpS1v2cFgc
a3INHveE9jgG7lKrprD4lQJWoyXPVgTl7FZ9lixfw/erwsvnJFgIknHKV9Tmy3LG
NBbk/3fFl1Qaio8Hg3/7f4jFtPlq5LXTE+KhKvIb7LWKTKPanddGweYmYDXiBF8j
d3mqnn9VSSR8+S1CTG2Oqz25ilHSXZ3H1L8tjVUgpLtVokdMNrVHNnGRZgt/lDFe
oeRtWN4Pz+XmJFii9uWrWWDFU9JzcQtUL1VzZx/ppv431zFdKTc0qMC7NSGgZGHe
jNw1eTqFuUeFTokJ3mHxfzvyZ7mrgdwF8YlNztgbxdZvNSHBt5JEhetA9/I0quly
03wVlGSv7JsLNKo23gBEtdx6Hiv+AMBErPmBBY+VVa7glAKlJWXAjzlwQS7O+AKG
fkWXsSGXug9k0yPwC8EipkRlVNgW6eqc262UjxpcWedYpjGnONlFVvJI1eFlvhod
jVKtCNDLHPe3fCCq1KkDvg4K2yU5DTAkoTowI/4Qa32CUnvRSvRwRy1JlvLMqt6J
yWQgcupm42CMo//nORMHrtB4RbNZPCkwiHdwUMU9DHC7+TJBw7AG9T1u2ZZRGkvW
R/0tZ3tW6hNbC9o8Wd5LXW31GsVph5EpJsgPIkujs7/a7QeQgJ7GILDUfmQ7w6KN
McVD1RpYf8cCEVtai5uevzX249J9gZ7ACdkh6ccUqRt7OYP9JmF1c9/rwPS9YHhZ
L3V6mF0rChzml98pjV986M/uHY8sNQjQ6jx5h023NA5yrElkgtKpuxHaiPotWPrw
TAXtto26+1OJHC9WEE2GpvDbtHsIR1EWGN3XWNu5P6EQBrc1sG3QPLOMylwS81qV
SWpZe/KKPTySiQzNtJi23Y6HQSqtq2D5L8tx1Y97/2mzrNaaAOaAdwxqC4HnFhe9
Mn5x4rJEjBedqbOpPOaqXE7opUwGGi36Xv6PoMcBoVty6lo2zDJgrGTghwuBjBKY
yohyNvLgBh93oukB6/BKX/NSeXRag0gvG/KyF8JCJOpBAkjWL3wNlPNToze8qwSQ
9zFe6UWe3qP7wfgxZBoMMZvtw3Va+RxLRwuJu97MAZI2vMXNJUco+hItygRcFBfV
sTLzyf6HBINa+wairwmPSlwLJR1/4qrccgLq7pyWvYShY9/JEUdCl8E9Qd9owKsW
C9tt0dvPb/szap4XcZuCxGDqopGeF2xRdEQpSYA7EQKug1ZAeEtR7KxP7PGg2/k6
bSg3vP987ybtvQSF6wslHHsbN1kTrG0z65MBKys0Dkkiy4cy5XolbmsNUYNBI5RC
4iw+L5f/PfHetU8ZpSmo+k92RC9wpcM3k2dT2tFZbBvuJ8MflQWoNBkwnB7rHNNv
ai2Av8eTIB1FJsc0sHmVTFwbkHItC8lG4bSlljMEcUkEwiljwPzZNuT8Unv9vUd2
/d7gGzHUIOO/vCLhEuyVfkVe5ZGU/6pJbhBkxwvDcQpeH9l8EV1y3bBdK3VFlVCq
JAByDp4rqxSJ9V5HmZfv5+5RzrGd6cLidd3uUBrLJsKz2tK1ytPS+o2RHA7lUWA0
OnYX30S5tSWi9nPVdBW+vud+3U5vdUbsw9+hKsXkIku6zDFTOoJ56JG47XKMaOgl
L8w55MACBHUPhK+vj8VDUhZ/tFcRwfBOIifu27D4rMqgCOyQCcDBkTp5jqgzw5vq
n0RRmwYbfVaobrmFJbaZEnE1+HKmL5JeVRSfsEVX97C5X8nrnZSu3DfPhmRY3Q9t
Ll7501zRTuDJ9WW+ldHLvkD+y74IrcT8xasuAYP5j3GDSyNh9V1Doge4+fiWZ1i/
FgkKjrE9QUATP06IP0Smenjl+T/wJeBMPZ/L+UiajeYXdrfBFjudMkPhihKnd0eI
ClNtzivMMRLadKc/J437HsIQ/ySidqpRe57O/ZAu0IbfefW3p7uxhleLxmCg0pmq
IZWB+DyyYLLYL+jTm1vA4uz0vSPWsKZRhETDMkxeF8koJKzAD4+c1l149TkfqGG+
PHyFFS+tNONHAYQ+wN6R2kS/ONk40CSh9VXZ/rEPn3V/CU8qa/Du9ma5eHAOUSiM
YaOv+7cUQYFbcY7hkUNVvI1dFPnxljXehiPvs33JgscG2UFA/LMit6Pn6bx2cY6f
PuPMMH1k68aj1Hm7dB42h03AsldYcaR4XAge2wEazaySajwmc9ggThXr/UtRlu7D
QGIQq+3SGF550BRVMRHvJCa/VTOEuEvsTe69JbrcSOJvLBcoaYIvF12N9apqd8uv
MlFRuqk/I/65nv4o4Z61bdi2XXuJx2gPbgjN1UBmvh1A+C6yL5yFgUvgzYDuOffU
8OLwVby2J91hwr0UgIgcjhi0JB0+LJPn4wGg6+jotlq0GPV7wr6jTybgm6E6R2+C
90i4Bg0S7Pq24RcVOMK/XwxrkAM/aT4HxTSgLtBLyULL/FCstKc/1dE0fQksu1Eh
2oBwH82ChbBIe0I95HbAlVxaF55QL+PR7ixmuvUVUkKxT3AEblxOjwUk82SayMJU
F1UbeGBHUTf4E1ajP48nGYgqNKZkkn2b0y+y50XTNrsDbh5I27fIBgKKvidzUM1c
0SAztTop7rpseUr3pNpzuN/KJjbZwqGGr4s1rXxolicyOMcx00VXaH58yM3bF/9D
L4eD+G+ahzB+0RMeibhnlIUKVA24ZTYgkorUTM/WcKkSquEcNLvZSZ0e4UG9EfHd
wcsPN2kmQz4xOowjrOAU5q34VLwvJaFWs7Krtvm9G4XZM6viOUtpDajNHUAhOlS+
FIObAiOB1hSi+rbK9qvGE5TFo2WlDDzwrEclAMIx7ZkOjmMWF4tcOLEIWhnPWDN/
8N9i//uMTvzfwsBGcg3clNiY5YhdHBidx/B/oRO7olt5fh5lc+YGu+3TyNMMczng
+fJe0bECc87Z7HqtYr0R6vGhBqOsMfGOhhFjJs8gh/ve7EmMuv0sidDE7D7ZPJpm
ypPhZFL2w6vfQ9ZaChta5uuc7ZH+Z/rdnSIM5nmHQomyH3y50e7mMZi6mA8nrWo3
LDkCoCjdEwlcJ5skZgX2Yq1LHhbdWH4GFfN0BP2TtT7XygiX7SRpn3bnTNR8dOYU
EQXwI6JBo42oAjbhJIwqa4vfjOtHccv5JqSolNRtdhAB9+JrUPhFdfiJMZFiJQfx
2M1qNtuTyTw5QxPmKz0jau//fkb4G3tQxmoEJ7Pk8SNwzexSD7m9TGK/aHLxKq2u
gk9SXfSjO16rbyG7Pgg/t/AWKjNGklh+eQNuiYCNadb7E6Bqd4ZrfFKa0YDHuXGE
mQov9tZon0o4GrUkZ1bPizVBmhmkQRb/aTSbZsPM2KuDYRnjDKoKQxLggbPDh2t1
Kbd1C8xVlnYIaaaBIvcHeLA8MtUwZtg09ThXAR2sk4rxyyqZjeIxD9ryN+WzYeF5
3wnsY9NH7/pJnvAvffbjhDvJeYBNO7wEvvwm5r3R20/aI61FTjKYm/IsR+lwONUH
wC81Xg22+x8Md47OcKMsElod5F2OcFNlfvLSiEzpQduI9wtt0AlE6Mvv5Gs3L3ij
pToLJmNX7OshIck7tuhFDg1/NPwafe4HJJgJR4B1cfx6/YyBFlPxKU9vF3ebAsxp
JwDb4/qPdXZX7tklxoeSbpgMX3UzPcBf9v+nCWzZ6Qaie9V3enMWoOezIo8mzMMs
70yOeIDofkUbTXD+rlCmPGgHe2W+gxVQe/LTMTisHg59kyANsmj46lTyjSju4KTs
FX1xfrIF4B8IRVJ50l5nN3mL0jRLk/n/3+ngIWrtWYWQlFoHXCqvgIjbbgkIiLxg
t/fwor70ndcZ8nQ53uKS/dQbx6vpfNmT4IwaGLNjzm7phsSSTZJWrCh0Lr+ASV2e
57fgInE0DNDi8oxhMVX+mvkYkJc6Zyvi4lA4LelhcSUA1njA+N0L7XXvpherFUpy
7+PBHYpcg6Af7HrZp2q+Iao549ZR8GvnKs3mWBc1qUcz9hapHoCufzWdP3xr3He8
jsHEstB9UBY27PoKUDxlhvBsyRcz3mkAwZZdw3pFozLYP/X+OhlOi4tLxFoqZlQ9
gLbXDuVtrK7Mf7ANgmqocqzNUwFlCJW4eB8tpTnGXEQ0od+i7xJ1ecqACRtDf+BR
FEXB8Nlxx3MtinwSPkMvWwLP1FE60t1qpbN8IadcEsLCkSbB4qVg1+uNtJR+zKBA
7cl+oPLekQlq+OJLU1INsKBwcSzenjevcNc59YVgTEkbkiYF5czMCz7hUMG65cI7
kNvMeJ9GJrrI3NPydHeq8ZaAhISGqk6EPgxZJBCk6MJmIKfSy51BfAjO1OfeLYlq
LjQHUOP+2n1t4QHUzmFmxqqcsjxEji4AtymTCZ0XcQU4rT99EZcbASnNjA0UlkSt
8Ioapks5FMOj2NjXUx7NjI4McX6FTQUOXCe0Pa3EPifCow08XCzxF8KoHEPZypEa
y8IzauBYxWSdVh5oFXAazaBr//cEApuGL2j7B2U6n4HJV6RERPtvLoNTeb32KQ0O
d5nDj06T58ATp2iH1zFcC0oRkrwtIYWgeFOQaISYM6O7rnX27L8X95CzjNEJpINN
xQo49SNKJNYDLSbAGmOVqyWPmSqXzkaYfRaLcDya5Rcn+6yRPT3zYFsPGHcQZ0Fp
RV0EiFFtUvY+pvEWkqHy0EVW0znGA5Fd5yLJ4rjOxUxV6gfoaB5vfQ4BpZUdBIQ7
w+awddpZYgfL+ScvikbP/iAK+8OaXPnrOpO4UAsSqkyX1x49gav2Bglp43NOYBSX
KkQhOp/gUfGwtUQiXBpX5Paze4DGHeXhdyY+vy08k7g+BUbn0Sm2gh/VRGEOd1lh
rOBV+joiR84K5bq4uxDw00eF37L61k2uYnCI2H96wUOmjdbQYe2FM+hplxVG/Ao9
ThFMe52VtYCpAPgT37y/k5tj+Zs0fVLJmiBOxEO6u+yr/434uvTZ9DbyDpu0ME9k
c/8us3txgyVfJaFDi6Q/mXzNAHwFOke1Cx6vFYuZ2DVeAzFxjPOJMU1c3XlOXNm4
qzWtRpcF/3nunGkMBmnWHLed8dBJvRrOlfQWyt7D8G8rg/HQOjKDgI39tgS2m4+k
+/indrJA6b9KZN/pMA/9w4CF5odAuxRFLDmllMbGDEs9jVfW1aLGxlV0o4X0rePJ
5pV4lUxj4wDD2gTRARX9Dvs8bghqYzJONf6jtsu/wm5HDs1Eg9wXsyl9mPrVeF9a
YQ5t/0FZWD6GLiQOu/xA/NkLoSfKNkFT6wA5cF+bi3FIikjkyLXiBBGCVFEgPoNi
jKeCSDVaqOOoaDoPZCCmCTZ0ziYXrRm3KC+Pc3GMFBAx50PkZA2VeKLZyRFyoy2g
xpeZqMHm+av4otaQ8G4or8VlhMHQ7bY/MVmYPwWXUz/X77fS3siaI34Q30A38s6y
cgjXZDvQfsGrQaUd73g+mHV5w1Qjkd1nHexvVqlZ+t1gY716yA1xorp52WnUQhUi
6C4FFyyHRucWOevB2g9WnzCJd2PJyl0CdM2pfPV0lRpK6DIHh/vEk+ErKzTFvZQB
Duz6kHF7Q0s/kFKJqb1+0NF2kVMpHF8tEtLBOvrKf2YGry0VtKcBWl0BFU+2Ecb6
ImtAAcwT8/dBC4qJT7rDdP6h1S99NlP2Mbz6HtWOlx9WmT3HWxDhFbL38DbZabBw
r7j3wOxXONsrMr6lm0V+o7rWppXdI7ij+Uqku5hMCgcs9qu3oO1I3cLorE/rjtuh
9KM8IKt+zD4dtrJNxzmnKs2+K0VV+hB3ZMUeZ1bCLAUIuWJ44SfZPAmHkSgiLHG8
+YAB7XR5KybWKfnvKugxs2fxv4f19rIoNAq8ReRmGeHN7jFKV0+BH5ZznWs7IGmv
qz3fq7NPorJAKPkYxgMFMT2gnX14MUlwi2X82h0ApPvScYWFquiDAHTWLChrfp32
T1F7c39fdq7OGLWr7NIAeqNh63IafGER7ac2C+IZ8C7pHUvB1NIxlCSWYv8KEyun
xJXI6O/N2P96eWWq12NNH9vHIvBsquSJP2jBLnBqIEGUyY2vUZoUQph5RyoVNOY9
sWAXQ8Z4bNP3dnc3YlCFYLuLN+X+M4ijWHPMaCDMJDkhqXB5V8XcvkNmpQno5bMU
I31LJUG8q0q0jankOMXE6hrDZC3j9kl53B93se6jst98Rk3TvLQpVHWATw61xppf
Bu2gmCxK/sStRmiDQHfN4a//YEPTLt3UJWgGNoB0OQD54kz4Mg0fdJEtFocIyD9b
oa2Y0JGeNNuwdXE3CUJ4TPcxoMo6nnyr/h4d2ckII1GeW30P1K7JZbWydkLnPwfl
pURj5opPZd+91fcGmn7rN/YiP38yqUEAzKVeacgLfQrQE9FkuuD+2ojZ22ar80fP
uPBWpexSE2XFRYCalOl5z4JlmTW12ctW1y7F1TgdUd/amfIXVX3l7Ln6WtsoYD+f
gtxtVH4QrNtvqUYNe3sTYJrRCPhW2ZzT4FmmQXO1HvQWJX2/Pp0Cgj/R4U6kX3AR
0SgoWuhGFC0sI7mZUm9CR3NKmqCTgut5aD7ISP+rAhItXyQcFmPjPPOhFzLircmw
wAeZegghZ5UGyYfOc+u9uQWJRdUteT4eo0yaPxsXhNtYyNlHNR8By2y5NdV9McHv
CYmhfbQnwBxoNw+yZHJKLo5pKqxBOO2J5Yv4n720KVYnBIWEfrVOpuWCnp9Du2nw
H85AQuVVlTjOhOUDUweqAZiVzXxkBtO3EElMnYhpr70VSL/42oV5fnl/ZlEUqkeu
K2O5MkVFwiW1N+kuMnCmAoP1gFG99DRiUxsLAGE9aX//BWIAsQGCJ4EqFm9LZRaG
+o+AHK739F7kmaDFCyiMTmSJtALQm1wUWFzRAKGUmYTnpYA1naFD9duQliEF5QOV
TYe1t6UH+2ZGG3siTW5oGqRuT5BvA9jOw6pzBu9vLjhYxGNhcCWIqwEwbvndBHeR
CB66+RhUr0X0izOx9QvKSu4iz2IVKlvQNL4vUiHZxwMTAu5W/K+JptxerGOf1G/h
v15U7eAFXpQGptc2bcJMjSH1YiulN7rt379KgH1lDVRHflYRGhrUBob4Kdb3G4D+
NeIHJOMGPSmktgoCnUuGGh+TLz8xbHiliHYpF2HoryZ53aWGqrHrIxFdTvx79Ays
W3arsdTPEviGmAMo4eUyiJ273oglVKWQDA4c0ziHQ8F+G88M4sfVTZQjajSYkFs2
KEooVf607RvYiY8VohE0oU3QYLSHHXGZe+g4uC5CpGfJB/pm1tweTJqKewlYg2h3
cRGx+FYCRlQ17fXptEPz8/uNJ5qdjRcj1W2pRpkh+EvZwubG72wiMoBvL8WEGxQJ
2fOMRCNwsMxNglrGIVtuRYPykVy1J+vunWB4TFm91rIAMxS9aFuh6xNBIx5sachN
8decoE/HNxOyXqlcVo6rbGZ2nVN/mFZfTDci5kC+Pu0a12A3dc6gqjkbkD/p4T4m
+S4wKHGdnzahMNJIKgRLZdcNEMGry1+3EKhYOtZEBQ3omeq50FJbe99feOfsjgNw
dM26pxCSPgAA5JkHlgu0SZu4CifiZyKjb3C1ojhYDc1/KIZ01u+zsZgurCVa9KbI
odwKDB+g6t2g8fJJ9r52+G4U3J9fiZCW8JBlCoKwBSfiY+sdg26CmXiPyw6sS/kK
WcJjbfebQosLXgkHHE37Z5WBecw5ryTIYU/P7LmQl53RqqPBDEFxgcCI0RxSNGbb
wiC88OBcEia366/voeNNLCGq8nxSaCKbdjFsgquPVHZQOoeWMClxLYBGwRG9lbSJ
v12RzyWRAnwL75BQ2icPRC/JPB94iZbhNVknkJ8H1tqjoskoZdPNaZ8710Bsj9k1
9sN8op81rOTYYtHOXNXW0W5sTsax2JiscUuOct2vShnZuvrrR9ZlJOWRYDGl06Ca
QBme9UOorqs10KcNaLxKhblBvviByp5Ed6oNlUCj1e4H3+1v5eDUcfmSnEfoljlX
0ozmvSaifJhH0hlCvGTpyKhvhFANB4f3eS3oMaZaNv2wD0oTblp0scJ20iOXXOZ9
otaH6DaTjDoAuVlt7fcLfPSn0WMdeaWlrLOeGejvfSS0ivn+FSekytiWyjqpXzrX
UL4gGrkMXBGCfiBOsGkbH3RB8gR3t1YhTh6smF5rfkE0t3Z4DCS30qWxaRwhuMzG
1n6LXurYjsdWF6k1ZCKQvDENw1B1orQc44MANJOkTf4eEPQD0LBUjbm7I2FNcM8m
V9oTcxKdw41H8p9meVTkIOj5EYGhnhxVw8hKSHFvJlT1QPRrarH7f3Oru40t+EFz
qgd00SxjJmNQxNGkUMyQETPNuRJKEprHwe+wsCNE2bg0IIzrIUEDq384pjk1kWdy
xotUdQptteRu4bwXoWd8Pxh9mqvr/2uGDuXlK3Lr0vdPW8KaafyDp1EgFVjO9UOS
Cz4ylp1TQJyDG7OdF1vliBpWSBIW801LKwZ4j5LrzP//gF5vnVyKzINfqdZKyFky
HEPX3GgJYKEjXRYW5mGFoejHP1bcOqWF1grVaIqEV6T04IqY+AND2Nljq+3Sfz8n
6C/vrPIp5C5lkyv9eCUQ+FslC0FaqT1mabEK3A7rVeSUBU4Bbk1Mh+U9vxDbkXFS
zhYHdEi/tbni1avABe1YHqggmAQIEa27r8pxPlceQK0EbC8VHIFpjBcu150L1VP5
W7opmsboBSHEKypellDhl+z+LKnCVL5vxgzSbywp3PdHRurwVrrkCPyALSX7kOnj
DNvP7Tyh0iAZH2AiYJNN8GSk0nPME2+iNaQjZjdSPTppQ3DUC+besPfoBkXARtNf
eZzkIM+C+psS8WUMvxQ9PD959BORdn3V/zGz21vljST5qtqeMZhOdC1PiNfAXpes
9O1iW5X1Ob0NJW8ALszeuKCjRtCiFz0HMZxKctKSlaoyr5o30CFv3mPVV1y7712+
hX1HP/AtKsX/t6+nMJ+g8azwfZlX64O9F7Udaj4NDzoCIuLX5XopVGyn1rxvxerG
sLjX3eo+NROKhbwNdEdWYWmZ+1oSWeckS7HEYZfpA0aUTybMyS6ntPAKLbEYPTu/
Ws5w2QQZuP/k2ojn9XyW5cGgo5y6BbFyJGwaSP/tVInVpnqEzwsTtf4vNoRVcHMM
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
h29pt6D8wHFUNkS2v4ij4o3fqJECyROETGNve1eKn/6RpsPQ9HQT325j5jJa9EjT
bkhV+ekVe3H8OwGPMLa7LnHznJBdJiuNzdO0Fbd0wHf9bcBc2qfCjYtqh2h36Zpz
/FGzgSYWMBHYDyGJ91ycZy5WmnLpCB8ckXIo4FUWYsU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27600)
q8ETMr/WBh8gfBAo/H6GDQlMjM9G1MhS22nGCJvY68qAN9iEP0bKIJEhZwdltpia
F10oWdWC1/h8Nr2KycPFql8C8zyK41jozy4E7CFI8IKMZl8z3TWTubSzw8xyujaq
XS4HyOnAUB403RI3AKLl47dEUxpmTtIagishoX87UmpGTv+JebZzDqUf/plsAlNJ
t9Yr0+9jGHl7i0u1NB1gHhHSCVuxB+uLd0A3SLWkVvFDNNjIfj1HuyVaPH+sI8mQ
iUtImRqw0NzNMIrzrvvGlR1RZ1bb1BQ42tg8/5slubT0thhwNeQxmL5tgWNdVWIp
XSP7sFHYDp1WFkUlsxwerUsKoU4wP6bqh2zzbcV2KNyDeElFR6Be1ZIRj0FCJF44
A68ETGc+VCYjmOMcy3BPfMI+Yzyh4H0VuxNfNqKgSz9IXaascqdU7mKVtEHADAnj
BZ/jE2tw4zp0Ip2NsrXSJgnVyBpu8n3JwuaXMq7e19k5YdW+b4hXHgb/C1XJeE62
cPkiDjQ1/HnQOlUad2J4MTNXowwIOTb28UpXc4cZ7tKxDaHB8nNEg6YcDT15giw1
uaqQibqKBRTLo6JMc5anKBL9sWRoO3wqvU8vvXI636G1DcJKmbDueUoVlE9h5fo6
9mIKYugJXXVgrCurXdV+FasAsFzri2nG4kwfGmzLreWhL03GM70F/RUuL4iod4tV
2FCkV/DRN4FfUtjJrYfYId+bi6spiZSarIyg46PSItnWstvd8BOAk9+MGGV24PNe
Kniat2AVzja70ZFALWpdRfiztYoynB1bjqa3qt7B6ojFloEmlww7frsz/fLArT+K
9oxf4ISBZ+k7qId4Lp83JtubSQcyWWbSVgekTT0kqg5LUuwt0WFp9KxmT0WUsYJy
p2JYj9MsFy3Mn3mFsEGcnVCzzn8aJjXcmMK56VTC7D+jr7FpfDkPVVFEAQ+grYvo
MJvRBM78SJ9NKC5R27PihlVmCJR++3mZvuvFovkQKcdMXm3CdOrcfvxV36WfZDyx
UNZWng0fH9JY7WkDZZsquPXo2J8JfDGjpzDyveanliNWPxMSVH/l88dX3uc+xR5z
/JXRKVGnnTfM7WTgVLm6dSE0akbhAUx7E0zF0zUghMJ9jYoGsruB9GS68Zh7NIg7
Mz2VL+WGjrnmcmEYk/PVJlTQJDm524ZIts43hVizF9HFVv8bPubqt5GTXjmff51x
7tk+9Ie9VQ7mIlao8MtXTlqkJhX0KraKkUG2RFap7somVcJ9+5qLIr6eK1J+/YKl
JW1RkF9+YSE8mkGbhcPLIT0M79kcPS/TXZzBedKgO6Jew4ZyA2JyPNTsCeIosPA6
xc5J0RbsuOzpuk/biWFHVb/fmGoAGap5Lhr77vKRv0UAHsnckRqEJBtRlY6P4NzL
6eRJXeL/EZoJZ6dsc2LwHub8cDu/Lip9K1MTqDy828EhV6exbEcdRJVReTwVYK8o
V5as44GpmG+RwJT/yY9gREHZIOiK8F9FJh9UVjogVuUdEhKXbGsNn4WoLV9UzzRg
O+CSdEmN8UcbVJBFl5biZGQlFiF3ZnFaNKSVSksziopgMLdaQvMDHaYVDmHbjs9j
W25rv6a7tKLkz0A2KSw3ta1gYVObV4kMbN7cmBZMYsODHdUTn0ma7OZSLTHAX2ho
o1n6PtUiT1CishFq55V95WSQ4GfS2+rYv4hvG2C5X2yJtHejn4A6ntcVtYawelyD
3B6sVt5c9KTTAc8Y8ayA3WI9/dS8XSiYxaI2S8o5tJ9x58LCRmv0j3pe/XI4TWrF
jQ6ryhnzyr9+/AdHWg2OhmQlQh4u/yxe+nUjwvjQ0zZSnav4F4vXqP1Q7oXgKrYr
AyyS583vBKTm8lWA/0hgNoG3VbJPYe1GqToHFGJY/wzSxXeO68wM8vFpGoBBLfJf
8fq4rPffEXRU/SULz8SWmN117aH2mAzBExU5nQUD4fS/XLRB0scS8DBCzq+ISZcu
wxnRbCUU532vfc3K3IgFVf2NHFT/t+oxTDtB/36rdtvriXzOsDq6jTfN9Skdk8sx
nrrT/Dp+ibKs+8Py+KwaMbOaEIf8KzBt3ecW/0FksK0TIaftv/duBsBx+8UtBi6A
ddWp4KHaCUneXMUmhSvFzQ5neGTAt9hDIoVTQkAWaqxmzZeiSeDURnoeJXcUS8DZ
KTT9qinhibTRP7KdZicdleVHwenGnvuRPDQW6/REWB3Upq5AVSSQxBqWHZYcCvOJ
ygwTN7ukRB18E+iZOASd9Ya5LXbIcAi2riJGYi2MwidXXg28nJYV5/dagPJKDWOl
BQmbgR8zUmMDVNhNzKx0ZdBd6wv0Xo8YterXbq0+LiFtuqTa7qXh+jXiICLYcRL8
7oKNIa4HH8emgCfS3qL2ITuT/82C4IR7YZZ/SYSwKPhNrn6GgE7hzYjN1NJZrj6O
roIGzeUl9Nu//jxUy7Gx2+UgM49CDKYnGqaSjjLyt4vLQJcTy9TYzXzjvRycQOwM
sF9Mz7u6jMHABruHl5num81sqEhs2Z2cFztBAGjhAH+/EyJr5E8DA9/JeB9NcP1P
1UvPoWTrzPezvQb2LTAAyUve4xARMNgotehtuBjk9hAbCZYVtJcf8S3L4IIjphz6
QGV8sjBE3weR1KRayhlsnf1XmVCqbnSQ2MAwdTI+/ICIJReyBX+ghfsI49ZnbHwf
+kZn1p9Kzzokkn7KTPvXF9wTmY8dogBkN7oIsg34Z4s4MPuq/RhVuPql0ti0wAsj
4WTXZa8SgPcKQIa/SOsWR1/qh4u6up2c/0HgKzU3Z0NTIyEJHLbFnRAIRvNz4L/K
AOOi0EWU0uyOzx6LAkqQS0pIkiAzziAJu8KY/YKkxfd7lP4ZWMLI5l5fQCG2fw8K
pCCuEHFzy2wXmjrH+U/b8teqHRl+GImlJmTiVU0phcudRlR46ii4mSjqcVVfOUxp
HZK+z78Cfw2cMb2Bu1KXiQQ9G11a7BBMbIjDdZJ8XUVmcTL+Tf4ApC5H6HZcqfY0
684xCwzdN7iS4DIq0U4d6F7+ahDSZrpXtjRzZb2NsbGAQpsGBgMPOMwVlxNzCMNy
I8WOUAYwc/WSVfA/x0WVlT+25LFDkupIgSznB3DQe9o00Gt/+wr2oOr9I8MB7l3E
QBNs9W6ZYps4c4IerQq3S82fcepgokjblLiRTJi/tHl1wtsA7U+2dsNZZLP4hra9
ZVrBjTzM+batY1YicC0rloQ/bXizYMNwfCo0Coujsg8cE/VdET09d2lqnSJ432l1
O4ovvcXweQLrj0vdFmSwEFLE55EmkTAthU9F1hHjk1oh03aTEzrKDMb7IpVkIsCC
rBcv87nG6rh/V3ijof22wjQvAVBTXCgCFIW/8c2Vbfsav39F0+x5nQOfD5q5Wjtd
xJUp3Nc03cznMhAyGyRUkMlcJb9LudvjpVh490g0DS3E+CE/aJjcmxRNCMXiuM/5
GrUx2e09w+eHNV14FY1bDRdz+wO4hK4YWYbL6nrjjEmt33TKRZtzx67iz2DG7V1u
/kHs5KsQLBJaarb56F4VlUPw9s/or8v7apgJMwB82p12LmtiPmRyehsOQpF2cEBm
FUDBpgGdFq56fDE60hzqWjI+lH2SJyDazkK5x/2EsgqHZXFLtLr8TshaPqAU+yiI
yK7x+qCgkXPTeqdVEi344fqbdfRyH8S3buyG1H53tl6/gWYL8mJPqptPS9uCLzxV
/e17sEQp/Aw4U4g/ENmux47zZPYfU9sUMn2ymlXEG3yUfeamB/yogHBsVxmHZhvO
C1p1/gbMYhtHlFc1a78qFEwcjWqtsA9ImGzjlGTHrwZ0KXuj5TQLz+NMHyvtEnWP
PRWY0MJ2RPM3YWKmCyg5EQpDbadzZAFCfApR60Rvwa5M7TwCNEf3b/69vgxzvPUO
KMEOsYkwjvMPQFAGzgcVVP8SwLH0gOxJ7gQlRsRmuFH7Ft54/VQWr1Va9QLuDqZC
jmFmY7tLcg71iD0VNN3+imnO6WG1kp18uqOLD1S4fUikP3sISMj40gAqDilYrV1q
SHvaYROduoQBvS51v7AlivxNScaH71e22+ffY7QsOJA3A3pvVRqhPFJTSc6JveUu
JgGldishcMjMLw63ga/ATJgajUXulWtpgHJNEM/ls4Gta03JRyu5SCpBcuHjgqN9
g5gkq2A/3fgqPRR1El8R+l5TmsI1MatB47oywqfBHNLZfXduQJqfUMDIicSsbkEx
XPOIreLiHlggaWggVVdTd7Swiur9EpAJ17FJBldpuIj0mlrVCPtHxjNMpcpFBP5K
Y7Y7ocpF/ym+4WMwaN4tbkmXy4UnwN3JyumSqgY1t5v55lcB5AJoLqos8u3C8F1L
VgGhr2lGhlmuDNJo4UilQ1/p6BNUASPiZaHMiDwhuR2pvHB+H/Jb4IRUN6t0KE8Y
X3dQUiASVEYEbK5HUI84WNIZVRQj4kBJv+QPHJVgHH/Gw4DWztP6ZQVy+So+v4eX
rKOFAM+yXosW7cvkK6CLLLPPlR0leOY+87SvYFfVpnmrLHFR5KLbHrafsZxRE1eS
ld5ABrdVr7RZYIunRmXaHhfs8mMdCCdTBPROrn+WjrNyfABtyhvWzkG9cJKp6gCs
KQ8CiJEosjDyRQSI1O3RoQeyTj4eNqtsQaGqYcebbpVRZkSh8FevCJGQgT5ZULzy
3t8U2dmBFLvH4C8+bmmWg/EP1dr/ldDfvddrBjKo3jycv/5BkRcy08TIuFll5Bvl
6Ok/h4wRjKce3feT+YSEHGuqTELRJ1x9Wxqo/kZ0/Uj59Wlpt13GnCnS1jYnwqaj
q+68Bj5MwYB5bUc+ga6+3g9OUls5Wl0TwXzDyga8NoTK4fWQuAe2E9zMqyaZIgUq
XL5zo/X2in8lwAU8gBP6LSevIRWYIlZ3zNpxEeMV1Rf2IZDX8g2TFO+dSmMYHpIR
itZXWugm6tjAaxpXKxq88nbeNr5OXRwlk2xYsX2fgoYVQGXDshIxxY5wLh+HTuED
Q7573hJUk4I+TScL+l0fyvyXTkU3zZSuAkxbp0L1IEt1S7426ngxZLGs512e1Wmz
vq0iGT7glIbDzRpxqIqQFs++nwi6MejUJIyHJbYRtUDEHdtq/yjuRkA/n8xA0UMc
+STTkAxNfi0NdNqESQtjOdBDxNeOGFua7k9Aqoqow2zfiz/DpHzZ61sIjnB26DzD
gQGTN1gxmIZBlX86rU0bTFcb7v4lFA4Y8k+/zYWB+aplac68vVqaFVKW5hbNEqwo
FBo4nE1Q4K1Z+khiRGmRSk8AoaaQQQZbHyf+z++jKHX9eOvPhBsmkGFbkhiHJUnT
M/WK/hs2g34lWEzNzhzjZWjK5+/QSp6QLO8qTVbpzSsix3SMj8oFhS93uvA3FVSo
3R3s1q8PxIq7zIgcmQC3aB4MT26WoAKKjo8gOeTaOphFTerLONPgN89NWd26OsHf
tetyc/Qog2e67Vg+dgsHA2uQqgisCTIA6d8ZqDB96CanzQkaug8OdR1bLEERd3YV
PxBkVjbBVN+ZxL0epHGqqjpU/Xj+xxnQ85ZlrTlIgOLhR6+iGcexf7BGUr7gmb76
VdQIGXiv46mOrxsQHUzxQpXBAlxHMqlkMeaqvPjpyZrgruOMee/dPUAv+dj3iQYG
Kx5Sjzd+4G0yrEKgZlHjgpicwfM+Lv3BQZ5GZJ+sDOva2pvWI3jIWLwliftH038+
dbyjA3Uzasj8PfdN8DX5G1Sw/wOCGUBfZiFzX9hjCgHdKJx2aGYZrWeMn/nl9NFx
/rXF5/FMK+NTdzGrwZRyFIjKbKGiIhk7Ttn6VocW2zBb+fSSDhyk3P+3yeNt/RHA
mswxFGIjSnHyMVuJXMMbtJiNhewFCsze59FCDDDrSzdG9M17JDoLys99quhwNPgX
jCv0vvMrsIHf8TctLDVzbJLAxQ60vWB1iSWYJZWuintsenggd2LIoQUUsb02RO0f
PWwRY6OwUgqQKaRWhSn2OAyGgILUQGgJ8HPpdoBf86IrZOkhjz7SlE5dD2ybeF61
7ABs2cwItelay669oNFarshKi2zsPj+iVklmmnYnbjaNgy3rKI4V6euVivLBs16h
yO3HvRS+WnfhOHgm0MGeEZ2O3532EHcfsHXm6Ss4pnnFqZK+GoD9VWuEuBwPIx2k
3zP/mG0tVmwAOdvHbQntemQobmc8Ty0zfnJojGrh4u/MWg8LpqP0ngtWVRcYduPT
3xs/HLU9ki6yHDAXrmr4F1dQuZzD1KabU1OKBIibfSSXHWDp9gzRvvEMHvuOFuBL
6TmOGcY6JX5hvpb/hkUlk/pOcGIb/1vHsDWCZeJUOKJndAbX1pYSZiOxm2RiVlSs
oECRZtzWEpQdHBvxr/gnmNuWpSficZYE66SSejhH/tQsZ+lO0gOKosvaAsQRlWY3
hq8UZOj9o51iFGJEJ78ZE15cL09WO9KzPJzGX8XWZbGLU6jJPlCC8tg+wN1N3R3t
nXLnXIs11f9ubhf5agELwHLnzOi08km+o4cVHNwUX3xa6ySGuZkXHNEqq4Ijjvjb
erXMcmhj4MlQhZ964TnTqKglIzU4SikqmUpteMFE1OBhakt7h9eZ5WtZvXI6j5Wg
OVfM64E4bkQdyw959CC4krjFvL7LZm8E40f1lnHoUq4u+hhK/vmnQH++ocrMfDQa
bI0OjMc1rUOwstrbSTlQtMKdp2xOUnXEq/k59hqqNuWAOJHWevizIwAt/VfDDQPq
bU11bcFr/bKusiywBQxRI4osTpO8azz57skgrhl45ROAj+qgsJ4TE37Y2feYbH0+
rceWopW83foMaVyLe68aExNwJbakTVRijwZzp44PhpUYIxm+0Jh5K4nl7eitjnoR
PbAWmEHw31Ly2k8iQSqADBkCq3/95eOR5kB6hgTJGmib1Ef/pqGy3Yzl06bS9kpY
tmlkWzXcO1iToQtsuJs0oCb1EE8uJPjnS9FlViLNxxqRRfgZ9Tuaot2SMrYNZtQ7
g5Riad6xtWBYEHbC3W5muhUBANbwiIF6atTlNT3vkid3f1b1672mDGH3HUqQ6gt6
NFZS8OKa7c7Z23TZkqbaZo8TvL7sW1zFMXmxJQaxwxtowdTU9OdBV1HgBlYGnqUN
f2X448zz/6qUqkV4wza9p+4mzs4zgMAdYPGYqMC+TOgBY1jlk8LHjJi9+fFgYo79
YsJ3y3Go68FCDoAmsOXjDWEg6T38R8uXOjJQHgGujovvEDbs6/g8pxzGJiOPbeWM
NHe5jSfLMHzq+XV/8VUboy8SmDlZN6FPHlvBtxsxYdCWzBbc7fm2RskamAdXQe6G
Bd6svMcd3XjkcevGsgwuFuJ/JSI0JWQJETNDET2lhfyYbaj+U3/+U66TJ5Xlg6Xk
L/vVPsvmG1JTmbQVL/HswV8j1mma6hI6L2iBmX4QyHLOWkYzTcZNUhg1qex22GEz
kLNyLLzh/gwT/FDn0SkzBIw3y2katQnRZBQPmfOxR5eJzbKXxah42lzGPtO2ScMv
vZf0LRX0gkcZGuH9eOAy7T9A1HR8CQOl47j+mMVa1tx94R8RomOWm6QHqZnAQSa7
Wcrw+uJVrBDYCqkYGjHWvlD67aVAN9HpzMzOyjYE/h6L6qq6s02hxnfmF39qBN2r
Q2DUrQqZ7pgoPon0/nev6kCZtOfIjZVtXI+HNajFsYPGXdzqoAmzNbgoB6Qf9r4U
Sw05GxByeoNOk0/OW4lZehqmvP5zQdGJ2n4fkjbQ6T4Ijo+bQilapQTuJBNg3erj
3yDs7+bWTMpSsPycB67xUr9ftr5qFJ3h3sS1jl9qxtksCfGj1rxytPR8IetsEMAV
FGmkV7lFUiVo4aEAZTXvDVZzhBh34oyDzjt6piwMRLL3owvtphlr70LyciBvATnO
6cH5Ryk7vyxYTYNQRaj0ggA7nMPZsO5pV3o1f9iU2yOMY+ZVkCa7il2/KIQg/jMy
ebocl8xIiDAAdPcICEoEmTqG6h42zLNg3VRC0e6uPMkyOvCK2hHIfObi8P3EMgwG
52Sisrf5dHKBfej3Z6xZQe+ZekteeQqEMiEcRipzACojofP3I7HoRfkVtQI0+4cy
O8f8ar1aNtUJcm612Lld6bf2ivtIr4aJXBZsRf416fn/as/4CtRWeyxbXufm3Jgq
5nFl2ZCQb4Gee9EL7kZhzFuES5kyd5b/JqyITVC7l6Bm632N1LW6q/ZK/DM/2ZFM
TaS4RF23mWikMQsZJOT9u5v5jbVdLMtj5y/nE0wNj5SL72WSna85Z5SWY8tUGYpN
VPhr2/0fnaZyc0SD41FfGK5h26QwX4AYJMF1Dp7S+TICxHxx/bqmJNtAX2lJwSjJ
aTVLVEqZNsAPOG9u8okCIykMDrJXT3MvzIOJOC8FNNpaLIopirSAcnYqgSD5EGba
FXsWbYu6XSX8vw7Ve+w8Ea3o3anygMM71RiqYkwW+Ph8X0bIxX//8oA6ZZ+KER2B
gtZahAE6ZDboUtaeid3JrcR6HAJwQxZQ2ndy75ZBv6EBMxxuwOB9VsKs3OaqiZyU
XkWiDVx7ognsEGbz2TYMkpgqNx/Nj6rJvhkzZ07O2IGzcI6joVMSk0Z8t0HDxqeN
m9bXDoTcBKLKiQkAGj5ieNtClRVJklDBBw5heVkGvjXQOherIXPyb+rJAQ5Bi9rz
2777nVm/BBrINabxVOG8+DeTygYHhMBE5KQ1XyfOLTAsDE6tKKZXcvwkApGvyjBe
UqbqpJGD9gP2k59ILpuDXM0HW4NurWE2rYxzm16YmWC1YQSYZwUqsMsJI2JcNHiD
g/zjgLvtHvJStTkk6vtvnoOMYGGOA3MbuP1rlQHmsTsnXJT9H3HHXo+S9McLiLA0
CjH/0bCkn6HcN/yJYH1xMbuqm1irCn/oov8iMg2tPIr47ksLOS1O37Nlcw4NFK2W
h8SNmBxjf3G03cyftPiDBTNKTOsMzA1omOgQqVI/szJwpkIi7RWNI6nFrijWZ8Q3
d7kyKDYytgyo8ZdOj3zTGa0za6AVkI3RDFNMHv7Kt8oC8QEU2z8Ql/DtC1GI963g
qdWAjNhdGkiFEr4/HUe8bdYealyYRPeFb+KgHnwM36Vjmzup693Ojxkfsa0qqgO+
TlvLIX8mVkbN+939nY7976wNNKuHpnl/3uZTgw02aEFaTgXi+IvWArLFj1byiA/r
zElBQAzOhXSwHUjTWNSUycpgVP4nBJMT7p8JYwNVUVD7ldxtQIc7Kt9O3b4giewu
azlkxvm0gKQ4YrhTvHHdhAh24c3uBtS+j0barUbZojTUCjZiiFwzu0u/JD1ZksjQ
Oclmk97hzpVjCFzck1lslrOVdubgP+hj+pTVwOcMmYJrij0wM42eyyHgcJbk96HC
nUr8pj/hGzJbO0JRKatowgsNXa/4VYhMbnPiU0mat60GYsD/bXJPHkfrbVfa/Syj
xphW6isovl/AUPtlasSR4WVmaCTBvZPmWoUQLgwdQZIlSxPEtBToUE8bZSwQEPA0
FVC25UeZmkHykDJleM7Uj6Y0+aaLK+1Qf0ZoFHOkx3uWgnfBXHIGOoFUBjd8WJxz
JfJgwXssC4+EqnUMVLwlURl64CquNV/5bxwAgQNzitXNZow/X8oS/9tCZnYl/gct
HKoGaECH1/4Gp+EzWCuqgyoKmv47JpCpNIQlqN03Wtm3sJ6t5MCNFQDJoT5nDc/3
X+7pXSO9bvTUinnb2SfdWfdYAIXVDpEaKQy1PNFup5Mpd4nDQpvOyiR3sxXAk1Fc
9ukNVHKRbPEsWLlYfVZvW9FYoGMx7WwuVn3HMMCH9zJfgOqNR8fEgadsCMvVBWZE
hruOhvVG+3nzhj1asiOMh1dsuzqfc9wyVQTbsHK4ShkxLm4TWeynK9oJx2WObJxb
9cb4+e6Nizr0VM4j3M3E1waY5lADbFMQjhnuzYUfdc9Sr1a5Oad++fF2gn7M2PVX
CMHX9AFNm99Jdm38tvqZ+8nrIaEFjfHXnXa4My4ZXmJA0TQ6ya/IJ1xJNXrDkVLs
9xNeWUElHAT7ngJH1vNODmOOxx4QHtzGdnYSmofgGteu3CiSv3iGRh2YrUg1i5jd
TcgFlGOPOzVps6NVNEpb1/6aE59WHYnvE5Juz1NfRAlwWFWoST4s7qfwuY5JaLgw
veOL0tkbHF7b3vj0njqTvjV+AfSKRwUFdzCA0clB88Y6ierNwzGisa/COk6PfP7d
wqDvL3+ChYBkeoRiSYA/gHzAB4P3T71vMVERVk6WbPbOBS6uL2nFqxRc3f9vjawA
PIHik8ruQQR4ElakmlDl7/qcP2cE46g3tT2MgRl25YQNTKFhHncxQ8agDF9a5wNQ
ujzyUECthlZNo0SG4S/vvnf7xNhLJRJoCYC8HqwI8EpGLtfN6Vamujplw2P97sgx
hk92vZE2vlNtkXwqcCg7HZJ2j7vv4nSUCcb9uuHlLVJSoxiIUp+Bob52Wul052dn
1zou+2kFfY3hzk89TwBrt+hyvA4j/05qnmsI2bDEdmG4KgoBVhw/jHC8TXIyza05
SjEGKNV1Ci0c1KVz/1KS2vq66VXeC01U307xS22oN6Qwe+9nfHFChlyvIa8+6GlJ
dT3ZfP3Rtad01BMfrOiQXqg37dYYLbfTCOWACHBRYFEEknk4rIpYr5hvkiZxTXvY
6mFclSd66mb+vzVou2+yUPDpIina9CrJeDBlDyMxOif4OcHAVWCR17ZpvpBSFuO+
giCAUO4PTIRvYsYr0aqPXwxtDrYQPWMYvYZcAzSu+5yylZiWR71vIFOVmWf9gtcc
AOfaq30Y6WU1FH5uF2OgGV/3EGMZWKQgAX/7ptGTcAn+YrpXTAn/1fTXRuU372ax
CFRx1eOaVW0SC0wvLGsLBn1BAMjA6BM0asbg10zpk4rEY1jEwc1mL3Gr8Ob7hf7+
oHM7y/C0nGVkkjWW74U/Ox3Mpj83VnX/jvsb46JWa463GRpNnUYzoidRQz/LaOtU
wU+QNm790LS47WAST8OI/NbqUcAzZ8dh1Z4p+j14u5eLpPmu/AvfiUlfWvtgRCdl
/Gc6q22wX1BWGmlxNhTVy16aK7wMjUD8NzQN7eHCeMJM9fG7enT2h5sEY+3NC2e+
BuS0gKTELB+F4rqRhawR1DxIlLHT7mYxgqjCnrluvcVtdWgbxq4FCXl7tYnz1QSH
22xrb7qATcEOcuz25Tr/SCZKwDSY/DQnBf5fq0v+tTjDmAOzLFVdq5XjZqCvgYNC
vJV/hfGuXrSvNj87HN0OpR30dTnYLAsVsE/Laz1kq7Lt4tJP1GKwRna/734bQvdo
EOAzMd39V7HeXEgYxZWgLSwGOsHp6+kR0tD8ahDG/TRLLltCy5BEG9NfB5ORHjxW
B9d+VmSFgLC/Xl5vL4C55u3QfMtgdr+rGsbIBGEJzIz3OxvNzZ2j5vQKx2yP5f1J
B9YHhx+1+eZjOAJKHkEEsK1kR0fycrzBnei5YIPFNhxxjrWxE/mP+GcMQ+Hoi68y
3EwYFZ9dufmBawzSPBSty+rwHidHBY0xKoPojs4XLFc62APfvtw1RwgGuhnpWy2G
C7BmI3F/tmP9Vq597UKBzrWutBmHeNsQTdFDbt9FxuLydyBgLRu7otJ6x9Xxmaaz
R1K6B3zKZvnKEt4qBJUwnz+/Sou6a6+f/eFlF7UsNjibFltLEHaQzEQVfYX9gk7k
iWRPUTDxk3Yyu+dSdfB86YLLOP1F48VJ2RhdpR28ZSYV8mAHjJluhon06MOdDruH
uMgzJcOCml9uz3WLBd9BQG2aP4VehrpwpPCk6oZHdhM0YlmkJgveQ3+lzofGovak
pHFcuX6NuuPIsI71sLfGV5LWSCf4eWUXdL5Es5PEVCVWe8w3eApD+jX1o+T8Fk+m
XWullLh26crXosOrIsS4IwAhlfL/9hEdpvEKvy6CFscb4tkeuSYCSvFhs1WuY7XQ
t0eX9Gc8n6P8/Siyoa7xA06+AAk9Zpf9LVbHc8B9Giy87WskgOFm+pFPxwJQXx9e
+/ASgPvCQfPRua/7GvJnUTm29/V5CBWWpiucvTS4DrUUqrgR5sNkToA7vadjs9Mj
qUrElcv0YxsvQLaP7r+ODFFUKGN4sfnYraxsnhSUBpLJ0rVnZeVZkJh9i0eQporb
AQc7VeajQgFLO+ToAfwdUXG3jpMXOhJsEP2PlIWUiolt8BwYXZIwgGyGe6ixk+Ck
82s6fQg8NmcAAN3MkncbCqNUPC3jruT5NoJMD/5uKFtWsTFI9OFSQHulMG1i5esm
uYwVjvWHfKSYHE5Ck9E9LnDzk3S/vu7uf6r3EKG9Byp4Gbl33g9DS60w3NZYyjcl
h7gp1FNphJgOxyi+q8S3QrZudT51Tg2NfqI79xS2tpZUeTGBdwHtkLljWQcRLzD3
91CO8kdLESfeOI8UAjL5jRuCxTJB2TNQ0Wi61i0v03mc0elc1NYjJepRxCq4BVTY
g1GSvzg5VDG3HUUsS4aXKHwlkIYWFDc3WFhsCvnkzKRI2cVnZ5GU2ozdqZE58WQg
FlaFXZfGNCcuFq07g3mzBNOjsclJ7TudqGiMEH3rbhaWd8X3yluvOBYTImQbUpKJ
zRJdRde9Kirptv2zPnTuYGc0Nb6qOxWJp3WuCUK6cIIMX9HwMQ1x+xnuVEPZMWQZ
p7pgqFhjExMJZiklTvuN2C48pFzFVDbvUoFTvprFeZzKNI0+qJOH81idWn1CyOXN
5bEXzReRCrcGxfQw3MhfF7Rg45iUOa8JTRkeW2zzq2+XOrwczDKkzOtI/XkT6pB8
XRba9eK8AK4ccPcNe4U0nZd2t0PRhImW/JHZXZ03d1Nzi1MRjHbLJQ9t+1/vI9FM
WvzvkmhwxjEwvwlkLzAwvZH/p3Iy8v/HTTbGVVqvyjKumjfessomWf4vvLvaFa55
IFSM3kS6fKynLFlGatEXk5vdUtvZsnPyvAURHW2HXev59+w+cM1gyYpvWAQQFKiO
sOOy+5WJKIuM6TgVDkbDKQUpoq3fdE5HweEy2Pn0gM/w+qq5nTpt2ortloa4OzCV
4fX6FYOlxr6vZYPRIHxHoKsYH7P3ofR5JfufOyrO3FaYOCp2Ve/G+U2IGhrozLdR
GdR+G/xx2GIplvDYJCbDy3LDyzA520opKGL/nEjZZyOWt2Z6pd5l+YOJ/f8i9ipi
FeLFMQue7Q8caqYLxhbdvNa7m5oEbRbZCtHH+rbnmU995eKfQKoogs/OqF0x9pPa
VyGTaxFgk4NTBY3z4cdedeJlfN+puWLxsq6OWBV4yisvNfJH8LbPrusGSYaPCd1t
s1ZSMorvrWSOgHkEoNuAoupIGZT7fxmGtmO1ZtUSzaBAeIUno7o7K+Zx3KOETJsa
FElJJcbyYcDmDyNTnJPMHhBagVh664sjn362kiiCcozKjPu7DLpm06bxrqLKjsEu
Ec2siptU1Ge0qb+q4JsWg1SC5K/dBCmSKCk94LhpOnMnpbRg8b3/Wrzkvo7MjiWI
jp7B3BikMiANHPR72NJS5u+XLR0kcQx1SbQ++oFUjx/1c7xQT/rIB7nYWQfVNbPB
Vl0NSWjtpF9C9HILe5pnNpZdOpHySm4CjQvnFsMds6RL2FYB1gVjY+2yNBbCEwWt
wKHr3+RgyWlXZMVhhVDrcsLFXO+KZtkAYWjkX3A6lJDc44hK4ag/XOraoPdGBFu3
4BW9Lp/J+INfxdWscY7YlnyQNbiBRQj5yTcamVbPO+gJHAhsJ8/dzb4sSCLkNcNc
vkvwfliclbxF5ogE68ZbOxe0dnT2OzP3O6fl4akFLtUF35LhjsAH/NZhvlaMTg6W
WxPcFEVgs0hKgGNVX8OgVDMbtFdqRRoWR8JQw7HX5PvouYSOh0bcWCBMrb6+jxln
JeH9n3Z2PIChBCx9UKWTnk8sZwkPY0Hl+IO8zCO56GJNSbkCEqdEOnxa1st/3D8u
5t7Su9yoqrCFocmsdkcXwRV8RiyEdl2udge8VEpiFz/jXW8ohkX9hxNLvUk4fW3W
ERL4Pb9r7hzXeJ4v6MJ9UnLSUhXtVsmg6qoXrGTyQ8qexh7vBQcqsbX3n39ADLaq
iwhPhxa2RhYmKnMGXmz8oEVK3kyo0qtl1CAcEjulROlYbgvSYNxsf+0qcskSmbf5
V+Dm3AAGJnJ3LWJIbsfxs2Ul1aKniY9CX+yP8lgip4led+MW9pAjKX9NrNi/srU1
dafx+zrOUAxOsrd/AvfMagYNU8gfBaYPN0PS3dP1yQZuxLMt95/AfhUoh0KI6/PK
dxm4yF0HfPYPFMR5HvtZ7f4HqrNQIHbbGpdL5uwcwFSZEEH0UHkLmVyXQax5Esov
Bi6zzI8YK/lys8N1mohoUCq0T3C7EqE9qUoHvI94d+nMVk7jc6BBYdMXMzLW8RNa
r8QFuk9VxKzliBOtAGTm3d6IZKBk8g48F/ub2TRS1x/LIcqZs+joyUoY26gPNxGt
dyXfM2UBzgWfKhDvNKK6T1eBCwkORkdDGF7IRayN9WYRW2tz64bkxlyzJE6tVbSn
6kMKIg1BFXj/GonEyLCW467U/fQ4CAB0y57yDhRmoa2IsrUd4stJfslUVaCJZNTu
RIlmaucKT3Wk9qNM4XIZa+3B0Eh3OnEo3xPBRn1t3a830a/eYBmsX+Ift5tIzziv
VcdkN4xe1/FtCRC4FVGg56XT3kGH0Yw03wKCSyAl5DkX68fjdwyulwLb4HczStWX
Rz92vSc16VpXQTOieFZxJRNdH89VMrSLBEu3tFJD+HFeS9OgWOGtjPDkS+pf8VnU
RG2E6z5hsZYKC4Tgy0m6RjRou/tWetK7IVz1ZW4cngc7jpDoNwiu0zNeJJaEi3pW
t8+4WVTdPlPcooFxi/nEPtmoqKAPl6GXMzl7Xw7MvSJ8C0aDFk2eA6yvQKX/G/MC
t1WQgkE76426+dttEspIaqum10WcPlj5IdmRFqznjMXneio2WcH+2yW1SSINugUi
usDU03kAGMdtGkBJ9rG7BQx883JeFmBYT3pj8IuxjD/11shDw96ACuDT56ORo9Kt
P7O6AI+nWGBrOIpuE4WxkNI5kCEVn/FOSVJix7YcHh44F0s8lq5w5Mapte8CB49V
4Mvo1+bY5GaqWz/CxtRxIGM3xftMmKhlrxoLNM31vVMO8VAlO2/IsovlEE/Nh22x
9YOu8Dc/Gqg/vJIawB5i52D3Llzr4UFrht1jV35PjgIAKfrPCPKGXTDHEBOFNtZZ
ptFjA14wdbT5vce1oSR+rJwLZ517R5pTZsy7NRPncX6Dm3vUL6uDH1CMptZ1gs/K
olyp/ilI7yZQ3XqvoBgea1RSXDAnETl4lUKcV9Fd6fh7IkAh/QAUzgVRe6fQxBIj
zj5y7SZKrezxZjyHVLGZEFKUSFoXTHrR+//aNDa9idbfs3s76Pa6nhrUYzdXGvLr
JsI3gQyXmdU3RNjhVZpn8tUmxIO9dOFydhbEQnGkzBuw+YbXT/3cfUicizyFpMWm
hfow87GYfbcGAihR2FBxBxn2cDLGeoiAVp7u7XU+uslQNqPKxuwZDCv3Zr97Lu1b
TvJtoMIjf0R8QqVR/P68j+c72S8jxFgsPbiPMAUqdmE5XxAq3Er+8gk3dcaxUJCT
zZDerawp2IsH2UYdf/o9avRcsLeuZktodnO7DBXQCUsUPSfkXm5jvwKmZez46Ww+
1dRMpKPOUpqbcOKp0JwgjV2c9djKxt0RqEGRnshZaSyw4N66f+jjGuRe+kvrf9MR
0/Z5y7A4QLw+1am5a8Yl/1xa06jLz9WZ28MT4TghbAqkse8q6ZwcEjZvJJgkGM1V
qg7XU+vt03ZPClh4r3DucQH0hEhd/U3mEt/rg/JwkpOc4qRsiv9htlbeN+Jd2KZF
e6yISo2F7Qb/RMYhd1Unjtf9HMoHkn48EL+3EpaCXxgbPcH3BHbwANvI0VupYTlZ
EXRViMFdHbaD8+XyJShm3MbkG6nDmH86fhTWzxuH48m6gnD7YuK2BWFlwVlInKeW
ThZLgJ2J4NodPourQ5ArtukUoU5N90bpSuezOsymTNR02ZiVzA1kkpQ7OZnspKgU
jdr5Sr3l9zhUs89mEsb6PC3UkuR5KBvaNr/zlp6+BuJKG4gF6muHbBljYkRg59yd
/UyPJu7DDFSFXRrtFDPcJN1dVDgfICNYR3xpSTG5MiFouw7ZK/v0xaVzVGBKbyK5
FR+NXHjtgUKqi8r9gBwTNKufI6cW9mO5iXzmX/DdpKPcx0EDSELUg47/2CgLuFfT
5HTuxYsLxV/Bxf0C/gB4TXHXTdQISTHBM0xTVeUcsMs7GUpp77/61vgdlUCLTsr6
AjUCLj4CxNPzHJ4NEgYATk3ABZ/uysIXw550zkpHGu5cjOfS3QX/9my4weoEaWq9
Cp8QMX9lYZDuT8WJBIirfJiY3B7y69wbLyBiwcgk7ayk2PPh7JNixLxMNJ8xjhdG
HfZrZMRKT2E6aR2WbZZVqJ/1zVcTFa7Cg93S/x25kDHQOXwn8f1mSZzmo2XMkYHc
ZN5I2X1zdefrlA8HrhpGgy+Rdtlg+pUGE4kCdkle78WDDZ9o3lNaaFVRNz/L8FwF
qikxlTtHiNujLg4ouWiKqdqlHsoAGJ/4sZUlWj4TiK3RDlpFoR6BNSCozV2kkMv9
b99MxAQlV2WA5KaxBkF+Nc72/KUxLrFpr3Y5/ohNl6u1l+6ttSGdK8Tculln9vwK
treTxRAZlDbn4OlolbV4Ru/wXIA0ISPoMadvMPtsEU1mw6C3rfreb1QZk/CIu/Cm
rvCk2/qheX9SlYHYi/rw38R+J59zB6gy1eZI5DTzZk9KZH5sfyozo+bAJzC0L23j
/Lo1JqdYQRxlFU0Pq+6Mjo61TrI4Utu+Q1RJQZV3TWPHfDJwvq/gE/juZg/Sgoqq
HxZVZIJfhHNMyK0kQTfEBeFyfuKne0yg5Q2s11+kY30jHtlTTU3WCDwIK3Ii6ArS
MWhqdLzCImluirxew+B0czhg9Q5a8d5OVsl43knN6FHTcK1dw3dtZGyao9wp/LSJ
tdYBVB0A8Rspi2pY493LI5P9Kg83x1ABC6HhF7MkdV4lRBEEc0qSajnlbncZVixC
LdLS5vFRWLZSG6gNilfcGi9v6NYgVvLAIFo+H3SfdghwPQV5Ier5EYH/HBDw6IHU
p1L6VnDk9tCZWDeerzVpGlt9T/dBjG/8MN5bGVMYo0TtBCazMdX4EDgU+uGisetf
iCQSbOZoXXioTX4JYQ03GaYFjR2OZkUFxmWxfF5Ft4iWYTRjarUMrIkRYU7sM71U
VE2EiVdlFtMmRCube+rsGY3eAJyvu6iOLiwQmHwCSooAzLmUfDFKWZl0gawGkvyt
0nQAgr+Ok2ZJlnQNk7NIntyrwNyL+qJPzAUlOPpbI2t2dHvsI0geZkZivf1XbofH
KO5VRlMy13pbEqGltPBOMT0rbfOegW4qDNrryRrdNPTeGkaQk4SlgYZ1xXkzwRXn
+SDE3qXATOZpom1A7+9q2XdpwtRPif+ukSbgymh16yX05WNLhhkEi9LAETRaec/u
XjhvAx7BNeJmuFYD1qbzNVN1AyrKitpi971zoSyOyvV3U6NgrQ+3bh9ekmd8upMv
08BGg69ZOvFQUc83fRHb4YtVAlAq7pyfjE3eNg1cFy2IpXCKJn0JJJMTOl1jTmY5
iqIkl489gipkrBi0h/aiedB4+a12AhjPggKsmFew2gq/sHXm9/LIaFH7AZkW+pC5
VnYbxxD0F0OmYM8ViTNngotTI+HqtblLqj49z6EzcdbaTca/wWuZXBtEELihilUy
gmxpImpcxsMFySJuVyF29oMyXfZqAkIRemb7vwlnm63B5copdwfrkdSslhhj73me
PISz0cFkQQkKrFSIemVqTbTBpwbBh142rwSwc9dGgS96aUGTpHtd3EUwJaXupIZK
YYyJYz12SNOxWcSKwLMNw01KTvQM8+3FesEdGvvesCkNmfBOAWr6z2x9l7yTxnBS
i0yzLfqA4vJfk89Scv/faqk3QRuk3iQI1CcfDgbN89zW2wV5qgVKez0dE2WHHO9C
kr8jwGfNydXey59RHg4UT48JlsD3OuPDuTbL4c09EAsBkEDsbC43Jqj1bEQpTiEf
He+FAAzzDQr/m1Ctr6OIHmEQp+UfkWNpg/82KZuF9ltYFX6B+AMqS+L8up2ujzkF
U3I/qPooZKlgjTXuc8X99SQOhnwlqwJtXNem31SB8vHZ9/D28XGR3o9Szad3GO7/
k8XF/AVnKt9+rgajXTvrPMrgaqV6+2K4u6+157U07sJA52yWudXpzR4goqBzjMSX
/f0VdzqThZkf0W/AGZtDEKEp0NXJDNM1W8k+jFKD2h8bF1YpZBXjcnM2f9rL3k3C
NbGoZgwr4q1pVeWGEYzsWkZ4ZdDNwGmaZ0z+hbRDaO1ScLkX0G7S7hH0lpHDU83E
IhdHI6GmF5GYXeViRUiov4IJ23hPl4tWALjEbMSWMrcPT8KEf6LjLrTsDhQD7G8e
xpb9YcHk3fxp+oJalO9Pq1RMkjiURyB1r+xHc0SjetToXFlV21CWitjafHHxZuQq
XL0oAe2GCQN6ehqcqqanqOtZPfMEcgmZiB6NPcPp5llFVn1LaHJGxYrVj/TR3xak
pstidfV/lON0G0Xb4YtYW5YAoVNjDeDpA9LnCHMN/95+ES7C5jeo1seL98xgJ+SJ
X2K1XZJg36X5tYqFUNwFH+kPYk1giPwxyLBmTBAn5eBrAMvNaVJvFrya153rIWo2
Y7/LhZqfsNjs9IrkeIpjAZqnFnZ7ZScSqZgV/fKv96sTkTcFxsztkXkBK8nWs30+
EMUYko/tYKo9I0nzeccrqNexDf7DjW5N84exdLCeL3lrU15qaXJhds1wCwBWnLDS
OR0yYPpuFBRPnEjinr8qcl9fF0cxQIo8o1afRQsDMTKTGYS5d75k6fKHW/GdMhmq
BGOpbKC/0zF2cFT9LB4NgPW+Z/CDJB5rc7TR7hxZR6MCqJXF2YnNClHmi4hcPIrD
zIy3pmFA3DpD7+t2Cjx8BLlTCuR3N/Tc21mi1b9+eD5B85Yx0dnM4RKHcMyHId60
pZmaX0lptiugrKWE8pa35RYXwNfEPAxdUz6A6P7UPbbUZpM3tdyBMEgGz6j5cC+U
EwcEIHcArkRIGrHDq2cvtRd03aZ8xOBmcsq114l6fqeHtkkPzgwWf5e+wHRKcyuk
YEvAadnKnt70Y0ODBwMKVbziErUxjIh0UWDdZAp50yfifSCq/pBzJU6kZDglEiXJ
+80Vhsx7s498pCwGzxfj7MjReO9RE7PACwrQzvU3dRihAesANsB+xm7wQzcoevpO
ikUbAaTtvwlz4vrqX2ojWL9swMS4bpr9MoEi8fAQ0TZxttZIKG6aj+kHjnw09Rmo
dI5u0+tgumdj/Sn0QizfE4PI2UDbcLQy1uA7pjWDLtZYwkyPmItbpgCDFIVgD4WN
DLBZ+Tvh52l0rLC38q3nt/jcVaf0521f1eMGkTN2Z8VroC/SYQdoewRhjC/YpQrm
SxuZvBYTqOekx0KWJ6UUxEv/TA9p/9Zn3rNNLJoeZnrDFKcDvLw0wRaIui0JzlW1
D8jMqyI9pvvP9WJLhXFnDUrWhDwvIT/wpOSk/bPay0TUcuRcVOtIrOdosnLsnuHX
GWmWUoRIA1gPhcH6cv3FOs82id5rV1eo9SAUoWnnR6FSKZTyF5TVXuR9glzZqe73
uW0dhTuPK6v/obc/7/CmvxrArLAc753aqIDWI0AbPWy/n5dFDzIp9MR8qQeDPj68
xLAid/iYx/uYybymUuh4sQxaw+QVRra7u2OD//O1BiyHmMn69uL2ebsH2pD0FNUM
1S8/qsgIKX5dRV2X0mGZil8v7FtJcDe2VMkT4cNmBCNZHI/MoS+afK73UkeqLgMh
QTRGw+JE+97FNfLwts9aQcpgn9jPek/g08CbLsSik1vtRO3ZbuhCMTDYwoxhdBid
fkgAeNDYc4sMDa4K2J9kLPl4gdUm74tBJzMPz4bmhhKN1nMktMU7AgTqhwbzqgwq
tQh3LIfRTu/Ss+LO1vgqnS1vIM/hcqGhhK5s43zDC6sJc5sncYkCPXd5lCusbv/B
u79ClzHKOFWwIwEgQpKDMnj9AsjgnnXS3/5YbMp+cgZo40Oa8IuheQZJBXTvd5au
AMiawZ4j2VTYrTJXQIidS2jDDzfHVjFD9o08OfUFXhrvVRJESz23mRucicpCPPhN
n4SubaXLBYQ73AUuDh7GKaiHlXV67UORhv7GjmeNCZIchXO/2zWHAv645eS66Tj6
pGOYCDu5YKiNEw/WbHOdkJ1KY1I1Qfv3NHgile8QKXt7CZEwTFHDLyWc9Zh6Z1gm
pTZfgf0d+GN053DwL3nXtJFvUpk2gllXMh024PZ1AVBjB5cUXGN49I+Yg2xkzZ9p
NC9NJjkF6kIJFwdsRzceXDuFGW6OCQRDS33IVaQWATScauaHhUSh6dA+1R0J+yP/
nWZ6wqNl3mwFLw5xw3V09j5oaGOMpd6FGZsppv/FhDv7VCpftyfCAS+nyJUSKKU8
WjUAXFOgnm93bIoVpJxR+duwvrNJFPxVvGmuKgRtFidT/taVtKortht+kLRyJzYa
bwGCXT8rBSn1Vsdg5nL+FsY3XI+6ANsJJBmGTW5MkOuGrh+9FbapVtU9lKeGr84J
3YLQdooZFVFg4TzTUxWVHKhgIeqhhSmmLtuv/TsHkkN5skJJFXGuhzykEzjCnWT8
JWfUEFR6TUSTQEeAagP0HmINjvmJZeeSdum3n0zQgkS2O6c7VheFgdmjMm1AIKwa
UNf8Cgf/X22KyJVlWyBXhEfg12CoNSaq3zwhqL2aBLF4vCabsmXi2IFcI5L1ZMON
HN+TpmbILgM6tj+4prVrLN652TCWe5qx9oc0r+f+G3aj93GH1vo6LwfSVuzrvf9q
pUGBoTOWBJpgFim4bnuxnCYm4A6Mi6KCrsmqtk+yqAgvlZVe6PCdJ2yh/VSduUB0
mVCcB4f/HEieny7py/Dtxxk61EkxdAWEOdNKXSbsKXSMsP5sjxjT5uj7mHZwKT80
tbb/4d6QbFSj1gqeroSRJMg/TUMXTA5z6tBsYCQRMsz2mCAnficKSBDyXztk2OeD
tgGusMRtatmqw7qxAxmqeseiNA3iNZQziPSbhSZp6xJIuID41poNzeFdC/egnoug
mbFxUYmG7LjmKvYWpiv4drRelixF1Jc96CP6yK3ZUmylCKffs5iqeGuCmkkybhEw
qc99DsyYsYklzfvlpB6g8R1ak2x2fcUZ7C14VKXvPnu/ejepz4JrOBO+clvTXM5Y
/F+75Ylez3Yy6urSfgl2GB6B8kbvNiCTKzdkO0ppBK4MCz4m1CSbAuohbXbiRO1Z
BMcGjiM2ops4s5OQY15PNxQBF2SIpeltLbzHcGR9Hy6nenF2B5R6jAkG5V9FraYF
vT6jXanq9Xk50j+sW470yEwt/NacFuIx3sUmcjZBAfSFmzonmlxRO9gkxfK6cxlk
j7E0kOva7extTxcbhaC+ATToVw3Nmy/a74UODW3s16MtQvvlIdivnyTi7eInausa
YyJgnO+BmDcUkUoiYNRNQKA7lbyRuoBQfKEpzlZczxQQReV8+iKQZuZgakE31O4/
tw2zkEx8Xjh9o98qGiMebAVLiEU+HbwG8xDNQ8zoz2f/LkSIaD80qb2+NVlOC4aA
cx+dqmjVBSEM22fbflkpYu8+g6b1401Eivy4Au97uQR9JNh3utZX9U8zGmtOo8cz
vYyD3eNU+1/QfGiO/uqWtgVOgbUH1tU1aBwqY7lhlk8q+BIlS59G1yNhIhhGXP4z
QNk5jKMpDtCsIFVvOLaYGvVFz+5becVcSY60ERriunjKYuBd2QteNQ/+SkUZJ1Q/
uTRJe9tIbze7UUd4+3lmqP0INO7hfhhlIUDQXj85Z9Lf+6SDIKCZkvu6oh/IIgR9
VoMOpQcuwMAVS8JYVP3e2qlCUAjR6GmZeiwHENW454JsVlci7Uxllgb8BlLxwcKm
jMG7M3w9Uc2AFMpS/1diyB2JG3yV07onZwwSUc8CdLlQwnxkfy7F3UZevdItvCgN
nyBZ3/dhLBeFuDMwj+ErZjvygio+wSY21PATJCdSeKeplGih/luRpAYDn6WBq7TZ
JFPef3n5kZSx4MCulm8QmM8XXzuQvjv0IQPyKo26E8u5CozZOfKaIzpHYBhxPW+g
WPKkmsW7jWD0miM/eVL5Pfq73haU5zeM8+HslGDDeCtrACuOuZqDZEv8UKC5X1bf
CQ3tUOiIsZ9MYdwz/j8qWlbw+plkAHMk7MHbFuY/bfmvKtTDAepbOO4JiH/8UZSR
8c1em5+vr1AUj/bL4upvSzr0h9klpvmitGVplktoS6j+y4sdlIzkcLmVz+dheXYv
nSVAtQRMJBA7QJoXbSQDkE5Hy4yQQRbtEJ7IXS6z38SD2MBOt3SB/tJ2FmDbmNka
iv2R5MV7sgYDIawTSPvMIGczgjHUCYuG9ADlMS0xddLIXz67nQhO5MbkAK4TegM8
yUXHd52w6Giy2yqavsoarejJnoB31mz8ONYBv4AwOuz1sS+84dKMTiWAADqXEdRG
W2yLo1cjkWDaltX6BWgKpY3gPiv28nYHfRWPhplPTkP56mKJDeKhcVETyGVkLIy8
GcwzLrgzuHHQlQqaYKxsgziXk1UbXQCsRt3xZwdcU1StN2ROS8Mza7XkW8Dor9V1
fyG6rXXq5QnGzRCXN67Q/ppHM0zYUgInOAGcOUNYV9+9cBfCM79CegNUpHgJzzJk
a4v/eZe9CMI0xfXkGwEUk5I59auE1QHHfIVm9zOYdjF2RKqTMFyxh4SdZ1NMEz7a
gY6KOlSEkjS1zye+EWMD7+qbNAPLN3ey0ei5AjJ9W20J524jqk05EoSDot0/8PJm
Of84odg2LnwDC7RAK3bGmSwAuzVeP16FzM8C5Nb7IZ1YM1Ew6GO3ov90otLCUUT6
Ob04spcduAfPxMDvMnTL6LcvR0XpdrbkaAZw22YqaRg4ukt6dBr/vFMzYyM/Vov0
zbHkpQsiFagShqfqVTa6m+Fmr+oJdraoO48PGUxVR04/2wUAqEeyU9GyHa+grEEE
fgZRQneAVEnzvgYsbzoWeYku282kYxHVcQGEGubCbQmZm+ika2hpyNn4rTGO1kOb
38xMjAx1lOA5mGJl9z4M3OQIgMmlAySqp3VUlrj5TT3PbxaEZr33En3+tUuna/QZ
KvoNw2JcPAsg6QqcXW7TRiN4rY/m+TkZIbOq/mtLWF2RnccFe2DiDlS9vHhbbxs3
Here5nX6iwRwdw8snlcjuH5wXKNifj49z54RQl1k8xPXdaPpDr2/vZFBqADKq9gB
CBvINcqQK3SatAj84gkJckqV3eaZ4S3ktMOmMNI5D2CLvflgRch462pk+EAZwign
/kt3gI/44iIQ+AqyzfYa0VBDRwmFMZXS9nuseikeTx/HdxmiCFEWU/h42Fl0krvo
NqqZnaovu7Dx9j0gz4pfIxyBvRU9kZX3YLbGSfJQUZjAUnQO28E3BNFiib1f0qnA
iSSQsd+UM1bXbOJDe38dr/B0o/XkE9ZdZgUJXV4P6MyMRPVELezeTkbQduEEnmgf
z8HuQc/EGqoVb/M+JqmypicOsQdcGjbEY8ciPIRuZaGK0hW8pnXVQMkkCDhVNlD4
C25pmNGjdjF+FtePlHpspmfPXuUqizt75/V1gtGn1R3Yu2cM/5FSEkQrU32sQ10C
kyJ24Mkq1FZkpyLIzMtDo7eoCrsGXamQPcfRUEuNP/RMhVoUSd30P6O62VMi9n7Q
NB/+eXHyk+JhiORa34DDq1nbX+4R3U0lzSCx45wBplIWqZQ6SKKnkrp8jgjqiEmV
osvhlHHbzZ0ahzCAjFjT5bPfVqXv4qjGLeczs+niQnWGgwcEgFkdVUiKiR6fvc7j
lPZXhIpLVEUdFd3UyAQLaP7iFZuuHigbkSf2YJ9Mt31dr8Iajkqxya4lMLfEEcrU
j4WKh+HWhkevdiHUGujoJ/FXkjEd1KmBQl1CokZJrDhNbFaGiSCHhj2GnCqmrvHl
kiIBILvJ1oy6L3EtXPs5IK1ro5GzfYygkiO6NKAwraodEtOHKhpFGTijkjm4bpQz
07BueO0iQ590Jb6e1Ql4AFCuu3uTcxq0gxIIqQJy0cdkmJ7RK7dmRW+pVaO9slzQ
LBSPtd2jbOEcjC9AeEcn4ptr5BLr0TqPYgK/t4EoeDA26mwBr2qomw0ZE+VDk5Pp
g5tCLwCGQvgLHb4+rIZayfOI8dzbZwcYZsfT7s7NVrFG/ye+LCoCYRLCLL06pEqG
W9U3AHqCQYL/LMrP8BJRD/fKzrJRm7js9npld5yW5lbvj/I61udtCdRC8+c5HEAo
Iz//Zz4tuK16PHLd4VYjlT2323MuG51N8Dn/78f3cN4IjOg2dL8C2YBXkyJRMLOF
yVHdD20KejCIF5YOgsLylA7dM0Dx18bPpQdRNwWOz4UrFKpiINdnNqULP7IiPjD7
fn2FZX7jKePmOpJHLNOBTH8Vx0ylfF8ppqOnOSKIOksM/kGRe+iQbc0bKUoEJExz
GwyoxmMCefS9zJeYiArKMSz3bFYtHGOyDrLjJOQ89rK38qi0AY2ZT+E43BOU9syn
uDuIvfPwpzGWGhD4K7OGYflbxhWotwuBmR1J2as43hdFFVkP3B6QJsnFIZarfKU4
qKT5yOKmsswAfGCnPow3wn6kqmtVmBqupN69hcVV6w0xbBRHk2aGAThDAfmwPPYY
OObsmk0jvjFzuWdIDCTBXhKKSmennfM7FKep0VCRv03DvVxtMU2p2DktzpEdxLRE
5fhPXwj0cNGhma0pOcbsJeqedi9rNA/ne8/21GycgrsmIvpaL4NH+PD6C4PtnE/5
uOGRl2azQqyjt2jvZQ4I4pXL6DBymo7SNEJqSy17+wP0sS6IB9opqBnSSw6quu9G
PTNZyY/SALWXj9OjGgkpgmopOy7HeBxeVLU6d/J7ZmRYG3kHkqHoADPgRfNi2Uk/
43AtHW0+lq6Uab3AQLkW27ITIROAHjytXdjeeKN+9b2aEcQ3YU8D8HGANmcv5YQp
WmvQXHmSzDEvrvxjASTZwv6Ip7HCKMWMX/UR5kZQBdX3MqmrYm8zVV8EebFQre5g
XOukVXtqQwyPY2cC3a/HA2/F4InK2L0PUzmaHGeMQJU1NYe88gn9ryq/oVzX6spW
l6RWOHC/WlcBWHFLFpdLE6FiYeE0ZE1wVtHXDvu3WxW8cWJgJyBWnHNEF/AANDyv
W+Oq538dCyA1Y0OMDiLhScYnzZTDVtkswi6lY9vjkOsvCHreCBwqbXiiRUZF+lGh
NNLRWD8QuVyLSggukINgAf/WW6f3Xkzq/oMTu6IwJI2dCzYAcO1YLkxNMCHbKKeb
/cgieGnrlrTxb50vtnsiPEY+AHhk6E23vCk5ahYN5WQnzHVoZUJoV0xLNSIL5nYS
6KpOFhJclwsUGYoDrOpEzVcsxe5GXj+ioLFwwB16LkUooBAAxwnIUI4RZ+CEo4o3
wC2F9HrZwWBuG9o6tF2sHW6ehiumQNxAYSa8JuyXZVs6u+QP2JZ/qo024CJEvua8
BmdC3D7rWHdMmTaPCuZHlKSmv5zQW0RN/Hvb8/B8v6I+TVM+onm9AygDCNxh2eRp
3fd0q8ZogDP9Vo0Kh2CBqlM8yqCB7ZcFlp6CWCnPCFQsEb/SJZCJkWTdZTgEXsu2
vZWW772Bnd6BSz1dzYyrWUUPyWuV+p2fE4AYDlaoaTI/zngM4K19CQ4n95rLM7dU
C3XKeYyNTP4BRj4FbQ8q8j8NToT1TDntkrdyJHcovGQxAl9xgC6qhpamgpFTK75i
0yajiGvTQ8t5VGvbit7KPSBZOELdF9haHJcl1nKus5bxNNMjk289Dv6RIFs1d0ce
H46QUoGsdDhWt4Pb3qHl2UH0RgOhvvzOzPtqPjpbxH+HE39yYc6vCY5C0MmoYTSt
iXGmoW6Uyf8cLOsAscFES7YnrwwtqXJ3i6e/fUmowmImMW/kGHpmOAo3LOJPCTB3
gspVMxH5SwQzQ1SgWZIBjG22gOTIL8jcgOOQMj4Clucx4Gy/eDOkkNYNUPjdFgPI
ZF9MBMOQ2CKtsSaLthUvZO8BsHPAH/WmXal22dL6xe28ThqG7c8Z3AkHD1Yn19Q3
ykrwZdvBQkn1cw1qRmIwzZf/bkfdtjwroiLAl0pPYazdu6C8Gchp0WzjAc686ehI
7LjuKpQW1woPlroQBX+j7k5J+n/FrjXvGR43VOCz9DJ77Et7Ff8YgAz/BTZYMU/P
8HoqqPSWa62vYPWod+INJBNAsq30SSNzGx2dnpjuYq3//9sysh/hjlR+wTAAg8J4
soS/QaG7C3GbqrWSfOsaeLEFevp58xLrATn/NEecBRWrgkR4xVijAYmyN/Z83+XN
936MA+wIl+l/NoKJGKQDwFazn12ysQ6TjbVdZ54qIRdfQDAufJnQdxKk78JMfE1x
dKKsW3LVcLvtRUYGJwvEecZtKL2IX8DZivCX9/AkbU6l+RqtV4TfpA9Xtrre57X3
tU/LZ3nyHJVh+z0a2Gc2sLjjnhzNQyYJSCOGCKKN4JVZLdXEEFZhev8LgS0ApDab
WbCI6DOLrr0qn8bmycPMkPTs/whNANrudFA8FrKnl4HT3JHRfJUTWtKGJ/Zn0nUz
WbM1cQpKIjLManpK/TlUfGznLXxZVGhgscGK2VANeOtwsR8uayXuDvLOjlswTvEK
9Q9CVvQgo8w8tg6tsVZDQJ1TeQnHCCAvWrxDmsYgW6pA38vg7J8kSB5pHVPWVmp7
Cc15lAtghSTt4BqOaLmL7QagJLJRFFyw/6tu/pzA1GQuxjWNehSu+z+43hsWb/Yt
Hil82w4PKng9mj9Z8zN7N/Fz5sY7oGpAP7NznPqLcXNDje7cNXVqx/Vdyd9gqYWI
RuEsvya0jIv08LTG1AnD0VkWk6Q6zdwmrQZXDeeNsqtwvJ4jpgpi4e3UhwHNfkLo
7ncRk2QqHaKWxhQ03QI4gf3G/oYnet5OsxWW45j1yU20l4cMezTovuXMaWSb8NUC
zfBzaLUdjiuFZLkAEc7U0oWSo3ea+pyWaSs4OBj7IrhPigF8hDy5mNQcjTtD81WK
+u/K2Yb/yfs14UICHliFbEmFJX+hSQxnVvuUAKUIVGcerK9jzvVOdwNu+Tt/5vvk
1k49ZkGapWa6Gf6unq0d53IXnVZUwJmP6B270zmTP/T5yJG3UtmJDzLsxGSlRT+0
wU9sBBbSr9I2fkKNCn8fcCwPuxWMCy9shdJIZK37SFjumDKmYMaDHEim/grt0X6D
4ZObhMA2u/et5c39MSwQ9Ku2euqqMPsjiOmmr7/8DtVL0WUHMDZROVSTmEkmf54Y
+tWFsTNzo5Y8KhJghjuueqBZKPA0b6y51dfzu2eZDTR8z6N90PcvlKMos271O382
KWBmlnfI/j/n6TPLJpjhGJAgm0gmBOUjVRNc/ygwg+AQtLKRln5TC+DhpuAAsF6Q
NNUeuW7KvZZBdrtKnPDLZkaAwb/mwnl2dLWTMPolQ/wiabMqOeUrxKGMcLX5iZ6I
8rF21q2+i9FhMKFa5sWHd0dn3Pe7fI2smyPL+4HXiqzpgi0jTfO1F9wE8Pqnjvyi
1KmudlhtUj2afeztv+M1Wa+HIOlSidNMPL3oqY7qaS8nDEKaW1oBuq9THV+1/UjB
7Kl1yBY8apLfaOOHRejjwqe7ObtzUs3L7AC2/Yj9v0XlIAn6zQ42+Xk03krbpSub
gqCBIpGFcI+i5NxAXb4YlSGP7hBZ6DiOBra5xqCVk1b/X/cJ2YRZPx3zDpa7WXtZ
QSdI5t6iFi+mqpRFAohoMDJ0n8FpTqbuwNQA68idPsamOf+mO8lDev5tWj1PIbKy
nGErk5EN7c+hl8rt/j3tucXk1hvA3n/t1dpJbzaHd0G3mgSyGoBTwo1jpoPko23/
fI4NPGM7fzS/T/PLrwpvEq1Ig7KgL6uYtJxyqGs7rNSgnOu7qUIkxyHBug6h4nEQ
m7YwJ65poJcAiCXnY3guGJYaOAS3zkSvsR0I99FqFbrTyYcennAKqg+WtlvUxBg7
WPpa8Cq/DWkv35I2xMzg93iJO0DPFmitFfUMlaUY0H8XVC9seSyatVN9YVGlT8hw
2pp1mfMetGhfSNPegLqzUgLGyI8yK/bmcwZ8blM/PAswIAHEwYL1rTBYBcXZtRxx
YuleeFJ/gmjCEDvyqE0o812mPnIG0H1kUmQSBA9ua3Yfe4af4rRrBcKZAE2gxQwD
5TvQ+5I8dBiBbUsrtWtHoCeTFZOULibPH5OqfUP0jlSnZVFMirNJMxXfO5gYWXtw
LgLCk5AOjkQhHBiIr5BHqlBeuHh3uqHNl4fKfP14MM94VKfDFzm4iiPb4YLLqjvv
gmRbC+0lg5TpBTgjtSgTQahKsryu7ftvIX0OvqArQoD1r77Iigsc6g6ihFhCwMaB
6aZb3YTnOyy/uDVGbtA43Tq8hIupAEIhiMQjbpPMpNmvWaPeb39wB2Td0o4nzsM4
VpujVi/OiQAaGGMUbgSGal0H16DDoSmIqlhtaUyWfUkGE0CxtsNTEBMQ8RNvoKWE
G6LGHFRRwSRwNYNRRyFlxf105n+bi0pdmhkFIJskClgdADHD3ZwiKfmtCGzSud4b
OQoc+7Kxzx8PKR32aDICsPgpCOqdNNfJ9KDm+HPImv9BC8zfYYDpbcgdgZVHSJIN
lezzXx3iN340SE5WSbS3srYfNUABElvzhRMv5hGVC4qpcQmea3tIfTFm8QQKJpYH
l7GSZkPvK30Ln2Ih7eB90xbUz/RhMlyw5zoWSmX66W0jRIXdoNzKWLmnqcy5rY7C
x0xZxTfGRoyds6BDlG5xfnBynze6kVTqJWdOgCluqeh7ZQ/oRPDkuuLJcUuzBaBR
w/Q77wXwWh7/2pD1BtZFB9kiQOJpAmN4EUrX3EBuZ+b9K1rIOy/673uNkEGt7afB
btiJAq9XDzqbhHf5eyBU2lT57PyTc+J6O4g3fE9HgWm1iKpHvQ62vzp+xZs8BoeO
hqIL0uu6pIUxc/Yg/lab8YqStu2W0GnkYzNN7vATfnXCvAQcdaWnezL+ULYCRxOM
JC3p4Qk1NCNH1MbtqDgfrvCa86vwy4rNRALwjvS27Vhaf0bd6f4NSJaB1DEdo17I
C1zStjL86+mfHaTbMr9IpNFMP6ZxMOysIs73EZGB0lTdJUogqQg0x4aYxrEdbUd8
6qiTI630N9SXqpM/Ba25t4GCW60B21j+R2VcqwwtdU1WCXQGLPRFFEmIufD2doyd
c8i5KVmFMF6Oz2OGWXzFGRBjgHNpXDIMDb/V5vzT+Ams94pv/IDvL1XhVPdmgOht
FxR/GJqSpJDp1Exbme5nKCObNcezj5pgbUIQEIoB1cBhBfv6Cjm+BlXnw2s/mVf5
6atHCCpIJ0ETKaVsTi5XrKYaXjMDrNnV8hqhbr2/6XpLYCBgbozbZwx4Rxp+25Jw
oud6IfLNz/Kn0V18Kgj61lQs2bFfpZd6rpQj1heWKMsE4hl20gzrzoquOgpOD2Cp
AvoJhCLWipfr4HvH0Dsf4ZmcfPdk3v63xzb6Gp09Eank0CQJsqc+gi6kvsgKc0ZQ
8KEDOHw1AsG7tmnsv3XayD5oPLNvY9nMWJ6Ep/dpqgvNnUnnJGLQ1OWctWy7jwlA
4Qidhc/PdePilt2bOy+92XDAVKmNdADLviELRNaLUrX1qGaNA6Y3mZj3S2x/hb67
dS9sd7uJ82MTTz8FFO3CABOfaXB/DkgC39WvlvomcQ7ZBPpZtckwRTs4lnaQXKym
eUtu3M+uWycjKcxdWVobICjbroA3eo5lv7fQHmlf+hOg695HtQM5KHYLImUjI4fo
ke8trLgGAGlebUgnPMG8flmkiCXkoPgiNaHfWXt8hHGnUPRaCYcsTcAGCwsuUn4f
CdGcwxZjxMaG6JTP+B2JszUaPlAc9n9xqzUDZfInjvG0jW8/P5BuBnm3N35cbYVj
6mhwvmvfjB+6/2LNOcYtOr1vzvp6plZZe8rYt2WedKgMIo9liJMO6+LdTl1CeL8I
zs0SscxwYDQ4HRwaNGT4yc3ETHeHC8sV09+1/3TDBt+a2+Kk+KbRahIKkp0Hcjh3
EsJqPmU/nN0pA033uZs/IyQjWmQlIjIcNJn1JO4eDq8POm03nQTZErfhcXPbH4uK
ee1tEQwsT1QQBeGhERSZ0oXm+y9Md05dAt50mSj73rsUhJLzb6a/rB2/Kqd/KqIS
qEIq1EyNYh/RQOLt9l9bOcKV9xelIMmcOrwSSopki8WQYRB8oobE7PFOW7VjCDp+
IKux6hq1SN7z680KZ5yMfUgXYJCNoUld3V7tnPavxxbYBE5RlXjit0OtJ2ogJ7oc
c8vE3doQMcBzQsKLb9SqSHYk4684Gef4UJtfjRo6AB0zPDF3o9pMxdxq+xTD4zaA
hrhyvLX9Tgxed456MXbjQJVThtoIw8yWZwUv52ZBdeJfdfBIfRN+CkwhpnXgBkx2
jmJhw+HSQd7Ps+Tyv+PAfdR+YtOn5DCb/cCcHEcXr5EdIXUfOoSAd0Cn49NljWiP
WJYN9076iU1Uf+BEInBjdiwDPJRBXCB9cg4F5isvM9VwFT66jR7Id11IlE2wPOCn
nhCRJRjIsn7zvE1X+3j2QnhSUcILsP5zQY31MgoNcL5++OkmU93EHfZVAoUf8Y9q
IAcIVO3q+HzYmkq2KmANhT3ATuv5OLv7b4Hh4XSHHEmNBME7OnpeTdfUXHzqhMd7
eryJmU3OMtjjbG7p+ihCn+9pX2OkYB1OqcGLj0n/Hb7zxCCMiXRvH5pVqBO4bkQd
3npMZ9kMcjkP9h1/impF/y74SoPWO60NTZOnlNnGE6OLeg1SpjfdQ4YQYW855vZ7
ebhUQdDBLXArB2a639X70ZaBGXcZo6xWuPcQIoCg1zGpML1kbAoIUBaUDlpMVDRF
7eZyShsoARl+LkvqFOHKso0aHo8mrMVmzasq0HGOYXaO6QwSNA+vixdgjqu9Azfv
/lIHQl3BpteMuCkUHRN60FtE2AeTFRuT4EIoI3THoxnqwkbCJ421qd6z2ALKiw+O
bv5S0bV5SgEMOwJhIGc/5I7dizjU1DPdBc5yK+nprcXBOPyyuzLuE/ea13NRHl5g
tv+EmKwu/XrkRiQfhi29a3ugMiXQTx3ElIbuaVLysE7kEgYOMR5sTJJ7l/ar/Bdz
EfQ1kSVye+/Ju/4LRGLJXO8QGTjpJ++G0Pp8ckQ9BmBHjmy3I5WtYrsBMAQf63lt
4TDIn/6wQe2xNJQDAQluatq6sUj5UPXw8P7xmRPsALClw9wl0Xo5tcZF66BYdpC3
cFkzJVSrGFNkcpshvQNIC7JH8uZAa9fDXw+MJh9Qayfx742wXVSu1z8Tzd6DW3AJ
P4rMESkb0aadnbF1tFv3mraRvXGJWgWHpprPFZimQx2CRRFv5o16/ukZMKgwgNCC
EqMEAz58zRDeAQNHootN+9t8F4wxfghwjRBXr0wKsBmo9dA6nSz2WYGOC93X2VZc
GuKjCA6JuLU6uCHASXAX6mX1nOTAEcC5i2Gl6mEEauMz0Eo50GRxuQ/ahAV0Kh0r
EmFE/9dMQAIkZAg9PUbxlqQ+GcUU9yrQLr9ZJbiu7BRsdzO++lFYn8Xj4V7nJzv+
iXi9PudrXqiRZlQ/IDLq3VFJIARwIzw1jHB5SndX1CR9mgiu4eELmcEQ0DLufXmg
ZJYRujBcmN/s4oICv3W1mJ4txt7FLE0/eLzBc7pVIjBVujyYy7borUWBwW+8l/oQ
n6bqnYuniH40m6c6s/H8VkDpfKnEdENwRJtMKcT/FuQsbIB2pWc8I131LDnIQC4f
FHKNBi4YHu9sRfqXS1J3IvHWRyT5w1l+//bHZTD8WDkK96jnPHW2tFU7bszp140o
tgBsSfQFNO68Y0X15no0iFxts00kHLoZOo/Db/R7vkmc+Auuc0nQT/6myNzg6+GL
4+wNABbUSPk9W4s/AxqyS6Hww5xlG4hoaMmsTcQYciU3ICK8kA86zOznBpd/bZZ1
rArxlXqzJAFanAWE99FWIemXHLEKet/bJDQzRFqBJnVAYJZmafcxTmrNsya0hDFC
0XrmQqOgk3p9m5sLUYxDlRrlhrIeuprvXDKmPiv3uDgQIU7kogmdu3yfbq+DA2F7
h3aRzTgM3LxXTUZEPGFfKtIub2b3eoHqRMVu9j6bZU7q68XkPCnyyxHSSjL32pVv
P+1rW5YWr4u4k7mJ7Ok106tuqvkUtf7BnodYaSuNvPpbpJpgzAbfhQgIlVgrF+9P
ZztFFbhyWQCX2E2Wu6ovR7cXCsdTZbd4XFp4uvUctASJGgWz1O7Kg6k0xS7HJeXR
bV3WZkO8RU1+cODSNhS4mPmrUgtnCyvFqrGASTQUhAfu8wYKN3wH6fw3+Jpb38Wa
e5sM4e1ONUcajGxGWykOGJIkW/stmZSPC/inayRl7WNjGgOVcIbpf+no0oFHCQbq
rd+Y1/aZl7aE+QrwruajGHuklB7tFK3NkIIq6H5jJStkNGJEa77D3Avcmrw5YUvs
V7MAjm8Lp4WqffTFEWtngrxnmwlsIIAGIjNpOAlvz9oHhtbNszuDfMwoJCylBNpV
B3GN6ZvQGyZl7dCwvpYnnuuyY0KBQc4HEZI3rTfftZsiKma8Z1cVSKzDyoROfUC6
MeGsiisjO+Ed4rcvMPaf8hLzo0v2Qeow1dzF54TDduuVUF9p6sO3Gu92qWui0p8e
XaP6LrWnTFwPIp7kYVj6z/E3xYs3xWVM/r2yFWxRce66aPX+DKhq1ihzvzLqD7Pg
kMFs1b3N9tAGiiPlEP5yFuDvt7c3I3zTYuSl0HBlj6AZgN0M0+6nnSIlZSfB6mDB
5zw/tlZfGV40xdwl+Xrq3njci4lN5xTa5vTFV/CqQdu2LimD5urGPldt+Wz1SuaH
3JUho37reyQMObs8M1cBSxYNAWKXvq63Tyw82RbApfRtdyl60gLSPp/b8btzh0qw
JJVbAtpH7jwI7/e2STOUE22RAlndCedmGX48sejD9lq/MvOKku3DpjRoCEO2Kb6P
VRRPtyqK1S/+SYd8dsOzDefe0oZv4a71utkoMpayq6wnFBsZPq+cHBx28vy4t/pn
5SRa/SMw4c5RjHuzI4S29aNWMiy8/eInrSBSgJWQEIzkLxzxzk59GZJm6GPJOBiS
Yjpk0nDUrQN97FLwxJTgzIKr4qFeaQsJgOggiZT14/NtDEtX5S0N+sWr06zJyQ7y
sXV2iMCiKiWUxR/jTwQkSFG1MRYbO9tRNKRm+IgNK826jPMFJTFkcZjkPKjBOQ00
qdSuRDoY0rvrcPJhwE9sBBpUr0rHRnXk/eRxDDj9DFyD05MZuwJucBz7GlVJy/fQ
8kj29xPiJCebNt0n1RuMZtj50wFgrTLfrlIwIbTcQ2ZHU4H6fqwiDVMXxdSpArSQ
c99CiBnjGf97NpsQVKk4ud66VQiaoZdrKzdSy9wPca7ajWf5OT5ATRWhcQsqBEPt
pR169N3T2aTcVE4Z2tm9UEg2trW5qvFSauXcS90zE04pO3j+mvVdDgzoDYJ2tdHz
iyZNtddko3Zdz+TJWY1Sbj0DElUzFoggABFHI63frCK28JDp3P2E86pKhSBaPtys
ZflW4IS72n6udDryUnTwHfvGU9G6rwEWepZPXUVp86K62aXKOyKQRxJI6aaQ4p0h
3t9Qr8cv+tYt0GmArdrQQeGFjTLytb/+tAl3t54jEjVbaRmoM/DV1qFlq/V6jMZv
XD7LMwJVbVTsK9yKv3yWnKPrfgvFkcjdWFBonxOOzIdIe/rhLMTJ7BUXnN2fZ55F
+xdjAWwbzfIZddZkX0S5YalU4IknXwIXfsUe/m8/aa82D9GHbAyooCAugKN55i/I
1PaUCdWuniKLIKS+0GrO+O+w/Lv5NQqOxkdPXKoIn54oOYmJzRmFJLXu3D+Ow/yS
OWxMeUCxZzuSb1HtZLR2GNtgwddGqsSYpgtd2ZztDkOF1DlyBOwE0JLpM/l6BAtW
EY3+ZKOgV8cJcZ+LkG+wdzJ5iQnbAlbgQtzUvGmEQxhiODbXrd1gRJPKyw6hssQO
zb3GTcT8yHEmoFAM5sAjkAvHNxjm2M5VKOKGMdSQEgSFXY4z8AnNcexn/gGt4d5D
xFcnmP1gJIRG4y6oqC850ZbKmVEZGEVxypKWKkz5I720CKlj0ZcQCy5XhPGZfjnX
YQbdCjXRdA+bLmfv8ktXzpfh2X2iP/vdTIHC5KnVvO1d2RQobLbvPtJw5jyuScPj
FKbCTY1nTOg4zVQNtbahtm5twK3A8kvp8CMbt2pa5VBABG7w/avNIHaXwM7SSEEu
JlEeppEOF0jxM9hkgFDkTozZpVFOvsol7M+uny4aNueDhkI2G0CgDqRMbJZvZ3R1
JqRl7mvB7nxryXSayReLyBSQe/xGQGtGzb0+HPknbfaRb8JvGBGi5dbWtwyeVpVm
O251yz4ho67uH5IHOvWcBCJ5bQALYc3Ix8vvxwucXU7nHymMgV08YHmX35VfYA7z
ioWC49e0sE/b872+FBYlH38PDvOk7OltnhZLkkSa+6pJKo8ehA/Z2LTQ83N7xmg/
5shykPNW7lPDUTzwgcCWwG6HRuNgw8VO1tOclGksD6f6S9Oy7Ua9BlOLNh+RY39E
nvx1Grev1w0queBDyL26BXVp/Xy6nHv6+sEL6rpJaI3ZXEobdSWVNR/gGQ1jIQJr
YCs+7fPiBHBOeVuhhD3WWY8O00x1G8MkkWER5YAsZ0oKYdc7p5Bq2c2VRDxosJ92
WbL3Zkaef1wwVNhosmGPnvAkbfHCoWho79Ryqxk6dEWCRm+Eh0sNCrCygpOy2Lez
sr29S0V0mROX7OtFoXilIVhnpZhWhrKxdpLmSdiFZnu/eM1jH2aE+vPUs6BYT5iJ
FGh5hRKaxr75OmdODqnGWB6ZVg8Crkdycxu4T61recC+R0v6uCLoOaFvoFC0Pycj
PDDgyEv3oK9FPFTW1RvqltiYiYfM9ouzdEgryJ4LA6fhT2Nk3Je0qFM8prWDkIUs
sQfzlVm1ZMMkKsCEQ6Ef0MyJHUBt0HiCxAoMGqSCSRaqBugDCvbhH5LJM5cXTtR8
nPaayizEEAGcZfkbWpspQ0DXRbJxg/JApW/G3Pu/2iQP1ET4SBmiCFa3RUCSC2o8
wa31xiEFQerkGEHX2OZHdS0cAKrDA0pXpfDHA8P/UVFfH7YSzAGgV10VBuCkhb5w
v43rPHPJF2WM5rLzpY1SVQ1nmwLZJobrk93Ov+/78NKGkDXNR60iH220O2HmsaWW
Yx8K5IygsZtnYM4SNqJ2ECh76bsql16AgQjVoZHLxBPrZgmn2NOY8a8ijPHLI8EB
HHbGNlT1woc6Q8vboxuw4dYqQYJY8lqOOLAhEr5QsLg/Z4xGh4inzN2qtla3teUs
pyY3pVQC3iJaI+Tv5haVEv1fdlL+enBcvtCZbJPZrkJClc8vVWbW/0JVB6ijHhq/
FIay78vr/XmreejaZxPyYUdoA3W7DftfXJ5ItqiuAJeBeUUv2U+kKCTQ6A3UhO8L
qtRtu666bHIAMBnALZou974r+eyEKj3IxeezxouN4cUJ/mlbBfvQr9AZZnAMLu1j
nNZiaxAy0SMl8aJ+Gq7JD8S37IAKeMRCUgtDOu/BfHrzY+aqb1gBUWDD8aGnQTnS
+UcMFMI1fG63zYG1xD3aJn1KIjAxRWQZjUICfIwuUKF75iqWMKo5q8TW9S6s8Nsm
IhjOFFB0L5+kaOkbYohYgmh1ZL49GOl4obBRPfvIwb0kh+iLcCdCT9y12xx3K6Ay
IRz28Sdwg5czP1GHLdbXydtdE50Y+MGurFqBBAg391D6ivuAv3kVQY82Jo2/KoXL
pyRI7AjO6Ra23SOyOsqRctBv7wNOmnvPafImTrmEXpCtoGU/nwIE9w1S6p3zjmVJ
aZ/KDpsQKiR/yNHtJRd2zkCf07rWle7+Hf4qqSqEkI+Fmrp/DYZtr3znMForJByI
+ftX8JAG1cwnTsd+90nPFiEPLmiVQ5k4IH6dllwuUbBfuSQm3F0nV0YV63hJDq5e
bh+clbmUsdmCdhqECqgHvW+OUQKiVGbWgSE0AqKz4LfU0VvleuqPv250+s3ErXm4
Soqy8ej5C//Jcrqdc5qmgg/l94fft6t9Qf0yfEsPpqDYIUczPLG2fX9nGjP3Nwp1
kSY7ffoeGquakdkJYY7d1U9rgug3hhTOWKx5ZXihOE+I2VZgS6ymJB0L9oQ83AbM
iec5uq61S8BVDSSdqU+cgCWSLQV8eKeYq8crPPhGjfabTu6tjArqDY8VFfZ/lpjD
GAPRk4cihpiZfRZfGCiRkUCMbDqlgHrwMWtbGeEEOYz+9OjkmntS4W/ZhrXMUVzO
TlCoAePlwONXbg75Gqqt0NFutYBHYtimMWWXXEJanwBqCLeyoYE62KZUp9haUR8Z
bZKBqOjk3iTtNWlNNMCFrdvaKhK4YgX1IUWWK0aS9L8m7LsOdeq2RCsu4Y4vNtU1
be+ms8OfUvdh2l41yKkuIOhii/liqhoNEZ8IRmz3KMKeExWZHEBckRvICFHEL+xc
OhAeYM9qRlIbPf3aNuNINK+5+NpGMVca9FkNS22D2/7+6KyD30s9eYemBySCMDE3
+xA2OP62G911lza/Pxx1GM2YeObcsVg5Z+UsB0JD1539YhYsnGRwNVjZQI8XtXzH
Z47r+K1rOyY4yfCFfeMOq2qbEpWNgS0HN1PcpWI8rb9nwHLUzD/vT2qip1bx7BVQ
Al+T0CmT8tO2um4q/ESvJfzE1DLeRHERw4CJ1kqQ98BDmNnj8W52xbmOFSYzm/xN
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
mrwQe1+XruQOyKbuj/fjiChaGpvuVBaXHIC3Qh79P81yJTCPGiKtNzNBZMR/3nZU
aDCSq+GPLBIms/vU/+DJ4gKlg1aRnseXI3ZGk36HRGgXy5I0BQr1hm335ZvDwghh
yu9sbK/8A2V6Ze00bT6CR9Ria7D9rl/5LiNVzsOks+4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12016)
WtFglepXvPpfeytXf5SZawJ1PPG+xBv9jXC64Q/iLu5yjSZE5T5jqrzOlQjFNhPY
EgQmDXo0CHxJPLX/8WsJHOtrD6d3qTVckb9eUbSDYW4UyrIhiOEFzVX598jrOwmu
GfN2tNvDDEeeJsUFKudPMXvd8Ap7p0hniBSNRGFjygp+btv2dlDCrgaBdeV8t9Kh
gMmvvN824jJS2jL3soa8ngrXICYELCL7IDkNa3Wd0/j2KlGIk3hr2cavV/p8gKMt
spHzOelqduOkp5NlEO3RGzfh4tv5p3EGtyGIhH2AozgER0IMhQIArLN0Vdz8jZIO
gdhgQARJlCyxCXPJCb27YFAO2sYDvWDa4GJsXSReDWBFdlaT+keY9aHJrFfosy2M
/MVK/Utd4j9zitmmsgE1gUnlCs8PSmIOA8ZVotjJidHQMkOUU3qCV4BhHIqVeUCx
BdpYKAHiDxdc0MGvB8h4DAoO0oSHgFyGIyon6tEXK1OlGN9xssqp064XXmj99ea2
GCabAAfunI6lpj8/JBQWZBKVJFHQkjhP2d8T68Azl0hZSBhcb0u/oA85EpuR+eL5
GG1nW+EPaT200W4fzz/ppzBmDqHE9XRGO7K+hX9+f599dsRnniNeJRB1GfV/CzEa
nSHf6BQe60jIIZ9X1HU2DRvSx++A/ZBJriZAXwPWfQL08eeepAj4jfid47N858vS
mG2cxgO8zopru8Evl2FmZKwHlit7HA4EL89qfrSDcEwSYWxacfHy13hTjOSsGG9l
f/S9eph8OnZkP3lzTqpEN29fLcSrkEPMBdQ08XVXztrsZRNSZ5s+djdWErFUBMTZ
Lp97Eo9a6l4QzRxVgaC6pqNU8dldDrmYsJBXpAqnMpJOXt7WbIADNr8kg0T5N0iH
fRsqy0EKsKUZvJLldVZjasufXpZnz6hT8iXEOqtUhipxht4WxQ7YUyGlTTqGQDRn
T+H6S6NO9zWczz9vB/8PNW/Ql/NdkHS8iYq7iDiVzS9otxIJvp8SIYIoICSUJHVv
4Dnl25H/xtcbQigkT/qkWKXNLbboZEnnupSlqU0z5ZaasIFk30Xp0IP15o4Xupck
vr8UZlpKEnTcy4R/PsD7hZo3JrAcwAhR7JEu9553Z6S/qsxM+DzH03mpgBJgKyM5
ou4OTolTwCuEjtrsruz3Wmd2MzVJbzvDOmA0VD74p8glcHZPvCeiz1QbyhSaieyj
mKJczOov+9k1lYuQ0/UFtwbNg6GukC60qpAZMdgQX79Qll3aCyNFkJyp9TnLJyds
4uesrj3uKM8DKBOZyXO80TO+9SbYuNW5E7VQRI5oHMg4YBy5kRl052Ts3wsCd7ZP
dKkrBgefLrNOpH2TzlCC0xb3JvI+zPSLkTu1xWZ0BldAkzePDttu5dGpO4nFtJ2U
+t3YTf8OZzscjgTiXZ5ajuIqnQ9CX1FM0IWAkP2ePPxKhqXIPJ9VZF2uhmZ11dcs
iSYA2BWIADFYb2wQvZHIpMnn7iXgGHR+0STNttqMtV8gbRCM6gcrzpT8wYvQ/GHW
F484W3tAAFz9LRWMEbIr7b0y5bMsAzq4oE3lWQJkxoqdJhOL7D0wpgG3gsST/DmU
k+tc8Tor0uIhjI4v8VHm9QGCMMv3oXcExN4w5xUcpmuYTkuWTbx2GJYAWnIxuuQT
1j+Bhx29qpApl7buTkguvr7X8uysELLJ01aprJtj9G1mMDiy+DDLJjVlsLI+l/hs
6dJ/gKM9AeGRoWdy1TW3bSxA8xsE/ZMY+xcyho8Zpo/6f7VMV9M4Jp3vH3lPBITB
Q5yiW3dmrNUih38nmBl7sudpY+W9lQyXNYQjKUVdUhKcEUF73JdiNKdo5goIr+nh
+ttY7ufrS8xzimTfMgk4PvwCtsjImNAtfW7c5053xAcqmxb5gl/P5IwDIKaC8bB6
H/c0pr8y1W2WuzajALMzIMZiXu2smvIPrtPK8Zw/Q26eaqH4l6VTjT+6BwQRINzr
pYQDe8APn5yddyf2MifkDkn0xJjPMx1v8SsIIGU1kctwdgi6kGIxXj92bmQvlWDz
atrKQAhwEVzsAxNuvn59hv+26Q7RDYndcBONW7y3QDybtQpnSWnxxFFLH2b8rfVz
JVerV6/rRjKt4R/v6+ImeFP1b+Ad5kcBayaVHtshx199QHpLTJ61YNqVJVQaHf1i
XePSpPVO28ApztJKHl6TohygjiujmMvTfzzdhQhV/FrQzoOGd/k4a2N313xBTk85
0LyIxwfxyd7/ggUE8Pd2PBaHnxX2IpDrOgjMSumpsjN/+PBXZntenwAQCm8iUNJ1
Oh+aNxAe4m8+6zLA0bwkrHqob38HmB6pEBACzNqyWNEszcKEoOZEFCSIiGAjTefM
oIOnL9flaeDG2Al4UZN52qau7Y+AzUFo8TO/jKDmDzl3tyIjqS1KeH9SNkGRsBwn
oca04Q7tFW/TYi8M4poAiQ2ekAiNw6nUS/X5C++pzhNks1ajIaS5G9qfZEkQJRQI
j6RbPFQRN4VTjdmkp7gNsIsxay+HP8tKSVIMDiX50D+BpWXBLQmW9Zkjrk1wVNQM
l2gp8pVSnG+Vqj0YeP74j1Im4SFsgMc7EhoyQCFe+wBE7RUXjYzos8/h74A7RmYD
FMfpuqB0ZQz7j8guQEZigKOVl3uunCPbt7DGpLtYlQP3UNIvOqf+GCVs0Me1IMIV
ZMr3jZejd1PMdyWSkdt2tD5RMhoXDLLt7j1lx2Xqfb4sDJa8a9jXOmch5Kp7sMbg
w/VALcojm9MDnQ08sHG/QlY+VLNsGzqF+tU2+SJ/rSkcBce9WFxyrSdE3M/iZ0QH
5OF74B1sq0iGyX2QHuayLl1bAUDe9VMa6QCgXWFrdpWFAzd9iPs2LGNSy4VG84ZG
QwkhJyksIOofdfTpcTK8S/HANnl590T+T+dz+3VlD3mNuuoe2/f3zyV+XNW2RuNF
CXhm/pY5p8hnc34OKFDcIvjzefCQzqROkJAb8Zs5DsMlicsQmRstxjlbifLAAHxi
h/icTR+NZYbfK4NJQcnFD9SHCNHXudeb/Io6hti8jJyGwmdMD/8ogd9MifCmwByw
RPvny2zgFxSISQqAVB5p3NonHcXO4PPY7ayNLSDPpf/SYGh2Z/VW4P5cMaXSlvBv
gYb8S/YkAX2irVmj/D3ubC+iIPrqhZTvXatSAc1ys53Nzf4SSE7VqMcKlP5mzHgJ
vgn7uXphCoLMo1A8i2CnL5gSoLhyRxeeG2aLSoYo3RrVRt+UrI7QVpTdmaFsLCBj
O2AXm3edsFnbCf6HTrMqkKAUx+FJmw2agX0dLerek71mf6KD599ROHIQr6zu1Egr
eoHB8o/b/IKzhTRq/hx0gEim+HjiP2NBOFSHAUfZzNaZ33R1FRhedWoh3PrYeScf
pNiKj43KBWMcAIcktDknKDc2GSu75mn8pNBKEryBhB6kGrjBbA7bU564YNb3y+J3
AAUncmAiAknM4+L4D5UVIbd+jNvustn+hzd9PGBRc/3R6miUe5O9mgpXHXQdi+vK
Z02UulYJdB1GHJirMFEwAWDGV285UO+sF7ULfyXe44BxngZwxShqTU4+BVlvJECk
kNSnfyACD7HTMNFun2mNQVNS5jVI21qO7+lUx7hcT52RRe20mmItZpv3+kD3k33e
P5htDBbgrdk98nAgnem7+eKOOxqRLYxqyOskmtewjWZch+BecVZ8nQvD6WmhxBCR
HwOY4FJd8S6e2Iub61GxTzmEI/SHjv+odDNCCT+PbCT0HXlR36boMHzV7xztRNAB
fear2BEJpGTBE7C7QiFTb8ox2bsictq51fjA7cINGLMH2DvbpaOCgp5BLYWsKGrv
28dIT+W1wxea+XWwGKxFM69ZVnIa6eRxj4WFVLlK8kvt979N+fLOdF3IuiH0yung
OLxIIG8ZKvYoPu9d7LfosN8YLrZ1BZRbu1HqlzveTnLuc8HCEg/S8JqLXKWDBWVZ
EO5QUa/OpE+FDK9iJpV9D3nl8HBFvAhEE3diFd/IvwynJRqGhFcJQXSPrGVP8QV+
03R7dr+LXCg/Ll9b+vDz/25aPp+5xli1mTiX9+6x7ci1fuanGkDWrpxyvKCt+rXV
I8ZLJGGHQsiuspbS8IgJomtZXPuWrfR/5qt+TfTYQHHSSrpuafAIazVQuJRJBKuh
z8htdWIFn/k2YDhdcO9/wKzUrUGD3sNZWNWsMDPTwiHSBF4jevOE0n4lryZG0eKx
jOA74lS4IG/Casl7Avkf3NzFmuGZeTCQXWVaXDLFnxesFgwTVC4KcE5hlka8ujRD
c9ExvZJN+j2RIhV3RD2D8W32S8tpv2zjJBF7l+BZ+LLIg3rTigk5ZFHbtO/F8fUb
/qJGDDqJYPRMH088WoHMacn+kWa4WxnLU0sQ5OaHS2BMtQQ2ZR9Ny5X0GWiZWNrd
gcKMC/UpY25/d5P55tZlLlnyME2MR3hoEok7dFrQxr2CfYvI6wg9SxwWlP3V2hi2
nfhJL9lbYcprCRuQpS9P2DlifTPsuadfsyTTTx4c7ihXQFOn34xEEl0gM80zlvr1
c2D90OUFRgThTxz0gd44qYq0NaAtT8hdU5jmGnInXt5BNCCfIQWsYQXN3X0Wwkhw
iIYXzR4fQmuUJEZSY28+5lpjRAK0Wf8Hjk+fNUdu1vA5fF9RMpk7twbHlE+MS2SA
DHis22oli0IiNbVhzkk6QoXvZ2Z/Boat+HlSWSLDJyFnMQ+ztk9IdRfefdtCNQ/Z
OFD/Hq4ZPQ5jJ3Wqcuv4FlZxVrPCxsyyWGZ3IhRZoE3vrIip64S5ZXCUSnzvOnL4
od7/J5P9lPaGOcjekJGzhAN5xwHizZ3AZHrfSeWoRv1ieWftTHtRGZgPWlwOh4Iv
4F7ZCknWy7ykgThqHcl0DpEKyN3OfVcD30diC4tx8WYdOMEtH4Rhk+yhUleorhIu
Y4S+wBBjhgEThr1MjxH3uHLtY+ds8oL7u/LH6HPqV119BCPZRhe1QgjJE3QVaORQ
AokJewpkGNw13LmCeSmvKsGYc7UQBBFDB5mFQbkd/b+KpXOh7Srr8OsorizSgh25
jzZQKbugZbGz2M812+ZT9F7kwXTgHQw3DPn8snDVakXrYXR+JW224hwnxpHw9jWT
vZzhu64Np+4Kay7jKEQEvbRfAkYIVe7KB2ujraIlkK5W7ckfmfjwvq3C2IN8yftw
GqeGuGu4nnHx0qSHqii5LZWWIKuqEK5mLFlifJsDS4aMeSiePf7CAWzeV8bL8Mf+
67zS+QRMx6cFVziSND8nU9qq9TF2wMYJs3Am4TUtHfaA1I1r6IjxTyR8rSSOwduT
B6qnN2ttl+9sj4ugiQGKuuvTmfXoM/U2N0AtYPgVvnVGhSaccK9ESRhMr6uyx5Hv
HgdjcoVHpBXWtaZmk6oNEMAWe+uu2uspy/UxriNUO1tct/H87bhPdyWrblKHWVU8
FPpvjaYX3u9dykzp0T9ifLzeADrZzUgaMx4Xm70dMxu6ImF2iDucpLidt7y+alXc
oSdmIpw1JPo6absJW3qWQ/yCaCPMv3XJgwM/qiHgEsTpOaPmcjpIybATFjkQBA2m
GADfryHRJGBM90uZpXNMtseB95DSiyOE+NALiFO13GbAuzuTkDuLGHNuei6f+Mwc
5Zttb3/L6bvo7m+/Lv2asHajo9H9cEnDRp6L+BOY0qSqtwnrNaDMdpeVapsXiZ99
fZoc6Y22nU0hLD4vK+bkqPPys9YONTU/lSLJZ/kkvtkLNGyqomfk79Bh53VEkaO7
6bQv6MyJqOSXQnIjvqUfFs7e5pyHXpVfrwQT/HUUQRsM9OSLKEH9L1R62fBQpgAX
AXv51+4M2rZHduBEwhucBB9OpNNbajjMV/WVPjXzWbGT7LhaHyvhw1cTyPlpbwdP
mQUzAnvg9YDa4N6ojfst26+2Xsbshkq3QZdcEnDRq2YSz9RHbFyuH1zXcx9Tfobo
BlF8puiIWFwlv/dzMX4X722014ixoHrJLC7Fx52KTXyEC9bV9yZRoSmJtC8e2l9v
viHM8/LpaL33ZrdHDLf/1AfMYaG8NM5+P8+K69Sr0oR57yDBTHJ/DfEmlBH9fHvl
jGgy7jt0cl4thMuvY09+joEzzeWp/XNTfWpxlBVwcyVtZn9Nn9eGp/mc2nKKbqVQ
eVHNPFDNwZl8jv4JEcYK0c9qdH00NxAedcDOzq1mWeiPyUYu6Ahbi8pWLpLLzScd
0X2PsO8/1h+UNqgg1FIbpilf/gHv88kEQLJVZdJjC/eVXK0pd9wJaPjxTczGfyHd
JZXX1DwCxjFKjyS59pBcaunQo0tQZuXe2cWrYtzgSFJZWIUZuPf5K6sZHSh4M0yy
x7neSsIB3yYACKvBSu1moAK6HHVjyyEDDQeLPe5AXTklPcFPvLPcBbx/AJ9nRmqL
oBpVbZ7TA1SYZMhDvzTkO3G5KXtzvF8zwN4e40yoJIKq4mraC8J+/2wlZ6av8+k9
9ogQK/44YGBrFR8OJ+7p2ZKtd7rSASS9I//jOMg+3oMXktaKGgFqTnmT923LH9+2
OLF3b0aSh2ZzSRJ3XCpmmecBhoxpUU+HKExSvoBVzy75mY8Xon07kgBodfikpJCu
Vf63pS4lzerbAcZSIreDKGPVXR2XfY9rucZutG+dqtk/vSYpQYOtDW2vbz6RTnkm
6Nl4j4vY/Q7gR0IZOX0uu5Fvw902Hcjx3GA4Y5puPjFT9Sy/8JnSPCYQh4GMarRE
2UOw8jmTqpT2l/ZQdYEflimxQWr9erOK/VShTgBJSGjdMEMzoRQwXh58Gm50Zrng
kz6hFBC/EM3FtLMHWqdm4q/q1RIYTRGR5rj/eO8vndS8vWz27E95LP7aGqli1rQ1
NoIoA7lF2bTTLaMSxKE/zvoAlhPkHGbBLJnyRlGMOgG09iMiHkzzjnkb1Qrml++3
k7vHJdtYVKA4vx7zcJx6j5qudY2D/n4cWfIr5Ef6TKgfpCFD9NRfQSEoTsj3zpJC
Rndcnxf34Uex8em7bGkv69mSFfKc0XsAi1Bge7W9pSxyx23pVvKEozLqvWpSrZeo
lF5u/r2irqZyeCuwaW7s7EwW//n05b92/AfifYajRn8IY1BBn+6btqms4WHm472A
kOk3C8eRLGJUjdQCObRrUAoeom7YyBH8GVVfGs/yIOhOBUrGHuhCqq7TDTC0GAG8
wiKKO/5gg78/63ackdGgQ3W8/PHzlxLeCAzEzfXKjlGczPfVwn1u3XYnFGS5k+UI
MZeU0KNwQy3q+S1YHHjOM2e5OyJfCyPDPz1Vd3l5Lmrijj+RIKoSK04tfuwGuDXo
xQ530MPtzDoPuMXjUtS9YaTOSv+wcPj7vA+HtyUSGS+b5cNloq9WpwWnDKIgfBdT
DS0fy6dYhvdWVqEXkjqVwWCRkY2NRzbt/xtgWrHJ3+PQs3/TWzK4UvSq/tlpKIWi
cRJ++XFJveJzpur9mRyJwkeNILH3oZsC9NN+MBp3/RqLU8jWeYotUtPsCfXJzcn7
OS8EFC2LYcW1UG7Z/0n/6Xpl+ssAuCVDhD3CojZmoxrjlbIA4to284P9j2AFN9DC
FLA+t2vap37RxAclX7dzefI/P1HQSlJEFcbUO2XXiiNvMSL+9w8MbZwTrt3DtlU0
tts8FK8qufLD6F6vMtjRDQr0lcHabfB8JvvBjCpTR9X9UEWZBE2C2medBN9SW2R5
6Rl1vQXVUxmXOJRox6B1/0BPUmvYyMaqPe+6WpiXVb29vYfIA4Cb/TbiSCBY5roJ
vrUuDQP7+GPptlqyYU22Pv+Vy3/qFA3CihLY04v7mnwjHFdTOPrkS/BMeXlf3Onv
s2cjDrnzNbtQrvZWGlLt/uRjMUqnqOjrwJ0GjgxqEO1VrFkdsYylkPBCteduSnZw
fW/WMm3DwLwFj7338ueZmmLhECtl5NswpEzXgFnFzH0g3BUagIWwVq4S4eJYOKcb
YOqjnItB3tv+UkYr3ZPrfHoSfHsHgsfQ1q/e6+NrjjI+9U/ZssOXBPOLl430RJbX
i4RhCBx+mul9I7Jiep9NMhgRp4P5FQlbVX3IweeHksyU7GJ/BxS83r7lcbRBm1g9
4yzVN7JMQsGXw1xoc3cBc1gQQ95VCxU/2bdxYlL+AlApR9zVXzPI7WPY9tY7gvoU
obopMEo109nJPwsSWQpAj3z9UO0OQ4M1m2QKwZksX8bxiy0nZ6jF5WyzAIArE/cl
z1HDo3hsN0e+aH/hP3152wENoZopgaxiFHKrSQavYIBmL5fcRdqCs6ffWSA33gCR
z5MObqEe68Z1oOP7+GpG0d2GVIMkFBECpzWv5VZo9ETGd7pOeZjnt8Wh83HJ8Ts0
8dLqAg83k7h+i8Krofv/mP185R1NI3p+BkGkjxQDHNjORWSEpWGDeiHIjB+jiOMD
jahpOl72GXkqalL/jS5al/u0Ui718A9oc1s+FPsDfnrM4FMZv678Hsl9My/Kg0hu
33dcwLlr9GwSOsd6yjNkpFO4tUrUyrxUl5eBIc12vgb1/YzaugGfrvrB1ZfpH/9H
WXZfAEr2WNfxNUlACsV30WGCrpRzM3njo9aT0XmEycBRFiXC2DRAgui9ZAgui0Cr
5dMqacuWYMJQeZmatJyLTHkGiP/tEqQEUhOkJXxCu2Hx+Wd5NQYTlf4agLHoHf/C
7vsKL1PMP0074q9rfrtrpomY6xKZflNsqD8lgpgiUAZYeBPhnJHhQxmUiI1G38e7
kTWalU7EmlJaIYHbDsjvgnovSP88CoKEbnMEPFwIpydZc/dPDASkcwNSe7J6Khfs
RUjpH564cNLQhjs+pOfZWj12Vqmc8EcQPMPvJLnxtPvSSmHLtCfVtKcygIOzHPJ5
/mZwx4+G3gQSJzTOC9Be2tcgXu+OrV7sXwBUu4q357GIIgfCVnGq87bRg5L6MrK+
EGK7/RPlNJc/RyUlmwEC1hRupFVQDcQgrq++LAqbXVkR8Z/zP8F7dffTpvKdwMs8
AUwezjJ250qZ8U4bOQ8WCR2fYJqUQZ2XQW/scQoCHPrcillKL7x+QS694YpcziDt
VxScK229SthZkECRUUYuf5eNcNeSfdXTTBEW+Y6IgO2FEZX7L3rwM9syNX9swmGE
vZe80NTl7lIpn1S2au0T/9+mWqSndumbzELsCN4GrczgleAlbGntIj3HZCKr47gv
YVvtdfr1yOckg6X3PVobWUCnEXU1E3tZ8div/9tzCRfzoigXa7JwMKiZPljdZ8LH
MtwT8eXOG732lvkIBJyvBfBeJSaqWTgW5HX2O9OiMa7Ke7SfhcdIBM5Bgt8HB4qJ
ngA20BYYH2o7kdlDfDeugAP05+7jw0zzkB4aH/yWJTU2hPdnqeZ9G6uTRcS+X0Qq
WsarkZLbSn/uokwn/m6JR1SLeQtW345DQRJz/5pnwRAzcb84JzMYagX06GvAzaLa
Nk7rMVMQCQqty9wntlI4R+nQMMzDOFW5E1Fj1vDUoouMrHmdBads/ZMUGGjoY1lJ
A5TCxETLwgrvHIEfRe89nY5ftXUKLmUEmZRNQDxEATWeNGu73zeglicwOk73UEJL
JhsjaNy3fou4H6lHCx0tuh0Pwx7EFxnnvpYx1w99E/jTT1usAp+MYf4blma2iFk7
SbjsG8z/1MlwO+wcWy5XRqAeqo2MDwvGqxDG/fufCIJy5kCe+OpnzL/qxF2vJ+EF
CwluseYCVvArDyTyEO8T5DPhdvJMyhNW7aWcMWn/+OweotgXWVDzYDI4ebkWzn6b
e5hC0nPPGdvKt+UfQb9vQ34uJNajO46VG6jtFQY1AOBlat5OFPQ5goBH2TiwpFyO
P+wpYi8iQ4EvSMCDQdsANn6mRS19N3tbZR6DOFES+RuXFxyZXR55HNEV1FKG3U51
JV+fepgDndHc0/2pcsJrUoTDSwySmt0ZTLmc78CiDcIN2nx74R+py57v36i+gZDO
u3KsBb5b/MFhMiuUxXJ93hZSM22q/6uCeboo7qy5N2V3Aw5zrv1lmjn5GmqGpFrW
VWXl1RKrxCJwctjcxSUuVi5mXvV6w49chv8qtbbNOHeOQ+aNqHwqZigyq7SszSQi
y4HdDV+/bD2cDkvthhPEFAcEqCNppwnjo2A0n9bF4RfAjsvNCufonhGItGeTID6d
QOtp2Sk24jtZMtG6OyPSYDp/0eYCJLTsehAJcPCJsPJ4epGzy/pcbIRz9Lw2XJn8
DaDyLv1bfQTGdbDjFX8T/r3VGgWFdfWwktGKhcwsdRmJVjVwn7+HHn0AEniN2HnA
WIKhfUwwBj6a5Q58tmWzOUxQhn2/oX9pkz0QG/SS2eBY6qonYqt9pQc1nAwjXSjU
gQSX7Ity35JZrfov31FV1gOnPjU712xnHvpz4Vax2R5YQCW7+dJHOHzCP9p6O3RZ
Hf1pYLcw+TqxyfqmPCnwOkYkuSP89SOg8vVqNvDpWhGhngF+wHk+vwX9nu08upQy
vpI65kGbBGjyiPBmal8/niWSe7A1FHV3vnhwIChkNoE4DV9g4pncCS/A6HEStClM
khjU0IeVOqLALZXBS/PCg7XZZCIzuRdHH6WwjRRRsRfC00/wrv23kKDT3VrOud89
AGXCCKAmBVHBzDN1nYeLgEjDxXaB/Kv0w9dB2axrklKL0Y1xpdReZcsOoOkChSJA
PVkkxxzYG+HLTuZ8y/sjSRTRcfgovaq7rCrtKVmwkTQjK+X8CGaaFXObrYmARbPg
OJIwx7MrKnhs2AKdzmI1warwHGgxBYBcmM9Wj+B3xwZ58L96bxhxRnKggxBsAdow
T6NcRJ5GAROgYyQE0UbYS/hh5geaJJqruZrcRL+usED9oX38i0oO5gFcLgZOegXf
QbaTabKMGv5nGGH/ydFSBCBkZzHXFEB/9eDfkqjhw9tv6eJ0uJaSWoy0fdMIVESw
5GpMck0FLjg9vOUxUczCcxIe5tSo71sHeQSsPSxlmoPjuDPYkOTGQOiA+zgTK2Tt
49SVWn5maroWtf+coCZUxY9slAQwy9d7SCxVW4a32LD/zpivXg2uBWgapUA5v8ox
ru0Snaic+HTBydQW8wCmgWeh7PYCOabRnEu44TjIg2xOLoGEApveh8mDlKT3LeFM
JYXtVM8gHkVlJZ52XILNm0eRxX6/eHTJ59wrjhRHJ+8RBEO/KZWdGJfKZirOkDiE
ud6B4xOGHSnpTQmvLyxAm7cm4o3WPUlZrmYR1tutezbHZM59HDMYQTJGetqM7p25
wZ2W7GFYm2stEUAd0Yd4dNDpUxWny2ZDVWJWI4cXEOZEYuX4sXvJlZaVuzZaRxE5
4ulmQlYXj/8eqvBjHCrKFPCuppgeND/GrEM9aRugrVAUhc5EtXeywebriXO5O2FK
1aULNP1cDsipBkEw7Pk6R2As20U7BZFCxWuvjKjVTQDBYaFxh2L/4icDWfgL0rlr
j+P7dQkgqqml/39z+4rbTmEMu0cWMH6ySqTRknhKo/VuiZ/qJHRY8VN/l+SQO29E
/XVzopsSEVrk6muK1yTmYpKg67aqeoENKka+3ByxyRDvm7OnFzV8SxeyM5r1mmiI
2ioIpChmDQXFjuD5N7+zdw1HsrzoHUN3P1ltWucaPdKGpsDzRPTSPhW6f0JFtrMK
rOD/2WFtJPWOtGuZReRmWEjGlUO5NqSeRu2wpxKGC573D/0szQQb2EDFKKio2dJo
QMNFMBPV0A0qZbgKFeeQH2jWygr3UwLucfLN+BfOA+2th1VsfgV8YyBiIc+395UH
gVJAom3MaFDlT3l60jWDpUC4IKSyx4ZP6MtQN7EtbEus+rrUWbNVPGOsR/akT08i
hKLp2p/cPdj5I+UVpqR4OoDkTNRKWeTG2iHCJnpHL1/XUSFIMVljo3xHKirJZh4C
76Nnz86yqs6H2HtRFwgpAXO485Lp3BKci04Jk3QN1sf8YY/O05ZI/Y+uj8bU3DWj
Ho84zoFka4rNDocUWiYpxMues+Xh54aLizDAAUtosNJteuHwxFXe57/mOaCVhRdH
d0rrqwBBlb23JHqfpctyQ3i+OqmLjJPWCLjaANcCPaIQ8OF7pUUuq9IowxT4Wqv0
J/PQLA9nVnZC1QTRJ92ReeteKYt4pls3a/ne+dvrrBO7LlLvU6S4Q8kzR1hYUlwT
Dj4TolgdHLoEIYHvE5x2pLG+iTE4H2NTd7cexo3biuVH+Y7+l5mpbp52ly1ij+rW
KEpfYO0TAWeFhbHKthc2RXg/HQTgyuRp9QC9vzMkSu51KOBA/PchO6u8tnoWcD+P
Z3dptscm4UtYH4qKLAcTrG88HV1xrq+8HlJig/QOk1Yz+gkU8zPYUK7L2tPCkUV2
LQKrtLLSKDViOrUkf2eFJuzfimqumQAo+DMLxYIKY1k4Wj7DmxSvlg/2/Uh4SeCu
SRQN6kq6CxnzdLS3fCRR0g3f0XKdCwWI6+4dXRB9AEWTDNDmXH8m55IqyttWEvx2
QY9bMxMi3urGp8m4GXJbmIR67wpx0x7JtijjbS7i0vo4jP1i6kQNhvQEwNFVDSID
CEx645G+sJkXhrR+lplAe2EYOKtDlPnFlxr44ELvDzQGkOwJRBy2TR1G6l5/ARCP
WTtyUDfn5XiSWZjqWWujCYeZ5qiwp+GBHRSBeTnp45xfJ8PBjpqjCol+9ZNEPhpF
yHPvTT2/5surwwgbeHVQT5IX9SYEVcURICBZ9jLQJNr0Vn3IUQVUck9GOriIhyjr
ooqId21tjCzVQWvlT7JSAqIX3KY5lZVvx4TXi4bkBtaSOBaU+vVNNsq3/bWgCoqF
xpA5xugiFC0gnWwe+taMXgtwuJAKKYWzZCcGFly4dJlcRyzp/JD30XX2rSVP6aCz
j+wdmWpCo/hFxNYE3vtLCQXCUq2cJKa0nqlqiriJOyQYQHZtR6Q/zp94Q2bqzx8H
kMnjUglYVxb752XusOP5pPBP9pM3QBDfm9CKunbLK88cy8Y7vSZrECM7IwizN5XG
vBcu6VQsfwsRiU0MYd9n+j7BgUmhGfDp4FXnAWFP8dTJVj2JlJBcs9VF+k4uhVDp
+MimX39QxZPHl7BoZohB5LF2NQxQbvJgRkJSkxC7evQZ0yQw+/eXdWdEzorHR/5e
GOkrZQaphX3Jn23BwFL8K1PIZilivV6zcAvzHXI5gJENwGRlMjkhgl/EeqscUQgv
FC/QBrmxB3/MCUbbZFYCaYRVl8O2vboWFydivpeHlM96fVYgHgjG5l2GSGcVM5Q+
EZ4UVgR0NjTO57OzMjKtsT0hvdNKAQN2BOQlUdkW37VWBVwynXCMh+Jes2hAbVM8
RNOVDNR4eQ6LegqIp3690RcknxO+dsD36dyI4c2dTruKShjj6IOaHE1sia5RhaUF
vjQByjEsV3XiYPp6qcX3NZ8RpFAy+FC2DqBkewpK8z7V3McbdSOiFVAV5eooRT0+
3T0lWgv+O9Ib2+aZ2hHON5wjWImfaMqnaGZ8MCoPj+mEi74Mp11Em/dos3sESU+n
rKdDLfx1ArKM6wFjz3lWfH44fofedBVLEYfAICnsxKjtzyYWl8wnmeD4E2lGYC5o
EskTPDeXGt4ZEVGX5swH1c67A9Jy3og+Vy83ghWUlVCPnX64Hm6kbNnFlX+/GHKm
iLSvhHNj+X4+OCLoED5apxcW0SPSq2VT4BDB6UPgqW5/wnFqcXx8SWCuZX/lNbuu
JodqzSbtWk81CYKIcyt1ruclxeWkFz55DuoZ6QFEd4EzGstdFWwyXl3fXnStAa4W
+0zXomZbhX3dgoioCzNipCGXG0g3DLZGCP9HZlPtrHlTPB03jmDznuuSuIWnnKkj
JfyFj6iNgba54FSGbh7GA0tRRXIV+IuWcEu+2utqADTpgGunT8jjHNltUBGPLc5x
CpeI4DeeJ/5usMqZVsE8IxSQ9UKgXtAe24n7oN//6xmEeutbfcnUrIDlTy+9Dfsm
mhr780KNY22lqmqQJCYNVifnioVv4Rgd778Vb5f6Qq10e4WPX9/1zbbWil24/PDx
+j4oPtX27O1YoSBZuEHxYAO0Ul15qHRKpq7X+m/gmD2T2UMw4lngYABbAmZsrAHk
6XQ3+zfzKm5AwqzdpvZQNtNK3mW/GBik9UyL6A9ybh1z2p8uVhNXvcdv1JUr21O/
2rB3Vn5mRU/S8R4yzsWKTvGQ/xW566RS45m6T3VSNIYsH9HrFzIzKVoB61lSUZXH
rMUVG3tEHtwQCSWLHM5I+dLA/4aIXT+6bqBgGrVprZqJkQXjzq17OUX/apcf45c8
4OLug3f8hOMJORZVP8UL58i3B6ysbEn+4fnUJLh+6XzWC++ne3SgpzY/2fftpuQe
i2JKfeqLfVzW2j3E7S1KBn3ZwhhzvpnofbayXAInkRTN9vtM1WdsbbkzZv9h55+F
6GZ4dSVVRjuRipQdNqvdLV6A3PUHbgJykOFf88jEskrnu7q0tpEtGBKM48uKAVc9
0eGJYVgFMb1ZpRO+R1zMuymemXFU5U+ytTcsAFQvKNXhHBPXeNxsTPivz8MkYYFp
AT3CnJybc8jK0YmhOt8sXbyarGVhNRsFBIEYE913g2drnM/iFfzDWu9wScemTqPp
aeA5aEpBFqwWJPz5EDI5FHGFN/DzQTumERvAFB4yTCJjDL3SKJ853t6OZbcfUloV
kgSiEJgjyP2cJsRdTL2pifNRJtyZw969IiHij1A9WyCIR0BeBoCxyWBFiEjFyIf3
i+kwK4oKPZrSqtRQ/lf+21NcL5lH2nEmAc3uEyq7GoP5WvqkvhrNaIyl5Ac4U2tU
jAZYA6WX+BpTpv9hlATs+2+mSGD+Rw25CMakZyfgXgKB2caDeuNFTFtyIqm5eEjj
Fvb3ajzkoxMmtW4P1+zL7r+6y8P0iXFONy2CAylhPylAoqkxgqggsxcqwZBsfggW
ubKF7IhqOq1sYnRFHPsPirFDxp6EbM672+lPZpnswSSt65YApNa2jA+On0t+rGHd
FxPcfII9kwvKtt66XspmeA7dZOoVHmhNLRgRfoR2bFVSccHP7CuQ29j/ioWpnBs5
JMiCQQZUGEse4JucGDJN2KRP1qAmgkf2VZ3SSvUO6r2AeJFKY1uu7KlJOJtoPLC8
3Hy0XMG93jM09VZvQoWPd6ixb2WwqxLaSwmdJqE730Tbiy+5CGAWig2HGSmsa/A1
g5UC2rRqxbIDC0IUxE5ojnSxihdwcJO0g+D2pm0s8V0VaumyOdHPyPvIt47ZZWkQ
TQpBs1fVCS51X/dO/HWDTUNtd2guoRe6As2NPScNgQcvavjLSXFcblpTto7JY7qA
r84l6I/ul9sQzHeEGDKS0YeXQcTCHKSv4p1ossnQY53RKzY6Qti2xgeAgyLPdg6x
O+nnlugxv5EvQGs6Qo/fq1advYGI/M2YaOIx355E1TJsdl0le8MT+XqgU9jzG6vR
s+ak+PzvH4+VU3yy3oVk1YUAo8RNQYYcPm9Dxl9jcw7oaxM3MxxA02nL0v8yeofp
VyAYT+hQ3ByFSlHAqkmZbkQAuejzab4x9kxQRkhfZp+4GbLfos7w4UCAcgFn5TDk
e/oqHlJbLXIpjFTvPD9BmqjqD0nEOP7wvmGOe3va1vxTul9CGOx5isH/uxmBKqyR
IUNUnpWBlEZv7c44V8ARvGmWKDSkCrbPBPbnx/hFjORrTj2/VzTKmkqc6qynQmo6
HOc7D0M6uLbKH766pkyNZ3HHDiZ9jXhTNhFhYPfPz33ndDrg7euTuBze2Vw4QBvh
EJxpMyIa2vHFHAAKn2hQy2Gha8ytot/Wp0Px81OKqBWRDYYyrkQK9Kojzhakh7og
W5vRyBAya0DY/CcvQ4PsfZ2p9mbxi47Pp6lDqygHy1y8WZLPLVAG7IU++RsShBMD
O/2xjHUMDP8UbjX7Lh9UHt6nmph+dZpZVqm9S441JzSlMecJ0TtQtCjI2GXuoq+p
F1hbvBqtaIExoeYI4LsH4Dpu7kFApJxPdLv2amXfbLnJQhMOq0XWCDoHXnbL25kF
7d/0Jc2Ef2vG04NeKugf9JLkPn7W51aO8hp2YZKUUZr6/DC46V5cjlJcYgQdRTwu
MlF+oZ8c6Os7tT9DqGKIfA==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hYUMDAMumlcZgtwEaB29bKwtzcNvBDZl9pxQck8WlWLiMWbIy4iyCPQ8djgOazZF
fQEWPsb2llGJAXDTmGeFsVIuuPMg7A9pR1c4V7qHBxsJPLEy4TYaWKF4NxhpcsKZ
zWQpQy5A4U3keiIv13RV3L/5pznw5JR3UtbcGhB8EC0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11392)
ELnv0IcMrCKSkm+Py7h1+4rQUf9j3eqUnu3YZcfDdAtkJP8kblGTOG8/epC9pJl/
EVM/HyO5oJvfeOUdUYIYL+tYY+EnTvG7DwBSyqC8NVYZTfseAHu3+93bVWOI5aS2
E8OVRIEahOzg6tfUfIGkIgG9qSt+b/C4w3QbQOslLiGm0d0RbofO+lEeeeeLjM8X
uH9jQRUJ4RrxTy6UT7TNn27UyAyXOR31u/kjqhcwZIF0C6UG1ZsMmNYqTsFMISO0
xs1jptcd4iUu5+6NBzlkjpaIdIt4YHLHvLW3IQv39N3a5EcHEc5aO759mkDnSEKb
WQlYN4fpyKrxT8ybesraWxuFmjVSR2vdFjSanoGA57ElMtT5spi0AvqUQhgcom+4
oF7HEWhnZoV2k8l0XMcMw0DJ4vnxFoLD/hJpYV2VlhZZVwzovsn8G++YNZgx3TGa
DEEvCxW0Xz8XaWYrJdky6YWp9QUs/5wzFpT8LxoOpZ2Vd2vQzhHpWi3DwFK042hw
g81RNz5lRhGfSbKLe9TPcx8Nv6GDFR96oh+UQGztVpfrtWxo/d0M8g5i0iuBPJE1
CXyC10cAds0GF8NDqOHgOBa/aw4BOZx86UN/sOdm67+AjxlxLgep7MbpzjjHBJ2W
6sR2YaUXA80qNd8zfZeYnkACvg3E1PJSlzby6Rx9gv3ruO6iIvIOT2HBUtQf44PI
MB9XLbGFyFfS04w3NslM5NZPoeIknEFS7uHoEN7/UiXw3tJgwoTSrdil8eq84lzd
EiIO9Q1z5XMFZshNd02bIx3heF4y4c9H3ZGzy9O3BE33G1YD1SnaOacNPP/8NZzV
e1rmSMtULuPAUmsNAvyS/fJGxiTot5BH17yt2F7K2R6jVtCgT+HqcwMfGfWh54BB
AjB/jED93xaHiijkjkLNzeBQdf08N7jqJ/YfT6VJdbPR/AWUcGtTvuqdYjuO82eb
Po5sAZkgvIdRIzugJjKvnJo9svVnjd70rVpIr6Z3S76NzfR60309e5JKZxFqvMqP
+tXHiCO9ZFMxQzl3rKQ5eFCFQpU7WWWc863+PCRs8Pv1+Ynte8lCTwFwEqvsBXsg
6SmHur9Yfuj5rb+hOqV1Irzv5rTwn0ZqNnAMcHMNxtK3oit+z+6Bso5GEFY7eKCu
QAY98Pfh1KW0ZkEAa1IRHqLU/pGo2c662ojdZv73xiZ0rUWZCuL4DBaAkz4loMSu
OXJHrxtOG0RdoewQMFfb7RYlkr+T14yxpX0h2ATHYo2tOC8Fg5qcUm+d+sD752kX
eTDNrrqHOi4hzQOv5mt/49yZo7CxugxCDb7NCc+H93K9ZXF+inKFyXCrz6eQto3Z
lAchen2X07b92+Nj1dpG5/WhknF/irDJ5kqaJfyHSlwb0Nkmpo1KJl2uXJ+fdSTg
+hAP8HGZrvDpSGdNj5fCkob78sLrPpJwfm3kut11cJ8oszD4IcRGdr3+B4+8bnw6
W/EowGALGjkb+RmpfYGVJUTNjVkGDtp/pxH7qsdANlb0eLqwXPOKKw0qOT6fcT4Q
CdQL8mfwN5YnCjJjVKag/KtM7oL/sO45ihCoh4uMDu3R4RwiAoReEzZ/2oYBvChA
UkK397WH0s9DxuA1e1X/F02viU1qf4zwI6tunMMn07ppqHwYjjrxjTCAVlRMBoKl
fvwOgWQkfTcc6dNjZYC9wMk13m0GblaMBAy+NpQ8zc7XM6oTWaLwRz3LbXq8ODfK
ZMd4cL0L4hNpm6Y08urIDMS5JQbNZqd6+ziuLKfSFHBz6F7c6+W/2kCQQOtfjCJM
+8I8XBtEqhtagAvrW5E7reFz2D6wKKpTTEaPcmaCrHMqN5d5Xz2sT7NzG2y2e389
ChmLqsTSDXFxq5oy584kKN9XPfqXhKfZIRn7Weauj9prt2XoCzaWsw1eG29YHOho
OY7ioXZkQvpTH517p+SsSR9YVxZcT4DnTKpnlhGhqYcfJEGfi3diW3cQVv4XP7rY
QF1w10g2V8N0GLRdzEJMxRt4J+OtBSyXUr71/Gre506sG3HkL6EqxhOkNMHfhc0b
T+XgmoXOh+qwi2+Vr6SBjeO8Ybf+kfINAepUJr3UEoBbl8B0Ta7utLYuOI+HyJkq
AoX/un6BMXfJTlcdsGP00wv6dqXCxBn67wdDGe83mWVDVCqbMM6edyJh2AHTl077
wAMNf+1Bte/so+F9QifR1FYdfWJW5QRDvW3HtA3YGkCyu1iwCPCyKR2kDwmux/3L
hzjv4Vn4ismPY8WykSdF35R1AliSNCY7dYCDD8avkOw8G6C96HMww09kfXrDHOBB
hIFsmpD2JwymM0dQPSCxO92EdcWi654tPS/Ry+7WSsHrjLygoFODuJY+dyT99tju
vpytvmEuu8K1i27wricJ4mIegoVJoWwKILsAn1hhvUTneiqhRhWbcRlYV7LPG4PH
v393XXEn/C3i6DpkOeLQ8taEt3CBC7FuOfl+geS27lqi2DwpyA8WzO4w7i960f1d
aVNzKC+1QMaEI63GPrXJZ92r77oUrVQtIJQxEAzzDmoJUhEODUM7jNKYvUPz7NdG
bZPE0XNytKcG7IUcIfV4523PqHSYQjaUcuwYPGAy5Jnnt7heSzYzQrrfCUu0/0nK
rm0Hr7iYyApqyHGBI70HkfaTqt20GJSt6+YLzovdHPnrV/YOi212+qMsa3GFNzPS
TdqvW8ieKaFipUG5sFEVrB/Cb/NQXxPPlAV/E3NM59yXdqDVJWQ6PtgC+Yqwq9Az
dguavPRgLGh9B3ASBLjLOi73VK4Tk1jqfT9afZcGgBPfb6iUk/6U9lyvEMj66KCc
MvqGt6pxhiHEe4Cq523PArbF9fFtWqTz+P8WJU2/oPdmRClOu8NMbiRSDrtvSqgC
LEQoyXQ0aC2EiP4MYSiRL1d+C5Gy10rhDKGhBXevyLRtUkGkfZoGNjtQJfwBaE+j
qgXewem5fA4GP0eDzAGpH72XxMvjFvcVzlw4yONvI9zHyAkiKAK5ZRAqgsl9QIRn
pf7oYeaUBS+Wm5NF+w0ol7WpPxyrqlPDHFlksT+eySK6wlevmZkiadlQ2eY0ZBzx
Oh7UtPFnK8oe+kc63WZbybHaVmEaPOsZIQcvZXw17RoiILc2kcaRnzKq6nZEVWeh
NH6jgI9KcdlLG2g1LC6y2O93pKGWUSAIBBeoc2R9Gdli4WLRMl6L1EXze/7U0MvW
BuwAPnFVaD6kiGD8BsM2XCf8Gg4vBEvOcXdXf2U7mxO8PV7kVfKz0cPTxbL9ju3T
6/yA3jAhnzP37LBVpbknhiLp9tEcrycPRknocqtciGDRaJmrUSyJYcJBl6Q53xe9
mk+qDirf1Ji1nW6b2RdFGOI20OZUebvA3NWa6wcZFoNuEQJ6CgBdxqaxIZNpee9B
uimIjt5wHSPUiNI7NRi4YUvkk19TT+zatkVfcsu5cgtzx83cYFIV84BQvV2M2tl3
5xf0BQ4sfEHVY++WUHq0MgKcdieQfP1KJBi3nArHYTKiaRn5fZ1k5sLVju+5d45u
NYF9V0HqJNetkTbZ+90gJE2Tug9XJVJEZ9kd9Mx2frxod9OytIdIWnXZSJCHHxmM
4/wiEz2+6UPxhxqG8I8Vv9XKObiPzuZ0UngaL5qQGSpA8VDicy2X9+ORNc5X5iDu
+7/gSx3v5Kq7peiBaBo+Huk2cuEAUue+vwJ2+A6V433svSsp3Ig+BZxF5VmUCE0Q
gXOFq5HDzO8p+pjIgBFx1Iiike/NM+IZamar7iE7ntXkcIBmFdTtotatPKWo+cGJ
zp0uHD0CkbADm91MzRTt3TZaVE6LEi2yAF+M/15SsBsvWIMjbnfBdcRKLKxvFT3R
gBJNFJFIqhWHz4K4UQZBchNPlcrxwmg1UA14qHk9qmHo/Rh5bK/shJ3v/iDOYp82
jFe4qzSysLfJvol3A9MvGI+NRe0XmfNjbCHSm+gayHFRyKpy/RHlPzj6ilQjrfOJ
6tjhD2Bt79jPU+oR2PpfBhsnSfdIkBd/il9B09/OirqSJtGoCqP3OKihUYoQK1n+
RTQUeHCCQxqJhqqfDMcXUb5Ax9+hmic3BhCnWBIgOh9kyKT3ZYC12K70OQI18Y6j
ReTouAzgNdOzxP3ar8l6N/Z0cXmMZkmEyp7YYf+I7nIF1NBX+WU0fTjXAhQZNqN2
yLz5jzqui5+xXoa+/q/kS+goljlyJ8JVeohqjPvCClgNZC6vo9qIQx5oEGyyb3O1
HIJvA15eGBoVMAmyKGX9Y031G8PnykVzTKhYnSll8W1dURvrsbGbw0W2/IBUUUeS
1zylqKaFNc5XIiSyqhEdWwjg2PoDX7WbjPsNskEALfjIx8v/Mm22vbrZvFYpXRi7
2M9q7NBc4DMsRrZ8YGwRRsTuzKKKf40mZ17VOASU4pLc1u8ZXf1Sjn0T/Jr1lUSX
gdpIzwkCF/L2ZkcP3s2JHvd64Gr7Uwt9FYkTOrVmBuBI6z7HNP8VhZJ1NQqOgd8D
0qHFCH0IrUIgaKsYIVNbncCImBc0U9kO3qqb3edrXqtbYJWrTEFTzp9er/2mw7xu
06V6yYgSWZom+g+0JUDhikuR01hoQQtPRS3ph0jgg8zy3jbVB/e9FijY+pOuc795
WkWkmj6UmDXjw1MXrTyhg4vLsQW+ofLg424WcijjsQ74Dr2k/CuvI+2tsPfmJxk2
Fso7RZsFj6/rdEyBhMcyFFVrPEOv0p4HzBw6QgOyXMnwutjF/tCzn2LBaAXv6dkw
dr1nPiIvIk/aakvNytiidG85lFY7+x5J9B1TZExbhyXu3+J5XWkOLRODen4HRDc/
g9h9lr2hLSwOY18K1QVSbbAQMMb66jnR6jbfsHpXSJrHEwI+mvERwkbSLWlsUqO1
5Pe2iIgjl8YGEfgNhhSy9mzWxT6Jpc09XZT95+UyxslhKOsoYDG01mpgPE8PrVI7
n7s0QrOzk/TJRCT/ldfpUDv4s79RTS5941nLsjDXcJsdhFLtD+VMz67C5bYsdbXc
e+7+FTOhDjdDEmQPiBi4MH3r99qRHTyOZBz2zA0kWBUtDzMVhnyOyZR/WxJdDlDq
4Gp2cR2pBaxrTeA8lTheSphaJz6KsjqmYAh6uvezDOSgkhOIPpqQu1jB92fHEurT
NH73De2vBsgvA8eoERa2FIlIRsazRX5IN0uRgO/tZpnVKBoXH9lA9E6NYM49cXcd
sxyflML8vELXra/3wHICuFO6xlwrVaHVhsntR3BEM5zYOigxgLz3HbTE/abSYJuA
28aAQXE0sOmG/BIszeimckBy37EzB3EC4XaKBszcveeBnF0e3Awl0sqckKjG8mss
5nOiygq+CmRFzdtaN8xAeyb2vqCrvOLUsVSnuoIH+GB3BkP5QRr9fl1yO+Ukuu/o
3qh/WPaykyyTR/Nl/4Fi2qjqkb+i8Z5d997wxq9B4pMwLYNc4pUtDXUtkS9caIwl
WqAGy8lpcG6z37bIAJk8sDEzoGqYM7XlJ8BlIwfwIscavUq337ROixBSZave2w1s
tcHNQrHjIPFcpAkuOIWDUURWL1kKt5T9N8LT+nYTlN7k9jP34gizIjj3l9913WhG
vnToc7SmWj+z+a8/SLRpdnDvVxgqYlcz24Vx+ptEFBoVuZKZ+Lfo8k0rKtdjWYGe
3nzCUSKUrC8Cde7QVcrn/Xn7JPwjN3DzvcbR1ELOWNcVuk3ss6b46JO2/uij1qej
cpML5qc+xjXZZwf8SCU2RJPv1Xsw0DtKqOiOV719wHGOJ2k0Z320D79VAkGGx7u6
u2HJChTcrwBVYE1n9htlRtI6edkEMc+u0Xh8XmxTRPRCa16KY6nW+yjxm+S8F91F
onQsBZjt9DCZRoLtg1H+fakRw76L/mF/G6r00vtdLlwGaEb3RAoVMk2e7Ld2bmEx
Pdet5r1Oq44ZaT4zyZgWn9uFEFB8gbU+jQV/u+NYraWzUwmBUXCjxdGQQ9FSjb4C
YVO1fC3K5ba2HUuD+8qHIGwYJ9rTPp3fCB7+Wd7fRa64diMpfUWZoy1YCNk42co6
prFwBGCUpMWkrE75FmmcZDhOi1ENReEf4f1hKpLu6AcJwfIsV4srt7K12cxYSZnj
5MVY1EzA764fAHOWWJaPkEZ9plmo5hgULGLTEASrlR16Rj6KkEMuzvKrdILsSQ6G
r/OwceIESiBQGXk0XJCBwvhkLLjSprrHL4fte9b7CiFk60G0+XoqvPWx1owtopGv
LfDRf9kG5gUhkLda+bk8FZPMnSOAQCCy2Gn1bC6OvwJPcSfJnTN5y/9vdiwajIIR
o6PJvx/krJ+WvaKaoKitk5Rb76kFsrFvNiIzYoB5IWQbtKqnWKgJG0CaolR6dTHe
/TIVw+fJb684M8WZ/Ml/IKIJKmz9KvKfr466niDqafRONRuoElexUI6sSPG1W/Sh
2Pe8JwqrwdGmnSRrjhUz3JF5hPT3SLJ6IAcbY8hXt8QqM5ctkDUgZactuilrxny+
EePGfg370V9JZoVJHsK3H5YmVawxTgN9/Wln3YMAFw4UK0uFIzmTfr0bNP86eKhz
xzZRLSJ2RomT7h4WvvOemOV8xzO4BkyOh1V5/7IU4YWD/NjCX+Zjala2Vd7ukJz/
HYWwFX4ENX5vES/XhjLf6C9iMRh4XqudyqzlYtqUFM6SmuXni8P8pXjn9e1nUL81
rmkxH7SbF1+EX+pFI/tKU0GyCC5qQdWbR3FjIm6zJDSzPjB3p23GyBWWzqAsqg8X
+B/KJpp8dZIDDkxAw9p27qkXqvJyQYpAwF5Jjj2aSE1GuxRDNsyuO3hReTZ52k5U
SBWXCkyooQ6OmjO2oSBJAmJ4AcvOobhKip6UMgT1Yz6htLTmovZbk1v/EJfLW4G6
A7ZWgH7idpHVsjNZaTeUOwuXkNWF0A9/MO7boDPN2TzvjRYovOqwP2gdhQzEamB2
W6WsoX36eyGnx8Lg7o8baYZ9oU1pLLffd+cRoH3IpMau8yEnpk3kr4+vYWKxiUlL
MkfRaxlykE66tWacs897jv0Lhcn38T4QGV/lR13FL7dhawFVCWTdpHLnx8XTYnRK
Lzu7DtLUgS9lCUNWJMotH6/XCYUWmttSs+YKP/Y1qMMulHMHzi1cRT93rRyB6gLR
N1VmuL/6DtXxxxYIlfP3qked2f8aE3dlHNiHnew0ComJ8A4BxfoDVwl2n8l/gL2U
HGMalWgqtb+mFQeVfN/gPYAq2jCl1a/M/rqQ8CfAGb49ZsI0QpZNDw+Xi68/vOW3
Pp2d5T4hXokqgArBGdrs/COPu4GnYy9BRyi99mSGbXuXvdiltkpnL73kZwWfK52B
ahnbK6gudr1sm43ptzxO0cqru4h8zrvZHtvA9TPiXW2nyEmiqzdeqoEpnZ8JImfV
gx2J/vz3dGys1bukPe32KNbelAo0ett2kFnEt4dBd45v3rM+o/h9DpgLoUlriULK
N/HHx8GHsSrMSipq+FFKcByS8g6LygHUOBVvmX3IM2f3Vv14KzMMjZGx/F/wQvAE
A8V+jn1YRMi84HPgUozTd6Oz8kKFQVadp+vLvx6zLCvpnNgKUASbK/DmVsVaxsqR
O3oYw65GjM0ZF4ErDpIReHCSNhJmrwc6QiptxnWJfSfiQWVC3CD27aYB/NI3cpxC
wqoj3SYX9jspQV/t3aY+S7Gygv6WhG8rTD4qM9ThzlnMk+bTwMR2PjN3NsBcdFjO
A+YHyAhnVq1x4YjW6enomuba1IuJ5Yhh5ZxK2l+6qwGXUB97FRWuc27VZPgI/5yS
NhBZj+udQBPya/DxEqw4ZlfC2Jc+7/7nCTaeBj6Gk+xnvNgwLXfBeoD1x5a+djKz
ElfkLXzkTqyxt/UJQ0ciTKc0abJDjg8dhr3e6ftbOmhSoUMs4HAwP/Oq2Gkzs8Qm
VJbH7Z8FknN8INHqGHJiSwBgVJRNEYCHmV7ckIj5laWBUwNK8BisRZXk4TKWlxg5
pgUSgs/s3FiqrDor0SV03hIJEFCTX8VFU0w0uH9CpdeWBYxKqmm5CvHqDFjU2ZWQ
vNvkzHSas+YulQqYNVC6CUY55hkLXJubZEZRGpdDWFZExML9V4hu4IgryKZVRZur
bVVHJGD242taxfYB3YMmMPcmMW7ddGl6S3LDaDdXSlYUvBmEjvWIjroU3dVpCeKu
8WAnd0gJW7hce4L9RVhhye8RU/BMyhiPnlFFEqrFpNUhTn4s6d03CgH9r1HiNSdB
zGkkJsWOLlT/FFuqqhFcl1paUjWMrHLYuP2LZ4A/AXRyJj/uCyJcGBTkzoBW/N6D
HOJgS5XpugvVfPDJQHnrchsNiRFF9Uv8PBgbfBrj+jaKGhuZg+8pCoBqtl98oPeq
yAokDGqA+oChx9wKV/pH//eW9zs1CJvegdq3tEqZupJCkLVnTNdPBZ/KsZOGnCHZ
RsONrxQY+syWy92i1ouKd8IzOFUGsa47kVBXJDO87RvH73aYq9oRzbvAr9VMPZ32
iQ3s/aXJU0RQ9RHSCU+1GXUn4liexh3sIFhK1BsEg4cL8IHmSkAX1RFHZABrqldG
xC//MkxOjx0KURn9Bpa0/KuNDeBxiM5KLnWC6WdUZLeDDMPtPSWDHJe9DBv23Gpw
qvvo1XOlTJzRdD1F7lUMDW7VguuSf18KjC8VQolD2ffTLnJUT9Vej1kkGPa0qjHY
VSMQnsI6bhF7t8vHRKACXmd+1bKAv/uNO9kwcdSsAcuRlZ4y05Bryzvg/7umNdsU
BvTVc1XVHI3SjsasgGehZXFK2MrkahgXd2nBHvLNuw/yBDXBbYHpxyK/f9UBoN4Y
Pnw6fTNKOwzKyDLs1VdzMxQ/dXTmubXRYzmSZeSuaHCOuO71looWQ2zehWrcyfIg
oIg4Z6t9B8j15zPtBHkp1YVYNpO32XtlB72FPQReERSDs41mY7jZrDlhtH1tEtim
xWwBWVKcOLn+oQwrCJvT1DzV48J0Wf+6Zr4A+sq+/1sVsMXDMPXcz4XV9YIZP28r
JZt4jZMAFbIBf6NPb+wsHUdJrW77p+61BkbMblIxjf1A+tdZ+E4mKUmcRNJx4znd
/4YjVSsouYnR2ufaZrHLw/0X3dWVZ/c8AlysvHxhfUbf97++IJMmboPcxrm2WQD6
8tBCQC01WrAMmQJtABY0uDQgw3sT+I3VOajCUQoB330C6XWk2vBbfrchGqMEnPwk
y5PtSEsv0C2gILAgMWOc5EyTr7LimaSNdNoL2AsVsxtztPG5HtAU45A75ox3x6rJ
HvquAkQ3h0DzPhQnPu1T1emgaU8GH1/cBdpnOy41OPJnEYwfzKfuM5awl6Sk7UW4
T5uzcjqfiEnH3S4kJRZMNtfl/w6pLhbm5BN6SOpvWrlGBvSBeG3v8cei5kKR7Wyb
A5sMP12Tlfjqq+dL8pNzdBt6SEggHjQ+ORU7knAkVZT+Ok8XMGGIFDFQt+GJ6lPC
MAZazLAOSBL1E1p+vSFU9ye2lXaF9VXDnQjeHwufSs4Y8NPaqNv0qSbcuiG+Z+Hn
UPKrhxazby3BE1Iub125Z+SZBhHnYQ7ciwRi04//kktJ2MaUvwaQFRqN8D+DClaP
kMG8803dYyc7AoqDhGB2xfnutPzqkNQc9VDvA0GAyKH0zb04v3wRRCAqc8pttfuy
3saumqdCu64+N/ofUi+G3Cq6HkK3vG1yuE8ljqee6qjS5PjAvB+lO+c0TFkL8p+A
2Dv6I0MIVdqMWireTL41LpYrXZW+wAcMBhAT5tgyswqu2dVCMUhGzXCWxFFrtkGs
ANmbjUs/w0JDjbOc5r6wm5tMXRtcFul4VGtBPzhI505hf1Y5DLbtwHOVb8lsx9B3
8ukq5MOhKdKWW9pXKWhnSIZqrrS/6OmlqxpW+SeGeRVfw0LsTj/z6mdMGuWay8B0
+k4qdFbTi+MVVJQ+rsXBUayjoJjlWuhqIsJ1/cpFzKxOOHrzwxpEpwV1E18tVXBy
vyOnz9uobXAkDu3t7y/0bqnEyu3GS1lKtgYfHoCb8P1JCUX1whY2v0ywXxchwWhO
dqiQXz565HDQWgyUh8/2YCM6rzkMUvmPUw5QdaeJrmIItenjutpA+oH5rwzHtopK
gewtV4Bkdy/XNndl6JhbVpvQR7n41XSV0MVOCIRNXUDdAOmYyxdUPkz2ktB0T6zA
F7PJzi9tTwNPYyrQ7x6YyPVI7oypQTRWT1ais/a/gw/gP1nTL7OWF4C8G9tiw44k
ZwwAXp9Q4zJaPdX7zpqaN4qKFJvxcKZXS9Sd2SpdLKlfsovpWjdb+VDpJnnsekdd
pGuxrlzBu2JhszHb22kUDXdlvzhxjXR/G4e6gJkPwCafTmLM/KhXCfsP+UsHyClK
X+kJwV8+WMdDM1fnuEVjqSyW+izaIHVKllnTH5DzO9ru5ewtjzpnc9OW2ZYSKj5U
RI98lvXLoLpDsNj8YleLvKeWHJcnd9euYrKhhtnxjGnmiNTz8hPxGxJ6L1432kwe
lwtT7Wy+Os8wqyym1EDfjcIH8KAZIOb26j3jkNccZF5dDwCP6fIkg1BqGxzV8WDv
Lj/YFIHMGNouzMJnurCTMkN7ZszHsOj2UM/xtpaypSbWz2xN5B4brVb6fx1l4yEz
tl/+WMD245i7YXlI2UrcsNV1VoIcE4rwIlExFioRem2cO6/ZNYvsOkC39eFozoxq
U+Zhu9KskcgqyPu/b0GleU9b5L/KGNiDHfOTLQpbxXPcZASb2lBiJLQu/S4rG8Aj
nsG3IEtc11Qfe36cv4ef1ADJRw8E3HncFHEwPLeZnN3clFOYydAbtx3uoFwLRtBO
kGTf+Lzp7xjTVxs4vipHXCbxTOIpTq/h3fRuBSuYkweHIUQsjJmxhG1k27a3pNKS
W+zV7z+PI+RPrOkC/i1O3Azwp7VUvGOI7mkjn3stm+bSxgFjMXyO91Frphns8cfG
rZ7VKgnKuKRRL18dqKeqOUYhcJQb+1hWxA8NdwCQ7LGcZVXrWdby7agxMWUl7Jxk
mlkwcRr8EeEFsj1mKyt54SWVtLtGcow4dkXc6PZ8fgbovi9mfxvTPDDFndsJpeT2
PB0ypgp499IKNID6MqivFeUvIRRFpbPxRQCyEPPWjVFBNSzZbGUm57iX3apDIJ1N
2vzjnNLFFNXZT22P2pEGdzRD+UiGw9habZV4R4HV/qQZLe2Hmad4L2emscc4WXvj
LTzhXmDsn1XCTFw2HpP5GzdaErOhbLwCZx5CoBbvEMWWnnWPmnetjJzX08cKsheR
xuT+cxC0V6Onk9KG/t9p9UQcFfo/Pozxpi4USJ7+d1OO2dhgWHR3Gi5enHxtIQ23
2In1KD/rChadVQb4pQ0OtewTDJWTDX7miUveu2XRhpIjP/B9M/H54h4+iLsL5bO6
RdnrfEwHBu5w2Gp5YtGgN+1rbkCJYQwRV4IKpVNEG5nm0ks2c66MWUrKJeMCkTAU
NRApiCkZEKj8vgqz7X7H8zu4naLhIyoYWVTT4xikb5+yAWz2hZfS5r7fCOhnsNDa
GaUXArbIEyMjAVzdyuoTAj6gwF+LZojoR8T3jtJbNApjKgEvPrdWyADRqsBH10mC
snocLBjllVeHEWpdC1LQECGyMmKdqkMnmSOO7uYo4ESgy/D1+F/b61bKuZgyIe3f
njv8HBefHbE55pcV9EJVCBGKnCaH10Mas2Bvbgz+HJE2gWDHnwdVM1cfvKpswHAv
I3YtpOrV+8KihssRrhQKlRd1EWh6Cmmq9hZN4SMO/ki3TC8Y5uB0MGchmYq92Zaw
kT9VWpmsNni3/pq3mpl8CMHZ0JZQYwtbHMNIevtfEd4o/CaJuvXJlZycYec08oCX
0r8QRa/ZPsnP+5YzyCmU2cVrABGawZAHmu6i76o6B7JFsZENt+3yd93Vw1oulEC5
m5houlvKchusw0l1sOd0apy5nP59BWAA55nU7qD+d0Xd6/pZEkRPdUGQ3iKUI1MQ
bwj1ybZ6Ig5ZLhvxk/E7QV0SRCqogWwnSSkECmwwHMqdBfVGAvvXs/khxuPQIIOl
FgrLGosQ376YK43m9af97V24bQDotGvWNxT4AdVViTaouin5RlPjH/SvK5mPkQK0
xE6WjwV/GHuqCYs/8FYVlfPBbRoobI3vWWBRAykpKB0Q8/EYSlY9qu+I6xM0TXyq
CUCCIaA7w4fvFUlV6WcEEZLssCa8CJMfZ6urflv2SmjsNNLffDZi8mOhuDFK6HCd
UlvaQRuR0WPg2JBHzedaHleqQNx+z6Ic9wBv4AMgBP1eFsK0+xp5iF5iZ4DPIVnO
cdDdn0LMK0GjJ4o2Rqz59GfdrB4RmYqCJXH9OC3zZLEq3vuZfTLZmcknJ2Ff2bZ/
z8jOZfEW9UEht5pDSs0cRFvUY6IQzUq64V7vN984f+NsNrdVPsOST7wI7m+V2N2+
v3MZReUFhCc7QhJ3+gqczgPacUduVb+IkqpCwsYOP0CSBEXnD1m0KYE8OWdfjrWC
71a9b08V4x0InEsh6ggBzbkWJQ6UXeOKG/gCK1EVJt0ndgtBnapsPOYSeOyll+ZN
l4sWcOh+r00CFcJ6XNcrkZwa5wR1ypTiuWkNGXMwvEuCLqhfZM3tt3iYzjI1u5mf
I2AadoWpAQNVeszoipviyXvwf5z1u+TsTJheRdzkGioCmbktzQDztoZf0RdzqYn5
0ycMo/UzsCH5NOfAXAx0QxvHvqRkah/WFCoJ6/5fOiur7ejZI+c6AYBc9DiA67Ij
m2B7YAZib5OXvbBXP+ToLBHuuaVXpkrIgUMMlDjO39jQ9pJqqDlOq0y/wO3y9vGH
+LowSmLUqT51iFU15ezy4+nUSw1gN6fBxmQIkTbzmRDABeXOq+7DvWcXQMcNBzIH
la9ke4oPxSLqzLykFQnw61yThHkCe1TRULYyOlxijeTAJbsEIs9Q/peFmRB3/Cl3
6awmNKEWYrwKzoXwzp9OnnbI/wAaqg5dNaJ23LA5E2dpVfxvfdiUEPUl9A1HrdU4
TKTfVcA0XREbftLylYb4PA4Tj0qApMR2mx5S1RvSG/sACV23lfgLpHSOibNj0SNz
WU+FWyfuxuV86rdDqw5vjLJK3twJpWBzwGFnkeVCOPiuoz7YmDMK3sg6DypAuGQc
GGGnUqOjBRMeEceij7CKbe2p9A07p7iR3+qZa78+DRk1OVuLG84/w9qYNvn9Gfjg
i2nsKsTx0aSih4Bevw6WfO4bItW4MBeofJKv0GyNckjd6NUTj7OrufwFrCu0YTNi
3Nsi938rEVCFTB0gDLmX0g4xQf/unG6JxKw/8DOiVXPBmstSQhVXHOu7625cofzx
h4sLr8t5nByloxjhGp/N3+1V1QGOnXEaZ/avjkCf/kdKa/we9gU/E6rtW/v7oQPF
YtGayvTlINL0tt0kq5TptrbPNHaWhuq2oJJsMPCSrJqHZlq7z/JniyCYBnKzab/P
EpvflOlLaUVPBM4yXZQKlmYAOFq1hOHye7ipjDDXczClFQTlZ3KxqCgHD45lOKow
HF0puBUThn1TIb1xHTR+s/AXmTndAY6Dm1gDP4je7uMB1pLevZ3vXkqPRU/tKM5q
LPWyghsqirpFx3tAT9r4ht4vQhgN1G/JY3DqUa1vq354ro9uKJAwWCLyN4Fdeko5
qI2OfZS880k29UCvkDJFBxH05YtUowC84lylPBzz6Rd7GUlZHtEjF62kULv62+zC
pRv65WkUpHd1cg5ilOds+D+QW6fn3OglL4Sg3iAm06stmoNe/mVbcEKlO27EouZT
RETsoWnBSo3VK8XINYPuuZnZMwbn7eWuT1Aams2J+0RD3+JGi43KQLobaePEs7wa
bjWvJxt+cOSpRs3jdLq/WvWv8qRCHpXTzHaS3G/GAunCVOJ/UKZV1+prRJB+l0mT
mTUAwK3sWTYMEl3FYaxMkfDmhXYjMtXhrsGGGM7Z595JykssyT4q0Z2W4oJ44BDk
Uw6oDgiWG5MdNfFgShsmzGWX61c0xxVk0FjG2ec3DJIBaqK1Svd2ZiLYB7ZmlHSs
BpiCRqjBtylhpsV3mmei5ydKUexb/0Cr9QlRqijXc2jp+bmc14cvEpKijxJydzpr
7gZfMLaPLgqdL9qbSvqEfczkUFu4STX4bR2sStZWJdsS3LOVn/49prCzPJKrrBUL
64jvuQ7h9dI0t7JvU8P8PmtrbpAATQ4v3pP1hbxhgXfUuZqZeH7/Xvbv+CMsjlt7
VhWYj6eflFXReYolyCwbCAIzGYtFFi5WUPJAbXe9zzS5R+yGlcR9U+KCiU/CWbX9
Gfp0mjfyNiPJiI/uXHoc8L8Tjyb+EyM7CEN+KwMa8Mf2yNUgUrT/gphgHs6/uRSb
YKue7yswNCxxlyJE7yMh15jGEzRWsYzk4U8wW/uIoC3EDuaCaGiL/Oa90oUhb86z
ettB1IIVE7byHiqv+EmNMRFsBeIojXQJdVxdov5Q4m19KoLQUivk8HuUglEs2+Rr
8GUK4AerybBYmOvsb2wgA721zse/8vwonGC7QIh+UOwLgYlNSsUFICh7nZrUfCjd
BqYffS/cdNGipLkspg8HLXHUa826gxxE0vEbuibBihNLjY9C0QspCWjzRgRTpi81
krQPrhDVKsq0WvPAvVJXDbytPTDiPLWPzQDxFaXL1VamjG5kD5LD7s1/sCMC5LZO
N91x4tSo1bhPBU2te0d95Ebmu68WIab5DrycX99bYPF54XzMyC0CQ7FglihjGmcQ
aibEfZdFwdaPghhQQCXoo+yckjvopYPZD1GVTXWOteB9FjEflOreEjwP5eRFo2XI
saapqP79LwirZqP0TnI7rzI+P2uOPTf+RolnkICMG2np+LCRPOU1UeDyXXVMiDvH
Rz8shTeKL/sOnGEHUC9iNrBVJ05dw0aoR7PCcO011goMzjAi0/vgw7PKw8fLcXIT
VZd3bI0HC9Huwu25NkCxWzwWh71hc0i1gZggXuSHJOvnI0gFOznjHp/SmBOLMZoB
MGX8NSto2koGqcO+im/IbTkHWQ2c+hCuDc5uFqIdsLciy3NgeX1dXS0yzxGocNdH
w/qh5E6tmqhaVG5YIXo0TK+59lu60eEzx2WRR+GfutdK0bUu9tsNUfz0/pP7dkTc
D5OnlTslWBCc268sHcIJn3gUfUQfbbxGz+N7X8u33L5vNJMzjJ+dtkP28FrhPngW
KJf0P6QAYfAxDza0/VpZpSt5DV49gxyk4rph+LjFJi0BmMlAgPNpeF7ITbDLzqGb
HCuW4hP96AHcRVofAUY0GA==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UUuE2awigsJifBFE12jvbCmo9LkkfVduLw6cZKZDVG9cGCTicNB2V3ij0LBcpoAG
iwsmbD10n0x0Z/ASK4gJ1+6dyDI88Tq6oE4sfft1PIkoCx0d9/PPt+JHV9bWVTEH
GHgaL6FjBXx99e7SAPkpiKUZPm+MkYiE9bi3yvtrMvw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5504)
o0bwulDFSodvVr7UyC9fLpjYLxwjwMfMrg3D9q+lHyFKrYxfpgYQPJfUf2GIQhFC
wxKxRFa0mY3MY8cF6P86LI+59OXB97vU1xs7Bgw74iaRE+gTTp74B2ZTa4xEMqh4
zlg/9ZHWLO2/GMSb2C5WeiOXi7XFpx3ef5q0VKZ+TxqwE1nA4jQ4/AcSEc7jQH+Y
9sxgjRbFDLvgFp5L7u/A2kQwDn79aexCncSr3wcXIuSYUeayKBr7r3I2bomCqy2e
9JrL5BzU3gRWE/EqcRwOgGFm6b2Vjkk+gJDR+4Uu5b5cUHKPkAGx3RFLBO5z8k0h
pb/9s1pOAR5/Qw0C7j5o2InrezoZQQ7QyaZuYodzwH/P+IKMb6MPw/VYrdnHQcOI
eD7ZpqMlqdnXoNCwNrQfYJbNOw7ajqnYfyz9PcZ+iD6ltvZvtVAoIMsZfJNcFjZ9
SQgUtM7oBPCGTlV4orX1fc98ykXettQBciC3zlTToIcx0FXAypXQFkmxKuADEGrE
p/6s7Dz+i5xRGwWEYAQjcMWSA490WkmH+xe5pgu69LZ8ewKEDBIVUDUNvgjxbeoE
YufktKVjWax78CU14mBqzKlImIcuTbKDMuf3DBx0hPEdeNAW1VFdfX4rTLHIAf4q
SuM4eX/wD7kof9JZSGDFBIs2sUAeWDMi5d9z0Tt4gHCWnk62cKzTE6OTOwDZNKvk
0sYgfSUaAcAQk4G3QMWNBmKy+eSIrhE6WjuYYzF6jucsMDz8roIKB9gWlgaOc3Xn
K51UCNQH7f6pmkqKKUHQ62XEbbfzWHpYE4xBRyJsCqibHrbg1M8hFfW7+/+PeGb/
Z5PJJ1Jz2HxB+CWW7hD0rewvcWo3aY0nyFsGKO2osXBchOH9F72p3efmqXIxqEfj
qLgODjuJLZhW14C6xkgAGhURIMV1TYMw5JdD2BblXct2DcmAZ6MDoxkHfbHVEVIk
GD0ICHdFQIQAHmCYN7qTgdqF3QAPVfbo3qBDlu1P2dNHxUmlWS0U5NSEPa9yGOkj
j0ENoz1CgqNHkWqq6R4/hLBAll3K+kw63Xe2IxX8GpYK/Xqd1uZ4sZ41jLO5dh2T
7Ik5WCfhjhOjwgz/i133Y/oTnlLl4fdKEUZthX9n5YTyM17JUNeiNbQulSLXiC2y
AIYePovk6JDrNmTlmLilR86CQviPnPWwDJV5LBbJ5WwqyhheACX1HbzT3IYiT78/
1N2tcidAIGhMtJVz9IL7RsD0y7Fis0jKs/fjUAuTCgkPh8wh1PMDeNDnJZPed0sp
FZrnF9i5XaqmjdKoTWY3R9kr/T/JpghmC+ledzBZAJFPz2Y+wIZ40YRYWRWaELZG
MWz2NGe7gnyFcD6SstAxrxOAbpdBIq7w7Z7KQ15THdGsb47Ud5TOkDm6ULJdhgYx
Sbd91Qoic5+3FRY06buBezEQULcdtW5U4IWWRCJMZt+L56DLiP5n3FCvMw1zPYkX
AMvkngsfiqG/TbpnC5EJAi7z1MH8CqDBHdHUWtRFGRi5wxN/VjAAFYovqgzyebIT
VqlsjPXzBV6r/JwDNm005CVst8I5kc/R0OupQpPDhjdET+aKwvHtdEGCWzzedT31
2mpdRC5Bb6Vqqoo6qfqHmSzA936nN+UmmhkMcdmF8Zv8r0cT77jGtLvYqn+jb7g9
MFpk1dsum4mtCkw4wmwroKtqeDJPmwTWuT1Ug4U+HZ7D6LVMc26rLNZD/MrUu0DR
md8OY7NiBn1Wl7tqBwS78OaPBKhKi8tNgvmw9VW+yNDfFdBqD70rlH6o1ug485QE
P1lb3GEHth1b6DWL0yyOZRZhab1Li/TBZ2Qla2F/XNfXMJDWjiKaQ/Ej5S8zyjuE
FMLnXrkHgU91CFkIKS8MB5x7BZcMo7XD/Qj+65fm5WPc5gSpWMEBwKgaEYnEWfxl
U81/O72mBGZcDcOrddAuV/HuQzZojjQAgj6qszO2tCVQVETui1Bcw2OvdzaUfqKZ
m74WW6BYwTxZtrM9VG/68K2Ii1oyAEg3aeoZTr8r5FlFRZwU7iK5oOYHROGSeS+P
7HfDZ+q0MJe/HTQ69JbBquxrdAyiAk2DILO1/5b83zgPYZGeY/+1tmKr1d75wRMd
KVPvG10GhOU/kWi2epQG+d0wYnKZkXJQI9Nd9CLZadUYMv7MMolyKP7QYUW2e8sf
IjFMrPAX68gtPZMlwPn+3aH+E4Av7q3R/0G3ajcU1BEu7wR4zbvWpXJQfQiyxPj8
pclmLQelY67UXndepeA2O/hzGkKGKTfZGh3+5iB1vHGF1vN2eTmDtBdQs+Tdkd9F
t16SNc+bjyynqCPnUKxA9JJ+xZ2R/56g9zqgJXdvNz/Dw00ytRpX6YgVYtOfMnAI
1lnDrcmyG4kubujQQhOw5Brw6EYpTpidmJqPdCSI5MXYaP5uGFlgznXfv4970SMG
74oeIQPZkjUyj3XoEijGBgJSBXXFdyGcGo+WGmvrmMn3w8mkZd9BVRIx77EWtaok
3CvB2yz+SNDPELsvKOBBqCG+7HCmB2V7Bt3WB0VZLHNwgTcWcjeDGQcN52dQJkjC
XXOiXFSAKuUWoPjjOeKzmzeqtvf83u/6ROizpOKmNkVoGzRpiWWI+oA1LKOirFit
RUQZTPFIRndt8pkTFS9Klo52ROmYztLuN7g1waCAquUpTfq5s/ePO9mx4Wk8WLVo
qBnj1wYO4SJtxvjnSwiilKuTdikD41G4gHs84uAnkybsJna4a/HaYCMvqhkgK7+b
B+h/q5TaxLF/0OnGIYfQe86ToKCXycuIaXY2rn7JPHTiiY11deV1+3SS3nCFglzq
/guK4uddg/GsIGy/61XGq1iokO3jfQIs63Ox1W1hbQTkxeE29yXu6+gnRdJBLLE6
/Q849QzBSm0p/rOtyD4f4sSQAHXUVMcbEntYP9UDy5vfLwXNltP0LV19pnBi23qi
OEh1Dv7euqUuWb9+wWo4TPT5YTv7eHH57LLYqhJ8aeB5WfgZtFiJ/dYW360epXOs
/D0PFZVvDEMK3z+tDw8V/pwMxRsosYmz+yaTyomm3PViAfKHqAlAgQZ8ZtS445nF
uJCIx80JLVwV+glHNJpvEJwZMhhngW5fbHiz9MldzHxQlmFMN6ntk/ZPlEYfT8Yr
i6gGsjD2AVKKOLhs+Z6+fqGp2S/fPzW42b1E8nd02GdopM+QfMJev/0mSKB3h/wc
lcYNGF530TDs4/QY4Ql8BF51rhqupwCwzO82+j+Sbort8Svo2eJWk8VYSMSve07y
mXlAZrY6iAAROuHSV1YC3Opg+6TmXvqjyAw9eC5/rluObRdL0SbLfjg554xJIPKg
tSz2OEJgjYJCUxJBrG+xI+ibpN2SKNASVB/JRWsTf6n3ZzQ97PvyxPW3xrUI27WC
Jq8N8n6J1AWbAxWrm+iPaw2Xm/AkoS8bpID9dqSaZzuQmOPimpws4VB84xemIaOJ
xms0e7wUpdn1BphPEd8YzjSWnbIuiqO9zm1SjF7j6UnYiV6btdwdNHyxslDDdLts
II1/RVZnKslDknWPLkw03x7kNj9L2Wfg+W2v1ujlYdVAWHkD2Q0iUAEVzYb+dgGa
eCu7BQOr91vAKnpafNmnQKyh+ne/w1Ymw8HGdNHoaEo8Em9xRnbhWjRNDQdW8e5D
JDxoj3qL6OlMXD8C0kOjkxmHHeVWUFs7JwQKks6fezBTlXi4rK7lkGCJ7nTRMnKv
S//AxU4YCuWavMA2y3fftXMGI9dZ39PoHQfDogKcqsoPnQTkDjg3OBOAleNyj9gP
2e/bc/X24a4SFOo2x2m+ZPE7OOxNoV9ExZ+wcNXVFBnDa5A6jXsbq0m5Ln5h4gbv
GJd1YPgaJN8GET/f5ge96YPvdJBlaaehBGFYd5kMpluHcCQ8tBMbmjgf6qWJCxui
riYc8hhj9tijf4Q+2xDNtwm2ysb4iClgv9nA/2GxYIwluLedMYRTUgX5glYKrhZ4
AX42Z672q67qmHA2lRkAk8IXuhzrKNGYpncCZ9OotLaikRSceQSRmP/cqcIgKp3g
nLxVwRoK8Y0zof+LJWVA/TH6LuFD2o6Bq8x9vv+DhFOc9qrX2KUPTy3r6cZIWz78
hOYkDhGCVY0R2bDerM8roUdj/SzlZyj/P1szKKbszT7iYhxhrBWMAwuhWSytzmov
Hd0jpFji5tWEipPbyywNdPYoQBL17vgJAAUxL8h2gXbReO6jFGW6jJQ8gbvYFuIs
b8e+ow2dOaku48mnXkjButC88mJ8JWvwzWjp9D/e4z34/hKc2VwtbhjV7hNMhCiW
T1Ab6YZlkTgf9eiTzXRW8PN3otYHSgudl5RIbgL5fGh0DbprVeioFlOwlXDmn04n
ohV9uSoRqW49Ruq+dOsRbdOgPZMZjadYXRtTJ2S+07tnGOoUo1HAtwfssB6C4N2f
zN+eFKmbiZqmp/aZBftglYrflraQLE8BRQW+Gggrlojq7p169Z97RVlao4WW29K+
86IuvPsh8YWaOaRCES7CNwkI6FENDkiO875w8juDy+AEvCyX91HeT+0wGiFzSppH
x7CceOKkN8csQ1s1eqU1SZW1oa+TizFJ4NXXNNNgC74GbM98fwtsVURTO1Z7qGNS
Fp97vJhQ1LaNIGMoMNXp+XXe59kExYoNIZNfTXhyEIij8V7Hdjr2kfElr8LO0f6F
omHzfW7vAoVKU3UIHRy11jhmrDkhA2wCGlRV0bFx5tijOec2lpT9I0O46G6JbLHw
NsDT5wlVZJ1JnRgqlVnzv8Ixod+H/U763xvndQLcsuc8SSipsM+PZQpDNdsu/8MQ
iDm56L1Y2vtmLQXtmqGGsevajxS4o2vUdoGUboGc4rHBrqYI6OLsYXchSiod05PW
SAigfFn7g6yk1gV2aq2mi4wDX5Mpf8G1izK9HKsvuovgwPVW0+/kLn+px6oFnk2f
MhIyka+HZYO7xxSq+zMmyo1hhuzY5ZOnnQhhROYEJ6n4covwCMcTH4PUkwYeSwpt
hFzEK6s7Nzrc/N3gEj8ezF9nRLq8GntClamHKofhU2YVqRaG44aa+Fwf057boFUz
10aiIFUOx9LMCJWgizr/Pa6a2NoPUAYumK8sN4odYBoNxUGzR+dQwhulafUNsCrX
Abzt2rZaNp/u8D0h6HKpyAAE7iIKZD8hfi/tNaTJFEk7PzRQUC62gzAeAOEgTPm1
M3PkTeZo/e1Mjv1hD/iSydCyXqugy26yftGOekMSOr+ntIFz4sbLM0IgOP+Ld9JL
mM/GcZjXLtW785u+gGrF792BqgiE+WtvbU/4uAfZjIBwVHzllimp2YQ6x+OmfF51
rKnJbv/epJsBgIIJhkk0gIE+2rYmr2IraFci6xr7RB+8763FtXtQqJZMdKocDerk
0WD8r5uW613jf7gZw+5nR4nqi7irXxcmjVQp772mWqxquItlMJ9dWA2bjJm7+GpG
RCY04uytPZwC4LWVw6txm4zvEEDCVZ72dXl90xnIqyudE2580oX51j5yEtSdY2fH
6XlSYnCqibik171YNe1XuHVpNfatCnz0uXWVzL+V0Tz4v6l3bHyFqJ5mq/sGL4ey
nXFwKcFZgJwWNfSBOX2+PXMn6l4/ToIqsP4ovaX4qnoFgbaOlQQPsVxkACO8qmP+
EZfhFDBOfTb6a+ku0+6gyHAKe8VYHepVOaf5kIvnW/Kpkm7o8sGlTggLrb5n2WOC
0oqOniYpyuuVeIcsZr1Mtk62yQ6fKTVjO74tVJ+SkWLMbG+6mLhIjydzGmbqayhL
iKcW1MhY8H4+qzYiulQMjFpNRqBa79upLxmNGG5X3cjiRHU6ZD6I4/BX7IEbgMrQ
MFg8cLAXcrWiUMOneEyCRdpUDXrJWfAAUMPgzH/8Yk57esZ5T9ZpCdtzAGc+F6S5
p2VV7AhFa0iazKZGiQhmbSVMraDGZM7DYOxgMeXoxmNM8oXi5VDT1tgQEsmKUpwg
2X+05WX+KJ7xxnX+Sbs9mbPad3baby25rGg5ImAhTflMyLrOKisBDy0TkGUlBx4q
/OKqIIBUo7fiys3S/WJZeXKQQ1kmWB63/gQfL8wnZxLfL/acUimO9daVWyxv3vMm
0QoS8/qyxnxrzSlbEqENdlPzhLRfDBmzAvOixQJAShebQhIO3Izc/fE0cEtembW7
AgN9uBpUqmbPZC4VpiLzltRQN/gHgJ1P1Mh6wYp/T7GnSWr0PSnFyJ8wy8A9z8zD
xN3HQktzI1z725Oasq8UWSXKh846tVFIOzfjkMI2viHjQHS+2yxpQD/RB4px7H69
V8bWmSatqSy9A56Bi1RR0QOWpVkOq4Ya8sCcs4ulCFxAJiCIQb0hUV290fmyZlBR
JaMF16Ao5WKExXQjlXXrmB44jzIziv8y+OxQoh9lhA8vTdXC9T89cjx+UdWPkQpI
VV4KjwnN5B1GqmVM8TmGHIbUXV+kLwn8km++ScNDVozDcuLupCz+TEG+8ndwfOmz
VpukK81wX0IrJ9WweQ8KrWEZitGjo1QMWa8bNhA3zcM9/IXu/ZM13j/ge9u5BuwF
rRsfOdeb76HRbBbzOOfwGoFg/sPtXKQl7UsXcEJaXReljDIVOhxfq178TxveJpOf
jut/D91gcSWkZmEx6mDMNqhvrU5YXl2B+EFX1t2ahgZnMYrLO9NQ8lMQXBUH1wM7
ENHLts4qSq4HtyBwCG0Xlo+6JdK/DnuyFkuf3FvXuAMMTNVhA2FMgiY4o7risJ24
9RewspTA12aOaAYZWVxUu5HRjIRZOaC4EynyBw2e+EbcMIm/ezRk7iyReKQXn/Uv
4hQIiAX4SxLezJ3hgB1oMLTZjes/YTV38SJEZ0ugWqzYu6qxzwcgqDU1WWONGwOs
CBGtJSd1FIiJAXCqT/YPwA2QANljznBwM05dJEV/TSIqmJr6/tJEKl5rtsS6JOp9
VQykjt61ZM2TiYqy0q6oD+9cSBkEi6FSmcQoDn6HiDylqPPpYyW9y0lnYZi8s03R
rYzohvN26h4TxCXqqR7JcRYDOL0ddA4eeWlYXZidjp7B4Y0F2xY0ujZLa5Nrp1W4
J7K8QO7OOCo7xPnRtPfhPPqy/mkxsbOdRucqmo3YurqwDS4K2A1bFWo8pu8F27Bf
3AfXC1B4itiS+ZDBON7iBEtcuudmHR56MZDeCT2TCI/5haMmK+Z/0GYHM9ott/z2
R4RElUt+NLUcCkMippq5nnroHe4H2WDVtLGWEDK7FzYraAe2o9V6qDukl77vS9cr
leDwaKGTvtu2yPXOdIB7iWQ8PPGUDUEbGDc/luM3Z70EAi3ZUYhFoJDQPcd1qKtp
Lhn+9FfSZ4b2nYGgoDSG0SOcTT7JPKajTiC9yxgENbQ=
`pragma protect end_protected

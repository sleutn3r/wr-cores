// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FOZzaoxBwD+iPSEDPftSarmmF2zw9/xU6K5Z2p35WjR9o85mCen09/c32hq0OgIM
HnbN2jfhgwQ/epZEgVNvd16pnrWhJEI3QykuHqz29bcBytXaTNzqmHxkxolp/BPI
zV+Po2ektQPbrqkbitSHMWdZRK51HmpcYwVU4qtqNEw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8144)
pzjOYFydJvbrS3AG7sOOPKmdSixDMXTEvIF+9AlHjlUEI6uoJitqMG478CVTXsUH
XDrQEPxkurSnZRAoxJplcFipKKcWznJvNAfc9fWskYnuwObMuCeVJtsiSItj6nYK
Rugk3afCtIKK821RvL3bbZj+vPcxRPG1R6EkgUoUfYwUyyuSShmPyZuOAyGj59Kb
w0YZtAgExfBYLquOvHuSz6MTz4+psHDEjvnqqwID7Hrj7fRZOJVwDvbF0pRmCsv2
xDUbam1YGcCvhdH++XhfDWePWGVPQ3V1TNMLxPtfLfcaT1NoTGmfNbmDFRezQ1xH
ALq7Y9yWnY4zgJWvHyXOk6F2dZF5tHn/5OCX8ukD0uy7K0eGpvNneqgrCYlAKVm1
HcxVFG+STCLfoqK8PZxA6WDvo25iNdSc8ELYYP5s7l1LQzbmW23UfffhaUlzjwpZ
WwQiKer5YVwV28fk76rp6K0FlWXnzPDYQDv/1y6hKRZbf+s/W3WNKlC/U9AJj7N4
qhpsShPqjsw7JIb+ewEMl0td6lBpfl9crapptsr4+XqoQptQzuce4+3LaxHZd3IL
z1sj6mt/6Qr+S9nr3oGWT5Ax7qvF7Hk4I3kWOwxB9e92Syi51c4Y7TgPrQ0eH8af
pyogYY6CKnOVxejOQnVC9nZY4Xa+v1+8O6XoSViY+1ayUlriL2mUXTQC0xA2AI4U
OLn46ceVCamYbiZ+k5dlktBar7Ny/XPrW5t+cd3uY5U6XCnlKnMWtYMjOThSRFai
YgzKekVPCcUnDimdvJioeSZ0Esk1autDClRwcyKlKnvxbT+wn6WeJtM846lHst4x
AL2wSS9Zh36iGp9skpBZgi3K3nxymUNI0fTGAdtLXM9rLlrIwm3l9E6hE3QgbF8R
0GUKW+bucKDkyXbiZ/jv7DDRBm1cBanp/2pS8ftcEkfYKxIfuws0F8CW1N5zqFu3
RBaFjpKPeOeLbpUl0qFc5fmMwS8OzRlMiSkvQGaDh/5H6NEtp8XrAuUvz2uWLgCQ
+CkduhmvfrHqFRlRNvTyyK9X55kGlfILHYQd64RTgqk5plCXzgtcs2H44o/QJOog
iYdxYXTG+HCWSrDvsadT6Uw5SO0YGwjFubJbj2pRtjss8/pxt/flloKcG1OWnAyc
NU6sm4KpxpTNesU76U6vPAD5VDlT5zTZEUEdecXXD0281xz+tTiZsTNEwsA5yRP7
fc5ia/w9mQYAGLmPUA/NmqRWIv7WT5iiuFYnkOCVo9R1ymKXIYPy++IqTh4I+4tO
FlHx5sBums6uGGYd58WVPRaoasZ5XVhwJrInWyamDewFrYfiakyzflofHxxTGYCv
k268GWxHjsZ7VzmL5QZs1IN8H9LnrwGkmWNMPCZs497DNL0mnDQrf5Wi0cUuSprj
P0b0EnWkTpV9Z3DzqgLG0qIE518U1+82Gcr6oxi8T6T1nnV45I5kcZZlqYHsOvrE
bQ33g5f2V3/BMvYKfRwd56d+jvR89kzQ2s94TS21tShu32jOAKYLi2oiLX8ThL6b
bF5C7P5gbWG2ea6xSzXze1uG4rRmO23hWRlWbbECQ1s7lwJInbcyFSnIkemu1226
q3qXam6VP/AV1ojwFYMMMhjZHKptPmL2YRlSWKgTeaU2jYtssY4y95uyx3tOXJxb
2NUAofKDB6a3o3Tzum+UAdJA1JFjmKWUqGjvYPOHoR7YkbTMeJenI38hZr3noxAR
GAeJ34ZhkYlwZ0+pCNDtTPWLUuOiz5ufhOM2k0tauzkJ2goYt9z3ioon7OXuTbF1
Hi9+q1Y7lzDcTuzagySRSUuMorsgwyJVZ45TC5GV+Pek35s3RxzSFDLXE3g73lY4
fbIYYg1wiV1Q/XxgACbEquwGh2vtdCPVLIgwm1lDBeH7FbXrE75kgUQfig3u8G8p
oX+lTFtyD+qdcdEKltH8VZMdY6HKH3VR+/vaan8TO3TP4yn8VHeMH+DjDwpY/grH
WLGlaUGihELqD9XAFq6I0jW6t71vbfqFN64jzeqHMT6mFKEc2T8Qrko2sewO+xiY
OAsHSG/qzpDbIVSJNvPYX0Nq723fgLi7z3wIcItBy/Zlm4xrf2kKSO7TOAb2RLv5
b1ZBEMqRatsDhq/e3xQCbvPWwXUl25vpeMe1Y7a+XYXigizVNH/40y2Rbd4EIUw6
/XMDGXDmhukaag1Dqya3IdMUOJuDtDOsSvvSy6Mggl++ZLJTd3HoSABJxgjfCgY6
z+xzw+5C0YWqzkERlgMKx5UXQEeJ2S0NdRu+ZqKcj2cf/PEdMqiqJ/Q5p3XJFafC
G+wqPTxH/GWJsadHHdANgHSKrG13d9d2Jm+CLIAgAuKIMAbJKaW3EMdVAEysVV0d
/mzIqyEP0TLwQGXMM1wf8SP3cd1aG2ZieYJp+3MronTU6Dv1ZmuAXgknokDzIG/H
b09XqysAfHhbRIkh6LZj2nDXkxp5/yIowlvI968R3GxaHw6iiDiki0tGRVAYypJk
j1GmTLySyfy/JzLfRZ/IjRpAU82XR2wgsMrKmG6A15E9idxdvghgB6By3TMSnexa
TnaI0j2A59PMZDXoDjA6TrIV20Ce8JuSjPKOhzo8jWVYV69b+f3EpDPR3DojrnfO
yhY3Zrdg4hQAyawKhv6+2GIhkFP2q+ItxVIWrjEhz/UV6C6X0RDbyHufTJ1+vRUB
Pj5GGcRwsEsaDr1snxHQuyImTfI20uiqO2Plh3kfYWcsFOtUzNG9uvp3vU/eJBqR
9xFpx6cbjT4EUfvxDM3pUQo1YHuYkOlrNS9ns8Bk68Kro9uGStuHOIp2CADpcjKv
Vh0dyGApatKS/8wlA+sLgywMMT5L55yOgrN9+juHHdadG7a94Y9WvNV8ccMFCQbu
ErARHnZ6L5Nwfv+HEsRrK/3oLoDQWXB3h/Ywl7jTvks02zSDNmpRoqdCjZWxxCHL
TQsvsA8mMi/SLazxyXATfueM8V5sUs9TNpUfmGq4QplpNqgRyxlrMVjzLj8VZDhA
5AzRZGjMGD8jxCQLTuaVFKw1XJgIEmgg7pkrZK2fj8xxkpuKNExfw8U/DMiQPLxm
UZX6EmlC7xP+0daGtksGshp+OTc3cYGi3ufmB4eADBBuk60jzfMqA8Gl8WNiQlXd
rdKxG2r8iN1s+BLT2WaC+uSrzqWFXY5+S/E3hOkLXmccYAqD9B+Bx8xmgWwbKcgN
rQDxMV+Yn3ndlOwNT3cBM7H2Mfez3B8ZOFTnFMm4eO03/usksKMWHZrh54Ck/b2l
bJwYOhF85Jqna0hdt9TahktzU8vjA8diFfXCgINcXOpAEJg/BqUemqnx0nWXUuWi
8ExzqUEd+ysiqBQbZzkJsIkMZ07hxMDOsBkY3NvTHqCf6ed+059WqcyXqJy8DS/3
SPwkNU0d0wOsv4wSXb9wS/aiNAlyJQCAJ0pnpxHrgLRlYdivc0+pASDLKo91PGmt
Mr2Mw3u9CElGZCAcglQ4PxKwFSWIGRmQIh3PVP3c3L2vgQP9kVOWPwetmqySkCfc
5cUU+o1lDQHrio/VdfVV4uA6J/LFqWfqaou84uyUI1MjLhZGUOFuky9SyWFOhHYR
hLu6X6Hnbed+nH6Fpj/SKIO+daTks9I+U2PWKcmw1bPiE88TUyI1x+aREC1NLw/c
NtoB30FlLyKPLQslYgTDiOKectXtuPUryYBQeYH6lf/aeF6B0q4PQr/R+SSYccOl
J36OoJogzEtAmXA6PjR7CzQ07ejZ5oT79OKdp23XmJafzJ3Dj9sy1HlS2VFvTtYS
dAzAM54UGUq1YMVwdHJ1XePjqTbrSe5bmMh/cJowLgj/R+Pw78aN2tZILwd/tkD+
2NSdoybTxNB0j5eYd6o0lsH05a+zLy1h0PWUHwAlkbdVqdxgAEUap89SHOLxHbgd
83l3f2P58A264jwOVw12mX8UiTzmMHKzTGOaDTiWSKz7WNFkjmS6Q98rHCp33zzE
I5aN0F58urlzQ+rkdckh7yKC4ujF0VP7rW8JF7IfnsSmEA3Dwz1zYoNHpTDKauXQ
+Z9zmlbu8xH4nurZjcWYTiJtwBxI73hOTDxPKLEiHfEb1RUtY+Ux+Ge0SSlHl6yw
OZxWvYBYcFL734EAibzGHhDYtVx+Sl6BtWki+uYwMfrdmtK0Iae1O6tFdbwuPMPX
KZHqL5sFsYaE7x9FCRGKF7LS4O+JcUQ975pEQq6GE+34P7agy6O6QUFGLE6fNjtL
oKML8LAwqN66EPYTI8nEn0/FAIeJCN9f7LDrJlKvGpCf3Hgu610Sey7yoJOJ2Om6
DC33R/pyjp/9bEBIZvj6L0Sh8MPLcfLF2I9RiqA+P/dbUlvpd2FhFqRagCRbxofR
ItQbK5D8qN/S7s59CEziG4cIyT+8Jm2sOpcF4BiFMM0H0pbwGEQm5j1BJaR01b28
pwA7sO/FHnuIlP+v+aW+ITvUB0MN15tlQSOsjbhLZoUuGbDffFf1RJ+aRJ3m73yG
qTaCC/gv3Ct+xXBzKIPzjgpJLV9jdybooYFCTAnvz2xCAy7dnfhON6abOQ20BgDL
ClWKdNpjWAaqXcHoE6neRak+ftMfYRuod4L0JGssu1V3l/orFPSrYGhRyMTN0gcY
WDfBOyxZ9XsN7roYYrUHmHZwvH+jQi7U9u3yhkFhlbWqs7UD1h8gGaJR8xtasZnK
J0ZLshmFManmOK9O0AKZBSN4IRH0C0eo2GsCetPHirMJd3QwXVVZ5mYp7/9BmvsA
Mh0Pvsfssp/BOv3PI1xTRRvjDXROqcrfZP8VzIO0CJY3O9FH3zpDzjhdtLbFFG0f
XmWchz5EMuMU3iMErBPnxiImScQoArxiUugutcFtXQz460+AJsNn8vKKcqtpkovQ
i83Ewc3tM/TKs5KT/XlJPktKH2UY2CL3Jw4vDkBpotnPfnx5cqb+Xg6XDRF51IZW
a/VY45rsxa34AVy73ip7DVxjUCr5M345TA0x/NP54S0Xt5uNvN8JofPK2tcpHubK
tSOHuFfazjoZEDg8/kkzywibgdeH2ZOJHkppdWl+kANWK/F7GXFpj6Zca+APuHfN
KCrCqHd0eojWa0P+4pB8BmtsXbWq1oLWXjDJGP4dyL+MXoshwIUmXkY8pEPaJpb/
ecYUp/+OeoKqNH5B1iltsNmcMzsVz5SqsxRozCWggvVRyKTZI33+nJdJnxDfPGJ6
irWk2fz2ySHG1/dnXVHHT2zPT6Es9Slwa8HoQYp7wtCyh0iDGBTYlpxEXOH9PtKB
frfHcuabenoZdGILtqp3CFyFXhdSfU3VedWmOCkkb5EjAGw6Yhr9QQatIhP4imTM
idpjtqIDrbu9cEpu7HNwnQR92O+ivnKqzPVAAB+Bf6+vlBE9tyU+R+TWBTw7oMno
uB2Bf+u7SjfASE2A1tr7K7wAM2ZSJXKWhu3ctrcQfUv1TdVt1ESRUvqXtiMUPtac
dl9N6jfmayiGPs8Jv2NyM2L+CcpgjsnF0qEF2mUqpzVtEe3aYDhZKA7RVXhbYizl
VeocUYJV+NeYJJTkHg+AsQ9wZHBc+LH2f6HFtdQ6xcmVM5UB5217U7RpPkd2W3uQ
Uo2/gAd3KdrpO7OBPFPxX6CtkIsqsTb6w8tvrTNc35aq6vjvZJjqtPrQKxdRPzEA
9rMOgK6nDy/g8zV50TlDENwAzdHqLEV0lyJJyEEPQfBvfZi/lef0z+lSAnFjohNe
quZnkyNU+6VJZ7hDxG1hmQn5IVcE0EOgxe8lNXkco3Os/4A8v1nyI8NM2JNu/FVV
Rxw+skXU78SpBmz8CHKbgItG1XmaNxG2Mvs3lmCVUqLrG2TBfdKZFyIfz0AFRP+T
AaZ4Z+rdr54+M/odDxD9TFUhKZx8Yvla7YrQ+2NPoWE5lWzdDpUdyqriNVNg3p4Y
9kM/3WC/p2FpzjyPTTO4P+nxm+Dj29/oxpQGpKLkyMaJMGXMuZf8b9qgogSqVpLd
La4Ke+5pHcfUkinW6yTwrEuNRrh7z02D24WqtNOwaFBDJN7knVOZ2A7oV4TWOurB
xtYmcbirXNYM9iZIP62U7EAFzOEa1DWkjKJauqbbLMDA7na9cOdwzUOqzG6DmIpC
2b85gQbpHeN8vQtCgwbhX7qCz7YsY1w54l3aawlg3492zeI/bXYv4siyVKg/oZW5
6qaygI38XXpaAgRA83fv+7URcWTS18ngweijz2Oqftu+yVh2GdOxkhGgpBASTVqd
h6v5GTB/RakuLRWcS53a5VxlvtVw2OkUUADa0579ZWsuF9CoEMNQobfrdErLzh5/
bxGat7B+67QmYB/67M/VCtHvQLTqrf4wzwX/+Zjet+MeHImEsweyr36L7m977klS
GUmfTnPfQFSUGI4LARcer8CAsOLCf9+OHNkGeoLeHhW3xajzt6Dzy7fbdCEPS0tz
pceJ8+JxFqTXLPIxa2wRiCXHmUG7iVDqQrEVSVEcP941tgszwkfg/WIJRAtRZb2N
k1/tUHG5Cibotro/iBzxguwL0UWm5cbA8c2352Ji5sPy1l4bSl71qQM8PQhbF71Q
apYXOsLY/N2/PYqnkPqY6N8Q0pU15kTo/Sci5LISZ223obv5m+xpKi39//aSV7JB
pSiWP0f25FdWujrJMysu2AtaC9YX0mINf5y22cVN5OjDtekDzN0DS62/1EfYmbb0
e2tdJGzin45Z9YPlBHgvHa1cF/pMdh6Ut8dVrXt2TWfqVYgv+gURQ2EJlk+OZ1cC
OQzW1bY7MjVUufkiPFEcAA2Qa6ZH3GmDaXoOLCkrl1cDKFiNb9YJGhf2tIj3mAgv
zCUyhIl2ulX9X6pzPxj7peumxhjK2FelqBTMVfp6agm6Tj4emriUKIpmQi57epb0
BezAuIbaWi01wXzlA1HQ8WUTvTy+SrpmZGQCh+ls/tLDjJ4PNCz0ecE8EgFBUtcp
K9o4eAaDvTcuvGZYjFJAvkD9IAmG3s+qldIo/lcP/lMeQCRpaD+8zKl57SKbrSlj
VnCUKnt7679mA+Gff6LCV2ZOc5T9u2KCQ65lYuDZUtkh8P3TX94tz0lO2OdOXFzy
SOsDngRjvU/7GwhPT9THEubbzWzTQf8udAEhpNEa9tTWQk4DCQVtSSFvgzmoy/Xi
6Zrosdj5k8zjmIU4J9SEQAA4AQXogxAqayVUsb7aslbTLQjAtWe2c9BH136YUl39
MjSfK/SI58AfDI273sd/xvVAhhz9CEOZkFR5m6iLEE/ivKxfCuzFPnxSoFVzltUk
mpOXUixLm7Ooi+EMIc0+5ah2IzbF80SlxyjSXRHYJoxiXbhSEcaJUdtKTJQU7hAy
sTo/Pk/t9pkw4oAMD+PU07uj6J4c512adkRDLPEfpe98t0Ekxbnfuhg6vPUY4HPo
MhuZPbG3Oh9/hBRS4CzEbnrkKPr0sGKdd2n22+dVe97pKm77mWrHBCfvCn2DfMTT
Z7KFUO3n5eimr/mKkfS2Mco6Pxj79zuXZiLYcJX4hG41irk3wm6lryAxBnDibhbW
gtW8XLTg9kW8rXGkG9hsC25rYvqoy/iZbJdW/a7G74LQNsCOpCLMJ6wIyjeM57Q4
6uEwUG1XRT55gSByN6Vj8jguRj0FoFcCaZDK5qjnmNkdxya/Cpm28UorZ6K1ufO/
eSDTZKO/GRvXbHnmoQIDongxWXHbRyxLBdPQun2vxwbcmakep7Z/boWuSx28OK6b
D2getzBqFHjcJaNGJnCAGNN/u6WXb09Pkm8/hvuZ/J2SRkkkHkkX7V7yKRxEnyWv
nO5jcJNvx0tRw1BNwV87sgP/V1NJDlwZ0XKkx3l0CNhwqPkZD1EpqpG8XqK62Svj
1Dxp4FRD+oJ8qXggZStLENFErxFayMsblKDD0PR1wFfjefziYsMdyulHug+d0qTd
FpCCJ/njyvvV7zbu7E4sK4aOIWw10PppOdp50LsAn6QEKHdE0D37WflvX9dhIqxl
SDw5aTMLB9jyYH4BdpMguyzHjm0sWZy4rdHApJN0TyCyfcymU7R/4IDEY7jUiB74
KXOlasrZlKxoULrSZpMzN4xz2lcjUdziKdNnn+ze9Pef+0HKhblRbf24cxUh6J41
/8BOA0ZNG7W+Bs4MsD0WjSRDiUd814Y+QMnx5Mf7kfLbI+tvPKeu8Q8GqFQaPH9e
PnEQjqbLYQ8uFGTGAB6Yc58WTm8roqCYjAfm4cj1NAGZRxPX5vpeHEWVpVmOBmb+
kupd+8+u4Y7Te8oLLPcxntB7dgurq+wO3DxlgSERZ9mi3lqwPqc6lNeQXY3XKwPS
41uzgzJMjjzCN60+hudN4FddqSATmcj7uOp/4NOFzLwzRk2FiQN34aakDWJTpPHM
ubdvRyVB98ilA1jumqpLaM/Nz7If8WBpTKwAa7Ziz/tvXvVDvWr19IXn5h+WFCko
Q9ZsS25z36CsPyyYiCdayh2Y4OT0IbpRV6fPQfKz4jZKBJv7Kb10VWUZISPyvn1y
P14NRyWXXHC6jMvAocWshEaIaIUrlLZ6X8JxoStSUfoignMyikY0AipGup+Ln1lw
iHKlvBBi7D3plTo+u6ux7FrGZF778hEfgAJu4W/zUDRjiK2WyYtSjZVeNMt5a4vU
O4irmY8KzoQVwRBnMcaUCLJK9VSp2MEFvBab56ltaU//2ULKEru8iDUUIX9LwdU4
Kd7pD1Po4MB6IRv6sFDlqTstcTZCkaYOPqWjLmuUo/6BsH7XPuIJDjExnNq4cYY9
Xy7ItAB0hwSF5f9hyWwO8ThdeIrd9bPxkUfJtlNpYFdIFDhj3rEjjpK5nhnSt+eX
2O2VYCXr38Sa1BKU6Udsf0XxCGVkQkgJoWDFoVqg+Fn5fZUW9ENB0rBr/uMDez2c
LJt8DzcT4VVcFy/7cx4pszkSu43yPao8gNkjEZwCEPSEMLuFEhBR/x2uj4S+hx1x
Amx9t4T37di82QeS8VwJihB0bE6LuZCngmdzq5VsrVmLp1X/kms/lLFOREwJ/nJX
I3URnfjKRU2NXp8jC+XwDtxAQB9ohKCbcgNuXPrGoq9UakVPpUdQ0nbP+U5VnHvP
bxbg9HyqNKx/ZXax2Djkx9q1jYvlLU7GCWNOL6ZasMH8f0pF4dDL4eyc4fPlcEks
SQDlKeEb4Fz9nSwKQfUaHFWIP0p0Y0+BYu4vmHYDaMvJCORcuj0PH4o7jyiOGrY6
oboho15jzNupy4Ep/6NT3r2RIFc9g0OwVdYVNqe8AF6FRfOieWOS+zguXRBGBXUG
qr6jDhcYVgCCyFjiCWy8KlVHDu1o4OgQf3bospwUSQMuJVzKY/7nbG/F9Ifn+rY0
sDki3IhhaG6AkJLZvKFoBH5vMFXBc7hN4LR0Kw+KXSXQwfODpJCFL+Cfl90Mb9Py
Bm5WyoLKSsv9Jg4b2Uf/XjfJ84VZE+SqbAzKw/WdOcOr3DzC+xD1+4njqNn02FEE
2uH2h45V2oP1kVvozG7eLMmRUhufCsbpoCkuVECkWAN6wOUeEHHpuMzjBN1WeFBR
6pqJ5i70Ol25YLtoWkXXqsQ+5t1CPUw1nlMihObX+hmsrzL5OvW3Sse2hUcJu/W7
6gizGetPDL3qqBw1a5AwOq67j8dYM7RvLE6dmayC5VL6NzBvvcm4rZ9v8zbbzJ2V
Yt2rmHkN9Oxrn4G5gHOMbuvSvRsP2P67tblffrhYITnppP7Wr45nGWuaKKHH63lE
75sZGHEQjoWJ3B5kQ867jbCW3zhJb9P1QNUQdGcmfophCpJchBdueRjYRO0gnLZY
ZAF0TUqiInO9CwJvnUOxsD91PCfWyiZ/sPdLn3QzXh+p4nfZ1GCMXr4AYu0Tfhy0
QP3wYTtLiQE0WZSjCHmCh5xbWJb8Xppbvxl3X2yOXz/nrkwVqS/H1sp3z+PrBcwj
Bo7Nj2J2BaX2SuwPwi2Kf/1B7CAKdGK81cGCxkEQgFcSSVWnpGsHUgahHOb0m5UD
+9d4xr3JmazHDtIS3zR9HlumPhQqyKhHeng+O1UmRze5zu/Y31RRy5gO7XRIocP6
y7nkMhECj1auAvEgGj217S0+0KG2NfHSGHd5u7/SqdAjJe8dRxqkOeYsGADyoHCX
/VMRuOq2Kish+4syzki/2LtBiAZwddnjK8IjU3cxcbTSjqbTMhCSAD1kkiVZihQq
xTluGa9+d5k4+5L8MDG1RGWY/WGleZU/7RQk+8VkaSUeyJAUvp+tsRi3xuvDTyc2
FqbwhegULCijhSi632mTA4yl1j0ZNv4/4Z49tdFMsopxYfEuhCvphBu1AOEE/8wK
3r1mwEf2iS0Hgtqw+qjjOMlM0+xlP9IDJ2Rh02ETM94wOweunEeeUdsXbKzRjPYk
qtRutL42n31HqBDOrId2mFBP93ONkspiaSmF4BAolDc99NSPzZzhCtRSyQLccbmy
1jpIrcRaTgHMdWJHN+FyYesRuwarfNNOmLkoOjRH6CRMO5WzHLmi6D9LVsb0XxTQ
qv9LwIbgLU1fAOS44Xp/FVPgIaH26ZeGnaeoLrhjIqvQvRarUG8gTXOWbuJ5GHmQ
hMfDcAL7+CBI4WMxVX4+erIbhotgPxi7UVfS0E5NkDIbP5kRhpB+jOKZ7AqOffgD
7igg1TfDSEW9Xcl9Z42aFuqPqVD8ox9wTTTbb1JIlVJsg9Lp1NkhSftIXFPUqJzJ
lpMR8qrDOZrw4PZSjrwiE5bK9IXMtdKPuOCaPaWtRKMU1oi7WwBmIZ4sbK/meQ58
DmVX97351aSb/0go6GpKMnDfWzFdZN5yVBPlOGMJcTmARzLvWxyYOArd9VA8YZ1Y
u+CXFBN1VKl4LTVMWJU2a45QQmRcrqtbtAqxD7h9i7t+Gm/fvyQpLqFIPDbd76p8
k2Wt/EAncBCMMJAv/QSdRXaDS5+kG8LyGqxVFe+O4Ic=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KVb0F/yMj6UAbNzcjlgo8R5Z3DZu6/7LI0OOLMuWIMUSU0Whjp+fvNOfo+mU9fJ/
s//07LADJJVkGASm/GEFk1v9YsFA9Efv1dgvMRBSIjtTQKMRbC73uQSjOc1P3OCM
1ePVtl8Sx8mWsAOnxp6DOYf1RofVJluGAeOP4877GNc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11168)
ET+haf9dp+cszjJlf+DRbQEuMCyppbJALmCwziMzex5haOqwJKxqwiIBFRR7AwJh
/lGHwqRI4AHduUHzM90WFbwE04pq+5hbIiDT+WBdQGRPmnSsUihg18F5gL4lBILW
lbdFSUUY/BKM7rWc/sVNxWDdKHhYxqHvw8T4pzL37hSNbWXt69gGiTrjgzT+oLVU
NYpal1exoL/LS7fUzClWUW8cPh1ko5YonV7u0F6/DFJ7p48TdhzNATt7FV0ULcwU
5oIDKhOjySwYONPfdwbt7I4MiQikBO8/boMuG0KwHwzxj0rbwPGkpZCJhLVHS6P0
kuT7btS+FyGuANxhWLFf5KYeChgRvG4fp/IKy8OWVvkp+KD7uNh5HQx+CYUpWtsU
OS5S7P4djxL29RLaWBX6/saAz8ZSXZxNCB7Qf0T8ZXJhhSE1K4gchmKgTHYENTlG
klbobnT8AgDjmnEQFD9c4w0iiafw8nk90D23jRdxM49QNo8xw0+5adn7+AbYCzqa
Qo745K3QNi2c/MhhGjZvtVM1Da8tsozJqZPNZBZR3/bBndQBh++4ahhUPRgS983m
fgf2xoAArymkLqasL8wq1dVGtqK/Gn9P8zLUH3JyGRZ6Yz74wsuxJ2Um8fb4Lh8d
MBsJVZ28sSg22giwIMMdgSGSd7sAHAJSLS6uYHCB9brU0ojL5C+AvJLNyc/nCScP
uy8Rx4FWSagKoVLJg/d/SXmaBLsD3yUFfmIzO6+3B1O+c/3xWtbXi5tGc94HqL1X
yGBu8DTgmz/5ic5fjx9Dn04ur9RYH22JjcOOOAZ+o1xLS7X+uXs7bpvACldhE9TK
zr/7ZYeArPseE+CjOWU0n90a51VCQWaSojPohENwVLDRi56pi4T19+UZwUmczG04
cUfGgMT7cST/DQpzSjvQlA/pY9wgmlhPrbLhi4Ma+zf4s7TQXPzA5oVp4rJgdTn9
wxqfmpdgPOpA724tY/17xmdnm5F1F4k7s33nrFVPJjDtMspoV1sh6XF1PCMBpqik
FP1MDZoaDm//qOj8h6JcEW3mHUIUOCvPDF60F6wPN5f7WkkXXS8s/Q78mOxJoQ9p
Mlbca62r7QaRvySMjU1lPwsnoAvUfcVBkqfgSjphFG1BXkRa37vnuCFXwZ1uHcWD
lbjhdvzeC+XwndFoWzamqtyUTPDd++4siGj4yGNfekMJLFF4TStsxu6D0TGR5fMK
5JqkZsQlPqYd6s+d6MRxMzuGWZAn6DzikqNsQxa6CQE7eTmloQzNx2KhFWrfTW/L
/zt/6Rsi+A9AlbKjfIIVVIp1HjYnENdeMTbNtDBL/x+Fbnu6T0B6jIaIjrRKDphZ
T1B//Xp55yXlirAN3VKZ2V7yHZmLQFdOr8V91AdEudKJX+fjOwsYxlvnL53I9E11
1W6J+txkda4fmKMfo9EBE2aJruWNJsxL0NWiedWl2U3VjsNei4QJ4tyriSg5+EKH
CQQf8tlOmm/SIxIvh09R+V9emHFb5sWTNcEZaCPImyjuo7ny19Lw1wDkrFl6u2Jq
srvFlWOuzdbkjyeKtgUrBpgq3q6XmYL5pXWlJiP1M9eigtCfSjY5cM/9c4uHRvSY
BpnzuiusGvheZVLLdmt90mwe3TqHaWTne9e8fJTupK2XWzz2aa+CmZ9FpiaVTTti
jPyFyUQcRx68vEPtuY+7RZLhnDAD94VkzyDmx54hm31atgapcAUhZ1ZFM8MYBHoD
A7cwUcmUCRPMS9DFGTypR+BRGKMGGbbONBLFlBpTgmi1OYBCDzrVLIm/KfLENYSJ
VvicjS0dh80R5jWZ7WB8aVeYNUWXJEb2byQLA+vw6z/h3vYm+zht3kIxFl6eH+ow
68MEUrmgeiWyndle0++94Pdw5bISKoQUkqwGQdIPsC5v4yv7yCp0Kf85748JLcte
mc3A+E6wgZwK9JGGP6KXUwo4z6KM27QYgBUKa6c3NbnarrmDu/WbMDjQCDhPKmW0
yKvW/BnlmBQJRGuffW9lP4GJ+fMutlueJ7h8RJ+1wNnScUkP6q1k6RYxZFpLkFn2
IT2HTiYRFGr6JVF2p6I6QUzQBWfbl3JhV9XoKGpZ9gQfNSDShwEkpBPW3/yzHxCd
e44DwbxiwQpv9brckGhqEjeeMU1l8FOrCSwcXiQvzHgP99f40MhR1K6wWYUzrDQi
7OXHHfI9OY9P8ns83zVxFmxTiKx6s9xZcZIsMGWlaDOAPJ8HxE0sV5Lj4d3DgMwP
rK7YFoNsjeTZb4si0LSuB0xh7tkckVCCD/UKmf9sXTawioizXRoA1Z4QFyeq2FIz
lbOcyRnhGkI5fL3sHM78LC+6QdcAHBHxOR4I/GqHjcanAPpOtAKx0cj7yokexVsx
OiOusjbDgix5zqiNQH5tqSPhwld2xPvktHrDvmxXwQCwobMx5jIUSBHsX02p/vFs
+sF+X61m9QI6S7N9hqaXAKhc1cNu8Tl/ZAyBYoZGbop3D9UDU1Be5YXbX5jYLOdg
kAVXS1afoBwnmt7v5fjmuZ6grWcw4oqLpMG/WxlMIOAwbZGvGFpQD5GFJf87I9th
Ae9dwwtQ1EgUZn0IyrOjkEB6bIjL9UY6QkA0kf1joO3ENL6iG+9C8lA6sh5NNrzI
KiHYG0ZLh4XL7vCMotED1OYXt2/0dpCKJHh1YkbUgHblu4+bcDMOWN3C1KfTtd5S
NEiVzmGFhp40/uS+efkBBmypTm11rdZCCMcKqnr1fvUkNmtEwXm72mEXoZpUG0KD
mtB5JhIRJe3yznFAwnYt1ys5KJj14Z4DhotJULQ0LmVE42j5aYI+DkbO5obbDqR/
ZHeLbS7361AboI8q2A+DTvrdTN1dha86Z/2gejyfLY9uXJ0KZVdSEfRlQJYjrV3M
4DUMCkI4vWVRibJQYIGOcCTS+cpZoOkfcPcHnX1tCZvPEXz9mGv7tmEB/ahiBeei
9JySeZXiF0YJlj+jzGYkz/VWRr4bFv9j4Lp4se+1Bvvk5bbm6wtpjfmlFuwBoJqE
EfU0XRTzhHacQgyZ7arFNKrpmA0eGA9GCcXVkbTDJylyy7RHZ8ZSph/2EXDMyv3G
o4xuOqzq/TB/UOn1ABO9FrhIpf19WN5soGrduRDGstg1ChPNEvaxRh7M461ln7sV
xLFTZjwsP9YXXf0OIxcFejRpHe4rqeDA+36ChvqyoIR2cVeY22/cyzI2pSkgDxQJ
vqhT2f8z1MSviGj7HGkRbRORURttbFiGxhyVRiOiEV3SKTsDDxJVIJU+FYzEIKOc
2rqgjd1HUrDq60HcG1KVQDldKHwwcUNZPtdg/hM8GsJqCgdkwq1C5a9ef4SY57Jl
QwnTok2UzqFmn2Ej9PUfC4wlDveWu6+jCWHaB+Z4U+P79mUZhjoDEguIDSET1iUW
BGUNOSkRSllJANhJJPmMPUBP7+/lH05j4BWpr+xdEHok91Wv4EFAz5V1QSUgfS8v
C1tbxjEemg9J5zP6ydO6CU9Nql1yYviFOYJhq3cwypy0N5o5XbQcaKtvVQm7BSJJ
fm2Y4ANkRTHzyqEIDtjiFj7lzAGSTClHLHfrCYD8L9dDNC44s4uIf1aLq4sZ0XF6
qin7PZe4px+6P/Sp4fHnBNrA+NgszI6vJHND9VZxZmtOCyXjOIGWCdrvBE6PWxat
Mcx6owWvBmqFd7/xtzoh2aibYskRGnMPgp9z/MJa8D16CTh7Kc1zHgzFKItRQ6hd
EE98YBbwk96frTKWo5EuxrqJUsmZYPQINR2OqhQiYF2PFuG7om850VSyKD8VJauK
8oooU1dO59CaVo7LlY+Z6aedFu3f4AySw+wbmxrAL6YZOYiDdClrfWdRHVpvwKjE
YgfD7VrG4R1nyELkXenvrYll0qa7Az4RbX1aMRVEmdy6vetAf8pb2T9z8tmOBXqs
94Xa7OwUlIMFYf0mmXqrxNhA3O3DhAsXtYgBC6MK/J9iDwNOOkGHq65Lx7YdU6x9
oN6kyDwLMXTrRzUyJFNwHyetIYcAo6HtKNYzCG19OWSxNtNdfm5RycKVUmE2zbeG
uywBj4/EQoUfg0hpEMFBWexazZpGRGdYMDnSkctVS8NlhnVM1c+1meRpha7l5p0I
ioJjj6e+H7rXbSOOi8Nl/GfwK1+BRYQE1WYDZTpXheWHIEqAZLzmZXSCkUH608qc
e4IXyFs+h/AWGSzqJ7GydBG0DOlfZsuc0gncD+HR3yXy/rBucacojEzzGgQnsQrT
VBw+OKMJ7GrA96XtBCyPAWelCTnhRGj2/JG9UF/fHqEywSPSb8zWszdjQWxYEmuK
qXWV2wX8MAbJgobwfVxVOhG8XA8VTdAZr7H+CTNv4OqzzrbIIz15CtxUrr5YKSS4
R3xrpTFDZKOAggp4mIpf9v+cmsyTlNihigTtu6uU0D4J1TE8dnprnF2rzcLKsAs6
rV3JzhpZNQaDFwZgb0dxiki9XW+ttfLgY4wipx9+nDkXE9OvCIj79TRIXUxLiMXx
kW6NGWlTuIB5Ai20/G+EXpEjLqAS/ZtcKvvhlUq9OjliR+CPaFwnZSflGAauWccq
w5q0thZ47i4GFPIN1CVW1WHk/W8njssBPC2zV7N9tBIFNhVEobO9WmvXJilUg0ig
7KUKB2nP+1AVLBtUID+qEEwt0Gu4egZ+Lsgoshi8N+Vo55wVX7Y9wb6LIVGqSpy9
gkMY8WAXcKtOsVQdWrV74rfGJ8yDT6ecrm0ecpBgjbq52tk7ABOY/nmxeEm/C+zL
QgAdrD4Z5BRai3ehE+WmiXv6NuOzXCp0QizoYi6cG+TA5nOIwfeWuXz5hvuKFk7X
aDDCf/C8H9XeJho+FIeI7Fll0JkdMwCY7DstoLgvZfh83j7vEqxCJ5hAcB9e/Jmz
FCpn/crdODi1RVpN6YIC28Suz7pMsT8Dgpp0c9dvCPm4zqCuLu69cyKz18aULZbl
93QiiTPdVBXo3xzMd22ELybXqIKs5lNTBnrUokpCY0Mx/4hkYXCEac/JGt8UFBDj
m6tVzOEjtj1CNyzXPfEU26Fb94GbyOjRheC6Fv8LcxP43zMPxGzLlsJgz+zbiIuc
0hxge4Bkp8fD6AmGXo00lP6Z2vfyWrET66rB8qF9Sr5VqxmR02Ztfxlr4D1Ka2m/
cGmwGhE8FsNslZJrLnzUK7hPdH8X/hix+h3HjaTStZQw/ecauAmZ5BZ7/QeCU6lo
RZRsCLd5N1EdzszvUY/MKnHpLNDRE4cQrIMh104yiVWalV5ZrTiEqBWzzF++mYnN
AcAG9XYvtpezjCucqb5it0HJBnvDMD49nAusIWRhRsvTNqzbLRVqW2KKFBMmDEUW
0fDAaNOce5TPitYN+QJGPDMcx08fWqPJVLQAbMRqPAvsq5wTkKXv9/m8M/RJr3PI
aUkwpHuV6PvrM+FL8ZYKbzgPg6lF9OWtTJwILhr5UN685qF/9aVulmrj1k99BHOs
glrcSHsm9BO0SZGTd0slbXSWqYFJjqEI9N3eHZZHWwnSHZTKSNEwElRL6G14nVhf
2JY8Cu5k4rwftrqFxZlZXaZmj1pLClfL4phn5xEksPAGRbX+90kgzIChUn/dyxA0
MzrnFMJxMMUca7NL3IiWvMyr0E2KYwyPx2IBSHrxgFhAAEL/q/NW5oKbWW+Jvfr8
nhqtfh8Wfu1ptKvjNkKidF3tBd3XOHIRV+qaZye1ztMNUe5GPEJkwj3Fb4edjHGj
ZBlUYfhP4qSKP1Fd/bL/bkHe8JUme9/H4FzJmFUBxhTHundhfOrNq4cV6nv2Wifv
nluUW8mwJEA4On9TGHJ96RlkZXupKDTp1wXOms4MgCVq6xyp7A0sDLdwS3RmYBWw
FKMWQ7Z3SoL8U4L7a+rX7Yu8S77OHEK3LTaOUIkM4em+sfeW3DxL0k9UMUJLoIwz
wbsKND/uibaTJhegKGcC5eu3TWDR7AmFjHnNHXQWvUQCIUfhh7sArcTRiM2B3ZYk
ZdnucSZaaPmfo9E2R7qP69x0grhdxRuwt0Ax8fmcsQ9q5qWzUrQl+SWr43Y7SgGI
73PzhmGfGpGXl5Q4oXkzRmDhUWDomof+aD/gY3A5MY0yn21te7de32jIGqINrl0D
rxL7h2zQYEGDhfC0Hrhmx4qASwTqTRV9rBEW5VU4mQqINEquJjdTBz5Mem6mwNC/
/Pf8Ot2yN3wlzeVgy+3IaOYpTRGtEXHVld3Fm3vbzwJqHIZut3Zl1mRSHgwbOHTR
Lgj5LwGBrOiSEq9b/eOBV9g5Aihw3DLOShTxOjV/xkpHRX3b5crIXJRbKpJyWd8o
AXx+Q90ZNDuBuQ8CRMkMbX7xFVl5G7VZaFkhEJe29UbxeUvkV7t85EE2iM0dcEYz
d4dDBuq4dOS/yOWfIlzoHJHaux/HpaI7AeE3aVCZYCf9n8djLeyH0alx9rTS4hZ7
EpddcmneChmZBBz/azr8d4b9ukzBrwZh26VNEKRrHqzGraMvg5Ls0F6vJ49hOfEr
9nOe+7fPy7IH9NFH81njO3q4goUYUW8odprkzBNSXlY94s6oPBTwyBdBi+Ud1nzD
ql4T+JeZonogQ29I4dJOJ5o75Cu0HjoMMEVsiId7GszoDnW9fUaNkbTqbpfL39rh
r6vwVuuUTjqkqqeGWkM/07kiaIxzFsuzV/eKWa/3I/EcbUq6jlWk2X68b0R25RZU
Q83NT3fXqQGenx0VzFOIdd2zYolfSD/XsCkdbgHRADEWX20Xpu0/cBm12aEb+rzb
/3KX+x0ncCZyZ66lD4kLdhqRifLrClk04i6nwQ2YT9HV24BPvKYKNYHcCQ+Tg4ZT
NKogVevkmDxm3rBGdBPdlbC5PjJQRpf2leh4iL/2nhUHvdmHDVMtH9+8n6ebtJ6a
dwyCDFf8gqBhnif8MMV+4OjcMqKoNnoP+f2XfdXTVYOdKjPbrOQaQnQMlkGJD3Dp
LjtPvt+PKAhw1cZlp2E77d8jdiuxL6XBXyQMvvx1gZF0TL2dXlwLkHE2ZiTU5pDp
V9tMYALhNRz2G3+VSA9mAhCU+rG1CY3TY0wd/aJOP9iPnC3/j+3t3hVZo2kgDhVQ
q6BUYMurtkDYZRcsSO9vTgak0A7pJ5V/YEp3x10goRcNiA3nlWd62Fotcmwtg0Lz
9zDFYTiScfXEAq/jaZWDtj/hrKuGlcsP0GgP67I1flgKuCkJ0g3PiJDyKHGz0EXH
42FNWeJPdkxKdNQg6FDwhAoVzjgJFJs6ehj5lO5i6nDWqSKfYiI8/CH401FGL00i
hfsdVgdw0NYOeyZi+L30zy6sMH2Ao9mrMlZYjPsICLDmYB/gsv1lOElCtyIvbg+v
KAsHRHR10yOje2CrxfCOdtlhI8rxRTkih2KxgSSJOVhftPLRUC5JffwZHHQE6D/3
iV68ZviHRdBmZGZMct2AgL184bma7TVH0DiNopJWJ2Ic2zUGg699mXCoXlrwGCUz
9LwLhJCcdY4K61eH+GI6EkZDw+3Ah/EKi5o5FliVIMt0Rkeh4NSSNRJq9KAr6ouL
XbEDbLGPsSChbeRlG7AY0bhfNH7vkAO9sh5nkzpN/J6jzm35I3EPdtgiw/bUTfKc
gSJMVktuaMzMdi+dLtWBYKxp5EvTlFHVwYUpdJCROSm2wUvFg0iWiW9cmvd93VlD
R6+XU0b3nKi7oNLMjMjk5ryIjpZ5p2fhoC5KCg5fSWOZuU/QGDRqlG63b2mqzliX
btTUftDxhotOWuyWDOk1VTbT8tNbIFOLsBQ6ngyTMBfPMUKwNajaoVrzXDDq8KlU
fySlbYwyWCoZHcLLeZxrJNSQTw/ylOFq5px4HQ6m7q+JbNAhz/k3TJkFGgN25VTH
yI6b3nEM/JzSWaBooVAzzXL1pCTEo3PRZKZHlR3WbmIhjguEEfGt/GgVz5MdLMRA
gkaBGBVjHtfqeSqxfoN7liFL/PaJUdxN3SZRXoDagtYJwxILXVZi+Rb7cl4SYLd2
6Buoimpvl7ysTxJZ9tzkBCOMPTZqa0Zt5N+OzoPRCNxaC5JpR3g6Uy5RQi+7nn+e
nPOP4/4uYN2tjtoenq7hMOaKH8wyPl8EvQBGZVzG9FubhcTkVRcQPzT1+939Aaq4
eso3Ip6exP72IZ2Bo9u5oyXiB1+Qt7hLn0tujhNmI7oL3e49gydvEBm4cfMdPm4L
/K4+tW+hVjDFAVdZ2Hc+EPjyxK/i8UK0zWGnthrCCTlkEeHh/rvbUZ4rApedGS8a
lJkJwZJXh+LePCpFHmTwSi4l88P6f5fqIlgkFG/5hygsMby12NASnz20cxk6592u
Ih9rrQGseRe/UmzVb7pH7gzHJzhc0CCfCK3mE4OTzRf04Mlas4bDRaJbuJx7NE/O
Y2YNqAxODeI2SffZl3cK9C08BLxQvzLurCiQlkMAwOKzKIDVHbJ9fvbbRthAaHrF
tkwxwpLVSV9KYEE5O1m3P0iy2EpoyZjBe/5MxCCbQhlEyNHqLypEEUc4cm8TGBk3
K4Hwl2QtrUnUdeoliuFbVaWgDTBCIdO4ZPToXb0cn7kcac5i9wrTcjMdUv2uRKR+
lgPokcoGAfUFnGQpgwiqhPiXQGjhbCNsgi5VDhzbEH3IelLeaXj/kihAnZ4YtSOb
Mt31wipzKm+3HLEYYlFsoC3176Ps+obU4rGjkeUt/jtHgrKSeyk8EUaFW0HUC/jI
em3p2d8mRo+7LLDfRgywWTWnKXjontrWa+v8NDthetwuGGtJMojJvA5uS0Qiqy+n
vl5hBD8Py1Nr7OrNwdbm4pSHKQPeiRvDu4viiYXuNLgDOlUsmyFqOTa/E0NRkwja
gcV1CtNCZalepPH3lmX7RO5UU4CF+/8oh8vH6wqP3AHixSMF7E9s0vNYISrYzDkg
eOzvizJ126xx5AFRsYsY2StyoigcK//pcnokWYD5qb7UANzTu5zTpuSV0a4LWgSG
WpObJwnw/moBihwH55BlnnGMMaoIPrc9qre9wyFiJaWfzi5xbjbBKmesmNmF3fhc
TGqJFex4hZb5CR59oKtT/3bQiChFUQfNziPE09DVw8Fp47BMkjGOPJINrq3PjCuL
XB+wqfyYWQk7lE1uWeIQwCzcF9Nwcsxlq0GP9UhwWm+kEC3NMjJAjt3IMtLc1lh2
JJldVNCNEUpU+XldaC5qeKGxRspcha+5vQCDyKx9wVlAcdM2c2kwRtJ4/YyfMVCl
aofkx0YjTn3k7VRILOCiNx4M70ncKxM/W1SsJPSXmdwY7muQCkC34AbUVcbEkw/o
i8je43w1kB1imD+RrO23nPTALQbuG2vET7MrCfBQWjnP2W+7fWkxpW8Dfd758uEd
X53jD+ARzn7BzVkRTZaaY6sRXDMnbKNLNqLlJhz4xlNAy0frJg4Eu1zg7JzzNki8
/v90YP5wx4IU6Tva+TX+/+8qGN5N22mNa+1DeMEMVdD1Hd5Px5N8pED4K4/03YUE
bfrk9QSGOUlVBAPcw8UP6tkpDXWG5jOk2Duu+UfigDnyj86Nj0pLGexAIBEWVEOB
krPl5POcIVnk1S34s/SwwzzdyTGobYpOkl7+A9SAsJGCEMLpdGEsSvuNQJZKMWyL
g9m1winYwVzmqdWZTIoT7CBPbBoCv1LOUdbRQg+41fY1Axe1x8lOpui2xP59ww/a
ug9VAKf5ez5T794XxBXrWbTHiroQjJ/MA8LT8+v1VDFd6W/iw40OzNtJYDcDF/38
LaYbGxY6itqteTRKq4edFz3ftJcT28vMjJFV0t9JLuosyvzOMpe+ryp0QsiQH2UU
LQx2HGwHSiEG3JbtTlyBr3Xs7UvHKrNbkLvDnpGq3Lyd85dzcI8mgPhxhCsXhr1Z
PBF5/Ou75wDh+hLgTfNEOzEh5S4RZBXq5BW7XZcPQLSOsygToeun8AE0LpcV44qf
yVALUKMJzFkliyCht4lz4BUwh7Yp5GcoWWnFgCLX+zWkAPEu0S399rYMFFoy1ZRi
GOnmbblo0FQOw0MDETsIPpmNO9z7UpnbFo61/8GpUOLNKkW2tJikR+UCz7le0Ad+
KBnlyVLVUNJIpTQzfJt1mcATn6FhZJBvy/ubxG6NupvnPULEcKtGR9oN2AyssQIR
3Ct4Sfp7Bq1E683c0/A9eMGBIo9j/J2GQDCesin63wfdMkfre81pjKqtJR37NM9M
0D1m+dbN5v/Vim6mFUlY3mJL4VRXUp+w1qRYTkgSFqOn3X8ZrXlq2kf3IBywFhay
mY3cSxA4iC8UDBdwRU5QH6fSb7ztkp9ZyKRVG5plP0K4UoKuQmP62XtjjQthC9Dm
b0vkdSTs9mBjhugPwR3OtjJBL/Czt6XBV7J/nBBNrNhK9vw9SBxCBlMgNTH6Q0hQ
bpM6gjsXnLQNO28cvSV93K0vnH2DvntSYjpa2WaI96p7n4GpWpizbw08kw6BkDqb
PLWsjcpr/zleO3MPcEV1gVzDW4EnFpOUXL2ZuVqFpv6XqYChPEVtyxg/ikp2imLG
TQX6wE9ICukv5iJPZ5Ao4Huyx9KXq0/lZ9Z9uIeQt2g68yvTAELwY8tkm7ZTZfvh
iWwv3V4k22q/S+HWe6WAmV5FT82b86BHuyuvaslcpe3dK3HeHc/hcptrGfTvfLMc
x25HznwMyV7+fmv8n8Y7R8c4JNilFbqEvTRfuRSe/yFPYeuVre1F1oEBlxCtf+Tu
0SYwJpwNl19qBv9blgx1QGTqsg0RTTyJOWiU+WijeedPzx0uZH2SwJ3L7M8/GYuE
TDzinm6qasN8natK+xIjB3DLXqu5L1Z6BvpEUrHYh5ypAhHw4Gt/YD2W/6jFmA+T
D2MBfKoyCIOEnNR3JRsvGBImSfPwvXvN0w4vhW/oiojskfme64K69apyxTpiw81u
bd9cYXcJ6XZ2zF2SDAVs1eLbPWuAweIpg4BL9w99Azflylm4y2nB58jankoHbsH1
ulw8wX15X2HdABTLgCMScswRG4EYC8jYOhxvGwm1h3MXGLs6NYxyKjrDH0Dpkh4U
6OCT/yaeAaM2y/VSYv1teAHtFFA4dIJJRVPTNJaKP0rWu6eeRQvHiktd4sbFKr1n
Dc9L3uRwA4RzVn3McKL9eSB/n8O2jT355Ly8Xg4tDCkIbcsuFMfRIGJWlLRA81Rn
hj+Bot3IU8u4/EYdmEjY9SnT9N3XgEqCb7fWfeCBoL0gJoTDXWHRFkKUK6huhc+V
LcWIImxtkIxNQCV2mfPuYZsg4/r/k4PzV6qRn8xdAn28nKotQXwnA/3xENXHY5ij
cxSeYh9q9AnoCZamXDvoZ2J7GfSm6L+GtA0LxB4Thf+Doa0YAIg6FFfWosHPPH62
21ZnWXWWqVMCqV1iuNeK91+uoiUHLq3QA3JtYUuqajXlH+iouHcHaomVEdAYD8zh
ujWvWoYsFbIgPeX1v15TpNzbe4xep7k94T/PHBtiD0tpFX95SFMYekIb1XWikOYg
wJPVTiDpLsq1eTgve7PrVkooLRP9sSrtqcYQD06Eb+/X2I/ruBSpgx0KuYRoITAG
D0EdcHkUXX+OK0llvhKebSi35mXExGD7rBpJ7+XmYP7Jz2x4jBMRIfLBDO2qGLv9
96DMB/ENXS6x6PPAsu15UQeMizfwF5tcgD+u2XyQdpBWPteUmB3B82RK1BpthMvn
MqXF/sWoe9ACDZDdQbeavHPdXF/3jHe1Bm5FRBu0OmNlawq0kdtdr51lf/vKg0fz
EAJdL/YDr7i5jEeYN5NfzbtU6rEVbaLrLuLmTmHS9ilL+JU0L0MnRKEGUr7qPICu
47TwbxO2dxDh2p68rV97Oc1j2b/B1iWB/a+RlGvQ7XAc/YQ9inhuOmWDeFn/2H+R
19LJTVT6ALAwU5kn3QnrjjKwzNjVDinIYcyHfT1aMkGmD5vnVvsa0VzkB2eEAJfF
YHzpEPcnm1WE42DIJJPqJ6WnY81wuuzFRKtuV91tZxW1wZUTCmRrvoNKi3TYt5mz
s06zSnCe8lpRHVZYoA617AqnjXJ5aXgiYTWkjicAFYyHTp7DrpIkaVPp8c70mImG
NGl6r5aAOmHTtYpW48RhCG9OGNgc4T4aRpH00yAYp3KDRA4u0DeoKYJ/XUvv9L6T
ZL7xFM11PSmtiJojHdQpX+p1NfesDR71qNzu29T2pPFl6h8x1bE2HDRJkKfutMaq
419QqnOWW7is5tnlIEC0XSBI79aJ/c2pYd0cr75kKhp1lR8MA6bQ8x/tEHdey0q7
Sk5rE7YVT1nVRQVytBTRmOZFYU39JualdJA8/fhD2YnDi6XI9WX7dpsKYdZVOg1e
D6Ik2P000zLX790Yw0xmHeYBBeVkKEHtfXCnkyoWipaczVW+maMmrs1ANKsavIJi
j72x11TVLOk0/8wxwH5OifQGi2djz8dYf9688MU85SB3Zx/Y42/K2NwwH6D1/wK+
7PcNt3ikfBQp2QvIB3CqJG3B9QhvG63IASjT3UxshGQ7SmLQm/xN80XCofQrpJps
tjEKY3q29fZRiQYOBXXs8CRRwzqo1lLdsyxvs2HgboREunYFFdJo/EF9qVde7sK2
cekDa04SE9ONz2ksaYRFToJ8J3Q4NOOJpDOj8EbVuRRyGtCeSjna7e4outWuejWw
0AGn9EOE1sfxFXLaHA4KwdKesAqud7WCgxHp/CidrWEDMehnpjwFpdZGG6xK6rLZ
r4XvuyFWi/wikiUfhewcM98bVCSZQoJvZ0pZo9po3FE7+nl9hrRYMBP2ay5Kye1Y
Ra/qGb7lN8gNz7S6FSDKGq3UhH/GCxCKnJGLuDm/YWuHzZDDC0Ojyngxce5LtY/J
O6zlh7322b7jrTrzVmjJAddUAN07Yfvaii+EgQU8rR77r/1/uxY0y6E07k2w3stg
GZqySQ6H2ZSF3BYsrJWg/0XWgzWEsb0bNwCrEsQQNyBCYisKbWF5u+dz5uaKU5If
YqGQw3MyD5Pnw57hgFwyKMvySEC4X0ZYmlrGJv5aC2A1uamNY2kh/rTCxi1tYPj9
jtNpjCzcZqHZP+LyO35zyXtg0iUGkjtwvnbuZLLWyH1QDIJwTI8yDinTE62ykVrQ
FsXQFkyAvx3UBWwWqs2BnYjeDyLqt2E6YjkexXCsLKbZXSJtjh711/+YF7oAMyfv
Fv5UabWwse1pJgojckdyh+TIvkKPtJLOnVqr8/pPgYgOFuDS6cIrro3GW5ZlrZN/
XklJo5lfmc6WsEn+JUohU9obqF72ch3JeobqTuRynRR+nO/hLDuGUCSOhU7q3Rxe
jutEf6dyXyZtMD+ZetNPxHQhAfQvPLgk6vTlbXozAvsNVpOi7QW3fbhBc3zn3Ugt
ekiIQtdrszRgoj5xE/YMbB0qcmitMFGnIKHDWLeM09J3N9w1QIGAfbc6bQuXhylX
b7alRo+DC0eN0SmheC1xPCF/xyR1Rx3sbMYSAqXCJ3a68kb3wAdDqu+XXQeGpzeR
jjeTiF3ELkUU2LRYPakoHucPHqFOcslBLo8th/fgSBMFawpfkuV7ba3nX0Ca0p0M
rGCE9mf8zPabVmZQ8nz2gNhdMm9XejDbCvun1pieCxrtyCTpq69g6pD/pgWjg7Oz
RTuIp/RAchy47wDcLPsmAoY0nRx653VLTQhS8mwNokHf4xj718DgR8JcIjewcBNb
qoh5KF6mXBMXKw+5sRjNiNrqxXKqC/d2+VZIr1lCjexsteNpD/ZTwrjUskSDfRqj
KemOJseIosOoRLw5GKgRcGFVcAxutrt8HDAISHKSJ8H6+WjaX3N0Uv5Je46pBHUQ
yJWnr1zztXIJPx/j05/t2yfgWV0DQkpmBPX2MSghG2qqB441i4uXIvD9vSnOS7zd
k5PfA+rPGTWhLc0EjMx+6KHiI7KEHs3g55UGQiVHqgufJvoDFKjDE7UsJyBMupfC
/AqixRMHBAZh77Gck5U7P2JxUWR3qmVmaYw8hV2K4MflZbE0y+ghwu/msG3mOXAL
+stWsyvt0gDt1dhy6dSFMq5HSf/7no4ZACMeBLHE5p2gKsJl6qxQeORTpDpRM0Dh
Gi6uiSZTKaWKOHS0IikZeSfCjk4tQWndqitPixFAMtdlMV5Mum7sPC/KyGKxEV8O
dV+1L1c3BrZKQEEOv+3GolquKUYy8p74Pnls+PEnsxgtW2Hp1mJE1F24phPqatFk
msSGdk7KCXNBhV+zFAwU4dp/3aem4negwB1mSI7wHXO3USWLGVwa8IRUZPczUFHy
IHXMwzBSthijMO7I+wkMyGqkCXFZsjAfSuQR7BNVllKKW+OjvdsQ0lPX96w7fPHU
X8G6vbOizrNJPm69aY3sDQyFkASNxp/IpXanGl9OO753QB8cQyFXIvFgk8gsLVZG
6vigv//Vg6WxBMu8f30MpITizJq9gLI/p1WwRo48+jln13YMznXukMH0B0oKhISB
BXHb/AmrOPwwHoFXF5DniuRCN2mCQUAWvcmgpcSV0xpg+Byrbh0c3SRdJYpGDW8j
geKxvFVjRGw4w11kEdpri56tBXlHtpQu6XtMop1hkCDtinX0AouXx4V0RwYDcQtF
6OZusA5cOjx2yOImGTRcmP8kTx6wtE3GhwPXyxyGM9Zpj4rxVQrb8prUdJx5ZuJw
j7/QIBmaLdphb0/w77jnRoLzIj2a98HpJ/d2KlYeuwlRlJyaV8BplIi/cbhdwGbP
jg4tzZm+4EPakNS7wW03fsOhFVPS2sztmuu5VUZUU7FhYuatf4Bg2AfGHaT7BrgJ
LNIqNrmZbpPpZWfjNPGMKvmXLtnPapF0NVusoCccNFa/kGZu3iuclNYgGliTPn81
0P6ttihMkvgePd9A6pZYOmWgJDbinJSwRqi4f0R22fVNYUibt3VBqVRmtOE8vz6q
5bzdKRU9iNISeTyQx7mgeTkBjZ2coKq+AIw2SRlfqpR3WwU7Cjtl8NH43qA/v/kB
3fAU1kvNf1LHq88GUKQ9uurmSenLcsaYFNrEqs2fces=
`pragma protect end_protected

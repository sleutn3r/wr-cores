// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:42 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JPAw5cjPCcQzQt9aHwq20INWEfLmu6k1ucK0KyVjYnUjEMaZpcnXxzicJtGK8g52
7poZMJEKEwHEC3X4qJMPzu4PtmXto9idsa7RnObP/POtTUIXsI5odnYhclZCDQbw
pZNGSDJIaFzH0qlJjCX51LqyglXcxjPczDWyXUtFx5M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 47808)
1/8i7IMRUTuapPxKxCjtL+/yURY1lfl4Z1RRvI9qOfqTemi9BtnICYnbeBkhVJBt
Hyz1iUrzRHhQUWS7Dc/ego2y1P7jdAmgO3yWkkdFoz2M9Egr1WcJ9sMWP5WDQFxD
NEk0PlfcWgICQgwEDNfTC+rzrivFctRvqI3F61KJyATRzXFPITYqiNn9foBa8Wna
2ZE+8WLjZhggkaKnI2PCXs1FIuFAah6ya4q1h5s0LubvGQZ/cQlAY8azM3Ezx04t
XV0n58RUyQpmwQiujznmQ5pP4c5ovp776QGiLXU5w3VIO6hW17bzcu/+9AdhFayR
lSdQnMfP6/3XN/lSK3GkPx3Z81dp8nqLQmVo5n12VAuLpP99dscCZkOtq6W4WJO8
TpnWpNFJd4ZfXqwLDa4buBrytOHTfWnL0KwyPuk33HxuPxKdidTjcGgDUrRuM5II
9u/jRbcSnnq4Y7KmTyRXp8xzbBepP9sHWTQyYm8YLjxvC8PAO2nqWvM6QvyXtNG+
7NknGltWWNDkbCxmpryDI3WvK62EN6L1blYxjcwOZRmzu0/pa/+l3QrfX4TV37Wb
g69ogk2iNotrHipSgKRl82olySzJ23JhArg1n5A3WGPBuqnXqg1/TSGDYE7s20VD
dYfYgKy+EFnwh7Djbv8PG6utL7HZO/esS5kMWhhVkT2w24vPP5/v/jvkeAZkS739
I7eRruZKZBz55jxj2MYtpnbdHJXOWR5tOO4eKSca3KtqwlpgICizqSZMZm8nVYPU
6SJ5DC+VWNFOQ17295GjqEc6yzsBJ70n4TpDepgsS13OtBtrMyQgY7kgtw5py5FO
a3jibRfjKaJp8MUwZUoIbjv4y3gL2EkcjNCp4IX+WQfxowmgQCF6RfUvuYqsSEv2
zblC3x4ijzmnPr8kAymakAlUg8tkgzD0knC7r7fRHhVqWNDvFZCUhdbl25WV1wZM
weWRxELNQqBegXWeZeozr7lIhfMHiqn9OdIqAsMnKEs+tTjtUk9th3BptCY4U5Px
2YQ/YcEEZNDWvh84gYZ/4ouGpsjV7QGHYCoFQp9bLlThOWjDPXrBFv01UalQuV89
mdyn0xfSMSVyWMGmv+tGmsB6WCGQXCj8eV/8Wy3ubxIDAagpzcyV4lVDY8/tqOBD
VBJ7TJ9nMAw4HUs3OAGWg32Pa6ElKT08jcGP1W3b+XVObPwgVI+ZHgXYAjzs+fve
z3Sujh8BFZ4MkByVNv2r/fGz9Eytl4kILw0G5LGbVFCfWfM48V0goaDWx/KzMkE1
VFjYDGD/J8PXm+D1FdvGGJMW5ezdgvmT2q5b99l2GCPTKZJkJJ7gJIZNh3UsDwHw
ukG0Y6KNmiT1n8KAvfEjkZz8LG75k/90SuOjEp33Djkh+GBaNERhO+P9BlvRxPxH
2bN0czOWB1IuXM0w8RoZfFtA9ePF7EZbXhwF7giQ1vcE14r8KNuFInPgfZNBh/tX
5dsCsb52rXkK6kM5uALpEpfMbGRzBi4Feyl6C/jTfGI6GpSukz809beS1ihF8fCs
trVyXlrDjnCCZ2Y+ZG+5LU8TmNXtZmScAjpq2VIZMlB2nCa1K5xbEkY/EJTt9dCt
qLx1Iam3hpvO1Syo8TAQblgS9ABuNjYWH6uNX+pZfbPnEb9UadaRcVzYueOcc6/e
8ssXhSKrRGuCukqxMpQqME0Lxf+WflIUPsJQ5Mq/CehOrmUmeen+JOzmADuI06fl
kJPuBTKftn8naKdSUVsfdBt5i4Cz86L+9DB9FX6kP74V7d84F7AMGLCn3gzsmTo0
nXvQ25no3W39lMysrrQ8hbFj0VES94kRbLXD0pYuJ5c2WSjHk7iCdNpuduPQ1kcb
kwDpfy5myxKsHyMJmvGUqVkHb7+/uPU2u2u/BjXlgZTGDdae8SaGLxG2LycDcDyE
ZM4LfiarEHkUtaDB8Ebm96cMf4nDTkEVARuiTcs+QhCyhq4PESrG0W3+F2NZRrh3
Q6ErOuN1JlGJWqzYBcT3u7mCfTDDV8Zd7RX4EnrBKy7/KKEyQHk7r7W9urjGh1DY
lNhph+p22L9shVegz5eQ1bdZMo7iq7NaZlXkiIsugwqC3qSdiCMCubz3Sr0h5zVp
N368hHj/6+II7as7QBUdNbx7YprKV8FEwVGsM3za5VBhf2S907czE3F88/s03g4j
kyKZzcpNxmv7AGjJV9L1mcIA4gLnO3fCG74rfONPa1msLG+lm5p7Lmzktwm/511N
sbfviI/6mywjyFp973TrVVwUTAB2rl/vQXgiB81Sz4OPmh9T5Gg197pfL3yPuXl+
nW8MFP7zNTjt7BxUPq1VbZLiCorlvtmNyRjMSHY0HsvHyJT3VCSk1AMuIFwRiwcY
So7asMMFeD7DFCfeHqcM4ZCibLZfdcF5PoH/Lv+q1y6u1YCr71C504Cdvxy/vOLP
GNQxgMGDEHfJWefKcjvLyr8glR9+sIkTzW+N1i9HeoNiV4zTFyPD5VKCH7wdyPVh
4mzr/Jq8WTV5fJkj7vlJRy0Kq7RWtTEBdeW+CU7Un05ufriEYylWsbyJc9Kj0SHq
rqY+UFPXkeKT83sWNxQKCX6iteRCy5jMNGaHPPOqE5IzUVnN1VpVTWQ+vyQqWWoA
A0stF/Xcvg9X1RN6v5VIeuON0abhR77h/2npO4CcFkFkhQnnryK3dgiIySaPlocc
+vneX6i74xB1QAMmFgNypyz10V9HHSfJGzZQqIQ3uMOLaxbwfrmLsgv6jFkDjGke
BwdxNfcrHSnYbQKwIgEE0K/pHCR+cLTY1NnKkYMr676IPh2Kg6TyApt+P3XCwxpX
idGZPfUtYnKfyKLZ4wtk/SoNzBlm2M7cmyF/NFpoOcsqMQ7XOJpU+pN89fYgFJry
VnKwi3evb6aS0wp2GAZ+iNqau+DwAcu+Et2Lhk8xCvcBkuJ9VAINkxIjE2eQHh8Z
Ts/3Cf7ZccFJdOjrksqeXxH8XMUeb9uehfx8+Tq/ncTqy+6k+URrXTjQt1/GMixH
+1Qbv33mvtucsPmVLLhGZFlyL3tgh9aNZRwOXy/054ZZT/56gR7/rKAwA6nwrV4S
kU8K4Sc1LqoXCXFcikNteLWqC6bx0eZvLNwozV/iwYGL5yoPnfSk1XslHuR85TJd
kdSaWfo5GwE2YoMbp3HjNNKujJ+e5n1ioQmS2DKZoA5RzubHXzKL71VqZRP6QT+Y
bAWBTTWHUgmGY4rB4eO4o+fHP1aB7qQAxgSNPukR1ZHBirl/Hgs2awH97Uy+6kAH
mVNxeThcTWtgkjplWbWvcNWDrrzHOkHZRcC5n9dGGKxCoX19Owp/+V+90umh+k84
cpsybz36glTlodVZoKSq6/Im6KgahhfR1R4IlGoumurzP45QMDTIEqxu64lyfGdT
VbgT9EpTYhsVaqDU6QQfAKVkTq6ue1fTC2tmnzvPuL83XOh0iPHAIWcuabq++qud
LyIXa2P2i496/09rIM0PecCij4dUC5OWXvooZZPOqHHZkjuYeUKk7Em0BXtLDfNp
X7GdJ/0aQNlHCSX21uOmdEA34zUeyUNAuHyoWPpUEzKF7FdX4YjDwbPf2iP/1cEk
VSgRrYFsk3KdRtoZEMvevMdJCey8nZJdQjr2xTwQ5BRSbkUz+xH5+FVsVWsK8CMX
pcHupj5DkqWSHzBny3VgKqLdPO9upyYEkbUVsLY9qEVAMxkqf7W7uScl1GrXRrPi
zWlbibNASrNav6so0AE8P4ur3hsBJxvoYFpma21b36zmWhgjYFGhDJsmA/Y0NuB8
rDTP3B3YZmcsxDXUcQNN9yIT8iqvRwGQtStWWANxkaQZwsHuD5n20kR5Ed87kB3n
rtzL3cu8xxY8FpKMQbLyqpaGoutfxgDT6i2PDoC2Woy4e7tOwrB0nWJhrP1hBcNi
OedUu5Iq332hlvRzOGfSM9yrHnWt+fhTQST2l1iKScJtEMtlzfqR7gWdLlTGPKAd
jc33K6QqHUfkMIYR5tm58ANOaZjyDojkk6IW6mbTKnPrN2vzFPhYdHkuTNcu82fc
NsZZ6UBarKgnvkme0wJOD7NCPo1oMH7Nwj4z2RoovWGmYDepPQVjOgkuGcOjE6An
bpGP9u0NwRTb25uq68JWgPRey6DimjPPyVM26vgesPigpjAqvLNkH2/nbYVR4Zic
LedCOGoQQMSRPg9BXSGpXtvartblcghfwvVu5WTFmJwx1UAYMjPmfGSJ60x4kIg3
4j29WGPqdNpGAGcdpuogSpTyAHmrNbIz+TpSbBbz+m4iZMGRoSiau0LYRWydwrz9
P+JxZP9PzkMEEMqayYFjKfEJxLFvt+/FK1gUELjrs0W8rQO61kVvtkgU3SICFIUM
UWd392FNT6CJNKV6tlG+HLwpfWnXy5TZBVlZMPHCJ1VYIp0nNIhB97zmaF1Nh9mT
b9hWSFvqedUK+csJ66kFaXn78xdgiROC1s3Jza9emGGFWpm5QzX1+HPymlZfvhmE
jzGKe+syWlnFEasnPTEoJU5dt0PFvM58Oovy7FvyCky3KWl00+JKBue2AwwMs5Ek
SrFoCYvPXXWvQm4uc8uP4rZOJnFpqDoymiOudGR98cfp1jtT7nu4SsTrCaIppW+d
H0uk3BzJbhNbNz71EMvuzK/W6FJQqIwHKRqenJ98H4LTAtRPegmUQUFCl0hhLUd0
ARLpqbgOXqusErcL3t3LSVpp+DV0i+xOjZdljCxIpSS5VB1FxG7civBJsDDGJWGE
wlbjbV73pR7GNoIjIN8lIq1C2hFimrfEmmMliTdVtyOSJl/9ONhymepuOk5puVbH
z9k+pMczSH/3EizlZvBV+kbFUUsBBGtfypNXZSkV71dck38vj/nq3lo1OgaKJj0x
Wz8xuT7K9ljyZZvo7D85YoO3FRqZ1DT8exBLhNFXDs0Mc5OTowXytNOZePYvYE2C
ta0hd1MtddX/ObTiltiCAr07D3SDeUQeISa5MnQK54gXgWfN99Onthguq+h5HkJp
RMm+KPG2vSurevV4A2PRmIIYTN1Pl/fBm7zJ7+R0mSGbKDQb9TUHC9/KOoztPJEU
Kwiazfl/S06turrmo/DZgzHOPyLvekrYgS1mHfMuFVayQYvIt+aUk/ZbG1ZqR1HO
Y8u9cqV0ovDVdWIiV309w2h+nN+7e9ea3P6d3jVRrSVAqA0eBUub35ti9ZSK3NC8
dmm/bvPYQUaD7qVn0CbApvICBO2A/vnMIuZ8Z0tNWELN1Ol4Mqq/jNq3zngTxia9
+EtpEkdIFfJFXlTXZbZ8UBD3dFUuD+qzO+mgSdLulYm8TlR+EsahFbcL1nDO036Z
nEHwSzltTizpH+wSfOjgQNQ7BgZea28TcpANYrIMRzVMVS7kGc1tbdy3HOk00Rni
Trk7MVPwSWdZbz/gHOYDvgRt/rS0N/2RAZ+KVw23OKKFBeQHKar7gG/r7JZ9edPQ
JBGjJb88c49OqZC7SgTmgUC2aHaoGiM345dRCtt0gdXx8cfNdaigUz/C3FqEdscQ
SyfbpDxlXIg0Uis+ndQf+G3KUtMpQwLzl/ZCbAG0a0qBnoqCYjV3zRiCzjWUDrAK
rmd3Cwq9paBBD/aBYtxMGt0IV4MSEX2qcQPWhDCRnXSLGL5KVSdDvrk+erOPybFZ
rJcURoFxBNrxJz7FudxjvhxDeJ9Ly4GBd0XWlac+KQGTIVTI0xEo8BtEDBAFFdGJ
dAuBVaqS8Y3WbKzDSTdSefwXMUOALVG2GDPWLOUcRry5zhjfXGgRT71XiusUxA3v
qbqsG7zDpuDuqBRpXrvTjhwELlaDOLiJmhw4N7wIAEDNX9/GTqWlySOULjad2Zuj
S4Mz2PqBPn7R3tEzvaAp+b1Tmvqqvk2Q1sYUvdKHpJxpgjufqgwlDt8IG7qy5vfA
Z8/5h6gDC9+zUlFT0qsy1eu1ZukAq5IC03ld51yZFUVyLDlYyu567+0BJrAod7Fq
5Lu3hDqBnfvrIhdH17BQSeT640Zf51zFW13mGeK9/+30AVZKzhKvP2MSrSyemZay
2f+FXIKOh7wcyQEGe3KgSWo0nojrYtfvu9+dF/3Qr3ZD1O3CBCnimo/FDx49btdk
n6wo1YWKJnKln8nQksTVQLusG9ZX2IS0xwQEgevBZzlw9nyZ+3no1mhulBwiVmGM
iHzhTx5BoLdjbocWcfSGfdFgKae8ul5XgiGywJFF3wTr49158Ka/TVvNJpCnbJ6I
wXPCdH55aPjac5IgWX+w2IOS8+SmsWuK/gWXr9sN39qI2m+hdNPHJs4rVfTBTEFC
GqCst/3WlKwtAT3W2aRG3MDUfSuDQ0i4StFeX7uUu/r73IKm+LHQzlfp9bN3jLc/
fSl84/xQn5iHi0pewlA9Y3pdV70c3zgQiGwofS9AVwAIWmVljw+a/bib45QNeaom
hA2G2E9YQ1OArfQ1YNgkB8Q1DYJyrPim/RBrURIa5fm5kWjDdX35cQ/ryQwMcA6K
kGuWt1MF6cUu53xreuaj3+K2F4zRemRWCejVVT5YyB056/6x+sW/LcwVe3a7eiBF
e9yemL2r+Cjj3BysO+5Cja6izZtawaCTgqcRZin9xdowLsh44Ef8yqM/UNKNSjsj
4Gf9hDDOxLpZvgwQGhpTfeMSAQ051Jsn88r89+ATA7jtBkZMPxc7Np+r2vjf9zMe
9KjF9gggpfzDTP8xIuEoLyreiHKkOzoppHZ+VGAwe1iF/PgQNObWIneJFF092Uho
o2LY9L0VkT/ovsKDTBLOaatIHHW9JojA2H5HMA/1+HB99YA9G9SdywTdYMYfnrGF
mz/KrDSCR9M/xvvkI6emg+xdx7C6WsFkGk6wFC5nJGLC7rOlNxg45M3U6Ef6Bwlw
WZNIMW9C8F3JGNjaTReJXPSZ6o7uSqWyCTHiA50Bo5UeUVwD5Jdq8Ag6uqPCZ28/
WwULIXo7UiIZc3ODkeRe0nubB/xhAyvMpv2wx/mCaV27n2YHyXFFQt63zYGrf2/l
DfkiUhGmAsh3FcK1ZMxCzGrcZolvVej/fuDXFNbZR1+bYwldrMUvK9pxc+MUEr9c
zdAnFvXEzclz8X7HtaCrvbi4yuA2gSv34sXGALDd3jBldRmyjlbpd/CZm6hTBDCV
+Zz6RGxZ4VkA3/TcFDKxtTfF1q6V+Ne9VU2yv4F2lCFYsZPYMMAqSiE3H8r9xOoJ
MwbdhqAypptTjGgOzl6N3hzDsxK0Jbv+zVEamYtAFE0/EArZVyNBU+PusVZMDhXv
SdCI2CDDp4Vtf+/fYjSl9ptycusXzjIwcJNRr8iS/3aUKT/hj+eyTSl+xHJhpge9
y4uEacBMw+Cks7ygoFXT+6JmRolyV0GxR5sRme52xA0NkTY3fX+JE8sJnR/pOlgK
v3//p6Lwey84AF99Lvv5I1VPAvL0+d3gxWXMcdmlWaTzXnsK1l+KiG+b3TApE8A3
Guet/pT7Artmbc6QPTk7D0wp5oH/Vatf3mtBKiueX+fhfdGFo7yyW4Zm0+DqgrGe
kc4etDU6X+12+ImGpWgti7x9fJgdU2UZQTSAGks55P2Y1/VMeJSeH2ayctejUjiD
ZUGAWbRPQmo1JvDFfDYslyAoHAbrjCN4R1FGkQMVF9OHkUi8lEKA0GWgKWDVWBcl
JjKAiM8zgy8+lj8IoqI4Y6puUQKbhLImKU/kzF0xKKzewQH0C8c2vHwqTnwRroDN
pFb4ShapJ15n1eoxLhMQ07/iHOCONUNUaN6bQAUr11jhGwyrJvZV4RmI1SOpNNq9
pzzwgxuMSArmPksallXmj30Y0zYGsItVucIXQgnfPX0vCtwJhLzwV46nEsi+Qu9E
DsktpuUYkGXKTf4IB33b39xJro4o7eoE8y8BgyJTYSMArGwvW9uS7rEEqMapiQe9
e4jVRzYoZ19gr5bNJVy0f2c0wZhS2kdactLhB4tmgD1veflzZSzjMXaVTDy8nwdl
aEmwjt8hjAnOX1Z7i1W/wal23euHI/7zm38OdzuwyP+iDb6wDR8H3Y47NsM8M6vl
T8xrj9E0NAvB1EdwDkuQPEmL03iPH6POTr76x7Hrr6kzwiI8nWSXeVYm9K8ILwUr
6vIyNIVJB0WqoXV/fiDGM4Om5xvYSfBAJyMb9XmYlzPchd99vsogxri3pWR4pYO3
uXrn7LFqW8tAmEUV9M6/5jlLQ9lA/xQIL9VGJvQfR+GBzgLDH4iYS4SUjPSEBH7h
MmGgz4rhgV6fJgkTgwWEp7A6eWYxNVhppY15muYeqUahzVJm87lxQ63CjXUrQDt1
0+74LYLBhE/pBQCIGDT2zaCjVs+Y5fSeaImcHTOUx9oS9hwrR/H7JW6UmpEk3p2w
q7fAoMxFF495+cuufIsze0OfWVv7w9EJZgTBaOe6vPvDxldrJJhPgvlPwFcbQaPe
6+tS0z9ACLQPye7TRpoU1a+iE7CMabE+d9ySdCQenftJZm0ekzCgVrjnQbXQXZQw
O2YCnqQ9NJgcYkPYO18LUZAArHd1LSGgybOBBDOQUkVPi39+iY/Fr+4C24af9eyZ
U+CcdOf326k8NFOODGeg/b9LQfzpjkkSDXCffFGGiOZ5n8eZaZoVqowlXZsYwES4
5HHcCOUXBKQ+4bf9+rpZXEcYOPN0F+4NUpt3S85GLtgCAbylGv1aCVY4me3gtX8n
agqbMkq7jDFK3tIdcKBLCgBVAJjNpO0rkfgI5y4t+z+GWBu7aEBJ5dM2bApKmHYm
ERqCRAXn4ysAfgZM5W2RHbWfVFXuBtpR2/bwNkiuzdGxi7vBN1BIUYWP43TkU9tb
TlhHKiNiOCjXPna28O0d0KLva8Hybhcb/GAZJ98Tm4JwypPOroXB8fUxBTVyqywZ
cIFry29IkQxJ1Hz1FIKecRfwYUAXixspHbFeGuP3H6J75W6/5PJ8LDQBjEys8XrI
02nj/CXDSmbh+9da8+z9bjrnICQFYE/n3TtdbeEHPwzYb0EY+lsNI8dM4ZCjf7zV
O1yxFJ/T01NFtVZA0kN+QgA4N1a+vapPbW5zdtjmRuJk+DlUC+MP0xgfMgISjNgD
6lrSQFGLAB8qCjSGiwZlnBNlx6tnPRTrxMyHo/VO+cP2a/IgDKnrXUlfOahbX5rZ
S7B3grGt0OxnjlUGTDNEQxhDUc3cz+bJgpjx6hQhSKpZyoZspHFJG33mVlDuWRbS
h7+7ZpUJyOGCqkFWcrEAIwg8LyEW0VlNxUyDc/hLPfoyvAsM4EddHQ02ZNdR9yxp
2chPfQysbPiGL3mKzwp910yRBmy1FibljKP2z/HCrujXbkLJaeMgE2xzqWWyjfno
MSG25RApuduzKBM/bb51mp3FYKSXLTtWBFkyFSKqcu/e91etnuaRg/B647gHz/v3
5Ja5z0O4tGOYiGeThdXjwGfzushVLCtowiDfhi5kGtXYWEJZFoRM1pcQ33udwtoh
VcVabXy1YhvNLEXUuDmGIyYa3rOGdWIs9nqn+V7ff3zAyNRykESE4a9Rc3gaagx3
RgxqHQbIvgbAE1xwoMqXaj6YrTvX9w8rdC/kZVwzNESpzUjFO0Tk/rIMvxOX/afK
xXM/GOJPjRPsaqIWMAU17NaHRyqulzBKvQrRiJrc9CxXuEXB3cZn+Y1cf6l7C4W4
pv4X4b1FgxZVD0yyppc5V86qGQCDAb9VwW6kKDB8426mSQN2f3CrHIXDR7W8/L80
GFOMPMg9N+ZbRvJ96i2ar+b+/JSetuJIZbq1TH9oFkEQo11PE2EPhcrh9GQqU25R
6wYevi5Fwz2RafvPuyEZuHf0GBU8rzG3lor4xVjqjUVOWC9xpuvbB2UAHu/+kAsZ
nx4KiqNUPzGkJh4Eekmaa2DhY7ONNRTuvJjjgyoWnC7WnCMveA2N+pnod7mVeMdY
OFmwUqQuu8aSOUzbWop228WQj/YarCBuz5v6vCEQXHujRpc3nSNdrkeneFNdsON/
+IP8tHGq7YXMUj9DbGPpYR1KOBEYN/xr/IcOIOS1nGJbsz1HjEclMBnVSXyKDfBj
gEE5SbXP8IuWrHO2EknutAaRA+ZQeL4ESGII8DIvCuCtYTDLawxni8lzM1R6+djU
Uz4uF6Sl58IvI7l8SGRzwWY3xA8Hgx2PPidRyVBil4zvr1G6J7i2MfaWa7YyjT1y
jDb026UsmSXIyevSpGQrvnDaEnIrogXgNg/5ouppGoAJvjzcPpcAau+17AjYoGFn
bD9MtlMpKdVqQGB4yQX/KpLvDQT+RqNS3EZEGUKaajzhxBTb9RSizx2MRBDtrfN2
nfLBSsEzIjudHcmGJXd3IDPgbYxBp8BuJACISuDCLwcNeb7xi1ZnW7QmT3zFRjNZ
xbTfcE3NRrF6eKxfDA7Os86wW0CTLWQ5pvZBiL0GzGkHoWW+8nOw7riI6kqmlJRg
3/PF2X+YJpnMYFw/JUXmIovWFR5r7puwU0UmOusY67dEmLJx5cWX8Ce9GV7zxbd+
kfBCp9UX8IdgxrWLaA58w4WknIGgUDpMlYFHS/InwVAUJ2UHcbu81T7cqTGBpjpR
iUuVw2AUmKuuvhmFYgyyMrvyaiLfcgJY5BRWgRYH1DWc52AavN0OQnTydLJKKAe+
h4M7noyadetcmVmbywdovYNzX3HCsVNipXW8jiRlLj9NauoHigXDiIC6lqgZJIhR
eZq6rfd8x9H5RM3omOS8BL7yTFZDkvJBAdC73jfR1id4srb+gdwamW3336YFnB08
ityjQ00GLE6diqcgmeZHGkIv28r6Lr7SzAOwL7wEoEeH7EVxYoUi8kvi+kYsiLRL
sxgW+hei4F7DnF0fKVylRv1V0V4YGqqkLZHx5Rhn5WXhYsIIxAMmba3KvvetYKKE
Itta78cdQN47cVGMOChBYQWZgb19g2+N78ck2wlOjIy/s/1Y9tml0v0jBrhVS5jY
kcfsGyjur41b43UJuoIu3UEXLEJMPppNvaxQYd6RgsZcL/eEQ7yDcXmgV+nwqg84
pg5n2qM2OQdHyRxDqwuRaTKordl3X5HQW1RHANFEW+etEScH5mn7/77Wt/0FHF6a
a5XnJgVaaRHuNWgfFYfgnXg5LWdesCslS8aZ7f8DK1cVyNHAscaKGnt30fg6ng0O
lQqeBjpMgu8uWX4P9632/y8c52ZxIm77VhF+ZPfTB+oII0CDPfH5GKBpW3vMM5bM
2jKLHkoHuyROStmG+/1rBkRw/PFPg6G1UBlyMe8vxyDGFLz64zF+hWvFRoYrzLNw
rmTehGjX8unOvBAsyS4B7C3ZRwL238/HSkIvsHJpj83tVFRoiTptvL00VKFUktgp
GdjcDF4YXdnLz6qQgi2hSRpCT/H6doeB8Q7QKC7z3Vf3te4oDnJLfk53DHLz8A2V
pwCUelzYubb4IR4jE4602KEa4umD1ReK4tScpsXPEQ29ZCClP+VO29Cb/D7Lb9zs
cjStTWZDnmKAKZjkz9VBBbogc4Co9XxJNRtdygrc572AB0pgB4YF0vqJkUAvo99Z
bbWMTlnor9M6/qSyw0vgGtckre4BJrXez/GbcPLW9qZDz0+Z0QrNqw0VS+BVPZzz
JhR8yZ13tk9o8kQrM5qSliktwFI5smYrE90ZK84YfT5294QrIzSLlJP/plPEi+Ca
TDC+cEVFFZSUzsx+OmIKnHNEIv4GmhDYLtb650iZkBzdZ5Nh2aes9+BQ5LWCD1A9
5V46C/Ovs5u3eCXxwUBNzpnDXGfCHwaaeQcDI9RVmCxbynWtFW6nFdzHgYx8W7T9
BxzKkWe9z9Dh7A+7FapR60c7TsJLvC4ZQRsUGguUd6abO3Orrk25thww4RXzWLUU
BpXJuU3azNGi0j8oOlfXC9bIY+3/6J/XmZHDNh/A8ej0Ndu7480OTH9bZeLCS6KE
PsRxkSrYqVnh6kscKokQWrs2Leh2PWXjLyCiJf7ULUuUiKp9G29RAl+5Gc9i1BKR
zEuvvhmxruwECg7h52lQxtxJkJDK+f3Tx3Fj4wpFdjUEOvYYkQaos0eyzudrRtCQ
nPeu7qxRnqtaDjb+WuVztgQLgcHPNvhIrldD2kDUHJv25rZtzAUgqEdkr7BBZfe9
Ud9EEp+qY4uOqOMdzBITzZi8y9ZfFvzO3Os6cRCarUnMBw8IohaQR69h8TGyz9Cc
KSo2IrNodWccyHSmy9ax6258f3gAcXoxWs5nCbEREPW89DrlUMbfB+Ypc+PF9aoV
Nj6o1NsDXRA94ibbg3Eev3SWwTMYXp+v30UIDWbqFXbdVDMTsuCos2MbKSp6Hj9D
ReimoxSO7nt/GeFClCE61yIB6RA72/LXeVCo1e6RosRsMIO30B0QSwp8DZ15BhsV
NkevzixrQU3DTofaqgpi3pS/n6MfJaaGDKBtsR81BPM8y8vLeVHc5wy1UcOlDVY3
USTZLkCBZ3tsJBKgUBRnrSV3RgDgsQry5eHz4iVUldMIRAbL/8IzW3faf1TsC/BJ
3X4AGqfGB6Gv3VkTnNcTaC/iBeMhS/ZC9ryIx7uQKpRLEkOfzXLqKASmBiiNlCCi
5CHajnSZYZZE+//Zb4JSvO6tzZgn5hCfX2Z5tPOnZVkjTc9KZyEb+vkMMZKMcX80
a/2NBxEZARF2pUCQr+wncf8pjfIOwX1OjabWSfRssiGbvanpWaUIyAULvCfv7031
XUFjyIJZWfHuNST1cGRqz0f1M+guVmhnIoYV+31qZtgbLiEDliT5hBNgcU7QGE1f
vYgspB1nA+sWpQaV0B2Y40LhpUl4OC5qFQTgeoQUiLeokBGjrKkcPKUcX2Wj16hh
re2E7u+jdwQtdQlDbXgn6qw4zNZGlXofKyLJs/U2ffDcKYwryS35vzfqqPhK+GST
R4xS9X8cDE1ojetY6P0McHFLdomYnUVgL87uetqCUXwqpY5cXP6Sq61lQkFepvFj
z6x7P41QlbOoFGNV5idV5HO3R5h140bL/1N0kj2ks8EvOpzgiMs/4ouR0ySi7Xp+
3L/ZWqYcs995b8elMR7RUmt9x2CmBm0ADn+53WLZg6ZTrVWKegnlYudcMdVcB4kv
8ezE3WKW1VHvGsSIU6qtlxV+KcF4xAkd9VGc0nAz5k8SE0TetMte3fA8kVfKhjP4
nFB9ghdopcfJkYxShLFllQNY6SPufSHFUx3tu1qBQb04Uf9W4efsjh91csWzUGSM
g88FVQ7IBwTheOIJ+WVDt0hTLt+eQKrHnDa66By+WWo7zrsxfUnZLG+AP1UHhdvJ
oRxpXrwSEh350ayu9dwyHuP+P5Hugyhxy0Zf6eRbSX1On3PNC3m4hw8UAxBfewXh
G+IZEhwgp+8O+O+x6N4bDG/xPu0RrY2xEZANZ3NVf2JQWsycjjUBUH6vMpenNGp+
40efQ+px3NX9Z6vfzd0PfurrckqPMtAa8TkbBPsxiE5PcLlQd2XqPXYkxYXXBJFH
9pkguKg7xLwxXP3kyflSTLrk4gw8jX0RsZDAxI7OlEQYzMsDB4Tb5WChWEnzFP61
GNAhzwnXJthNBvITo06vIN27dJsxsj9uFnubLUbzqbwNwA2vcotcOdDKjQ1+Zk97
W8I7WxiTTY7lUtiLL1Tc2VX+qLWw1mG2elOL6cR3faN7V6nBqwB08for3adY78t/
k/zsq4wJ3Hhm9BSYE2G3IhRE87AZwbbSrGlN/tHRNEGZTpfWhZsiEd1z6tcFiFPZ
bcOOwD6cwCB5xkNWg2Lc20xJx45wNFP/cjzZwPgMtZwks4WaGa7FC/O8RIcq27oV
fQIPH3NKNa4O7CXAxYrdJmusoxsW7q+zqBtzroAM4aMuE6RLkp3poQQGDogUmAUv
3CukuOfYcsMDck7Dyh70jzsf63ukFUTyo4NR39WPqmVOtF67M/hKn+t2y4Up+j09
FysnHXfi0tlbrO41R2Dmus+Fo203GShS3bMuh/WlyBsC+6RZeNgaMbKMvQCtLLIM
dwcAfS4j3ZkSveJ0otszzm8+MXz+XW5XAtbQq1/Fs5bfN4JjqG/ToA/3UnxCE31E
lmqaZ1TCB5xdycDe5Z7oU/wD7FAmJDeoWgeB+xwJvFd2W6F2SrUGCEIHELOAMeZC
IK5uWif/El+GbdcWcTvzNmgg2uqrZGxLVSfcHHbtJkhyhRZ89YbXrfm6umRUm5G5
r8uTcxNBfLeoeYzJcJ7Sk7nOXJtDK6C2E8JKH7KcdRYcw5pqfh7VwV8jEaYOQy+d
5//BYAzXtU+yCQ8dnc0kYkl/jVoy0btAwUdoYdyVCKna0dP4fOdflISUpLT0CPPP
uKCziiHpBm3dBriUTLS0BfLakaYTSjRkOhTXv2FV2vi1+fKIlbMMAYVJ1rLpxHzJ
zAv/pUprz4yNg7xER1TBNHiZvUoTRRW4ZoKq5Ko2h4XtO2ldp9I7VCPLUWZ9+KOE
riTDEhl3UsMS+I8NCPJWooXdebgKyjRW+50HuaSwhwS2TE4Dta5laqbrTQ/Ji+Tt
WoRf8mlD/m2wdYMjyfghiGbHu0LpLGOJAEJ+finsks4aCzAXTQlZOKSuvEhgnccS
riIvfoVySWL6y1UjI5kWg3TNQegWxxbOKs/ll4TrviO2ROAq/DA8JGPFwnqIB6qY
SDhgrNP67TKkJJrXMgAN/yar/s6dKLkXXuq/hgbB1K/VDnlRHDZbZxJDF6mYRXl+
uAasgnrfYYnEXfxE/M7ymBdeMtG1140kt2yc1uiUVdG89R9EDtgPEg7bUn/M/68G
yFBM0UesjKB5IrKcy9yr0n4rO2LpSIhE0jX+o/grTruMbGvrSlXc79Myia7VvTgJ
JnHxOf3Zm0XsO2h4vvMYP6yoOwMwdQhZQsBCPvRNt0o/ldXeal4fwG45LlkOkgUX
0dgrzhdu3zZrqFynFE8eaJ/278SrGShBulp3dOnsZOP9H3X9acYEtaB4YnOVFR+W
3Qd0j36oc01eAFRRvSKHQqt67nhiYS60ozh6MbmwC9zspRzQak2NvF5W/adTgBIg
gZTqWpyUFkmM4tnsWXXXLRr4Ge0v/qAkCtvYSSKK+WUlzzPNsAXJ2zotVbx6/LU+
AeDTzYFSBT2YMx4QXSF0NGvyPguMF4p9bnbUPYEQUMU8sud28T8IqadLw46AqUDx
E2j2XrTzX3fB0ZYGLa9BXfzD8kpOSW1r0J9y2kpQJ7rLqve1kaChZSd6rnpnvIC+
tu9/ZIAfxHbT1+8cyJFIeB4RNkBeiq21v6i/Ivcbv0+zDC2wZ/8B+mcLL+SJEQkW
8NAxrBsT04+sae3XxkierzIAFfZfXQRMiEJd0qGz57Sh6/rr9ALEqiKHvHuiPKS4
2O97hgV684clTCQpWhhiPfmRSeVKDJHUD1qgBr6o0hyUF9K36HYT3DcqZUnH4vLB
moopaJhg1qGZZlo4gP7QtB3nqS/pwqXSbAFoBx4E7NGe/JaHzbXv+zTmgla9su47
S5FR9S8ByakNsKDHyEkK7hkmOchPONPg+qS40zZutTlcfxCru6FH3zh4GUyH8VHx
S2gga0mqHuvJx79EFZS6mk63dVRFBhVx40iGAFu6x3c7OzkgC+UOGiaOE3rHoM5U
tCCP0M9zuqtnFR3jFzx7r6sVRfRtiRp03FDJvHbyxYoGLwAeEs4dkS4Bb4idSKx0
VuwXhJ+LJeKj6WxfXvggJ6q499r4JT+EbiHA/fzw6BR3qVWbjA7PuU9Hhs/tTQMm
2oljjXoKh9bh9cbrO8JiTpZMIl8aREzidF2p2SmmFJqPQaSE8Q3a303NeqY4kthR
sOuzUYehG+eWeyB3LGbOidYolFm8maoQqqyQixz5kMJuI0TxoK2L1tiSUKu1c8tx
bninuPRtZCjky+fqbsXcYUyf5Et18Fr4rNuVl+WcT+6hIfNcXvyI/8FsnsUsSSqv
zEGtxmTwb22FvRFjTpTyO9PkRYZDClZWeK2v0SSQKS/oA4cz+IUdx3A05lzgCHZB
jjS56z45EHWHavlQKWnWzAQxMDiQO/GGDt8gKBB4El28fGtiyVj8CvUJCyOcLNlo
wFOGynQn62tgx6Mi8fd8sv31V9PgJNkAhwgWRDkZ6Xub4bQ+7VgnzMw48YO9hDoO
OEFv6lhPtVSF6GVUvT4Pq0ldQXJSl790eZuMtJw+X785m9kaxgzZU7cyEZx40Afz
Eu6PzOh9iGTA3um8vNY4FXJnrGLCUMZEAnvoTHNvnHNXf+m4vvwZfiJNxsg46w7S
18EbaLBoJmBK5SpEraF7kcwmoZ8Nf2DaqsvAH+L6zYD7CPR2CFR3UqyZWrbFyFOK
ePjt1MiyyotFEbUpRuLM+JHmgc2GXaGiqlRFbAdpMmlXGncyZm6HUKXyV5c/dYXu
0nkLB8rhBPXW/2n0u4BkElt8QDnH2+XNtiyzmaD7BzCAr+WsrhlEtQMk/s9Ux7ka
TSGbL3y0dxakwOt1pRQcsK87Izg9o1DLoVzSIaDopq4bm9VmWm1lByXwjVoWtWVH
nJfUcwlU5Wy12sUFUYtgbQO6fM0MdmYomVD1/cQ/vnKovdOZy9GP/+h7Oy1t+EBu
2nWywy50niJOAYPErIzC3BZN1n468bWv7wMvGo8LrJEbA2r2KOINsj+4LkRn5R4I
ElhWu9xxe5vJxBjkHGHCWJsFSLNC2bZbXDGxWoiBojuaSwohf1PjpCq9M1L9UQnI
B85A2GJcIVSTf3c33TBQwTX45eVv8SIhhQQFsNwme/KusthPA594dA5xhlKFvRI4
VXPn83JftFAh4WaSe5yAMAm3sPUGuTpzXFv9/fkdOjV+iWVc+A/SlstRAzmhNUQM
aTAX0EgRmUUcavFAOSJobxt+D8tEjDcgF3osbwhUTEE4RugJUK4BqF3XCEvQkQw6
HUlQZoIF+l1jtDDTTW4swPvtk3LxShiOXPkLavWFcVO8ur4eyQx2DBEXG6a6G3t+
GpGgyIIDgejJugF+cpKYxNmO6/0DSCBJ5Qc2uQhbVb3VRroF2saJTM3F2pSHDWOd
geglVstzLwbDIxie7rLS9EZq9uQKRhN8MnzFyiyM17PWLWFkwyRYo6rQaJTchsn5
QEJZv8WfqNYtgV3hZKco/Wt/HWoo8VQSNbPoZyZbo/IFjZZaPDnozpA0reFJswVV
AHWs7VZsqVzpEW9WSmarNn8y+y8c17qIpVZhjT/HsHb1dQ36nPgsMJv7Ns7W0xS8
eMECwpkEFN40/9BtRm/LCVyIM284ORzCNqgWGR/s2vrbicUauoVxx5MC7zYgmuun
XzOWp0fEQUyVk02HCIJhRNnZ3jS2s1gjsG4OtQ0e4ywSlObnYjWxj5hGUB/N238s
JkpxMT122QAyiKPEiwQ+qIIwf6/wDc8nu+BX/TRvirh8dGsRg1lDbUx3HqK7k7tn
8C8PFkTavn4NnjrP2cXmuXSLYawwEwLDDP5HC3uqxgsOyWbX5dvUl8qOoz4nKShZ
IuWDfZSebJiBTPbhjPeveYZjWfYyn8yNg2kh+B5BRj2oEPXY3xoyZbT4LDGmL+su
4kurjNCJEDgoEZC8s/L6Y2OsRg3r9wh4kTodsp7E4rcdoN/agDHhE3Gbb+5g9Bym
/ercctCABJg3mjZDF6xg4rjgCmgxZgZyN7LSdTPyMqIDrg4oh6grD8XzETYXTkit
sP8gJ3WfEYizPN9gOgKELI5ntOVNe/LR3KSMSP8q2RMU9szEzpP/6zTr7pEckmd1
qvm2lE7OvytaNpgjFkkX7Nn0/Ih2aUeKUxZT9I/ewC7oBmHxtl10J5ih+Fr4oawW
A64/YypzyWxn6o91WScu4IvelA3onuulgXFGLbWya4lDo8T8tQa5GQY8l1F9jSPQ
TFDbHXZrqQRWXcHfM/2hHEeZpZmdZksWtplL1Vd1XRzAzGS/j2p5sfMhqDLdJ0rh
uAmPQN7+2iN+63JTb7Rmrn+J8TRLrEW1DtY85Hbk1Qtl++XMpO28Re3PbSNkKpPf
YLYSPKr2aYYkqunmktMlsXThEQmK+PJv9QldOn5WLhaqh9lzLipOxDRUKBuujQPB
8ZF/Mxzjx/IlkaIuP/F+v1CO5ESHgz0SF7W0EwX3/WvCdB6n9qrcJ+CMZ5yfubXj
gfurUPQR9XEI0qBjO3OqE30rZ2ydg3jHqNVrGGyjfXc1t3Yg/Z/mMxDyh7nslqGO
B+7xUuQgyyt17jVAZ3MfsQpHGQYE8IIrOepkg6WJFhHE3UCcC67Dfz35IHWAj6pm
n3O+nkPhATStyRT5q0QAHd6ElrO8RAVjXhWIuHMDfoywDE21YeBQhlhGxRIuvZip
XLIxqFrsY0Img0ubbfa6VDD8c5fyJ8BnVrrtzGl5snCvsjieq6jVQ9QfVG9iezgj
Zt1D3XzqJOJO697StZmLUfE4O/lRqUZLm/m9si8hu29Jk0xjxNYBDmYTZWy/jGIC
vBMQ9n+vbxgLz9UkPge06IPaRpEcYCMWLwAtflErLEryGShrtoDp6ez5E8gSPSwv
csnk+BfjLh6qbAgF0vjc6bhcVI6X+AwFPTqe74P5yfTTcm1zE05V18U8eiI5aXpZ
rTsUTqlLVMASZVTgZRpiYUnzfQSDyXX7xMq6l145rnCH8nzlyvaUsaEcslh22jcH
NJHfjYSWbdQ2oqLeubwBCnXELRrzExuU/TruRV//MzCOfzwt7QCXtiWNwI9Kaqzx
mWzJiYSm08+33qYlyALKmISzeBSU8E1ZGR48jNOnOir1q+neR9wWvj9VQMIoewDf
fab293gN2tzu/uT+ufRalrRRs4ON9XJnvx0CrbOs4YbMy4YMSbPN5vDh4W6pqm3q
NI8FYA0SLtH+5/TH7pUIvT3EXtujfaEGtkBTzOusuSdOSzRVBPtEJjdxRJfkrwMw
OJ9f1Me+8brU/HqZrWKNikNHLE1iyl40ZsfiJahX5uS7FQwbDKGfSUzA3aten2nN
Zi6ur20dng7jrgNwFIkkt2RFr7COivyOuqb/4hzyVNV5IIOJdcvkXqj9OfTjRbWC
jq43VijU5hkp98zomTf20jUcaiFmXjCectuPn/S+xINLxO+DHfpfWXLSu6yaov2l
nV+FO5o9GevOjVEkjvYO1vTbCwGL0krMYjhdja7SgJqsXIQ8coLkoaM4XpyE2aNM
Va1ImSa/hpF7jg7kxR+W5aURD+M42FYVns4ZS540JNM+h0Xci6dk1Y+A0MAVoSpU
2J+Xw4wjyDPIhC5goBwN6rIhkltOM49Uqe7FsPLW2dZveDwfMTJVO92fCuGPf4pK
qqEgNitwVhmnS73MUQ3WdNSfXv97Wk/xIdr+Im3FQyyghVFHR3GVcf5I42s3bw6d
+DHbI0Y3pNBRBMlTjDYeO5FAqT6tG7Th6MT9BF+42w+wKmQYkY6qBL7gxm2jLscY
zUWM6dojpRtqHwrut5D2ttQ1acs/h141qEfA/s9CEWsne/pBWSPRMt1Vt+iwyn68
CDdSYD3AKHVIVcFC0ed/1zRogqWCKLGQXJIIqXhSrXCIxLXwuK44M1flsFpBFQK+
RkaGJvf55B86ywce/w4o+8CHAsowxFO7pzN2g+TxFFiPB+M7gOTI3ixDOopBd5NP
o5kPZhGbd7UD4hzBMjnXEK1ihZMCLkytOMkxb6rR75s2Oh5myj2Y2Zh5hHjPYRwV
VftqObdrKtKABT6y70PbC1trN4gHAu8PgdxvGzy16AOUPpGVSoaEXkKgdBrWQH4v
/febIKv+aCRzEE5fEL04sJNngCjbALFYBeuZOwFbKkFzq0fKP1RDIV7Ql2dmsE9g
eClVlJBMUj/Z52YwUr9hmJvtjqKWWFwJzsNpHCvrhJDPUlnsIV0K0dH+aXUzR7XC
rejgcmGCl0xl6U1Op/JWxSHW2SGulGCfvgeREJp9P5ku1aI6D3jBACxwg+qhOPRA
5WzpwbxzHGBd4KWd+HZlFBOGpf+tsjhRj3ujdivdhmqiHD2g8Yq/viSad5fVOIr9
xePNR6Zb8lbx/fST3/47N3o+Fj6gaBcWAGQtfb4oe+v3JoTKNFLbziKha65sA+OG
ipVJ0Mfb2Xp7u4yEtPI2eXArjY4hT1eAhleG5ht3l9wsnja4EeeYUnCmh1BMx3bD
IKz1WFZOXHb2ur4vSUPRrQQ80Tv/H4BsW94NW6h/H+X/BdeSIicpdJXvfIcW8uqR
8tirIFW5jYPbf3YUUh29eU9LI96kqSOOWR6wCsxAJUchY+vScARt/R3u112yfxoX
Am80H7X9406QOT/xBu6qUgo8vSZqzVScOOUcdEtcqzLzU1e28O3lWTRPnyX72XLN
MpKU9yMBfKQOCkG+/zBl+aboCnU/s1DAh/W28Iv/BwB3ND6qbWRzHzFHhasHGsHX
B7cpR2s4PHvJIUn6bmt+tN/4bsTMIX/S0eK49fxFMlO1c3oWXcRyzJU9quUezeI/
VWz5KzT2jG+t3VW/k1APXztkj1DzHq7bHv7V00fBwOFim3/6ou5Z/lMtrwSAidT6
MLeJWH5NKG1Z4RUFWpy8ci2MBD6Y8juhoBtpOPWioS4r2ppdUpwGcqy81r4sgMVN
l4gT1J6ff+XabXStXzyV2VIlkzhMEh/GhWDJQNeIWXrcYuDx8G1H9pUJpY/c+386
AXVa1w7U8ZyUPYMAdWSNnGB+nLScqDtJBNG+rKEZJP8QODAa70R6O+aPaMTFAy+W
aZSLEu2io3yo8nx6XAJP8BLfv/ZhfWLhhJPT/OkUrANX1/dcDo4W5DhG8YLx4yOc
41rTkz5abLfQrta6nk9PcMODXr4fI2CAce2KeUVME3ouVwkzr+zjz81YAWbF8fou
WiDpGnNzIBy/2JdOXh3B6jfhGLnBhXPEZ+dAWhevTsxaiqYx3ZCnJBsGSl6rPh7c
JcKbPJfV3knXxhUbhdq88GDQRivDnRoICF84dehgUWE6NklxlbQTdfaReIIxzHy0
7b0n2HrTI1YbRVMV3M/VsyF9j4Jwnf96umeRJNXd5PNj0DT33IGu52wz7y6VA2MY
4JZw/iI4D+q9hP+8/XEF07WaAdwUaPiT5880U6GnxVeiJ4cic0IVAhSdX77n0jpv
7ldUqE7y+IfmsFP0Yiu/reFTtnMy39cM5r7g8a2lnDrqb8nQeUYP7UAK0mq3iwkb
gH/HcrAR5iltTMXFl5WeAep3NcKnhy8JXpRogC1LzjnA8CWZuqiawH4d138qHXsX
DyPXup/DuInRHZfYNcrvyY1Gns9wDPI9YDrvgZ2b9YZ9ipeGHLBj60ullL3pBpWK
Q1gzJfhJrTWLQIL0SEokaAkd3dYR9TCVN/A3YhZSGY7ppIuMREJFqQTJTxYyUU0X
kOXruY+kZMNEhhcyw8zKRTU3nP8FUD2bXzvOL5k64R2BQvtDeRo9djv/GtDJF3+t
9AyZXa6867oGqpubVMLlhmn5vwtFt04U+K2Oxbxb/Q9MXGDBX7wmR8t0uZVznYLe
RWIsqblJYU5x8LbJjizl3mGofeztwZ4aKp4lUnFjzKRpFflLfnpylX5IyzawF5a0
bTmpzyi4lmhFKcwFa0hmKJLipjSqwMJs/cC4sE8nnbfjWslX9NJE33fjfxjuFxon
t0Yq2PX00L5wRZ2VCsYgy9PkR50OPKmmpenPMSHv0ZF06e3IfwarrZrBZXWufBm5
lg1CqoyJC/1SnSgYsblXGwMLdAAxWFmK6Pj/Cj2Y3YahP9C/3wEvSHvudxhWv+OA
a2azvV6ziGGA7saxdbOy/JlKNaETRb0ESb32PIrWzeHT01tyNc8byn/30/nEKWcu
yOxJuCUh109kTyv0Aq6NkRXeKlfSwzLU5Mnottu5XINzUxvkSgU9TsLBaqsx0JHi
E+HYc7fpIYCU/Pgf+cy4J9Q23beIt26IOtqvXC/o688bCM/H4Fn7j0GARc+Rss3X
sJTyAt/fNnL+puqOHJ8DFC+u0rpBRAbmHVV1m6ynq2XNR/i3fh6ojsb/jymP0xGZ
DZh+wgGnHXExkWaFwvfTE9gg46FgYZJDLnD5YrGPVSJe0/RSPawF3KRYZVxMdwFX
tAA8RsY4BVhfI07ppiJeblZVg0mlvztZdJmmqOJp+VuHF+f284fTIOrQgZbaTIQs
cCh8YXBkldVgHu41caeOSx1wAsJ4sR8u5h3MVpiCnzuY1A7LBXAl6vYYcEMcCmrk
tp6f5oi/0u7/fYVl+faoFul8NoZDVrFRIEbr6orwTLgcRvCSwJnZrswZgqyuvm36
Y2X2rejKnP/Lo1QTlYuFGptcFB9bAVQwwv8hYIaOgylR3h/wAAg0+ID6IiBN1WV0
6NLeewOQOdwWGkMDMeLOPk7e8BTUmwvwMlHf8uFuGrcDHWredGQxZw0jc2fakYxJ
jy2Fe0pxvseZQpqdvPUg8xcuQPl9yTYc39QRI+eYE5+sikHpaAJVdJm+hPs2jXsy
5OMKY2qUlk9f0u83bfMSYtRcszbUuRj5Oav8fLxQ/KyG2JN9KhzH/MjcCI5vlkMg
IkCbKiib40rPLkf9P8ZApodDukS7zgNVG9hdQCTmPVho76zNM31qIRAcuVgSRTOa
jPWAk/vibBgO4vwlzZkuopA1/FLVkDt452Ik0yW251moZMcUikG7I94ziSN1BmOE
n+Si1xpHdgzApl+fHIptXwVLkVZnG55FU9iNI8kO5J3H16iz/kROpOxQnSU8r5YF
oLBtoy6C5FsbtcbpDGUO3qk6UokHTRai2BHHKNl2NodxgHCi/57WW2VoAk1kq4tw
zLCO/IP0x2/kdhefybXOSROIkb4u4HBLrlhGVanokX+Coj9K750R7Nn6E5OE1MVN
SHFiTQ8IUjNGLGQKmVjAb8ZdXAv+7iOrLX84J92mvwRVt7wrXt8U4vwkWC44xSz5
b5WjbAWkfYm1Grb36XmJoJ8q2uqgTaJ5cImK7vR2vSooHFo0aA4i3RC2e+Y26/Yg
3aVcjsrv5lOIiA1EHJSHpFxtV4h+BS7D3hbM1tTpMQFpmptabLriKkdiQszUfekA
vX9zR86cT3dxUqWfBHMJUpq/ytq34EvrP00T24GRFwSva2k5iqiAfrlCvw20iWJD
DIq5kKNYjxkgk837xbqPVkQj+NCV8Ht5xHY73ka7GQcEAXv80OZF6TvUrdwYEayM
OSBkQluNXBTlfw1+uROTxo2p0qLlOgpVKqMBGAUhKIfLzWDnkOsi8Ge+N/a/pKGw
dsmTPrZBvagG+6CzQ/wmZ1jfwduLsSZTN7919VesS4Yr/x6bW5xOeLTDZAuXmuag
H1cWzAlxPCty8dNR7phM3p4ngu4yEoef/Z4XDWsFdKeYXvIqmi5JmTR0NXc4OOYc
O5nkGaOl9RIa42h3zPQtg1iTDe+55LzAEs3pIpd/o6JZ6Ru2nBrVVyzv6t0AwWVn
gZr6KRtR7cDDjUYIu6lizVbeeyo+fswRPzMpQoxf8V86rXI8TgtyiznRK1FeCfNl
wIs2jNIQkonkUYpx4zuuURrHxK+pmfzQeB+4sD6GaBEZ3yUABKSOlkor8ZwjopHQ
VlfRs/yVyOth9K0vJhw1v+O3QeHUFaJ8bptwlfff+jzllNFb1D8HwJU+Jy2PsXhB
uaPgrlIPxg/kLmqwB/pqA6qDUFie82k95sTnzurbs8nle3WBk+iOrvxEJek7xBLi
ntpwBUU/nM0v/+YAMUY7IJR6ojsQulRpFhbGlugX48FVvKg/xCXfcr961VMk3hyB
Mq/Vwjiaslf9oU72fqO5/iFBVLKDw3Xu5iPSFiml92Zdn1y6+SV6rqbQesHTdL3/
jxybUZf1ItAyCYY9miiaoxTgKsytYWTiCqs+9FJEknCQCTk7Wx0xdNo0eHOwZaJo
xxBJxGwspAwiXa3Roa6vU/1Ax1SDs6OhzP1w+hhgVhxTIjNbG7JrMQnRhqljfYQm
1T+z12KhukcsK3QdWkBI+sGnroctf0W9EDdtTjai4VA4fiDKBRGhzwWC2r1dMTBr
l5sah6uHYNEufs5yxqx2zAIuNZV6LQS4WF7Tq60w6QiYw6ZDIf9adi+4wHNwoHyc
aDATU7GSTuitIxSrUK0yoAxbaoaDuE1kJK1iLjOPG2pusfrrbxrsZm2zWoBbTwoU
9PkrDVQ+bnCqr6ZFOm2EekMx/qKPGhODKs+3Ai7C1iOJ2pGGkySv8CjPrNt6rqRF
NqIr9exMlLSVrSib3s+Rbn5MoowHiJMQsO/FkK2k7gjhXmsyIg1w2PBFWwaSqeMa
h+QF6gLoGwJrEQoSr09/4jMXy7Qyj+taG3OUx96c6oqonuDW+EdXiaGLcSCcm6Lc
qcWJGYSnFjiCPaRGFppOgVKdKG1FsOgTHWoLXd4/8uopnQOZQ8ToxnKFQncD3B95
9QTcZJQpLaFtL5JRS2WnDkdYdflY1x1k+k/948MqVUz7z6YwgkxQD/gQi+AGENJ7
T7Vghgq9Umf4GuQK4ZY/Y6clcKfaakHYPtVR5j4dyBOWRWloJRAoY273/qOUkzCY
KJqcxGBUB57lWNNlbFumK7K5m6rsV1wcAxr9os0uW9X3k66uaX3F3l9Z7lYBkPEB
Pc3x95NCxqm5b9xCNczuE7ioBUqxgipMqOEMJtdKCX3NyNNqV32drcEcsMA5/jRk
JjbttFEM51ge7BAlLyYFK2rxUMLS/TlbxsLmRZwGOMP0ZhVQZQmyFLIn//VElJMA
JwLbxO3N33xIE9ejalTIKzcA64I+Bm6tc2qPlwWdgk14XrN677OB63G2pjE3ra3O
cKLgPgzAXb1hTS3qzeY5xH5DxIRSyTkkXpzKQ5yH8kXSemvbOtK0uWk3/j5cOpEZ
9805iraVhtS6CwW2mESVEECwpkvThwEMDDuFHwj6aC8eUrPTHfRm7GIzzpyjzI3x
RBBlbhJokUfCoTW4SafKa+VY+/SU8ziVxve4XdIV0sqbm0R4AH/8EtEWdqLyIBCx
zm0GX2EGX5hikCtiyBVTU5+xlSRSsKL3F8UIJTh9ldaG1wFJWQemO1YRWIuC9lc1
zeFcqnxTA9BbB6s/zmPbc6f1TBkkR0mvqOTiJxa8SQciJnyyJXY8DkF+7pp/OnBg
BmwlFDazkVWwv2KfFI7jTp5e+ROVpG0oFzGpdy/ion5VTyhfcI8oyQc3rkOat3o8
ZyW79tT8RIgKpxTnV5MSxHya3mi/0JWVbwOcseHGz+JEy37Z2DqJloEudkQNyw4M
F7TMtWAhA4bPr8Ht+ssIBgI/gQTkevndvnqPRGQLiBaJJl0JLsQL3L3Z3lMNIQj1
dg15P5/Y73E3uoGTk9+5dnbdl2mSvPtqYHwlzgS4KEcoqWzSBMnk5AIt/4wdjlEi
GY7cFoGIgC1gX5vh37mr9QkKFJucKqj070O6Tx91jO60JDpVeW9Cy+GNthOghZY/
e8d/8f8a0/h4xI6PBq5+eBsDNRG9wX0Is4nJyOyOT8as+bctJ8j79T+bh5GvNaNA
ZoPUj4gPJMdMfwj9HsTF1v64GCXIwN63f2QVk4Do8waRGDhp21uoB11MWt8ojMe3
9thMyzP9vKnTASrMW5KdN/1FEFE/KX9WJk0FUsx1MgvgrUDAa1zUa/pGisDC2FPd
vo1qw4g2EXUI6ZHJUXFGFilVx83GwgtfnCvAFqfNTXbD4j8W0UdfJCa5s8PH4uCb
uQoS3VYgPht3kpQPO9y4HvuRyIOfqcNR3BQa5pY2EHeMH7T5b5GBOx45JJg3LKTb
/psWjykyY0OjFuUh/pC2wRvKPGxqwpTY/pEUvrCo8omR4Rk5RCjf6jFSuuADuF/d
0JmTM5XFdmXLwejighTSBuHv9ERmtZud/60JiRG22d1MtVsoWXY4nV3jQJUMIx/X
9x4mTWmfHGFLtQKGXwlcf4Ysv5eRSadIwLQvoCxW9IDrtbS2thpRQXtyqOX1ZDZ0
rdB7uJUAduouxhxw3aSZEE6hQQwvHNTmTGjnf5mIndl/FUThc5IE3fTHw1tMEcXf
zx2aaPKG/qeANhe94G/TWKM7siMJgW2IiA52EO54klRY7hKi0pY6bsAFuXG4YzT0
Pxt/PwQtItNUroBvjksVbK4QM3DqYTNvCBaDoa1KhkGjzc4lEjkb2HOjJr1qiM7O
GNYyL0vHxgLI8HdkvlUG4fA5Rw4rIeVYRCDHP7ifgf9wXFf3BODrUg7vbeOyPKr9
0tQwMaCFUVhnbrjktAslFqeuwub6TC9kK3Rkyp3EhUr8ANEZDu643EJ2cA+3Wz2j
PRqaAfcLjMvbZW8bI5qQsx/+qnJqMFVRx1h1h63saWpI5ouDj9EcL3+dbg+bWO5/
jdiOitUi1jR5vgxNRLkwr98sfmrnHBAlR4QFjU25vwzmiWC3hZzQ3dQlyu8iK4UG
u85cIkDbnXOelXjeMEz2Cw0CRto7KWslOEdW2ZV/cH2r/cu6fdGON6aLfND7zOM6
5FcTxgLczCpRNoL6g0s1BwiAc473/7ax0ysT4th0Q/I/S0aI1WNO3Tnti6MT1yD7
LIVIZucbaEYrdwczFFK/gQDyuqef+mvXvrVkCOo9ctLJ/0uU6l8StZTFNYNbpKOL
X4SwiKHOBj9ugsjxbPvadITdekasSjhGXlqONbcCvE0j8OLsPRU+ZTBeR+fUBmkX
cFQzhqOvv5N3UebtZcPOifuPBhJjTyCT9uOhbpdLGlB+b3j3/g8encj9GfHU+7oc
9bF5IKdcXppyqNN+g1XQaFYSBDm+zSD51FSGzjQ8qW9GOemRlBeyYbZiqcwZ80ex
CFRlUYNt9IOA1FP4N+lCWirbSUPVB1DCaX9zDQYlXZT2yfTuvK1F+bsp1oem1VHy
c9LXsAr0VJ9LZZF30FmclVpeNte+aU6vvl4YyhMdPUyRYD0BB5LX3c/9O0j5xqoo
IPr/M+AqH7lOBAqPAPmEIZXnTC6Kkrdo2nOPfMXZaSHAnlYxCca7txIvvS2q8MCK
8yjTHoqen6FN+qmx3jdREYrbi+RPfPhoAUuULmBsh+tgZmbP8yiV/ukZE56T/H7Y
pUBl211mB+BwTb6MXK8COb/juyfSyGZfD0mPR8c+KfHvCnIGRmOpjDbKQ0toyaRc
YXH7JwZ/95k5xChm2k1E5yaur1zXAdi21Lb2nJdyE0OPpgQYvYotX14viBnOrs8y
45ip+Rjoikc4HnyE68af7E1B7hbBPnk6JAyga6KNVgKkTZLqKvDDWzFUpBrgxCOR
s9pu95Rt654ojFp9TmkQuUzyUk2+AQ14wyq6a4RWNqphIfTJCMr8iiXDct/ELUi4
lgIA8BvPNefaAQAo4aYRXGIkpWrpYay/yRBst6ZFxDhqkclRt4pucDpL2Ot8WUPw
HRsuVnzykyJ8ZpoOd2ahjdYFPKHHmkrbK0QvkhobwcF6djcYidmRhN+40UtbnZDu
iHx+v2lbfOa4/lbYZOXnyDhHtrQcBycQWgs/1pJ/KLu5yYHYk28lkVL2OBATCqhl
44DIIVQoLxc2aWDrEH4WpZ8BTdzUTRlGdu8N4u621F2IpMR5e7ZBX0ByqAzbGxu6
Y6bAntCT34F1+hb30dQKZ4Z9Bg0yNrO9MR8lKtjm5TfQcYCsCrLjSniSUtoewFAo
w/StrHdk9rgLbEIwvIiYzy2odLmFiGFHL7ljsgSskq9adecRavffYNpNz2CVBq83
2fxf6U07+a+BngmNimSNtZWtxA+KiGMbQURKL6XDSGQs7jWHVdrRfQ7qdLR3zZ1J
tIExlipGPrMnsJFLjqrO+vB3CtV0nxIQNQu06jEtKzpSVR80xWMPAJLdWjGoVibG
EzOEqEqA3uiSok5tq63TvaZWZ/MjVa3/vXnym32G6q/k2oj9Jw2MATJMEhXzJk4V
m5NY+tK6tsy1oYxJetgWtwLnKxRRB70B9B1K2tME3T6g1WcDFLnfXwuP1BeNmx8/
ynpE8flJbBrXQXKLYj99YwMNtZQ0XpQCWa2GdVscJsHYX+IWdUnJU26Vo3xxkaei
KHQHzRRUef54SdyrLQUdJ6/OUXGTmL71QB6GhOqJleT3Kb8qjUOkHKDxy5+2Dw00
ztC87K3Gsm5ThY1mIGXXk1J8izLq/wq1/eNgNEgWhK2uIvzvnP5hHn6U/cUUThqk
0zHIL3v8VK1GctlFRsE52PQ6k/G6o0IVAu+m99dgsMzHtmLTN6KwHVbnIz3DHkI4
ljQsCtNL1QKj28O8Og54qeXQMdg1Z/Iq15YLZ/Q2xb6XVw3EjFP8qpD6+pxbiMhe
O+1EYEqqspKaR9aqoDntOpKOIEaUJ5ubX7mMTYYQqSjq0HDT5OaYc0nw3dt7+3s7
3r7rp+R/QkxTmrL2DUj6OAkezmVfZsKlL7TgjNBs+nacNYZOswdEDqPEI+IWGJyp
k2C0yUmMB2VAtpQE4HM0+j1a8Msviv+7brc/U6gmeGOC1If6VtamQXvI5gOeV5qH
DLrhvTRa3hKCj3TUpz2YZ+Ew1oSVzK7aWI7munuuq/3IgQgAwJPtGjBtTXJYx246
Va4WvaulA/9FOsShhGzK5n0r0M5rJ1bH0YyG2ISy/DEA2oN4LARtNUiajXp5tS1+
qRxzaSZhawR1SiCorUl/f3H1z52S0mJaQLFlKbNK7gpNgXhQrnAZABg4dl68FQkJ
x2NvhlwNuyQdkhXlk3jjW8wPCcLM3r/yPSlwc5+X+doJ0Mh74PxA1RVAhrphossX
HBxhBPfQGy6uS22iOieUEkx7owFgVN94ogDJg2WQZvK/WT5A86GdAGSY07puKPR0
bAcqCb+WlrYbvnorSigEBR+b0q3/8YgvywmfaGLCjFAxiiZOq31Et7wcEt9yypID
JCKdq7dnylST3jC/yQFFPPk9lnt3xbG4FowalfhmYdTL9s1giW8rQTBoWy5t45r3
hh6ZN+o9zBYk6PRhHE6yDFaKCfcPBMgSCRlUtzPsoeJArWze6f5d8s8ikrSWRI8E
uNGMGEbqR+GkqCeKDXhWsfH08b1ZrA8LZEPv4QlA7HLONYheCZ41QUiLI+Fzrho0
BmQfv2mhTWrjXhwmxyfwwhkTnSzT8TiF/jOjrhXQMJ46OLRb4pELCXaDbKMokt72
v2VsI2zaFVjudQLxzLSJGzHRqtTZZI9u+I4ZmeSdv3QNMLxLhSAjHlpMTIXADj6p
8IsVxw4lI6q/5iS1jZJ9/ZJtlEuwY6svaCVuu9JylD9w2l7LcYHnEaDVTP+iYIVS
mx/hg3NlutEUG36bS+KIFsM+F+5NeGoQbf4MmSRsHJwaGEuzTNzL1u/njhT/p7HE
jxu4gOHp7dXV9UJu/660MKvzQ55wPYxTOQSZiYBn/nrNn9otqxb3JRsw5pZtzgIL
vnZCMzwQf0zUbmmimx+U709C0V+j+t365aTCFUeVBVlyk+7BLJiKi+DvvPQmAwdR
/npr2qeYCjr0eEMgrwT01E/AlDpKt8WL/m3f5unfsIvBCroJAUyx210fEwqgEFIF
rpGOXBNN2qWBgVElAs4KsyJp6vnMVQ1E/g1WF1srr6xoW2hYsg/bzbVBZe3bCMMo
5HtmzMQkKv0I82BMbp1v6aRDcRpX/VBhR00EHZpMnkdrqUjW90f50U13CzXUCCLn
TxEuHjHAmEzxvwopt5D80EQiTJXsJ6lBc/CauxS10MktVZ3FFYpuPoneV5WxZeRC
F4GevVNiAYNO/xLcKsbk87Xd8Z442AARu3+VfY3IER3iEXhTjIeur4zY+e6Z30XA
6YmR0hJ57k6p2XkK1YpqltzSSVnmMwaNAo90sFS5Zov9eqZk/0mVm6UYD7bFkAG/
Jtvl2Jma4h993sbjN/9y8GydOAda094DOgt/OOWBdQ5QfJtWb0WS8klKmer8gEWt
Dtjk4wzVR3MfvJh19EK/tahXWHQedF8dYck/tRKBzLIiAQuMfl9J7I1fr8aj3M+N
sxCh3+UgpK2Bbuax0YIxpLJsRW5wqfeVjh5pN7Uh/cQd/M3uBAobxkHz4DD6Kvio
15wFH2mgrUCYwcrILQNRJJhmA8CgIOpy7gDo8de7Lrry8JbF/NmnvX3CRi08cFny
6WsAzL/RVIixxCWRdtOOxmdpJA5405mfkFht5laZdOG7njsKwunhrt4n8F6IYfmz
LrnIbw60PVXgw+xuXVdDP+GB36scTyTmLOE5RWxs7gMLc/2S6Wh88lQnDMRCCNDt
RWK1p8RjKFL+q3igCBaRAEIFS9UkvHe82rn6rg8vLKGp9ZGn/8s8JNkLWCRwvp/u
OctOj0lJdxlxOrRdKpEnl4n6OFlXilpZEJUbiJQEorTM7awR0X37wKCwolUQu4El
cftZm50vArzhRLCPHfeCPtqfy4J/36ZLcKz7wj7pR1SM8kaBgUEAzL5VstbIdanp
QgcUsI5nNfxwH1MlTYl21tQR/OqKyLyMj1FeNWXNIN0U3/9OPPB8HRQSo3DAjWiG
wtysaSejYxiVUvKVtpT1/hqJYFwlh1TA5dT+xrI3H9vJlv+STFwPCtbMc4AW6sWZ
a6uBx1ztzL1kB2yADub82znXLe02KnWNPZGkA1XQxWdT5BfMiWR7PATu5sSpFlVs
aXd9L3oQkeP1pPXCf9DwpbrKBLLZbG48wGwUdNM4hCJvzJiEeMl3T7d2e8Jfpz1h
7YsSu6lF8bPAnVJjMEv6uHe2mVCQD280wG5bikt33iSPCG43IACfLx6ZPLQQ8lN1
6UEQx6m58m7YoeocKDHhpnPoPlgKz3xW1rQhKMRLNaV75QbDWrSb4kNnzzeJjTZJ
QwAWbWRheFusqtsRduP/BA1Ke20TSc6T0LloJT2k7okMNYMaUEymg431gudIbjTe
1xHYfP5QLkLLevwIw6HgLGel7OA+PnAeXc6LdMRu7rbmYhTlnZkNRyiDlV7mWMPY
vHEGs1rL8S2wHyxtuekpiWo2MGaF54TQZGKN/f77J5MNx1FM9Px0KbfBxefPx6lK
KqNOinr5lS08CalPV1r99OCW+xp0lAULRJLlWqOhijkqdWVmOKNwxuavNWno6uDZ
ITERbUIBIC5ug7fs3wyXWL/Onmc69IQk9oJ7kWLiGdo+V8udVWXSgzHzzZ33D7vO
gLNakX756XTbzn2TZzAg1FcXd16zNG+/U37S95rEJnkNkElNYh/DFtfTVt02dWlQ
VgBzILSU28wtYJJNIn2xzpdp/3vmZ2SGgWpUgL3kpO8UrjIeRlSFnqoPA6Jy2uqj
FmFWLR1urTFZXtBTeleXn05KBeKHTq5ui+cIS3IeDDLdh63IcDTb90449z4sXPO1
mVFgyOIMih8B/AcQsPTA8r3+3ulO4oMC/1BmmQ6BB76IpVa1G6d2/0tlw9rXr6S7
SZNbl7AzPsaDThmUqIC98vjSaPxc9KqSLzIxxjQu6dFOifeHcjWnz37luvUamkfr
5ieY/pG/5C4r7BsObYejXvGTPm/9g3s+4qav+L8muTBDC8GslU+8kv4e/xS4sZx1
Ff1OG1hH+ZvHQ5uStkEKjLYrOyQYXfTr5byeu1/1FlR045yLuVa6lZ4tH123HACM
CfHATTNnkkNugpReyCVqdbhNfbrW23ySkWFn9b9j4TrS4pv4GGhBDEedR8DxYgjg
BJ4Es06sjye84Xkumi5Q9BaqldjovrDE4Tb/5OcwsQ5KTw3ogNn7Yrd9NGlOc2Nk
FxI6+3W6Yhmm1VAYUmVzD5ys5sPGS2oQtXKJx4RO+abXkuPWhwu0TpotJd+TENbl
jf9SsN/cwFtzIyti8L+8s3L+4kUCTq0ZGXLC1Vmauhi22XevMyXb2a26on8QiSGf
JrgszKzRUN+4nXrgGAgBpKNmneLoWkx7EA8k8FY1JF80Vhz6mTwaiijjImdHkAW6
h1TbXYcK1S8SEIPV8htfR3ysBg4GKRwjc6bDER8ABJPd0JhC+z9N58uPGhmvA3nq
tzu8K62KszYT6PAUOUM8hufiUOUV++FQC1mw2VGSvzvqT0zf+X5xJktwl9wkaFw4
4IYd5a3NFexvvbjPROYKodePSvz8hZzEl9fjhemzXepMXpTfQ5msgxznBvshTQuz
8nU4FSDgGdegtGOd+LiJF8bOJ/6l97DseTx7k5MuArHm6ANivh0UN0gWIHmGFadD
c1VSVS1BbJK4an6reU3am2JIv8v2RCp5l8mP+X1cvgaU16JQk5z6iiua5adjsl0L
7869CqtjT1qbqK6t/vn5OEfTI+R2FKWudi0J4CVJsMQsOooawNgm2Otvx+6qzhtz
G1C0N6iP/CEMPCrPRyqCeJgjda5a7RDpLVb4ApWKz70g2u7LN0WisyN6x3fmZwn3
iRvqO8WK12gxL39bf1AUBjUuOj99SjPMg/tIcO4CrcyrJC5pahIYY5m1hTyDtscp
aCZ5p2W0vjuL9moSugfWi4JIK66FRf6uK1dO8N3EcoDy93jOrimMT8cOx4LJr5cU
UzpoBrSN8kc7J6ZgEdD+QaOgi63nWXTNYEN1zqQnqqD1hQfy5aazJkQ3HD/pPOW6
2rlAeXwThOBlXwUlUzjQCi7kY68OtVDnIX3MXOLwv0F+CkMS/Exvn8jR15g03U9Z
gvkdPRIYQK4c9/x6TR2oVrnzJKPOk3z0wrf4fVyccvTYqKSHhiYpaq4bKlaYSHCz
nqsOwxvhMD6t85aQpKJizm4+NCB4H+RzeQmcLC4Gm0sP0GIPVO0jrEGqOtaA+R8L
dmwyfnHNtiBw43dgEgRv90y9Hy6S7yy4MUGYvgYaIhER5tGfv7nNViwf9fmLUoKF
ePA7r6W40TM+hqNmgn6P7B0zYtKxZsgJd6xKFW9mT2f4AfVZf+MlwFKOVDy+rfra
rMML6BrPthwU49cmi1HfIeNCvce9s5tLSqmxAgMm0Svd8JICpN+L7HzY+bOu3bt1
8DeRtD97Kb9zxeRZEFLdwXcKeQZivLrcy13oBmSNjhdg2wUSk/UyPDKTX8pfAsus
Ac7GJS4+6iBjlSyZ9S6UZJm+c+Myf1gBrr0G2dYY4DuGg52/yV3/hyE/QtJ5Uxmg
TLQC04bHSlVnss8t2qMF+HiSACL6+v/E2PevFv07pqf9QqJlpd3gR0ycOHKvDAO7
Sx3xM+fJQP3cMJcR2OxS0CnG05yf4K+2Ns2qJiHzbVnW13vdbCrCTiHkVX3dEAWQ
WzNAcw8U8RLK/X2jHyM72+0mj8uB9b1u6XqiROWQ4YMVtkFp2p9vfeQlUQ5rbwup
mUMZMdcpqZI1pDuDflv1tlHBghKbeTjVHx1pWcCiCg3z77SXCDp04vN3wQ3yG31y
begEFZ2IuMBfK6xcxspyZwWMn0DCX+hPIQwK2HPiT9yyqzYup0jsAJYc86MPG6Ef
CX5ADSgpqutjAU24u45Vrk8S9H7m0mmKxuLMtAXK+FrQjTSb6BbYGwk9CErL6afX
MvzT6cEB1LJ5dpwaYKy3Di2FdUSzVhPFWNE4IW2QJ31DIqE+05NZpmz6FYCQ0j5s
MtZ0pigOZ2eQr3xGpVB3D7mrmE1h/8d+irQU4tApEbx+nxYLs6+8SeIsirZgP8ql
pCLQ1vkBpcaBU56XVfzezmkNDD62WlNp1kdiFwvx1kvDxn6KYuqhiS7k2TAM6p+x
HBJpshduOU+lxrXcZHpjD3jzhZuiR3uMDOV8MORLd4SAFpGwKFqR+xXr4cFNKmuO
fSgOz0gxXyVNQT9oPlVFhBGfH5mdqb+6mflfnPTJnZ6lP/vStIe8VFdmM2/EXSJm
mApT2PQWSND/rx0tkwUfEZprLaAuCcefnLw/r+2O2y+zWc2afiTuhT/LZMdO6ImI
FZy9qe7uuDcmYJxd5UU3VUGHA+nrhZ7NYr8gGOO8ohH1RNByJjYrIquTpk2Rtuwe
Sd2liwOrtsIO9VTz8kYzKrgOEnZ0XzXU4xDXUkn/D+edLYNsf37OCfEg/NPkjCyf
zMihtPbu0n1ZjrnO1o1CP3kU43tqLKlAcdssCxXmG/+RMuykqU93/ER8O4w9Q4tm
yla3EhpGcVhefGPQlEjw1Wih/7CUgA/xevjgSSrRCpCMGcYNSPIpCheZnX5tJhYc
4TZ33FwAMe0XbgJ1bTh4KcAy6cyyTLBlaBrw9dWHQJK2qYeSApCupbrc5gek9VjN
gLGx0QbZHin472baY3pEfQml/xqhpWiXfALxENi27k4qXXEcVJPMYemXPzXz1qpX
dzdwVU0QFwa4ZMaoBnA4j/HriuFjYPuMvsZuCw28QsrW3lahhVj24h3rsO4vELgf
qVtf8nHRVHX6FPsH2TCBvR2j6eWotAVBt+dxEso4K9G84BBk3eLxGv2+86u2ZP55
spu5MQZtKUQRbWyMrsY+R/+3O6XRDikMxtoIeIN9QdP1UuCamuPB8VB0ePwLolV0
nPigJNtxatqKnx8tQsczDbHqBCMrd5kXhHSKv3/H0G2ANG5HrVVCVIBdGapk4/DX
2u6J2sLQO0Cnm+YktatWGyAReKGnDVxfrHk+YGe3KsaSjF7XTKWndmDSLrhdSCei
ZOlRGdNfrvBrnvi79ngbWSgP9JaYPlQRH8mwNIdsSz4qq4N6hZDwQxTR+OCeSR6i
T7DLjTD9yO1eNmgSazrLQvfmwPLTg5ZkkHu5KXYznoXDBhMyomzfJj9x2ZN1hDaY
cSAKyF4B2RL1gN9/5vL8BgyykI/9R8w26y82ytaf8ChGRw4Jau1mWMlu8CjEYmlU
mEPZR/atY4kUIz11+cPntlE0VDhYZgc7Rf6nkZrFJ7Lgw6webBB4BTcdYzWtMCiA
MjoBGx+/vfX+C/PEmLDnexng6PLEnbIlTu0RzavTDX9DwweV2u82r8VnfhQBaEJN
y2dR3AGS7A/8I5ZskBUgSOptAmXGTgM2K9HEjRVTtSMfeow+HXWhd0ZHjwMfQrCu
HykI2+je1iE4P5cA4GwCAsBAghnyvJorYQkGAAaIF6QkBkDiiTCG0mOnrNOuxzef
1+ceVTavbwMnPD4TblvRVHAFkN4y0+rBtJSil5ULeNZ36Cfte5HcyGmwm5Qedb00
h0mydA24bzp/e/Qz6Hnnx5yBH1P1gQ2s69qbq8cHUfQim2MzgFQOF+2rpQlBS0EN
e+VlegBoCBTK5XSxNbphbrRNPxNHQBAVVWAerLa8voMQLBzNQyZRFRqRudzIpljT
d7qk8YxSZleGwMJatytZcxOXHrMyr+RWcL4xY3NcNXwPE2lk7yIMV1//S6Q0RPVG
7gulSJ4kj3na1GVL6R86nA0T2TXNMpTZTEW/MeEKcCt0V1hZZdqls4x9YJU8l0KU
9kY1yYN8J6Qs5+QtzWbhq64FX02Riv+eoJ4M56PoGKLtZf17lTzDFRR8PMBFJRbE
c5suvNOvv5DxbEvsmd6bVDhZSd9RB8P9A6+HZxFAGe8Bv+d+8zTctKO3+qO+3VeS
UCAJt2B+vE5I4ybXBy+iqEm76bSPX4u0F0Oq9QcwGeeoK0bVJENlp4gPTcuZEv0D
foa3ztmEgT6tEgbtidzYTtZZm2KrmNP0wBK64F6a+7JHUtBeOoXKGWHjCtXcJ6T7
b9SyT658k0ry9Ya7L+SSSez2RwtfFCOQ+ZHVIWSxld0WnAiVCBgCsx4LDxTY+Kp/
E3adnj1HbaJICDQp1r1VwxIe8JBg443ystjO/013VXsu1M2WBX/29Z3CqJv21iYY
BfsJ1ip6ni4rtuvkJoOdu+sLD0iY1+JxQL0+LfpeF1ptx81FQfjmH4OKWfjwf3pS
+nFL9kltOd4aUzm9vLP6JbhJNQ9RFtr5+F2pTbkJQ7iWN1EOASG38QOJ5TWnbb/i
hW4eqXU2B52OgOPkeBO9MYt4SxKb6kyPrmy6uradfjwQN46iu5VZl/UtC8P5DgJz
xHzaM5e4tG6S1TwJ+xNFH3bRhmIwkZlUtiRU8a13oSLvVOLSaUdc4vNQArj4SNRT
6NhDFiGbtNdUicAMLguX/vRyoW906xp3hIPsLtSnwvJ6Gn9ys+GZtne7fymQDMGy
RJw4doOORO2ank228M8q2j/6GX5tl1qHCblN08+ikVVQvY5L33IkxG0B4f/dFFOM
VCkSIdY+l5dHAqhYrA7Jo5Ut1orvZKk7RPPEsEyWenRCdc1Wvrwixz925tSU3FHs
mNpjm+I2iychlZADTHL+5dAgyRAO8S5ctqR71A23Aq6AnAU6eDbhtZRzhcMr+Y0J
AsC8EupsXp6O5X3qEnlZo/i9fVxfEOdE2izLrV5+lANTrE/uSWXWX2o1BSK0J3Fm
SNkCx22YAZROUOAo3bX8QKtNqQIIq0wRAqiFw4EaQY9r6PFIdpsMT95S7JS5oFsb
WhS0a+9h4YG+z6a4zwkMNIp352TPdfoArPUT3/KM2yqONvOVOHLG8pOrgFMCRRkg
m9k8OOoOFcWynsgnYkOcGcireomAV6sOLjEz7AbUFY3uxQYnZ+4hlbP3ntt3Ejwa
ViNWu28nrEDtwI6yHCvdDmdAYaEDKk8VK43m0xpPb16OVWw5qoLdSinPhRTA2zP6
SDaTLZAKmJ7EFKM57dw+yqvZ7/w+WrF0hh+34U4cZzla3BKZpl6pH2z69j6iD+Bo
KRHqqT8vdGXTUqPvaKUWc7m4oMDebXvKeKhaH2NmnoHRhhkOyyWmvkfxUsJ87tmH
3m9pG2Q22dxTYR1Zc5V+hbmoDluTcEpBh9o4Ngb6cDjONfAgpa8yFs3rVukDn9vS
4qOQ0aEeqGDeeQ6q06ViLSpQuwtO/cORo1oe0WzFcxgD1xP03viUQ61WB+HmuuhK
dVEJCApsiD0lzMRAbhFUfurzWR0+V8qRZk6xnNALSrNpfjabZs0TfXjbvfcnI9ge
ZQKME3r/4pDLfbjS6pPcy3Dpk0oly/KOWGawNsVGTAZwYTBMqeL/HClC80+e6dmg
UcOAZmvaK/jwXQLdkyVfByPiAbgstwJVUpPu1rKUEzQWnPM80+2ZVH2gaMW+Lnp1
WrVtRf6yHLP4veb/9Bp3d4FLhfcq5wF4QdrWYSepXJwl+DdRqihdaIY/Fk6A2C+j
SzymEqFo0nXj3hZjDWsl2YMTKdcu7h24W/CGM/hsKve4MzONR9P9pZsw2eLUv4ik
QfJY/Jkej+gyx5BdRgElzVFUJVpROyBrVCfnc1Zwa+w1yq4zJyg7gBcAm0nHNr2K
9GeuTOUeJ+b0S6gI7R84SYJxJ3I1+I7qkhUTXox9jGLCnwil8CExVAIHGLEuo+W7
pgncsrNmvNyNkGkL+fFZgEJTpxqKlqk0c0gIGaB3Ez8jWI9rPRhKHoqQEP13lVLV
rZWwfgj6jp7T8GZljSlV/RwPRAZ3iW7F0F9Wv/tbDSaDv/srOmPAM3ooiwXYxGZw
s/eTre4BosU50BaxK3a5b5IPokpOHOixB8aQYTDWCL4xyHc9bDjI3WJ/G1O818yv
UYKVLwz2ekTgZfiaL5KeGqBWZnEVE50WpTt/MT4u5ZF/QFFmnHtH1tHjTJYh5t2n
ow0NFMOAtLGlCy+5/zwQ8EsCoc5ZI3dd4f4imfIKcn5c6nvqed9egwK+LMvWAQt6
bEGn0sJPyzCwvixZJdwHWtjkRuHZI+AELolJogFpvqdSNkYYoDr6tlWG4elcWWr3
gSl9c+6zPR+W1Y6deqHkZwpDNYiWYzHC0ixggS1jTg/EYCOAxOX7u0tJrRe+KB+W
7hIwsU2zuFs/PgrxVG5uhrOr28FS9qI/hUB+fi+ylRZ/EtkS+7V2bUugWgNr2gFk
T5r1dRex1MCI+SCFegdTwHQ+16qlE3CuSthRKQKQI4GQPjtnpydwPlLC8piT9H/N
ucfFrFquMur5OqlbphSv1t+Rw6lXSugDSkws7eUc5xtAPw7T8LhgGpJuzR7fBu5H
3JACATqQ8xN1UVt+P0Gyi680sZs1mQa7XFWprrZgS1otzQgdkEdOR+PuhtGsc0H4
RfInj9ivxfPwcH/pIpjbMWhd05SEbuWFnWQmVnsrH12a/T8Bb7eMvLKUPBD/n/Gt
imOsxFW0oRvy0v1IxAL2MmELS1ZVIUdKOq3n4QqzV9J1yxfQWf8XY+RUhBZCV6tz
3hJpysGXDlCxpstdebEDQMRQn4Wgz/x3aNr3TVuy10lOqwBiDHjueoEdtVlabyyO
X0NWnTo2T555crbj2dyYPLbYmSCYMJhX7XK6ejQt5BemK7D65oiDmCuiD7LvlDvG
yaaeA9I89o9hOL68XV67BKxTE6SyaF8VJ6In925eoIGMDlQVBZ91ln96bCaIXXyq
qmRgKW6w4IvI5Tjnv3tYodJ1Y8+Nu4dRK3fj1vzEyiHadUSkrSQfEPpQrm+YffUS
c7G76SpQX4uGilnInmPVJJIwG0PcrJkv7o85g05q3IW6R+9pw7bT33tNxGiLQkUm
ry+pEqaHinxYEP76qOO3FhHzd+AddDZ73oRjjVw23UCTeryQsj31TOPcKv51bjXQ
3yh1FugotgDQTKw09PPmKaaicipQ7axU/pYEFy3ZMmA27EbiXXqkfNS8pbWAkt3N
SqHUwww7/PL1bEdsFt6U5JOi6NfcJtDa4qmPgpJVjqulG2+8mUmPxyuCE5RJIZp3
cikafjX8AbWIh3g58BB5vQNiLzx8M5Sp/dISCAn3Y8993VEWmXNgUYtNVE9s1Iwz
3BKBQp44I+VTkm0M82YVqIrt/gLjgnQqwOJe0PqXAJ8hckstbEKeACnZW22eKipY
FNYsLrSA/fk8e7ndDzUH7oK9g84M+Efuc1nPurWlGpHQ5H9xnnC4Cg92leQy3Jcz
zhlnj3alC86bKetpwLzZDjDay5CaprMn1fY5k9zCnTMuJfo71m3QRiHgy+t5zfmf
q1u6jyfZfo3h7mbyYerQFPLjOzTeLWDRhejcyXO4GXakW6JTizX+tfREKY8s4Ek+
a/bG0ipHCgJ6YE1yFJTzv3ISSFNFdlKhq82z/BxM3dp+GSzYvbhijdMGs5snd0pT
XhD3+q1T4cqv5+v73e3t2jwvhOQt+mXpKCHx1z1kcwGwjQYRDmgy/OO/ih3lMwZw
woQizBocWC7FjtDcGSUV3kIhDN/rTDEQPjki+g5EGi/M5yUY/q4wphbic+BEvFV2
h2JGNBWW5hgKCoIINm3ql60cxM9FloFY4aT0yLCObXet2Asst/v0lbT8f0u9FeNp
WXmmPwf7/JIiPLMXpiQ5+9tUAPda/1AQHvYshVMcmsGWmx6l/cVLsuBv1t6dUplV
8hhoA2SMVWekstVLBukMeKkG05gBlEEAUKIkuDX37VeFhbv+oX1B4lR91kQTAtva
sZh6Q1d64Z3CPMBhPn998UdsL2Nk3tuEt5uw+OkMo2Lkty5RjPnpf0gs9g1JSzka
d6Jjyvx4dElgWlv3m/vp/mS5qYV9T86U5k0Bd5fHjvDJvEekUOzyy6AqkjTVjDco
mWXZUlpTrhYddyAqlt8goJPwLC03aEUfUXBQEaL9ptlcI6fHTCnJWCunDWqdVYtD
zqx/VxzuguPXL0651wc5y+SeOFyGahxRbOWABTdXJfN0gidiOv0FbY/8hWXsJcr/
tTLegcUj5HzKrSZt71WHv/jU8XGALcf3QApCUMQxIthyJn3CPMxt+MiUP6JsXqtN
KHwRnBh1BSbDVZSk8G870ql4hdk4lJb2XVyruDp9g7LrhYMRnvV5APXCNp4+qhzm
xHfiBzA0Iozeqflofq+Yn94kd3iUBqtoq0xdhi7/4EifGhLkZiVIrYXJi6CWNZCo
zEkGUrEYQpeiHwJtJ+7hBSgzOiaW0B2K+BvtXIit2yrWLdRQYhVEq0dIEKjm6iSl
KwBAhKkXW7GliF0gjsqWT9f2co0w4kp2q2UgAShwB2X2WaB/Hakihmu/0w0UGgF0
6mJrctzXZdJIwCA+qPYDIIaATOI0Rv9nlspvKN44Q4uuBXMu9OXwiscv/giDd1OJ
H80Zy+8Sg0Dj5wDgDPU3y9xwjVZVXjq7FxAHMMI/x2bJXLkOBYrCAgN1PhMFZHz0
f9lSNaAVXIrI6Th6uGFFIP8mQ6nKKI73OgZIZB1G76eTgQ1yheBAOUliFACixCiA
DVzKpXlu2gSgTF/S41L8DHaLoDtRq11L32PJcqeqFRlchTVqCtBVT2BzBFEKCtjo
xIpnlca0+UVIf38gcZIjcJ4liUKqLsy3/9M7rpWHAs+I+r0LjUxhC0sSk/qonp3Y
0x8yI9bzPvP+OmNUS4KvmVYMHUUTzQdeozRHUJHcCHQZ9bbhDGMlT8YuA8n8yV6Q
jn02uuShz0Epbuo+OqMEkkd5OQdagH7xKSL+OIN1CsSFNq5QhmMeZPxOWGgoSCY6
QSz1yRiZdaRyw7s6X1kIbHRRJvXy+MmJhClQ60FJTa1ap+12iiuij+NsvfpmjxaV
m4aljUK7DsQiwXqyRdW3/2Fg6uX1tY3x6lX4Tt+pIJGE/ZRvVLzi8bI7dhIR9a+q
TmwNqq09ah/v86ekN9i2CYJwPpRHvvHV9Cg/J0+b5zH0/OzHmBD4mtaY4qEAqbHd
f7ZnZg7CiM4fEmzNOyNaHWZY8BITdTWXcS41S0gD8vr32iEyEQktTdEnqEpraFog
lK3asYVJ9fCVEeS0bi7zvSFXDTaGktFQH7Idf6f8K494mby9AWE2dwdyPnZ1wwN9
YQekiZw/K9OsVdiNwHjjYP/X6i27B+6/GMLo3HZfw3BMeqVVCn77fR2j6SCZth+x
IfuHMucsFr1JeRQMW+ZqtQLdJjrALk0ehrfit7Eqv6dAdN8YJs3bExTaJIEXhVjr
gSItcDtgZ/mXdEF/6PfBqVxejit2Od/3L3RkUXE+rEvOv7BVF1HNGVrOCFzT2h6K
SWFxWW/TmSinlz710+X2EWBBZ6apxEYqv3qMMEDc0N0u7Z3uyOdBbbq8izjhBXjj
k8+APA6Tb+FKBG4TWC2tmQamosksHmoWKkCsKcjOQeVzjuCJDjYNTMot5VA2ziNB
OJtKY6irdeAOwgNMS+h6upw5+PV5YvI5QV872QhaEqXR0q/6o3HRik06/JiHTdiQ
fye/fCA6aYLDU5O71Fj79dmaRzGAMvTTSqQXqfHMCJmOcp37gnFhP1T1dlK4AsQi
d0J7LhrMVGFTtVLvKdpeqK1V4z8Tl94F/gtiE5fkxywaJVpLevQhxzuKzwDkm501
aN5kjuPEqnyrsZ0ZJs6iz4L3k12j8hSi8oslMnBWGEfBe9GNmXvNzOSVtotnddXg
lbBCnAvcFkKnQmBx29kOaFGdFDe9x8iEgvLXAwPRD5xNc74ThyD/roUj3nelpKL6
OdGePXsntSPf659Y5NX0g9Rd7zpFMAQ7t3DAIMATP3KbFNbaPtzsNwj4A6Q5RRyj
WTMkGYFuMIpOGKMioGi1e34l63mnDtlLp5+GYFpJSsyzcHXqAAwrflvuCyZsgsSV
pfGTSCpDwt8dm48YTYdbEEAwswFD+bkWgTKFP9O8H35YdXpErwR4/o8E+3mz6q+h
ofMFCmFxcOa24ffwhhMX709iC2H5AzIK8KFbK0jxBVYSsOZyXR5jJ6pbsNSn9NgJ
lJMsWe5eF+mTKId18SmZDmSYPftXvBOA7+j45inyGHrXHrTumk79XhJQRhmcwdkP
u2lDnDq2IP9nBLYhLNw5/NaHUzp3QhOyuGfbaFTFv47YrLK9hQ4d0vtxEZtIi8oi
l3TOav8maRV/KVmv6whAccZWvKlSp5hqujQbXtURJWSJipJCgrYhZIOoXE2VEnet
324o40vwv7e2bdvl9V2QXo9qfFvD7OtwmJrFw+9GM8yA+6XyA/K4UNhQYBSVQx/6
qh8iV4mym8I9q7mdX5SsVB+v+edg2pvitDpKZBk9fA3o3BTm92FEEraAM2LDTLzt
lUUxZ6Y0A7U23dEC5GoCYLGtS6cm6PMkHAvYnBDTaB/QLYVw63xbEsKZOpYYICPx
BvR2qcVtYPa8P/1gBSBLu9PvwaB+fJrudALLgQf/EQzVb/HC0/JUiydl5bv6lym7
LVyb5FNTsTE4lo+1fOtHLwRd5Vq/lsslEvD6VNBaSU3AUBy2K5vSzN2NvnGXNPfb
FBMM8+Jpv0uf7URERVhD/rRcKBUO/X9Gtg2VpslJSrxsYfIwrneCfETL9IT1gyIE
xFkv/BGzjueOlf+Hjq1pEfhB97yPEQMqsYeaBv5IX+kLuI0mNRbjVTrHDwG9mRrU
BRWmHcVN/JMpFfCzL6vvkOEMmBul8axO3CAfPj37hJpX/rVpagQdgwiVO48fpkV5
gm32GhrIkuY1RFvM2uT+HTihqS2ECOdRYk/WLUzPxioTH73vEJTk0vbcDN5OwqnM
CDkWRiMdBmtq6UCxCnjm8suE+Pr2fN/gm3unN9uk+waThbd5ZMhs6EptJqEHRBoE
wMFjcBWBxgvs2fs5sQZxSIpbGhfnSl92R2QKiAILOxwx75lLAw3T4VEP9gR2nPsc
TBtuIx8p3OiAEVkPHdM1lMBUXpsSQrD1dXnRl1nYlygjQ97VO9HihhVJdRjYpfTQ
XDs63kdgo8oaYIU3DA3ohM8jr88NUeDyo6EQu+yfCOVkHmQx526wuhliA81Oi23W
N+B3KdVMFy68VUWafxoJoPLqEuf+zAjkPXso/g+KhNrMzh51V5oT3q/sa7Mofpik
sgESylmhE2CsnZtDjlvlOYs6c7vYqkY0zFHx3X0wnwiLb9d45lgvM/T7yqMw69Iz
Vr2QvAoMmMsPM4mV6O+7JPZqd7fAM4r0UadBAOMVb2xv/mMR7NRQhOHTGvtOuQ+J
eelP6KB6wel6jL4qHJk7PO6KOkxCOyDpKrDk65R9VkITkvuawq2A6JN5BikNIJCi
27TOV5Z8i3TDhtoW1mFgNJQvfhezr68rBgetxNN7kbIYmNuHYq8I5ic3JyLKIWap
paOr3ab6EdukHeLENU4Lae9Yg63nXIKCug9q0oIlrCU3UODlStjZPNTMessh8hSw
gmyV20wRiDGgsh5BUs/dYlN3XqaPuhjPYlfardUdktmrJ2cJfdomDenB0iCHKyvG
u17TubCONkOnBxSo5RHyk0qmP9ovSEMR4iVygnzUaXlrNnTo+NejsqQR4DVq7XFw
RrLzd/XSYPLKsBRV6Xpc0Vf91oDYdFYjo9apDLWOq1w2OkhHhzum2hRanPo9kIvu
h5JIx8cbHhO+wHqKnj+honCtEAsrP4SExDSKs5TDcfkehkqSNoF0r/hO72/zENbA
AkQpy7eiyWbzy2yPEgNsohu4A/SOqTnKGOTBjnpk+h5eplombB+tIQ6sOijUNVtP
Se4mHZcVrwR7wymtRQJEdScEU7jP+OR26Hr9dv4CG09Llumn5p1cQOIkmk8nCD66
e4uQZ/hpjKjTRtrNcf+gKbVkhx6MWYgpnE6ZKCM5W0YzicELGZBW0Z4CMXEIKrbd
q8/2biBk5NMA5MyYJVXo62bIZlAK2FWB4DVlDhAEkAv0WuGjnEK6loduJ48k9drX
J7ZuzguJlQRrIWdozINurXEqyPqLeNu1N9fqBCm01EIYa7NwKcH9/d2FDyGoXbaj
FByJgJSx7z4ok0srXYGZO2J/j2fkfM6ZCngEBVnyZE2f3/8lnyQDTOwM2789HtBG
OljTHvrkrht207UeVpiQbWC0KxmeQ6cyDY24cqlscdZVULZ6ngPmtXSBXPOUh8BO
BC040Ua7pYVKVzk6kKr2uYUh7eYX+Cozdn34+ehrh5C78oOLzJWaaJCAnMh0nZHP
sN1b4JNpGXAvRgvcxOOyXVeqaOBxRj8G/wTIyfqD5L0uxaxP+DNr/sgzxkhIiBcz
uesynPYhByaimbBR2EpLchC9M8fqy49sdmYgDkSd1LaBm/2E3XnW+vmgGQoOpjXo
WHlnNblFNJoIVuZE4tY2BEsdpDmX586X5V2U2P85tJtSAxU1IN811AOTJUh00BGC
eX96osWsGDZc/Ae4j0AKX/llTKsnnI+c3wzbbgrljNbkRUQris/KecH/LPN5IEFL
6IcUg239Wq+9qB281XooO38bp+snymcEPK/mw2eqCg/jevpeEz8Pv5P6PASC//WT
sOzPVW/94PyEXlZhXsF5YNHRPGVcnRBsgnQRVakYrAG3atJBmm5Ms0UsVIyXIONq
eWYA+uvllJU2+go9he3z9Y1zUMWIloCwA7AYvVkQxkjq0hbHf4Qz3d10zBeCOrbu
A5plP/ght5IA1rOgekkBiL+hEFFi0tXr5wr8dT1cXTziRbk1Tlcfdqqva5W6tg/d
Lg0OouQPKGBkinuPYPwgTd3hB5NKa5hu776dUyoALToBbpyZze3mkQPVUxZbUK5B
eEyIYW4TncMcsipEAE4gHUJzZV1bQlhz0tnMvsPubvJkdNIt19wlunB0LpqGzLGP
0WFFZocyewwN9DH8CMTMCo5Spvqt3fIcdKzx0Is8Y6ToOfqhTmzux3V4jldaeoDw
TZcp4u0qTVyiICo7lJ01e+A2JhDrtzTQuxPj+EmJ0a2K6w0WbTeHMkyHFk2/yG9+
Mts8QdJQbrBfqcFLJ1MQAZ2r+e/9coY7n91c1RaSeoqdC89zo/DSIZDa25BUuXXD
hvbvkBmYk6GYJlq4ulJWyBp+3BR18cjNqtMqj5VxH9b6ihQHm4sIw7DVgZx4zxFC
nWT4lPlqqcdJMUa5RYehCqyO/FScjXV1VUJyhgVceTloMFczWfiApRxvw14mRq5/
CZr9il9gOLAAUuzZqASOZx0a3BKZNJIEk4Kct6+4Z2y1tMDLE8K81ohYXAucl6uu
A5UrXM/7KHP9nabQOeTrgKXxlhzPB6tLcNow6uunxV2KrZ3pcge2eoARe4LFgVh1
t9af8XhQtxjxK9/dUjwIgki7XBqpzZGDt/S1T2jOv5ePTDzm4UwxAvYgduSaX/Qi
0P8eSIOR4G19FrKiLC5fbBYC+so7TjASd/xEeUtSIFMMwqucTvXLQ3bGSGyc8gH8
IseK5N/u1ELbxS0mbcNvjup8Z9RtPDxN4t99/IiGoyXqwt7vMzRpulfy+ecebbZy
7v9DMCl9doJvVSFkpn98hydaCsrzVDOIoBH0XIoA6dv2Bi0tBfOqXcBlRP0v36to
Hu+gGlmSPNLCuOVgIFenxnGArGiSDYN46BzlaQnws5CoYZv3YjP/xfJXQQGhbr8M
lMqf55mE57Y58uFT4IfWGUNfWSeubrK/vA+J6RM5eRfTeQKKRTCPeSLKARorlMI+
i4XNNv2fZpWw7YQv/LzIpVH9L4n5Lw3Mkg/6H7GrmYarBJjIXkU3cH2Bu6QMe9Pd
m6gDS/KeMBQJjnByh8++5vezWbEX2xVBzSlkVHhJR/G3sJhFDKJz3TOvB+hUkRxB
2WiCGixB+Wo5mV5taRXf/dhR/c68B5dJZLcw3nqb5dUn+zq+6BOrFwoyvEncFcyB
GBvlWuawhZbVx/38SlWzrvUG858ynKlMBjmEAG9VEF+MsMLRv63RAG7+eiH3/Z7c
FB18p1m06Q6jmKHOhEENmi7axboCUHq4EYWErcZExoENkC1ql47Q9e7tGTaeqXV5
ydR2dMDTVDNF8hHhgc2GvdBXG0bg1HCQWjK1gX9LdwpaaVvNm5VoiZC2L/OrokyZ
Pa9e3I3gaqitw7+SPnBiAxytTNxvMP+Rq0QVXIqnTt94MnKcB3BjLyaETIWaf1gz
DnHwNYLoSCv1P9b7WjBt9DYbWc57UwQ2xLHYaosgDkSk7X35XNtrY0CqQXwy2BNm
naFAiHiH+6n0LcKWgHRgnnfn16oaQOzbsRFY1hzfkwhfCBU4vHsjK//OTabY4G5n
KS9MQ/JAhw+yNlJRtQD7+1hbbIeO792toTshE5oYAmFqgbFIW6jTOnffUg5QKOzJ
4WYA/XIBw7tTDaxKALe8R662iL0ozVQAtPnqOT+aCBAw3DPUDC3DYlEwY0ufzUBG
glT9BNr4yRoQ59NatTATGXMJzn+hbf+JMd8Ee5gK7xIhXk/DLc9tZ4V610Shc6L9
sIsMLWkW79sChv0hdfwdS9+0bzGAvCFA6A3UBiGJJCe9qkqSDm+puxoqaG731D9f
z2ez4t1LV207Co+ee32Cp+RbglGZe8lhKssXENvP/iOC/5gZX2lk746NxjhyHQuW
eqW/MK9lOpvu68F/WUrJa7iK8WegieIgvqEHDVc9PR5dM3VzY5dkswL4Ie4RCTEU
NZoXk/Tutr2RBV8uiBczihwSM2IOcsuYkj8j0etk+Kp+OaW/fibERqpINH2D/W3J
5bZkMsAKKcIZcgknWQ/AYYUzwN77WnrYKVHWo54L345HyMW1o9SB9nONDZK6mPB0
XBaCeYTRyAx5hcwD/HISthWrdCbeHcmObbqAvQI9IQ27D17FeZwRsWSy91lOulen
r59w78FABIWF1P6q6Gv9x1XkbrOSm/0H59GBhZ3OKKwFfgW0xuYPg/rSjIvg5/OZ
zZcXVs/DRvHM9dCGCtMVlReOAL4I7paYI0JGAJES13yXvpdrJQXKPVFRugDaEaWi
0HPB5dTb2SsCo7e2ipnQwL+/X6wSw5sttwKTMPaW735GLroQMAhm29pWErVo3mIy
fwTELZe/8egOrWqTJVfeUFElS5QBEgghaRi0dM39G5xaGbY1JIbhS3OMNmgkDaRI
qGy6yTUPZaVWPnYjPf7YxQIH28Toomr8fdASUJ+9vw4Nqgfjp7DRXIuK+Y1ELfOC
MPlv+lPdVEwU7TMt310bpU2bAln/1vsHeejPbIFmAcZ3VQiatGx0Bq7eu+ccBuHt
NuZ8QGTrBcZxOLKGwulaQI0i8vEhi0a7anQH6RRx+eI8xTF/NH1h9DpwnTFY5w9d
iEDQvfGnK/LDDKQWkq1GAYMsfHF+wq4DZnRIKwXoTQalZisu62Axga0B30pqwWjJ
9fnGFPn4daTjmmdbS7+BxEfcS889CSow7I5C78IPnruNUqBu175RKL9OlphVv4Gm
39TTWpbwraFKjBmnztB4pwbRuYvGFL81jtcjeBQP8yXW7mx4w4XjkgWlDb+xf140
ks3agvBGcNfDp+Mxe80bxZ2YY6dhmAwJIpboeuTPv/DYpavdwddrDHgXlK4dZ5+i
HxBAgo5t8OSBoPE8FcKCI5NjvTDY/AhQybD4m18++6I69D9aDBPH7H4eMl+UKCNt
6vexdRYlyIzlzj8qx7xJ1ycFkQWSY2v4/z2bad0t93l2YxbOkOqJN+5/BjANxTTv
0K9vrPE0DFANlpxTTGdBGxP+t3vppQChkeiDf+jeEiA0XtvoM9mAMcIrq6y/HaLj
CjzlqLviORtkT9HYL8vT8OJhBBsNUZFY2r2FOFlSYo0mum8RO2DMPNiGbFfUziIe
yXXSJQTb2Q2Ow/DnzDJn7QoQMFuMghOBJS1jbx8qktEVLIbqNntdjPuhxS4eElwC
/ajWAw+I40xxRoyNAUW9u33RQ5m2RT9+QmzDh+fsLFLOJ8cHc8+QOmD74m9Yj9HF
vWO+qX4itTZfOv9VfTQoU+EMnulgEVGXoURkEfobjTHK6eil025ACPwN0oFiIxEb
pljjWTU4Cj4uzdNPx7vuhEa9uIezieVWN7+w02twzBWqZ1in1DI+1Ux2spNFtWRi
1dZoooMJ71X93/MRC5az5w9P+W3a1Zwax7BFJTFsnTlGyHXOBu+YtSYOkcRlDobD
36QBmhZbJqoqdWyWivbNKBJSrWoi5CSWl45v35iygN74LS+5GxYeFlgC6f8P5VEU
qAwR11oV9plHXgypVm1ZMi8kQQtP3nJYMp6a9WqphZehEOqCyC94I2rWDqEhczl6
kZeJ7U7STxYxG/bqKMOd/d3AgmT0a2BGRFTTmpBdEEV4DKLnFjuOnjDFpQTFTiXX
5N3H2Lz/7UpxmMwptopaP0FBEcdt/LDVA+zwOMrvW8462khFa0Rr06gkrbW2uCr7
RqoYWQ4uqYde9SbuYVuzw7E8mjZUwSzhHQwgMGsG2U0u2ZUyFCLhaZtrKQt6cSeh
+TS5sQ0IGkNwTn7S4A95K6feVi3gX55VgA+E0WBFfZGrr3S/t78ELxMVJctvH7pN
UjXoT7hKYSYy3mWWSQerMtt4N1oXSMgKrO28UpyuzuGztsETdOElV299CI/VjanC
3pjQHmVoPt6j7LlI6VwK/qFdA0vo2eZGKfTdzUHtu1Z233aeC85bwCZqL1WcYYhg
kd9g4rjZmWbf7NO8k7+S5u1RdkjKmBJxqM7i4w2Vrnf1Dlhlo6iMLP2kU3vVc76W
GqsJVOBlmpKhfXDjvAT3B9UBoDPvwt7CLaqBV/e8FuKB4Gv3o/DZ/8mHrzFiQXK1
mMls6nmQhLck48LUvmBMD9rSC7v8vExBoSLNgqDzbPew4GjJfSwAy3FQaKyWdtfl
NtvzfklZeMPmD2+8nqbCO2kpPzRpnfG7fija4NOGVZAyiVEzd32nzKZ3Vp+plDDG
paFAG0rWW7tJAmw2GKq2ru2M4n8L2M0PgQTVkJW84dyN4Sxe8hn2CSsnmkjMuN3K
Va16qaoy3tkB83C2Q4spaLUw2WmAW5rMlkeNSXoWvzZLpAc5oyahitXC8UPRRw5R
D23kgVWrVCYijlfAcwzWqyoVp+VWRdgONRpNrB1NcfOr/YVBPLwSZhdouCIENWjC
e0Y8sOu8S9hEGR4oPCsqSa85S+1UQT2Pg4o9Yt4i3gg7He3n0ATLOFmU03dOQI/j
2WgjrlSojKVDe+BtYpYM+FrVgLNlTmse9GghH+8lRN5GP7GGPH3NdFVIG2W73t/B
yobWCtygnIfpCTy+H9T5vbc2totfrN6lQ45D6wzHgFYM/z6iHW82em9Q0uVmY8Hb
ItnPIJ0MREbzpc70fLcxHOhRLLAXFyO5nHi6TEq2D0GGgt9A2tESYXLJq05r1smG
B//e2Ju28yQJEdJLLykaEFMNmLwOGEp1VCS5feGWEtWlxu/rtSfz2lnyDc2nnRvj
/4SoLRXXoddeKnNWXQRo7hGdTlePelFJAjjkwWjowF6CsdcU4KpSz/YEurc6gD/b
0+VO/URjuc8To5rmFZepqgfdWMHirnO/b0DLjE+knDCVaV57iwwU9TUX4P6uezxH
Ce59pgHRNw3eqzjQbZVGKdRnsyJ0jj/4NQrhvjyJvrTglZP5bUy71HmKSogufbt9
3RBHgv9FqetLYGpIgW++nkykeosCX8ctgZ/V9O8TSB3qxIucGBgpS4WnwOwqcOfN
yBpwFDkORZ6/iSVHSMzkAkgUBpzkdlWsYDKjD/C6j7xBsOEKXDolhssVPyXUuC7Z
99kE7nYpnME5bvrjljYbWrDD1vcoI3vYxnIWI21QjYY+FIyob4VI/X6baM/AQm56
RScJT7XXx/KG/dSSWFxyXFXLbkcd9w7UCDrpWB2wKdrq3iabJVt6hkOgTI5lPjYf
sltxP8h6vZsUj2IBZ8mu9+/7ZgtktakQljmQgqbCbA/Aincz2glzivG2ysj2C9gS
FfzNTahnklCTTy5nFGNeGpcIFoJmTfeb6QZV9a5kgkrF4NkDcOMHHHFh62I0QsED
IsFZ8J3R03RsLuqKWvmccgahx5xCJgp3pwZe3v7KOI016jjmwExOaRA4V99K4vRm
CrodFGjYual5karkF1a9mFd+BAIRP789nbs5w6y3PymS5LmUBrHPHlkyNx8U6ZlG
bPMADAJ4jBvNVavh/2As68ICWglNEy9XiVZBpxBzlf4nPeCssmjaQK+B2jFEsEMK
1taCKJUnrC4c/xskoyMlKD49mC2oEP8zKXCMFDNgaPDPQYCrBUG+Oo8fAIzimezq
eareW74tjlrrt9/q+kfywjQE8l2V9abNHYKJyOZSxb+qypYeb6FU8Cv/6k0NCnMg
CTTxhA0DEXUk745dJCdGZVq8GiaQOGeVTJcfaoUog8liel7O+TYdyHN75qjqZHYu
j/TUezYCF/Gjev2uL0EIQCobn+++RdLfDMou6qDY5yOx+seL4Zktz+WNJiNdivP1
5J0c7vsF4N3qIEWuW/OzYISzYDuGARdp3kOCVYAfw0B6SwT2Q3zKFIimvZV0F7zb
NZaYSEvXhQg58cuoPdQF5poixkZu56wYCQaZAb+U8pTbjjWiKzjBNFpdrjyX4yM6
rvAEP+rVSdPbOTSJ80ljOWPCUDYyUeuwETXONZpXXEWZewRruVQQberXJdLXTAF1
fUcOYUUli8Lw5MomdvujErUdYNpTpuVoU1qCDyoz8tLDouMOzPNdWVjRSx3UH9vW
ttrM7p9wFkC3TRiQ4+AMUpS0W+4LJUy3NpFMVdQy8eXZQHNwFdJut4LuSXCqJJUX
bpLmGrIflf8XltLjj3UvrICIPvIygpq8KhMQb2m+ZPd/qL5w0Etayd/elDTEunbc
NODK+mY686ElUQlrDQeA6n+J94lNVp9KwBIYENQe35qud+RJDqH19PPwj8cSq/BZ
/VubltvY1oRcEoJcoW43aTw4zNI1bp/yjODGvphalSLU/NLvHF6RyR9N75fSFLYP
GSdUC3t7s08kkWGZv0YGl+/AOVU2QaF9w6WPbyFLQec9KGIQTihQdxHU4z+tdWTT
QE1wT1WA5NnQd9nSH8Zu4/Q/sMMEdCzupxZ7NczIMYA+eEvi0WOJE99/avX20QWP
DZabzFcpvG8zpF9GQyv4GGRn7xBHa8ACNv5CGUhS7Tgc1Mf4kDQJDcuM46I5/Esc
k4uFwXzp9KerQ5eup28hPqeQVUAKam/kQUPqxieX94Tn1ireJjsvI0fwlt0zzHAq
FkTc4jG0AaBY3B+Nvy5HWKKGD3+cLMOx1ncS6qd3HtieavzLq6Z2JdiTJPGeZ1Yn
JAyXVRNQTfiJ10b/vtGNKSmD49kg+HibqXkMaTQl7MTyGYwj7viANCUOV6wz6csc
lSaZn+WsM9AZeDKEMSyaEpVNezAgtN+9fyzv00wfR6yWh0V3ePLwNxam6LHlepvh
OqHKvGD/6rXPjzyCpH+V/Si526B6v0B7y+KWQlg3TKJdE206MUZMpAfw9rTkK4BC
inGejdrj12x4L22mM9tr5V7RuJD5AwD2gNSo5T0j9ytvHKxSl4pT07McfNCX5rr1
UUshjjx1PNc6S4SgxEBj8Y/vmF8nUgoPD7Jkie3bfE2UTd2cFdrpOrZJgiHKnfpQ
7uDyYjqXSZtmSjaryzUBu1zfP4PnBvHSisVnSVfURRceW9zGPa0lXkHOgLAr2vdJ
uz1XizSd/yxM5ci5+QwHZMgkMVWaodwAtnXXsd0nkSOW+e3CZ7nHmhoWea6iwzuR
UFQa110odmnM3Q4h6RnP4MaMaUOH8Sfm7DLXmoop6ldWqgMytgD80GOMtfgmS1pl
X55QejGklSZGj5GgH0qGXCVKbHqwgCexYe8m1U8AZyOpKnO37irvBxOvjIF+KDwu
a2Bs1y1ZOkAfWslzB8MMDVEStLSDKn1R9q2ND79xmrE6tv+kWziBINPG66yF8ZaY
4wQ7xmeXt9b8X+hcro4cyrymumuQJSwXvcwcBZS0fa93X8olWiMIKXF9UFvnYI77
TltM6V2DI2HbDYg/Q//ZyKhE8mYd83tftTYEQh6IBQdQGxLZZsxtzTlMailMtkWt
08INYV/HmK4L85L+MMQCG93Eq1hxs9pvfu8AlRz4zbadT/EhhrE86+dJfeOeiUOm
4W8totigeXxXunObihEMmmlqJUhDHADDSpn52kO24xaVevXpv6hh2IsGTWOK2S1V
PMo3/uV4mKClhK4DKKoWo+gJDsjgUnjkY3V+NgzzJHSFfDN9aI0lox37j6d85BDU
eorkq4yNJ7hqZSIT8eoyuTViDAojI8xAmiGi8j9dtEhdUzsBAiRim/UFn54iJ3j8
hXd+mnQWcir82Mm75SGS4A+CrfrPBgURBOGV1w+1JFPORWYQpNWlqyA7gQCvmbbh
d118vjxStvawKW2KmRfz27R2YUDgOheZNSH2Ltan5qTvQ9BvUCTguBebNE1z3tin
IoGWY/32zJDnRt5/h5btZVtK9mZiikjMiVD89eTUkCPBB8s0aQ/DwENvZ++BtNvZ
rw8EOvvPuzPaTcBhjVwEe4fAL3vwj3gWt1R7bQ1hraWLfyyKAuN3AaHWycsuKGTv
ToQ1He4Lo+TWRxk62pZopsAzMVlw1bvF3mc6BcicummHXAjKcnwf2tzzUHK08bkU
pk7YASfm2n88OGNF1MJ+ruRtFBMvLxNZ7dNqjq9qZFFEhhU4fTeCsxkI9wGnGU2G
DqM9FUFqtaOJV2uaVK3zbKirfCwR2zaCYHTPcqKmu9Il1gHovCO/xj0I6g/OmnA0
MYj+Un9zJg/lITaOd4Ojo3KeN5/s2wMrwu3kcof+VnnWyhq4PqyWfjoKR8QhUYeQ
qqE6kwRGfA4KMA68BvOmAFCi/63EsGIxYC31xFdodFtbb2pAdkHTB0VtZ8uIa0JZ
9NpvKzt5z5jcp46wb2woLprliQ2QzoPywB1I6Rn/vO1NRFDi8NmlDvM0c5tUoQZ1
mpMeoQTvBYEgtKfx7ZL8aOavgH4fEXwfYe/zBfsQ8yjwmSXqXbu255jonsX0FTHB
ND5tIYtsqwSLAEzIdxzjrNd4+q08/70qgTHjj92AVwRU2UAZ3tWXBp5ONpwCd141
FGPKApO6ZfxxQ8ZxhrfUdyFeOE4Td9QegTM+BJb9SrFapOmcumDddMKesG3cmPGP
JwFBglmW6heJ7r7/bWFj5a/t+BnkLc0cyjsfe4w1zSf8NBPs30tjJiQTjjlsRN87
Z6l+Hmp9hjqaxZAszmwEm4wPOwCVdj7++lyNskLmWilKZIchl/bxHBTCM6UCF7yW
bUngZSiwY6ltrmTcvPxN6/WNEgbWyP8AhsUqYdn1ldX4hrnxu0uZ8uQPJcsOWVtY
sfEGZ1XrueJMwq/EVwkwU1++TuOmg686C6RBYVRYi+JKOm2mXww3Rx1s3737Iopn
6xy7WEe658AZCo7J/7dlN0tJrofpVM/nkmhv8fVYY58C/8sYDhcUo6ly5Y1Xh3KK
iASBoky1GKy8JKMz0pM4Yz7SDYEKw00eA1BWhu0ZiN2/X5WS9oHDn0lh8PF0YnsY
F4NsEPyY3L0A31d+6l6eq6ZtaiCZ5ese5lgbVUrnsHn642Bgv/8T4Rtby2DS1Rs/
05xMxhCT+saQc1rB80iM2q7MtoFcwSqXOEochlwoS4q4pUKw04jgR+4xJNqbLCfU
bGP7IhZqFmdIR+StokF7CR429tA8v/CukagD9Ojj0UaDDHcZ4bzj1eMfaE40myHy
voZ2zOxVM/2tnogylWweXQBCiQRpKPlk9axgVF9NWoBYewqw4XrMafpFtF+OM0zO
SlnQWc+3KgbY0KGhZccGSFHNhUiPKr/p42tQCdv2EJRDiJ/9L6P2fNhJ87jYGj3y
ywpQeY7ImzqyGtk2IfCjUeZ5163B8gjx52QIO89iupre1c7XTr9eP7HKhFJKuV37
1kvKZ1vENmEHbUFhX0uxtil/rxYdPXUfjZLJmt6DXL8cTHBCGlynTXvMTi6UkmvD
U6Qt5BJK7maZA47e8n4y2KHZ+PXHuwxgfWdBLhLbke9wfSMaqRwsXj9VUigWaPdK
lRg/pI8PIsoSVwWFXsuJnMGgVrkXIi8aTh0/pl3yt9Fb+TEU/LS88SYufDm2yjEA
mnxcs/1WcQbWjXzf+MsDKmvDktPDyCpJdTqmsjPSldXx3Q41R/UNoF3V+algMBxe
HSIQ8tArnV1F/c5xky46OIXXe0qIc8Z4ITshxVR5N8DxNNaY0Awh8MuYRvmB9xEc
Pz9AZSY163eylqC5xInfKRU1HIgqaE1AZ/9LPUr2c5L12/YU9WKXvAhNH1Q9louc
d67i8ehkbN898+T6O0grYA1FfJFP9xPY8/WDbpX5YDxXKKbZJ2/BhAV+ntjjpULs
cACL6FlyPuMyFoYJd1jTNerOsQgTfULE0jX5A10o7tzjuD3lPR5fThWNRXUCRZhP
x+wRe8u7Eis9J39x7elZWzanj/29+CxPeSyGrCbho/5UKa4VyN+FdfCSqUusK8Ce
nCOQMXtosUYAjXvrBiupkqmV8YY0DglbPJRUryUCFPa1K4r3TuptxD8GTPUn3lM1
IuHSNss5OquTRhS3dRTNL+ztzthJlHd6ZaYtWC99778Qh5F9NNKiz6a5zJTrs0sM
/RpVOyHSdNERnMIuXUSqkfkM8d9BFbsUDyNHFIUY0frHw4Ev8d7Fx5D64Qy+kmla
BfrkKDbZbhY+h//qK37tWemw/L/9M52B1wo1N10R81xSeoCkySQea7LYo77gx4rR
bbppRXylQ42Wnj3yfEuEtZj9FPFOzAPJD7O3ysKeNBQOHQ+qD9KANh6/R99sN+Si
8Rkz0oRFYvmo0EbT2cJP+vF63msKdBGr+G4IWPNmZ0ruP7FrBahDFrR8M7qJBUBr
G6AzxXyMskkOKMXi+o0pKRHYugNbug2Sy/a4Wwnts++d698uoLZVRT9CfKaZNT6B
BYjLywQ/Xlj1oBwIqWZuNVo+cu6H0XLje0WIjX140No+rwmkEaYOa10Vb7u8zyr7
gjSxtwjwBqPIGEG6kEZ8vAhfpt0m0aoOCdeXNPLRypeNUuPOmLfe6EiQaprM7eBK
Mmne2MbcuHCwnn3Asn0qbYc/US/TRIK91e9suZcOvt64+W4qs04t/BhIPRaSFw5A
oA1w5Kbbh8JWciB0oteG7WLo+/nRCM0FWIHIz3nfGEZH9Xi4B0M1RX4yQ7hsPB3e
xJ+Z1atyIxwwJPxG4cZR1R3eKYb7rUDBAlvoEc/VdvPBdmfat7caxXzu/U3ZHdIe
6POkqhdpnfc8g24AUC8e+nPzq+KclN1IKB9ReS7RcB7AeOzxxbwMjgtRhzl879Uj
l3o7RuBXpvoy30F7S8nneztWgI9w9W8WFEiJRRVAl14Dv0sKRYt4TLdZkWtuqAvq
Ros3bVJP1VtTcJEKCIwLXo9f00U2WY2WXYrNuewvi2AJvrlNOBsgQ2A0BAW1BZ1F
lFgv2QLrpGVmABhGmPPkX8QDge/YR+4aEg4KveFoecOPB8UhLPYtlV/2wmUKhfZ/
vTpuOKwU6+pkpOmhaQ45qgVxCOTtiYrt+L34sDINeqxumidZcAj9hNHd2M5M9ymb
Gpsu+VKkwEmGyt0/6lsuPCZX04Gmr4HRuMxegTS1X8Qkat+Y+kNm25qKwLghG4F6
BoDP+mz+HQcTb9elqwyjFQM3KgGxGZCVfyFFfoe6i9hxPSksCCaZzPW5wKqTZ/5Q
QETQMwF/BGTKGaOmlPf2+KFD4RXfdP0Oeru1FL1+F7LXXYCZPQ45vx06/ov8xTJh
/ku5W5cu9xdNMiSmy9h4gPFi73KIQku8pcKzL+BowZES1JgqeqOqY8hFt4TRB/dL
T18DbF1Wm/mu4uMjgaxuK7U8PGaVqbtDdFeU1Xmw2e4FdCjpNksI3DNMaTQurCnb
037n7zXFE1G3eglBjEJCKdJYfGMIgZp6pAW07LQmQuMWewsmtL2Q/kFcda9TRuRp
blSGChVXCk3KUimr3Z48oxaeFb5lV5qKJDzAmj174om2q8fhgNb9zwt8GKmMBbey
2Pr4yYoSZMZB/8Wn8J6PyHKbAaYaHTD8C9YENE0ZyNn3UHkFg9dzKMPrQySKAmvc
NRuiU7ZI6Bce65yQW0597IXRRFTXuGbIQQyxx6pZqbSAgm7IzcukcCjrB6S0h6mT
0sq7sbMGMJDKUA0e8THghi2chnhnGG/vJWxjUJqXTLiNDdSGazTEUUgbwvIkLVlU
N9yPKM6MaPqpmCFlxZomkZkzQQy2BetKmdAxGDtQUv5EZ7Qykn4aqOcNxM6d1Kov
2yl2nVdD2EBuNmBnjbcERm/JvzB6eU2mHbbRAM25MuxjbrXSlNnoRlsc9tzD83+0
ZKsqcBo/G9jjqaLjnKLXAB9d3HQ3wdNJagr9f6fLIrg30MkDiEh4hvo7kzoBPnOi
84DYYX3sFk/S2N27S1PzFsDTtzCM/daA0+Hpazm+flkhcdxWQQFpiCdImDE7pQt3
NYHxT89EHd6kWNYotxFuMY23StsRrAqlWimF8ykLwJt4p+h7H9FZUz/x/3p8Sip7
IvmiRL8QaGgE09n2McxQ258TkZ1q3HeUJqSxfQoSnUSTPsOIS98r944BHH7+cePA
r9rkb+RqZjF61MUSxzjc5bG96IHxMyXdk9vmb/76spzYwhinyZRSTURKO1sr34ea
JdWUBhEVWAufMVSM2nCCXmrHKeQdVe6atgrG1HHA5X7ZBj7+L3qSreiCYBZz2nlH
y4BPlhhupKEtP/G7uo9qlgYMcCyygINbo+W5Ycgz8nlzFOzcVlWwIJjH7q8sVOKh
9vc+3mSwtpIK3SygXvkzEUVeidn2I3QHkznCiMm4+mp+Et8nelAEF6wnsp3djhBz
4RG3Xgf6bs/KyETFdlA4lwty1LmWy5AxvHjmdSwlxqwYEsXzdPe7XlG6xEfmK/Mo
oDCHQ2knzSmtcfOqT0WWPcYajdt/5FJxAEUb/sn9opZxm7Bc7YSbxoQnySE8pBkR
ldBtBxcCfdq8KL0QbDhIkVj2QQ1vh7qI4XwSvzqibmiOZVyXOmdWcNVRxi1tI5py
EYZPDiyaL2L9jFlE3OSJDNM9oVxcTGTaRTs8y8g6ZDe/kmiYX5hFgj0CZoBYDc2H
Z8lWxyCPbiEGbLDzf3NvvTDOA8NHdoufoHJvAeHhaK7/1rP8DsBpfZYXk/Jdbb3y
3w3GQdci3BmZ5Fa4Ke0qnctzT0aio09i3DcWW6ghhTuZmqxG/m+re00P+/lyxHP+
E+4oKMyeP2ZE8w0IxbRm+pLvX3eW8vzUJ092pyO42zk8kAVda7F4X3EWCnxtWEUz
1/hoblctxii4ZkT2TdHChloizSI81bVZt4ig9noiEk8G8MhxSm1vKEWPpH/FPvr5
wtkqSpBXEweW8eROWewCUOe17Tql/DF0wZTVBS0+v4qOCP8Y4pmgTBXgtZv1jqFW
I300r8qU1AZds08JPx+4WeSE+XINUvE+TfiacWeRhbN++Ait/39i1kXSoEFZU50U
btU8cm6JawH8ePZcTksnlaUaM/ZHF72cjsxWDFE4ofp6mHO5JhQ4keSFhPrDfMPJ
7pzNoFhPoQWUrsU3pw1XhoRFjENa8e+gbYteOxkAspo596PHmdNxXqRSVXvkBfwT
yJCqs4girWc3e+JTFKweeeas1qQefx4cv1Cv+n11oKoKV2QQyoWAeVGxX5SI3Fop
6TXMrecbqNA0prcJ02FqXZHiu8sGCpTMXtbVYA2ITQHNBdeb9rY9XbmvB11rak8J
Dk3j1b6biSVq3+79zK+QNb3WliJRMFiUEO1RUErqwYukOit4uTkhiFvjG0k34sxv
Fjn95kD5ElecCSBV7MvT27Exa2dtNhpZk0PkKDyflLNuWMH3Czq/3l32PaPBGra0
TLitNBIxMpx8UElR5jhCh7x786JmGwFYKQTFOm0eoK+nXzKYMrnTKYk/HGuuKu/5
HbrhFsMWoqTbd0L5gHa8QUJoBtcaF6Oe37DNhmjX18rk0pQaKcD9/RJ/J8SppDoz
F4KQeUDBmgX648tYZp0eDS/vqexI3Hjil98/2ESyz8V//ZOAVJJBnMeCtpnOx4vJ
5cb5qfEA35HRCotxQA8L5NgxGNSiNTy3nUVOECgnjuayFH3W1uKP7ojdSYe7IZ9n
NqZaYW7WzjXm3vFJ1xZMFOnnQF2SLPapfXmTu0IeamVbo64WB5zn4f6fbzEAgDHK
j7uCrxnXnolP2G4N5PQ76RS5jF1ZJ4Hcds0s5uC4z9aTE9Lu1gmtzcJJVo0JqxGC
4naV28JEfYeF4bw7HkiN1vRV9ZOpXgau/b3FWlxmRua5O9sR4nGbL5uB3U/P2ITn
jytTf+RSymJsI2lfdN47LxmXO6QXwiapkL+jWxvX9kSqyY9BLJokj3RY+fzfEY5b
xpPCJATYOXOOvoABD0BEbbzqEA6m2MDABXaG6HbQECnVzzzauVXNvi5R5yYScv4X
ShXgb759lucM7+HaKt61oOF2BwV7awcx2VYQWTJF5TjvuPmsLk7h7LV7z28WYLE7
7KvhTLxKcdYreqt57pFzzmNyLAwy7AbCpHO0d0PYr35KVwDAKEC8WYK4hjYI1wc9
ZIEGJgrKlWvbP0bFXTBMxqqcCPBn8nLlzj4uoHPjWBp7BGWGN7TpIGjFxCpUDrzU
kepAC/3XlIIU9iM17Ag/Ed08YNZB8qzxY7Bib77iEpyOHCu3+SLRKzvb7lbV4XZ5
TMgC6kI/dP/qqM9SHGW6T4M4ACcigmjRKQscZ2GtA+7Ul8d3/k9M9vq9nM5LpiXt
KIfisghsy6SBYtO70MIPgz/9+PNx13KVALTWTVKca50dHXH60gRxtx734GBPf3y0
Za+GMPrbs6k1R4+DzBLZZjhhgayBHJ5JG+r9pl4yfDoVwixHiCAiWlvU4cjxEULQ
ZV37sxha1NOOxJZbZYaBJK/VdLLGvnrhFByqEB3Q3aTNziXSX84khBzohZ06vCau
KQYN/860u/nIVlvuF6+7elNvzPj8AJ/v9qI85Ww/94lbhEromWpIOVzxKprBtqo9
zQXCp7lg1eGDbeMdflKoRC7N42hnXo79cJiZuk0tf49WRvC+4byKfnYI4XwMwzaU
Uf9L/dHPg5Et5n84FX3wAOzPL7PMTcHELPGc4PdoVGbWZ20BCbCY0bAQxQghpJcN
69EA/G8PdcWrD8mdnYWQnfzuHTOSrvG/sRrG6fJP+5Y9j6RNENJZJ23NBe9Zsn1J
6qO6GJxdV4Exa/fuLlxFJA/JQ7ri8jQF/zuuCaHiBmeg/auTO1n6aluWA5DfVP82
WvNYU77wi9Y7OvDefnRtQicnNPBPy7Wb3EiqalNlTWavBUD6Rpb0PKUM0otiLnVV
pXKSwDb8zKkahO7g2o1PxYTAL5aazvfK4iJ6iMi/0AWWYVJ+8fbv6VoApoVFNedD
t/cdVEOBlVFdVXh5vAzHN4Bf+7mb+LuFEQeO/KAvWzUJzqPhdRP7Fj/xMCSmcrNz
U+aiwdLhvAMLriGIfJZU/hiAIIIkDSySyyQhhTxexP5yKKXqDZf/vl51HDDAyu8E
/mZzwSR0TeHrTkIB80DX4Ko88u+y3vfTc+Uw6m76FeFWbQ6VTyVbGDEwbQV9Lu7m
bsQFFSI1qsKE4dQ7wLgFsP0fz4tbfJdqQ2JN9PofOGxiOIWR9pnQflge4Wb+z6s/
1fp7dJvhwt6rzX9fYcmIWUbAYUJZdmTbZlc7CeFip7/o5PWbTcuXKk98URSc1Gp6
dLoQ1PfoCrex4Ch0Xy+8hTnq0ZXWtblD78PVdzVgMPTsj9M78trj5JKDQ9tTbaLE
005d6TZ+o7pUkcZd0zJjf2tblO6mFx9PFb9z3cVQ6wLQ9CDqR4ssEEeTv6zuhI7y
9T6JZaxPKNCVj9fyFYFa31Afqj8i1j0OtDppiXi73XQdi0hdfn66VpzreO095ls7
8hxaLJs2QuXCZnr0XQczq4lIwyWPWqkxdGfSJvhgJWwyqqBTfx0S/XCylzdMVL4c
ECjcqJoYOSBsHds6TvTM2jhjG/OuW0JWz99I8fXveA6CwvbyNH8sxhuV1lrkvnvL
vj9clr6UAexfPcRzvkRQNku2udC+sHlgSFsqe2L6DK8dreV6AQpkKLgYivctjXb8
hx4asajxODlHWP0ipKSKKGrMOgOvgnw8+moMMBGT6VgzgsPXg872nnQ2jXkJxtT3
C65cgLGDlbn5aTHFzXjkk9wBIFU6kFbwQVbTHi92MjuhZuZUScfRK9cUaeJ+5D2G
mNuvWvLARIgY5HgLJj6HN+h3zcVm0lnsOMIe+I1VZ8S88XFtjBghoAB/Nt0Wn34L
vh8QpLDPrXTPuhLz9j8NvSLoy+IYLLhbYfxAKfQHrjnSp8q6mjTZRXH7L/xQ+4z6
40bPf9vAgdGJMfcvZjMwGiqJC/ROYCnJF7Ss50F4T1U1Hn9Jgxc8yGKQofKefxbk
naUPTTYJajTxaQO7SZTPIQLs01yblFVipRwDP55YH1KEshIU3CJXdj+KSQovKUQZ
R2xv8LUJw8H4tcfGG+ruT13m15eSqlZ8YZB0A6t8d7dOA70RqApQ1dCDfUCQaQM+
32O6jYpjVZoguPjG93PBL9JzTwXbU0rTglnSHppvz3r2FucDyfkbwLV61OeEdoHl
25EK7eJHYTjUoOktb7nxdziRZDJl0SEQRNLLtLt9mmptJStjFAEbsJR2I8VU8tL6
udFMyzbwTaSjwCIzHg12O6KnpVAusW8aVvn7/4Cx711aFQF5EDo2IKtesu9rgVc2
S2Djh3MNL03Z2zO3wnZpN/SJT7NWaJQcZLL8xsW/V7uwlrodynrH14NYwUkwkwJr
1Yc3V7BBp9wYEeLmh6h/CC/zj61dFC1TG29FjsMFgOIDMekz7rkuYX9Fzuals1DD
gzlM9OfhS1V8tyJeSb6dz/hVzDTpEaS+1sqyFLmWxDZvaFTye6HjWWCM54Df5+Zu
LC9K7ndeCgPTacS4dIzVKVYtH9SxuTHWIbI7Xm7gxl4pEurLDA1oDjvBYvkisLyC
bmo+iIPRSVvZ5dDMf4Nzrww5gwWG2tSl/B/o9LpGwESvqODIl6SHW7lwJDSveewo
yqxkxvyxpeW9z3ZlOUkv/CHTQBzjzO0uzGBd0SH55hEY34fhbB4qsJjba0PWxKF5
q7U119wcFdu9BBUuvZ1hoZ/MZek2hP/DBl+JNVKkYiPaijJWBtMCWUZ66c+k+79Y
id7He2hYD01RGdT1bv/WJoSMpvcm2JFBiRoLzDqI9gNSzK0OIjZutT7Mu7Co7PPj
kcDDc+zZFEuhMdtMnNbRgUEEP9XtFHEBvSVdMcrx67QnKZeY+AxbQmR2e4DeihOg
FQFWx2x3/Qr7saddfeoI0TA8PP6mOcV8dpuCTotnLt0f6MYgFunzIt//i3pADcM+
7i2ziUXj37i+DN5Zd0HnxLI8Ce82Dtbb5kXCug4oO5P2LSn9UEiVI9BttziM2/1K
3Mpby2HC32TJ5XE8KqkP2qYNtYqWogU4EW9cZ2HSiCNkvSvS577vUti4kI2j1Sun
ubvMd+USwC5voehVmIVYnThZ/QjPg8VpE0vuJ4tx4Sfd7pDWaPyO+o3n5h+YsYwq
+gfpMAPwhecmIGGHwJPVSG0zeHlTMHUsm6b6qlSb1gUdlRfWxqLlxM2yPc/VHQLM
MEDWaWq4RW4RANpy/GHm69XKH8cMjoIPQKiTcsE+LIuhImQG3wVkYUtx99eTFHbr
YJo6c4qAJo6dywwB8tFJZie+BQnZQqivsALk+MXdkDgvQOxdRhkMFOuEA9E7AgL5
iyqwvc5d6TTSoFRJp1EtpGZ6+JVJcarvndIVDv0saq1Ls/lVuotbb6leTuhPhL9r
ziSIUYqForgW11RGNPSdvrjfkUDYYJNNeZajg2ISs+MpFAQ+cnaC0VFPjtobkmAA
TKEeRr70RG6Rw6Sw1gepjccXt/uzvyPtnmpNIEFlD/U8jGNk2iHHIwk8yc2iqPZI
vTtjnf8JnXUmMk/Ft1gZjOQknUqDsXxb+/ttyAq99HUZ3GqnhlbvvbVUem8nQzeL
rMH94LWEvqmQp+4wdyyt9zNeDukofnnlRS9Q9SMDo7a5Cx15EfDIjyQlSjhoC2Wb
FOqD9B919az657eeQMDHdluavQcefUfHb8hK0SEUYC8bw8KHknB8otcj1aAw7cTt
AXMgcdZWWiWDtUaNBinMlx42z80J06bzw+3bUyyyypRLk+j55ifkYTtonOV5NUR7
Db0Vz+sm3umAaBe6CDXT9PK+Rf3De9bBYqp5SvKRJth2pPZf+bUkopbNT6ZPDU8i
rpoPi8URbs0NF0tHKqeBabd6Jh+M1D+PKm4KJE0Z7hC/f3WAe/Lxd5g4eCSKzVpp
42BUCalbfsvkGDelrTzKCjLjkpgbvzcp/krh4fONrfpt3gfefxDg5QYSVTF1YQfi
qi6B6l/AYxvx9n/Mlryavi5Xys0D1PZbmRAiZ0j9tts335PdbmpTvZC5ttj4UcXS
NqQYzB0cy7LD99vOjMM/68oCEw9eo28mNRzF/WmfzZ/R3Oi9tx2GRY4rH2LJYOhn
YLYteOq5eE7rdZciCcoGqZ0MSrXrML+I27zYMOwKZFi/m2NjocNPbXG/jcVxzKeZ
ZtS0FUvGkpRJmn0PZw3FqPl3ic9dJDw76AYPrjIvfFW1xpx04HZI1HAvLufnsj4U
paWf9a/zX/Vbp2YR1eMD0+mnqSx+iY2LXfk3gO24jQz9MJ1mqOqdg2CdFDXCyd2p
EjHUr3G1V93zz361lPN3qt8p4t4roc1AyBIVVAEf1YLYL1be/F7d8n2v1YYraVXx
2no6BVIwDwx8Qma2yttjPbwvKE+cj/ZK9EZ0jaB1Lz75YLEXG2VNotQ+pghweJ7C
5z3I6yRFh2DFcmHcuAIGNBScAelA5/n9QZLASfNTLZ9QgqnuyEf8zURbDFFKH/yo
3TGuwTrxJVircHrXZpvjiWwhwQcuaIvNt5wQtW8TWI8EnhP/Z+Bwjjer3/fVNLIG
Wh/KKAaYOrIjepCSk2gDKgsqD5pHJnEEI74HvEWv22b47LvriP6hfOnEw//LUvii
VisM3QSmNQXtTVs5Ye2WKePtXYYnuxk/8O3aX5QeC+q97L/X/SVvBlSwscvaMt7T
0CbhQdKN6Lo1Oll2mcs24TJcYw/N/Th2ZTtpIhEtIs2uUKXGsXe/qfAREh3GCvGj
J3BJRKjAwqpgvTXkw2NbZoH8oeH++BtAqirNoNb3X5hGe73mX+ehJE69yiLvHxWC
GVoRnog1r9wQNjuDWJrXiIwRt5jn728ZMppSUHUCjS+cLIKdevDGWhqHu6qnwMCU
wa8R0PZ9v9nB1FkfOmuRgqCmOWeGNkBcJWMoWIFo4YEA1uY3ew8NIaHPXUYONeR+
DBU0ZUVdI5gmh0uQMoDUK8r/TbEb1nPGHV3CK0UZSUrgXz9cmxnE3d5sSLeZRsHY
87Ti7o3QKKMzxewUC7GxIxtEKG40ODyvtJxGhCQJd29pm6Kd9TNTINFdlMqXbKrC
OqP7jXpeVQC6jid8VM6oaIiXwHG9DOVTAnPGUZSTMT5dUzZQPKtf7CLDog1WhlbC
Wb2f/Yk7bqq+t9y6pgKjfqHCXOcjYvQRbv15h53jzdEAl6mEp+0cDWkpqtN5/q+6
Xq3L/ve7NWBzywtUq2v4sfp5IYk9R56YqnOZy6GVyPrQdu5AAavbdQfxjLLMXXyG
EuGAz9pjWT6SD3u8tH6uiHvJ/5RERf4Hns1lYL+QyvVmXgbJB7WI9qNQ20H9W4rQ
R5K9FFXyGbyR9Dhv88Oo2MZjUKAbP5f0WwahYkw2DiZq3YtHs4zfOL6xXOQN1jTD
78T7UaN5Fu0MyOns0GiSYWUkv23sNdg9Nb7PoQtgDZIU6trKHV0v/HJF3s6Hwgu0
uSKI/7Ne1qrjoxwY9pk1WHYlY/T0frDdzdoHiX0EgbEMo0ofvRS9ZaEEVoGPXFIl
pudHj0m69+f20ZTrO9sYiNLGCDzEI9TOBqZnclz15KLfEXnt5KtzYnPSEUwUaD2k
0Ib1jIsbyd3GN8pTSSdSSl/KRhfitPy2saXcQrFbsGv3Sy6IRsydW8biA0Foe4kZ
+bUdZKkZ2oLV2ePhgN7xaenuITyW+1GMNj+ytXAzKn1syMaYGN1j7rA/af7lPiOY
3JbWGgfWT93BywuxoBK0the6+CgRbB2kRYyHwtftFOFgV8LhxffcLEyQnb/LcjNO
q6uSeJZYTRGNm8PQvxoUI5xkjcvvIz6GmsO5KcBz2tuUCgqyngTjMSGQkPRkTaBq
KiXiW3aysUJmOrN2A8Gvi9gRuq8N5nAR5aaofWjlF7MwoJk3l/Su2fKmkaiPFl7V
niHRDFxhvpRQh12GNDKokRz4oqZhO8CH3EqRmVQ7WdtzNOKbjHf1LSw11edzIyPs
R/SQW12mcVLpW/52STCdYn27sLK2EvAAzXmXtQJSBJ9N+4AGpCUhP+GwKs8GFxyG
8b2zkmXIXK9jjsd7wO5Ed8ZN8v9lpfs/9nigjlR+sNMZ84j4Mtk8a9MCmp3fhhd7
SzI8H0AlFhhyV2T5xxI+xv45VlaKeoKF6nYoroY/bNxVFBOk3wRrG8jojBaRThU5
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LqEjD8dqvjTDRPXw68pLW/OGMUQSfo36kt1pFKJaEsyrRE1lidJqDkrhWX7+eR1v
+vnr3GSMDtpTfoZpi2fUpvvV8jOqVo9C0LCVWLyGNQStvT605X7zhjrihbMTV5LL
E1duDneA+S6C1BoU+S4frVfsXCL/NkCQl4KnUrOdYJU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5088)
hTTHfsFdzmTj8MtFwxkq38W5A8J0bohePuNLZU+p2QXf6vX5i0P88aYPAGb7sa5w
7gWAaboYV92RfUFVWwFWV8gz9zk7J5LaL4lDzv9lXRT3N2J1VDYJtiibBjIVnEWt
E6A9lv+kous8/SVxo6MNguG/anY88QplU8DOBDwVHHxwFAX4ml1b6kPwPdlqDOcI
2XlTUnph+4Ap071eSIKX9oMvH8o0akd3pKptPp0DASFMSNGimFagri4HPOvkTC+B
DmBp6ssVY0g9piL0oVjUKiVSRh6iMq1zQWA2Mm1nsUdhN2TzhwDlUTrYluDIHw6j
eHb04PirenjGrhwk3dzHSYXJ0pcsGSUJZzseWHfT0b/h2lNpvVBin1hwaV6p9LLc
Df4HG0tiVbEmRQQiViLxirU9Xddxhs5XRWVot6L7ar+tj2vFq6kKol+B/NhuOgLZ
DNEszQT58UKRlNnCrKLZNKwbLwQxhpXs+JXek3JbUF9XkVgWSuxkVME9xuov2Cst
cukyBaZfWOhDUEitzp9VNsCd9PHF2Nhip71DoT12+Iz0sDHPq7y3U9BN07HAR5Ju
s/LE3H2ok1E5vbg/U30KVQEkz0pEn9Tb11EX9jQINFVB8y0DtIWJJnFQzIvx0MNw
EZBvXkfHZvL38P3sZna6ovxjzCssdzicKFBC4OjBTdZLciijvmPxKo8ufVO2teLk
h6NDes3OGLpBw/+cmvYnrT/kzkNMzDOnI7Hd9zbdR45bdmxSn/U9+RV0g/S/7ECt
QVSkUmWTCuZLRX/R2dR+KVKZYaEODX7NqhiHD7pmprT0sV0/fcPLehKTOOVTuP58
7P98UHVV+WhAKh6TPf3svzlLzVD23P403R3xV4OnosWFEZv1ndciW2zfQZHNx+NH
hBS0VL2PxzS8JeJNNf6Yi36nTmU+MqVyrCzprhdtIvoPR9GI8QbU4fqIKZf0J3U/
RNc/tiwKGdkZqCN7Zo4/Fyl8tG29eWyYmWrAKMHEpwMjbPu1uryOYmaX+kY/Y0Fu
mgp609WAYbV52MwdU22pLXFKPJ/JTbWbLdKr9/k1pB4YzdylBdBTpgC8tJXNeEjx
EPQTegU0wYMXxEUzN3iPkyI+YN83o4h26oWML5C9PMDwrpXIg1oxjQZdh5DxP4aU
VqQjWd0y1oEnbOTNwBHiCzZieBSGIKFCdG15XupNkt0lkf/Hd1L40dtKq/8A6HQ+
2JhFG73PQ1+P02XtKCBF3wSUQlFsRr6F2DxDPhRUfgDnAHxxr+YkQSc035dca5ru
T/KO5gcx4PpRQ9bON39REMdDWj2fQ1NvSzkOKMlTpZ3KlJ3fUDnhZqaHr1wRm20G
kowThLRLKWIW0VNTZQ1EsQRyBRMOB1UEPdEJcyBLG3VmEdMQ+R1S84pKLdfidjZ/
+6nesVS1GtT1Ds5yBb2mIxufqsSYTi8fLhPD29IwGEqfDjTrrto9ZyCMaJ/D+ul1
n7o5olHSGfS3neAikbsvKdHb77bImWVIbm2QWWd1rT6TqSXo/MPFTrcqre2S+eFI
z4oIplATFQ25Id5U+s8sa8qjjS8WHEdgEtG8DheSgxexffSkeX0TaYrE0wAJZGT2
DwvrGl3rBb2fj0yL/koHRTiI0ljRNpLLBUCcxGyqlvSugJ1KwdCAGdGobzb69Wmb
YMr+K+ZXayuT08vCdj5evtvYkDRBY5uyiqNTU88AgUYUEs8LFv4W1KSrAu4WhT0Q
4EQ9B42BX/sc313ro04f8I2f970aZaa1puTbmENli+2lnEWG7Xg4Yf0lDBfHdNZA
IGitfBIyXI4mvdxFQUgN+8Kfn+oKT/JV5+ag0SQxp7ofJOUTqMkVczyFQ6FO9Le4
dCTxCEDYVMolgZ/epADhKqqpGEEUsvlNlv0uBx2NZIhkfAZ3zHbVb0I1ItROjXbc
1MpWKlTzIWHece1dOXzQM+5SvZL8FJKAVZDQWo3UURjGvbk+q7xHRI1nai3m3EPe
LFAhSOVQSmrlcOvnGbhQ/UQ/vpxOixe2YFhowAE3qD2i9KyOEukBo2/QmCjlUU5d
xRZBaJKggg7BUt0GQEEa/TblMdw/Ycar2N1rVb96JvXkf0OkbNKwEdl9vzZr3lLc
4khpbIklm29y5qNiCgz5t3LFWOOtQnFFoT5WSFSd2Ye4xEhV/8JK/CsODGl8EFDh
DmubvCGZh6Hi6p+ZkYVX1AveXHdso2gIMZEK0vPBRG4N6Dmv7jzWf87RXEfqvteR
ykJGlYTvHQKA6F4yg+ygU5/2B/jyw9eOAkjQvvsy7uCAqf4l8K/WHpGITOcrHT2V
qXZNdLZLa4iLwzUZd5FOy4szDVe2CMCJwRUNfnksIYEVou31V4+FGVPrgnqdUrA2
VdzeePa3EJWomxSvDNuo/IosvG9nFvGymdtLpL5kF7ciKR0aQE/3ceuLf3OceiQ9
5W1lHOrVJVY+NqKHiA9ixCxwxj70GgHzaxz8nS/3Y3dU1S8Dbl1tPBt/89CMPtEI
BuRxhYUvtKqo6zLzQ25Q9vTypesVW+5vptf9/w0RJKJXu47gScWWyLs3OT8Q1exd
GJ94iFu5Kufs/xLIjpEVz/NRfny2c85L2HULg/Dy9DBe6g2OEJ/kBst2rjlcjru/
kh/qPF0oB0eJphLT2jzEaA65YkuobgztWpFi3vhWcAWY7yZMjIzjNdespFBaYbV6
0lBMxD/vaXPBAJ6kRImCZs482wrhxHkt5oCZo0pafmujfZY2wcqcLC8iyS4MZ/AT
Mobe6WNXhj0PAxpdmL3grLpSSZvsTYpnIYZClCaJfuxRxJ3M7tb4WZneGH5T9T7t
n09DjSYPE7ptvpTnf431HfnFup3Zqcl2rc5pPD1wT7h7yKLNoYy9bZA/4YwCS+Ak
YNYE8d5wtBrgZz7hetUrf7psmqekrFH3HIxnn/JhTiifrhIhC9lqyHA1NaENDNgg
jhjyXavrdI3YysuEH4zjU5FdusBO8e4WYoFpmaefaG2cCCCZdFqLcCe/GtMHvJ4H
LTKBEysQNtl8yCcDY+hIMWd8S5/yZLakH85HnsyHoHa5+2C4mcECr/qXTi6/H0Sd
SA1AVs1Agl34/G7aQk0v5ZTXD0INs5sg2kEx2mgu3w0KUyrANZKTzdVtlYcMOk1q
U/BYHYOdaYdY9MNXgcSmRA+ODBqD1Wei7/QXv0aOPre0R+hWHjSRvEWmQQP9vTF4
5S0CGo8n9sNy+GgKct56MAF7ZCnZxFuUqw6Ql2nV6AU/QMCuIQt56VfNJaquI4Gz
oqOUG9Cp0powamRgLV5vIbSANDbWnhU73QSCWqPmjQ0Tlo77a7b5QIWBAISAhCeY
c8B2MEo6y+7Pq9tibOtvHLmdcJbIAjXDtt5cP48NHqHD7I/eTq4EDy4plNPaoMBL
A8fQjk7noLc//pzm1nxqs885zlYiWS00Zi7s/icthH+BVtyS+fXhGWscbOTAf1tf
Br1rmXGWO7HQJ5MPF1pHcTTm5z9qc7V0+u5Ws6FB0zAWNOsXT7sco3xyEfNOWUs7
U7q4fLMFeOM0k4oTN8MuDzdI6eSsMHJX04d/fakieGNAatl2jURPebw1uY355IQv
1Xkr84Tub+LPdYGR+4L8QuZ66IlJMKPG8tZkVd8HGsPjU852mSI57tX8TR24VNfm
IAsAEnmpQfj/ddh8BSn8G6Y/SUjqjp9bUXaoEqi54aDkMRNgoq3UNHAV9ReePzOz
DQtwTn4f3EFeqzzn5vAmZidO8/WdocbzUR6j2pz1G7GNEnDqkKchpsb2fkmY4WpQ
dSfvTA+3mZL1p4ACVNm4yJvoRJRz0sgBiO7bT0hTJ63HHhRYE/a5VXCNz6uL1r2T
AfhTUvPW+Ojsiu3MazlwnHH23yT+4CwahxuSDqooABdRQ7XoHvmFog95I8EbBRKP
Ux89+EKiccRLGMi2XwnHPtXbVUT6ytm4Fw8oZFawSneGnZQY3E/+1cCv3J5iMsGG
AtpTOXj1aKd9+bC/78PlUVAUWO+lV3M4SFJfI2MKoAXbhdU5vzhoUtRgH2bzmHqL
WUs5OUgCYYaER1dc/pIOSRbYVAIpI4QJmd9ZGibJildZ2FKfxs0mbQY8E9KJp1+O
S45mLOgBHTsEq9j0ZMEUqYqZS0ZznoKWQe9YYy9G6/2+mUa63s84HfyskKbjyGCw
vSGsXTcbcWRxJzdiEeIOAmVGJYobJiT9PsEEZjyA3pu1kxsUXS22VB/IQLsa0TQa
rq3GR7atiT8w0m+ByQRpx8ZvwDSxWd/lhAfbLy8zxEfpZyoxtT8j1mZ6sgE063iq
gwF32yffaXWEYMpnjc78CBz4bsZ+BLYPeYyfjmIpINi7ihxAqNwrHlDiI7qFfvLn
ASQPr7lfFMYBRJ0lt4Bx0noMtNj9Y55a1j09QOLWWVYyUCwXLyenjkHAWHkBemaY
XJPoIuXiIET18LRkVzEgbLUGeAQlxD2w6gn3OFjrriOU//sEIW+e/am/Jl2RxLY8
8tWWySuJnkSj4ZcY5DXhFERbF3Rqbgtg/SrMIskMwKPbJrhldH5Cqc3kGFK4KnfO
fxSf3sNgU4Lc1+g5qYPCPZPN9cGZKYGdj6PHjsMVs389URIufvXoAoiDFRCITCEU
EfFy9/FEtjaAKoWlUnv2JN2nFH3PNhHd5NIxkGb/n+o/4bV431pbubZZu20Xs0sk
YKZmoA4rK5e9yAhbullBsfJVYlRS9oIZ33jYQXawJMEclDkmoQG7Myh/9NxfJeun
m6LFiFLwfUFXyGgjp0H+Rvu9xHQ1QRqQDPDDXlezq1MRjYVb0KyLZzePH9LOm8vG
QHaAcbChPLDjOg2Flh3XYrDZkq7LFsZAjsMOQHvLzFeEydjH5dCxAQz/OHrUUhR0
NpewfEL/Y24wIZi8iBukPZiiv0UYUAEOULplhxyjm/XQovuVQnsdBK+jbZCY0Ml3
++AvQFZrGw55K1JtgyG5nNmr2+7bg4JquzEuLhAB7Pty6i+sA0AydEMWoOvs7NxT
MU4O/cLxANSbfnJdUx9vvYBCUEsZdH77jW0+Qwflksjpfcg3/fdqYty74ZVd5AQU
sHoBcORMWmPIhPO1+idgKE5MTYytEXsKNjRZwAmSc5Pgh3IdYhBqBvNpd90m9g0G
gQ8OvTa8r5x979ieWPTpr+oAxzTNnuCmcpiQqlk0Etn9x19hNE5Y8y81cHBcl25S
shWUZSnNyj7xNICKk5BAgf+JtBsq1/dbK+wsQ2dBjUq7fu+kgjzuEmk6Z1nLJnfd
z20jDBClaIn3dL3iD+yVZOFlGdqvhgkSKXbH5N9cW/iD/VYLvHoHDs5mK8hNl0HQ
WhTGfBZSLM+yEU8Rfy2C2egWCmbmqcQlPzzeAqj/EGAAlk9byI1qtSjDS1oQLDbM
UEnMZNjgRzGEj3kCJKzATXwy7xqbhLaNr1RmNbKvM2Nv7j1QnieDs/Ts8fOZNXqW
C2/B/qpdR8aOBEwCav2IQT37tk7lMvXpRhswV1/2dt0xLPMxNiHp1eO894Ku3VdD
vOiqrLErRr2tslj0EX6BAUD+xRLw01yoMF6Pra+cVgb0VBCXlJws0joI0yjptrnQ
cAYymZsj64flPM/bsCi6Dq0l8rgwmUMs0qCopKnCACsxAmSNXBP4X2B0Kau59epD
74MP+T1izWY+g2FTwlI+6izULJfA8d3wSLi4BlM4dMM1PTUi3fbiBOX0P7QtxLKq
nLDIQVlouI63iksdANPo0Eudnvr/Fqz6xAQq0/6BNsceCQ9eIrylTh80Xwqt/cqa
QVC1wDzhGT7Cm47/fYltGwxmROCQeOXWxac6No/rRpc2MPK/HFRxUky07u7VRebF
XeAU3uBfMD6z/+tMsJGxvlOPVXMbcQ13EzOCTsOiCKNE1qACvD+Q4bt1wUgxY0tj
rv9t6EDwf72aqFx1xyWUn9pXZFnyIpa2FWmAi0/0+Ckr53gckfIlC+skvwe1TAVi
pOhagR8F3XrPYtldNTxgUs4zZxhbPL/GN20MqqIElHNeDoA0my9f9ftA3Vm2IL+D
cRebn1Vz7rvHK8y5L3FunywO8pG2IN/Pc41O7rfQZ4pzitUcOi/kNSOYWu3ehYCa
I9GrxtweARG9+gbszq5VutQZVgrT0Em4GT84H4606cPLuRlTWtHj8eM+nUaZOBtP
lBurTVz2upRQXlrnl/mIHE9nzPPKhyHkzMomT/kOR6AjhE4S7R+i9y8T3HhzRW2H
vu/XNoRyxMsLvMuKChz2Z0ntzqZLXZLh+dT5YfHGEy7Ay6DvGisJsMvlljNXO4dg
T4jg4PKomICMzJh0HBunFtslaWdcqXnVHThLvRLQTjxSKUWsH8Fx97mWbW9YW1kS
6MyLbtyESxPJKdpnxD0hdQfhWtIxDahlR0AADgMi84NuG1jOf4GHoBqtjocI8uzI
9bUENcQzgpJ0k6DKZglGwVUsbVt/f7W9ci3UldtUyOPfE9b+m0UNqWJ5LFfbzjw1
cvzkiMgdH8Yq7IJ+DgZ2Umcq2Un3GjMKYeTdijgaDyOZvXDMFLi1YIMaqvdlrwiG
3Wfa75hQBLVU3NdexUxIOvS6yWsGOlDmWgC0kn7K2OxO4wjEKGYoXJ/CdLvSba/S
ZciIeorcW0LahY0p4v88MwAa5Wa/W22R8QVL1W2ziK0HyDyTYa0+BOLpGLGHjWDk
/bhBRmCdDApMA/thkBMPLkPHB73K83QTQXQV8cuzkX5vXAkl79T7eaO+Ljyq9Q5E
ujVVe+Gn3hm23oyzfd1bYmMGNJ3n9sVG5Ree0UgZlxwXySn6vAjTYIJ1wLNnemLw
`pragma protect end_protected

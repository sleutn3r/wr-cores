// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TvzWWudsD/Emhziu8wxLFAryompQIzOSSW6dBb0SvF/2CRKbe5nXgbiZetSF8Mnp
wJI4/y1JNmYoxOR2JMqD1cqgTB09QzkcJcrUWMa5RQFL1RxVgyKtq9ht/XvS4BcJ
6legrpqEJjxTkG3YrRtPpHs5JQbDmXlwPC2aqVKOf2I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7376)
0l+Tu6JlGtyjlKvDFJgp0ZxAp6KiXgygvcPJZYsu20IwcH01smi6kuoJ9zzyjLJ0
wAHkKBJmXQSzj4+L9Hh5dGK8eyx/rlAWe+Nijg68r2TFfCJMNH/u79kDpcylv2V3
rOspAiUvPCE293JyL/bfd9iNPcGaneRtBu1zuL5Kp3wCFjbxckMZY3cuS2v0o160
6tyLIdeIazKM94BGuwGu4s9aL86ynyfR42fP/orLUUf5mMKyoq0N3wH2jVlPsqVJ
HK7SHNlC9cunX+oMdu7Gnaqv6mjVGFYrULCyLWDC40X0/8uzILjqbNr/rww4qn4F
RMWD9ADaKvqUBgmXrxoVfWQri8Hct8XE+dmOmSs7oTMY4jLxQdpjeMBGZDHTzID5
1XejJtrs+1SAG1eJCHQrEDSHJNDXhNH8CUsdJK5GVTORKFyxRPhTh/Ke6Tug5J71
bA7fVxt8Q7/WlDFv1r24VptdFgkLsRjhhBFxFF7wexuBd7u1PG0S+R6SGD8xz1em
RP7t46q1vNjYPxasjnzkRRsJDLWdylytlDHoxiOsv5HfZaPZ0c7G8DAvk3a3p+cX
nxjitgoKmHN4couoxzFXrSQchUnlxwAyD0nI3HtUXhJxVN2POKVOKlCp2GOy87CZ
lDnrW607g4EXwIkwiie29+fvBN/bKSWfzntDblLmRPLyb0W9LmuBogEjaYUfxE58
3vR0zuU57+TaVrnLlRMmo3qBWQ7all6WLPbR0lwxMrbbuO/N/dEo3LLfJvfvw1bM
P4xLXUwGyN1dBveU29RN4PyQwccn8VPa16fiCdjwd1oP/aq+/00wLwBSlSfo3OW2
q/LS06PmwVdPJyzZQncDmmKL92rYfBmVGRfgIwqlz0jC0i8Ha/qonRNOYB5bow0s
o50fRQY547xKwI0rnPKpmweIuJBV1qSJybFKE4L7rWS7BzR3u45f+4S8Ri6YoJ+t
FUlkUXt739tAGGY+dG/HdbA9MQycezSf1yhlv3UXGT3gAvHLJMpzMxocImBcfcGp
jrK5JfCPlFSiPCRLKpzKoN16oWB7DeoW9t0ZgPEBWAJN8PClXbQ7fVeyWW650H1e
qnInnQhikqNkK1/xKYBwDNsCnEMXzKWdnWEmOKMBFKrsThoFfROXHUzfRpc4zaCK
nF7PHfxfRwLVah5bF9KwElMNxpGwN+rcHlObs9qR5o/iPSJxkl0yVnii6bWqO670
jHnvly2uV9ZcSpwomCxzpXr0h8u7dgFuvknxZO8axuU56Pq9sSZSE7fMq+HRI3Pa
Y2cph2s9k4JWkJy5TzgeMxW7wUatZ4AjOPx1z7AKtNpZzoN6X4E098wBfJIn+xna
j4kHpRRLh0xQ0XOO1UIMIdrCArv/10H507enVTmM5k74rrYXI/rOfo9ZZn+M72b8
Sf64QfxW9n0428pV4ZXHpdIVUCoDZtoYP3AjhUa346hAtYsabG+Lwf5cGrFDKSlX
w4KcTh/vDIO7nlSb0xsmO+liKPpDYPdneY+5QytIlHl8mrNr1d+r0JDPeiddXttG
lCEVRq8/NqDvxZPanJBlLZdgWeKgjpz5rfOz/lPMhWOc8r733K0Qw2DZzBL/SJRo
jRE2aCynCf70nZGMLFMg161TYQmRNDdaiF+jlxC8RlqJ6P6YvNSBlebUkjaouS5S
AVN38OWhPSFSeWG7csyOk4Ckl9GEyRt9JH3uIecaEANfkK6fNYhlyYvVpv6h+Y6b
6vyTLu1nWnOEvsXKquGM88PO5ckf1lezQZDJOyb2/13YYhBo4zliazJ2i4q/pw0m
7pz4DpW6WBSGhf5/TtavGOkbS1O6YvocfbxpxbuoU+Tn/R5jvjWOIgfJqx+1z2bF
x/rk/xh/UkGdi6rJfrntBxg0qyZSw05VSiA90W26O8KhNbl/WcG4AH0qBFVurOA6
thSmAliHn7kpuiLB5b2mCt2Lshyh0dEwv9HfHcGhbrmY8JSscHqGQ1od9IfBtbRC
+TFytXam6E7XJpOV7tBj+piBkz+7u9JItmiG86w8f2hNE3cGecnikvbCZ+XeSdMR
X8w77BPh905f43IWm/E7rNCpGiBlxJJb/vn29a9JAkfKK2jUntUwrepNeGw3vcJN
UfzwUjbraJuh1clXCDfRokzkJcNU1k308MKq3NqQDdvW+CdKXvGPJ/8FhfRf6nEn
IzLd6Bf75Rdbfhwr/etQuJRAmDpOGlTomp5CFbZECAA0nMNsYK1+al9sHOmoNiUW
R6L+pFgnazHyh7aEEmRSaMJs/siRtbMZmQ3DY7+x8Pm6KV4JHak0MWwd+5qddSwj
Y2MrHcsFHb94cJkABMbQGTN1G5VXFEn0ijLh6Ftcydv1RYtAJksoU93P0Wyzh+aW
8h6rrKxKYEDIDvnQMMj7vs/tpJ3a9zAtn2t9tHKA9rf3cPhkERacqgTrkqsvm8Vy
2gWgmr7N12pd2nsBXJuYS3SwniE703Vd9KkWpDD12zIPSbB9hBx0bZdpHbjzFJab
dVOhE6UqJyBR6vUfg4tidEGFV2qB4FOAC6bJhSBA+w3TEmyzQjvagOC/Td/9m/tm
X38sSgNtwVXIUg+/LuthaGaPxysQJ2Q0TXSmEn0gXxzQzf1+jqoan3fSys6IEn89
v41YlcJOMz2+RcQZKiwhSmcaqb0dzkGfT0xPDWW45wATXxKzje0fvHrSL4KqA3VA
UaT3WhJa4OSNWiEMWxXMOhQSGq72jlWvcRzShDEeWyc/nUa1hY71JYUB+87cDfdy
KSYBZuwGCWdAlkMJrGFDDHAAEODg2YN51rHB1JpFeJ3S+wiWovjm8yBXFkaw41Q3
c0uAanqy12RumUz9WEdGcLJD1O4EjwXam7e0u90fec/LC+Z1QodreILfU0UAuRjU
mImZfFrbhf23hMDxWOd//OtmL25reYrzWYuqfJGIZmDZ99hfBtYijzCUGSb7/EH9
d8J1RVrlHreRHzKUSaFWpBxyIJHGpm9C68gdT4FHOeR0+rQb8g6AQANArzjakZhU
r4VNo2Isa1Bd4VNTXiB0TN7S2+0wE8wqh7KTKXx3p5d7o4N/dS399AldZVCFb1E/
G1F9bkoP1amoDdebNf7tqBUcU5RdvX7dsXND8vpW2byq79t1MchkhjTCKxrfhB5G
03jMHW2AkPArzuGyKCcilayUUAnpeahvjU1va2CbSAmVMThYhlazZh3693Tnt3sa
C9NfYOu4nAO3Nbij3tLqBi8sgfaD3Xv4Mt6qFUUeydklaKK8yEiezFj6YRpaa+mB
ejpBWw6u8KY8i8XuFN5Ene+6lk+G+gFWwhfeAc1fqNyFvHQJD8KnFfJvQaLlBS8U
2e2st4F6SVYDCvoH2psMvj2ibovSgmKwPD/OGBzhLD2sL7SQ9SZe92E9Q9JzgVQ6
krGNBkT4WGzwY5ULpHnV2xGDw63SfFdIFFbn9BzktTEOEan37kwwlIi4XvIZbdDy
UZwJ4zievgK9w+8CuDvpRvtoHvTyvPGYMkJqu+5YGZmH23aNlKgMGATOGc22Qcx3
4zxbSVz9tyqnzSNGOBJKatB7z6YSAnlTkQwBdRA0MU/FZfSE2oFKpr5a3z1gmEwS
EEyJbGEVX2+t0QK8vM+M6RJevdWAQVAEHD1DUMqAxo+gGvK+mWqn+elJCh2M5KvW
lFlCwm1YfCQ/y0xg9NftTEPBnms4Wp9pyMT04J+kmfmlfItxsfSd1BBna3T7fbn7
EyHSZ9b6Uwpncgc7/Hbx5ZCijND4b8w2CV3kt91Lh8G79UEBTnJL2x21czKK30K0
7LBiM9LQfbGU5AJHgV/eC2Xd1Aw4CyTMc9mD7hQt6hm4eUS8lXOCTlt2qcVidhea
9fqJWVQbmp3mcP+3dwQFcd3UFtJU/aNFP3hcHxEkswhi4v0LdznQgPvEgvFZOSbl
s0FBhMbdaqVosPlFAoHXh7rHfRtuU+1CAjxync6Zt6oMRr+Cu5v4RFU1YdoHFnZZ
LSS3vZVUqg8++MF9VmGRvvlHYAyATQ3AE+0CtzkNFuUYu2pIlDnvTDnU5nbunNrA
bG+iHmHsCr5lxrrNPw89p8Bwq6c04FoiZz2wCLXT/xhd1IHLR04aIIry2SKb42BL
qBeEqNDMbh4mCukrZDZnOTi3hzRnf0JzYFvLEndKolBC9g+6X5JbmdkQeEJklVPH
xwakkQ6TZFy5SAFGLsSAvJA4M49+c0dkp5TIkVeLWm8FTaB+NJa+c4DyW4gHKobR
6oaEKjzXlt7Wawhl0RnG+zOiGIvD0nilxpTQ1/zYSKqyvBe/DoTVRgv6qUOPAkUr
Y16YmYJLTyJNnZ7b23lWay/dAHhMzCepcSbxcJj17IiImuYHOVHUYFbEwV20LwkM
aHd2mX12fjJgDcSYObk1/CZIuSligoMfaIqifrP1nAbG554piNYQdesnt62V+hFf
FCO5sRcRuPMvSVsIgYIQ81WowkfLNcQMSfLMwQRQebmomOeC79YZQa14euT0J1Fl
WDsRKD9fa/IYNJk3ZsU/XCskd1rOyIwUiv3Ar5Ys6yJ57DE2+JwD37WVssWs2XxM
hLlPhuFMbGZiOXu2hQPXctpltl5pdbgO36wUT6ip3rP75RWlXEOwGJW1tbBcFIWy
OMlCfRRsEv7MCHqhpugEog62XgFxCoQAtAgmHg5V2zSeJYYq1AnFjtg5PquHj/iW
W0+11byPM06L1QnqCI/U56OzAMNyhZP1kABPtsObeiJeDv0OpflorqLtArWGuWzy
OzGzV78AUxSZ1X0J7Js1HNZbCtGH3m3Kyvi7O7TqWIG2x+oQPxxRpU0KhzMA/Lba
cQKmo5y+IDv8zTKPy+g547C4qjyAIICZORXDaPDXcm45Qn613qGeR3KGLsneU8ny
NJBBQddQHSBvgXTUeRmARuOjKWRkWv0urx07ARFxYRyhCitMcwtXr2kCe9uh2r2J
cZfOhm+gcWLCwaIzlB/fqzeRJ4d3M2CgvZ5mlLI1TGSIn3WMt0zh6DxNLtPgY2s1
PA6AcrD5xwOX4rJss6d3aJp65Hqg3cfjQ6FOO1Pz6HWLamqrFO4IDSpStuy5ifNe
jidloVNDO+9yzgM4GtWIEgY2Wfon4GHom9bnB8F633IyLaBshGC2FpOyL7KjyfZB
1tZ+nKyngySUSdGH7rccJiq5DMdJFHPbK3nkVIGFZkzGA4JI81gujTKupYXyDbLO
oQmCYfgovwszPUtGH0SOXCyVI81DDunpvrvA8i+XZUN6p789qdUR8BJ6nq2UMzcR
gVZdVgmn7GgO28+GWHOnk+WDpbcnWS9+NFf3TE3DlYwFzZKWqPI3b0+DaxLeV8EG
kYAMXK39tCupuUMi8y+fmQWJJJYnX4DXlyZmrhZr/Y+vb9Sa7KkW10fWcg2R7Jn+
XVrczkpVRJ0LeGshBRpx2Lsyg5lAQDKxMpcxW9r2fHfSzyikD34nDIPh/1uqLsVI
D8mZhwkRCVglD7/3/2gVwFmgIP7szmNzd7eX+lwDH800Z0In1rr588nMHmpsuOY4
V63BUv1DOmxqvisF6k/7WHFib60CLeMLSfGmVarnwgi6gk2ooP+KNP2EDKHaLRAK
l3MhNZ0kW3mv/7XvSGW9XoyjGVQHslQJAvdQyXzvIZqpF0q05+34wJ+av4zU+3Kv
pFMr3aNN9jc09P9sxZDV4dvKLs1Pyl5jPY8VGnQBTC7geU32e69se70QxPgHFTf3
Mid4UgXDAErB3OsZO5MlOk9M1i4y0KyvNYwN4M6H6eSC5Um2aDD1prd703jshrSP
SyrBJzKeCBkLQ+GJD7Zxc++sI+SBXLGfQCzYNDrG9w/sFrKPVj9CG0X933WwtsGE
5zeyFy3/o4Z9LckQ0b2C8TxtUd2tKUxSUi5aYD5iNq5cAFVXt575DB5GaeItJjSB
zTEbd6lB3iYSFUJpxeQl6he+HgYXPrn3fNTTmL6JBwUjCrV7gGopelEAv8N06Ui2
4Pdyt0Ip30gs8FjXvIOMJp4PR1/UL9r+jNm8XBtwlwd0l8z/R71JGwZ2dfd3qPir
scpPTbzJIBITzBnsdWD78UyWTEAUIJlX62Nbr9HWjENgJwt8O2mRparVwHeeAZBh
mqidSOkS4h54gWNr6e05uLJ4JjzgNNYux8oOQFRMumNubW+ePnx/zgFUMThr+9a4
WsD7RrlFs81TDdgmu06EGDdExmhp8mOGYjgG7aT6hz33fkzB0qIraLHOSzzLsHao
qmIUZ11BcfL2vuuLHxxvttFgF7Tn2zbMEpsjCRJ48+P6BMXif6uNBJHXBvSY2Mmz
0vvFx+TgE4zi0F5BfjJVe/NMT8l4jKeTVUm0EOxgDL3Y7N4zNj5MqPORuJrVLWk1
1Nr+biGsKlKISrSZpxYBDTtFjiCGbMn9EssueKSwbNinaLWt2mZUq32/ytlKZ8E1
txZCiAjyX/q1SlL4h8TCAug9daHffbQnQ2L93VeqWRcF1yguX93ShSSRzPopx3z6
BAxTan1epn82dIikOw/hrTTgsp7R6EzZUXMMMYY6v1sbltOt0Yj3yE2u+TJ1AYj3
qJ4T/dqWUvEE5taaWZGxzgW/kTo3apU5Gn0GhCN1UC75ZUELw8wcVVnT9Rxj7zw7
CTZnf3tmxntihcdLLwQrSYZlsu1AxMRReH2ipLMpJMa5ym3b8+U77HRXRFFkthaQ
Fl08eq7X7IZfaPZ/HkKkw6M6/wovSFNVlABiZ/RdR8fLr3gbztvg1rwAZKWZ78GR
aJ/+cykD6mo0xJ2ife8kK9yQxRa65Bwy1sNRoxLYziSrc9fjde/WjNHU1q6sISFD
mB0cZv34OaV6V7uU38ZQeYpGoT1p0r3Ff43OwV19E1w9fkTayDujWpqIUjrugP8m
ES6LVaabV2wlyw0rdtGU7HE90YmvROudvYbOsWDlgDqdeQY/rErS5+pORvBsuOPr
l1I86dre7ztK/A1cXeHq5PRQ22BmFJYLzPwMBYvuvubseXNQiwqrvAT2WgYS/fX4
JbLEi7BPH9u3lrB6ioVUc10ZTcgBs1HzXLmnnvjgAAH33/A2dFohHtX8bWl/v51b
mOilL4x/D++L703eqU2u+TWP2Aq6JyuXMHTzv+jiYxH4xyE6E3oLgYOd62OxCBJd
6x8Tnej0h8cnM+FdRSlP7wELTADdd2MNCCHhV+0R59JIXoWdVeh/tA7vs12+io7Z
qVEFDwCmY1+QmyiTiYAjfyx3oCYP3QP/O0ZgLGjgu/Vr9+qxqHVfTAk4fzdifnip
pzSgT7NdUu5mdfHoEoaP5JHevwzSocjDQstgUVKLBOY12sLQn9fjBAyJT0aRYQGc
xBI+Eu6x+5ruyeBjMsXWZtKFZC12KzBi8nN9MRo2Lcw27qBromG+F7mFGcPUdgVW
XLksEeb3Q19yE1j7Uy9Ym20nZlN+c+ebH1yoI2NlUjMfKbvqiuUpVF3LXB8sEN4R
8kS1zglmJ5Qxw39G1w8Kv5ATLYGN5OHfHynK3+prCFygS2slwvkdl0ahtqAPqGJO
m96bdmhKSmNgwETUkhe7sJHY+AJgWXmm+LR7fUXX8qvBVxijYA/n48IVrbs6pOZo
ksnXSYC9kgzPrpFzXXnj6vAQGv68r2bsGsO97hFLV5S/rQjKwmLZjRPhFT5DORwW
YcfFM2WpwpWHrfETyUv1rnWrkt5owSBj9ee5KF0kOSM/7I+34f0L0uOpJwFb5eWj
RqFD8j8ePvGs0EFRnu1BT7mCDrmxIJ6pJkJmAlHL4zcINReiHzxhB7j+2+Cp78a0
bK1U+STW1mpM6KTyGUV5WPs6hVSQoI7kRSXIzedeER/rTGiJGRipM2PXVPxmFwyN
roWqAYOZtPIMZsgRiZTVYU5V6RrFYf215cYFKlhLqD1x0sAb0uNWoTmKkR23E1Xv
IfC8Ebv+27yMVC2OZQKBKmSeFiTbC2FUVDBlTgSAdshgcTBNFD2p6boOcfOv/VFm
TGaonwYiVTyrBbqq1ENg40vbX9KkOzctUuJwRzOzOnRZhPaw7udZ6CzpcejAtKbw
L9IbLKq+7ET3w8YqjLPyMAgjDZIg540ylbEyEnGQ+TN9xuTCzUQBSlA+/nKJR6dI
kayrfKBTvQvfRlILH8HrFO8/0WBvR1zQoinyyNY+Fk2MHy+6D76SFoITUuuYq7pU
vsmeQptsSeUmny7nsnBXloBtw7K2Zvx/EgFAtD1fR5tF1vkIOiIa9pp2jgUcZFl1
0F6oSQ3nkgxZ/dQ1D7wyzXQDpunlFv9gFPUMXwMxlG6vvqWcg3aFkaC+wa51v/QO
cIM0Q84MNoaSJCJPWByUZ1mbjgTFitToENGNnimwGLTTTJR/6NrSlqgEQOSJo5BP
FoohxOD8srwxbRGRtd1VUXjiLE2QrjIfuWCmmU5CxLKrLGKhGrp3YXKJ073yFEtt
fE0i2/f479FX1bb7SS3eXwhUl760sJ7SkY29OWtNHxQy7yD3NEiPlj6l4j55924R
skrm6iqIhTrTzn1Pbf5j7p3S+VKj1WB+VQreQHcMhVOqgrtPQ3MIuqMhZzSLEqC6
TUKJCOG1/6TeQrfxsWF3nD7C2gf0TVqpdgj7ZfFmvQiT9bfKWXAgRw+T43dpy8z6
KnQnChRMKnxlhMCT0ss5PcaczbDezJ7a2eqoEEPxwhXSe45d92MrJaKL7XBnVGl7
bPHu9XjXg8SAN4eBLmywouURwCHnC6wWb69V5tyvZzZcYexVXTbzpMOTGrgWsUdg
Nc9Okhl+FnAWt7ystPMqmRXdA42tiVA2VEfdn53f5c8iqle08VDuuLEjMhgjnbla
aciIOFk3oTta5MqXa5vhwdRnM3rglWUwW1vL6YE6duGsKKYW+j7wBaLkLKKpsSD4
AjgHu8AXHO83DwZHIvBgHUGTXTuLlS5h8fftZE0UKQusLbwMeOGob4IgJK3cQfVd
ZagJoEpJW0MhQ9WlLEL2QTHLgQTQxuZtrBs3QcM83qTiIwzzKv4UZcRK7iWYB5Ab
jZEqJYQ7sNr2ovfNM7JeWd0sIbFwTAV7uff5aRkC7aUbZHVwMkA1QZiPD2vNB34I
4X4ezYUEfJTm2pdDQ9nOlIdLJfhJl5ahpuPCrapRAVM5oFoNMEraUeFfGcMqKK1g
8JoYDjp1zE3Mbx67oq6WMAqZFhg4l9Cbl5pp/PDy0WJSxl2KI4xXDVbzY8o4pRX1
Q/Mbu0cPtqIM/4RGkFoOSbM1qW2kiNDF9BWQEzOW65qPO2dngaE1biw2Xg7hKKgs
4d4PB5x/ppbiae7AH9v151N/gBbFTwvqb9iOZlXQQg043Ca45VC7fNzin/ss6r3p
C+CSS5+R/5XrIqh2/29VKxWwTy2noxykgIH3Gp02MeuNBY04cHPPP1vkn7dSBbfk
WuX/GJ0wqyzTbJL1+66Sr4rx3AjrGeY4iDAcw16ys9bqnzujhGr1MKO+jtnHBf8a
s26uyON/ZhRmqQoQMNFKXNrFaQQlm4wiep/X1xi2M6JEq0xZ5oPUeg+q0bY+Sy3J
D+Mds8uy7aIMEiaO3iJiy50Iwhhj/9PEcgBS/ovUwVHSFfyXnhaWcUUvWWoV0Xtx
MkjW6/XGQyuIBtdHf4QrwfQhSDKouqacw3jsy757R7Cp08AcTtxhrYS9YJEYNidv
r7usxEU1vSb2NfNaVc21PpGSAL8cL774krWePcAfMqL4iLrgRztaKE/vKv33DY9f
Z8YigxL/+0r5J69r6nJw+pez9MYliw+02/mCMmUDLUAhZysGnaPB+HziThtGlotx
EzwS56strUSv3gZq5P0HO2hhbZ0ccXd/uAhvXlVgw43rTNzVqrPJkgar64N49yuL
0rOiMHo9EP+XPMQYNUjqHPhIgxc78aHduqarVnQAvvM=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J0SOBBvRg253DV2+sJw194cN0iP/yJqVCvEvghONYagXtXOK01UHH10EHzE+e5AG
edkkVsfWsf2hQySuDPSUj3tvoEq/+ifDTTaf+se4Nku/XACZQ4F5mXOuUt5PI1hP
7kYlYXOfrnd2AmHy+3ehf9PUIExFraD0+NVemdJbDO4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
rOlcEj4d2hk63M/9ePH0z9KI+HyCDXu5DhcrXtosX8DJ+W4Z6HgzACad6Ep9foot
oXMlCDH0vmWtbvi31qehL3A18n6W3fumBBNXfZzV4JZqDODKPj1oQUjRRIPrUj/Y
Dx6e9c0UDU/Mz5q1evn7YHHfC7XjagGZktnUNdULNKy9HoIRtwnTt9nVpewA4Aay
PwPJOyagvXBf8gapa2oxyfS9NvhKf7vTfPPWwN6KbNiLOstiUCzmFTZtB0xujAgP
VjNFS4gk6ctdlguRg/QWKkgDg+lripvy2UAx0SQBPzVxKWKWwJbTmwSI4torFXVR
WDYutPfIZd7AnFRUiDmIkCiIKfNdNVO2jU+p/3GlcpblQg9L2BzxJ4908KVN0yQI
EtVX/c41f9eLXvRCqe+AGRhGT+3GNT+i4BUZ6vZogi64sKRo0MEPooRjYYUHHyl/
qdDeEGeXrKCzvQw3GwtxS+ce8gwKmdxWQGeVrbIOlZlMinvE9TjNHEvT0ZFG5AEP
0Olq9BQ0aetUMy8YwLdDnD8sRiGmgPX0oeaDt5QwMYfvzdqQE4sExT2eIoHBVFSg
mt8MTPTb/qNu2YZfs8FR8ky4z9/F2ArhGwlHlQW5+OcLNkgH8SkWOjpNwPh5eDcl
5n6Qp5eRFWBYLDwt57idr3roo7Rdogici0cn7Y2ViZG8KhkoIXxK2tyzf/Uq4/Ug
D8lbms/0L0eDQJ92HS/hxEaXVsO+6JbCSVTxIQiyDRgUpUEomorxuDvuagkOuM0r
c7CP6UxaI7YuveF2H4VL/6JACX5ILcDw22UNTxLKaadYSpIq64ySJO1HvQ/wfD9J
pGs/E8d9Uw8P165Ycm1YDvP7kV4Dqg3OCwFxEPWqsmntiSsccDaoLPQ13muJAtZi
YNSjWDa2Dr2V/Og510A+1gkTgy9K7qn8kvZp4DEkTjzJU0OF3oTO8WVMsXnhXDp+
VILLpK181kc8/uXbDyN5KknAwYsSj47iP4Db8Xdul1DZ3sRMy8zf57/jdw/CLz2S
PPiXy/F8jQx+5waOBExlmym9RvArKlfeLTgDENHZQ9th7SWdOuqQ0i/KX38eMBj9
fJRmcpEwdWdI6wvuIYS99cNPFudN25Jw0f6hTCna0NkntsmzFo8EcH5R25eGypFV
ZynFVYKONJntI3rfMXdY9Zlb6+mH6zXciF+K/bHB7wQPaMq3jkaRgar1N0PxvD2W
72TSJPAYeKOeDLz4gQVtXc1bNQf3tJATc+LxDxou1dIDl8yJzk8c6OYkS9T/t79C
jfhQV2lNxirQAfcJuO6cf9i8dXOmpuWA+lbg02cYobtH0cj5rcLZWhUai3fxacEl
3eve4CsHRpJr/MEU/MAgWRtAitrN244n8XVhxXAgywEZJ4eM5vH20hI5N4lRBjfv
kYj98eehtYWAgkc05g9aYQgxX95f9JdzpFvRpHJIImXzkX9GRmmUHVq6Z0EAT8Oj
G6KlaV69CG9fN3y6l4nv/ykUdJaeB4crJa1nYckTIAFmpSN4Ux7eSyDs+Pem+5mG
GNT3aJO8rf69uZx7789/DXvDAp+SXcIP8x+5IVHGrnrOgtUvMO1m34AA6Ij3vEa9
Jfe9SSeNHv9DeRAJTwBj4gSajwNpQAbHz+bq08kGQSxPD45ym/3Thwdq7zw3aeB7
EYfMYqmv7fM22dv6XtP4KXDVRYTPEJJeyT8J0P6JwxetjIXM9JULsUemAVd+s7E7
MrGZ9OoRl/Hgb2NxvNK+e9Hdhb87aKg70kKwCJ6XhNJ01dwMcmPuKHlL/jwo22C4
RMgvJUdFo0e+jFfqjZJPg6JwZeHKFGcY6tfKgMAFkGsE12ld8HI9NekhHUjkvD/x
RFEJNjslNFkthErtmkEyKjwBFY5aV8Npq3K7XRUWI1notWfBngWLL4FbMbTvi1H+
KwyfkhXA3/NWIkEe7cl9z39DkHdibC6YD9aVRMEkLUrUuGVtOfvVBDluiHarWFaC
EKjpN9UY3NzMfzxRfh68nPhTO6kJ5bFTLr9PcJFjU1qO4GoL8LoHYF5izdZ3g7n2
NALo1zzcbivNDMkaBXdgmrme2FHpgNjNR6MX3p9VgwYgPcZdU9bIsaPU1t8GXTLB
ShQBPUMj4ae41+ncKfMmHdkZtLTuA8NEMAsmQ7oAxnzjcTjESZQhn45MbSEDPWbw
t0N+grF8FDiZ+9cR8Gr1knN3jRbQnFAvNW+0EtpTQEx9Ev4YDQXC+eRZSrf0pUiC
9SL28wdpHbFN9VNQRo0TKzR8/oXKxUdrAAHoTs1aEWdpPLCddXxn5cz7H/+ZMWEn
/sFG2DC8uCHmlPBezY8xBnpzKnpHdF4JR0kW8LcTKxTh2gyyRSP4SpABGxo/FvE7
b2ihVyGZM5Qa10aLIKSEnkf2INZSFnCnM1XOxMSiKapU7k8yVEHUE3g7dWNk4F2h
nK0Vjryq+Z6kTnTKHAuQf6JaOe+F//lyaWvfydjnlfYqEBUcezK+e7tw3U67vsrU
qpg3+12WwhwYFjf3ra1Q0hgG3jroGELvxXV1UNzVr/EajaWEvPBl+0Y6y8uHsJHN
tO1sGhzaYZXn3zijnNL+Jwk8ira6vLGz2BFH6GGAWNF5legy8IOl/GDsZ9LDCf0v
9TCtDHGxvm4qRJlykS32fGwHNeG9MEZza+1yjuOfwcOTsOmfJDVBu9aA6/c4uSeH
32g3WN2A9dFkv0fu5ACHHU4+KdtDdvqxE1wt5voMG0TlnwkBRv6k50NgbHGG7qqL
RMkCL0rqIwEK6WgAxVmRT5FcEbzbUyKSoMLrJNYTiHbvkVDrOfK0zMe+sAPgZAN0
I5EAIxlHzAlWHFdQOP48RMeqlLoBNUy6Jq+Rj9CrCMk0plSQZaTCAc6OFjU+Okj4
SDGnJLjhP/jPBBOTEJE99HgCGQ88nZt3LiT/QLsbxv7a5rZ9hiNEunDCDUExF+OZ
HUL08iOtWFIka9lPjsxVT0Ben3TMDExP6rqUU+grSghVoBlGAdozrwz71aNaOna/
qVE+bjM3CQBzhtCWDaUgUvWYoNX5HzLQ2Bkzke2V3KxC2szixU6E1RDrWdxlPNqn
HFxj98XUiSMmZ78e6w9b9iy88Me7KfmAvmveUFh70Ed+UNvay11VCLos2Pf50kt8
cHfILgI7DhKzzmK4Xb8pTP23uFhAYfxyh0AUUk61WfP2bkawZWfX2PqATw/Qfnks
oBqwSSxLoLlW2II4EyJrpjmDTEwjFHGmVKRFy1Uuank9DHL8Yi3BVwyqnSWzQVeY
Q4rVBkaxGV6pwoMyefCHrcnpSuzruJQrEx9LV3O5d/MLQOT1kV7QYszb5A9kERga
3rr7oNkvGiEionRxNb4o5eXvgrqwSB5kHIetCfdTp1dIuq4crWDELOXY38eKRAGA
ay3lDrEwpid+nKbQe06nLn1h5rRztowSYShTamYkNB+AsX8Zld7yu9Of2jMDIey5
ev8Za37bO639dMOcdgvnHeF9RW6Frs1LIESVLF34n/TOsydFueW5mf1AfPDXR8IL
R+4253/8OL6NHXU0yxv5gXkLRX8WQQt2ek+uw0+zyk23rT482cKcJAlFlJ7X6jCE
XKFFUYSIV9Xbo6my2QzAgp8f8oYRkrbTH+Kr/jvIU6RpNWh6ykkAYoijLeIdzJXA
df6tY/hZgelmHbsoy7ddX7Kn9AsjCzfPfJXKVsmL4yVSh/EJwqGBg5YSxr1rNXZ7
bvAJ/zRTaMrB64I5N7sTiZ62lS1SALRY/zkJfLAZFhwoNyW3nlmlRYVEYyL2SSN1
q9pKdPKERlaD3RVXhZ/28H+t/Ire/ZkW8e0VOHeB8+59UNn+tD7vhCEyeDgIdk+P
a1EnDXUmprzkST5PKwqlUhPhRXFTebnkl5ro8i+4lqOW2d0P1Qu1UXMX/rBAfyu9
5pSywHsSoXFAUbL7atwyxnfdsrkD0YlQOGbResjl5wjAq5iloMX+Zw8fHPo5rpQy
CQ9jhvcmrYgDZ33L2y3nA0T8ZHY1aDOFcKd11bxAxP3E45gshLfp3bCbVWKIwNEr
qU7Hrq25e6ZGgtMx9HqUgHCmd975E9frxwmwPj3deA5aCn6pCVLnmkspY5qqk1lB
OUeghGaX1c21rKm6r8gBILf5TAJxSx4puG0OPTANPAPJ+9NM8Sfn/VaXY3JiWccD
dsq9uXR2pvlrwNt9ACMHp6ibT3vM3YM1wtVg8sFiydvWcSvh83XSpWYuB5gA3FXf
7AOd9tfwI+1gOrWU7J8p+BSOg7KBblZomg8Vg2KEGjQ03jGJu/WqFJDNRuoAq45e
MqcKv+Rsozy0yNUbQaGWAzrW9rpyXaSY92MtE7ua0wsoptbCjk37e3y5GzgpedK1
mLhfbLgPaPS4bFZFaoUJbgljNYqK2mTAyZJwZV4vsGo9/+Ydm0tXgbkaCtRJrLAU
Aepc/duinecHiM+KfjLa6KM8db8xrcFn9b03eFEMGk45x0zOjy9o9FLtZb2UYlQw
OBcOGiq3IzJORXMjKgI2OSwF025OBxD6kEVcRdoGCNtxg3bE9trqPiKoby2X6CF/
K49YfPbA1ISS4WTPZjfI6Gc/l2pLNev6aMZNTb1mwodi1Mif5c6zVBPsJgqO+/bT
g1BFArB4fiI7Bri9Dg7cBXKJK1GXx+rFaz1bIr7rbMcSfW+cy0od4zxcZZpgV1IC
zXel2F2WRbnVyjpppVjneDndAw1RoiJ7XyZCQSNM+WXze0Tl9Qh+QHoVOwLnx1j7
kvX3g/XfyGDIHCuqTD3NgeIbzcy2jaqtCx0aq9q8Dd+EAGOEgzzgpGiWC6mqTO+i
VMTwh1FSQJnsX35MH4Q5k6DAUH6mhYveU888tk2QpdlPby1E2DJIrOgFXqxkvFiA
sNr0zj9EQ4QyMhr9HyDb8KZ0+rc4nCYxMuNr+LVsmBSMzZgxGAJY17h86hwBGMWw
386sZ4K2DgZ6+skwcQZCiXGXjak9yUznh5CZa0YoUMP7synopqvG1/4LjIRJczQ7
YDpSUKat+3x6Y7xYfvRHC/cV53C0hqoElCBFNZXNwVOn0Gcq94p6EcvC1R3YUF/b
gpZQX8qEme+sG3uhdR/GxRIFFO8n9EsilEzM9gix0p/tPu6a0kUnddt7OqE11fnj
BtePeaBskyw4Exk82cBnIID6QsS1oTz7LQX0hQjOVmDfYu8Sxhw37Q3ejqX89JO6
jLnI/sNxsMVXGWrMg4vcEDWc8C40YWrZRWgCY3T05rnmWqqZokn7v6ZWthG5Mori
Hj0t815CoZjJ4tYDgOXvAIyC1h0+/KWjwBqmpt7SUppqUzkAEfTSasHLBTN0xYtI
zXWuQjOnp5T/8z6mWPOY18FyQ8qsMLlhmpq0F8FVfVsxEwZjO/CPqEkoOGpbi19b
hDJaehE5FfIx3aaEFFYdZlOvmDYPBeHqNeVXcSPobG90M+XusQiDlJ8AGECLmASq
+ceo2QOgDEfj0XmIVgSWqZk85A06tAa6PLBsvZgrsfhPCOqQ0+KNYFUjhvcRct1q
hk7lm2B4QWqB5TDhNQI9DyT/zp3jj8dvbuJydt5mKWCmtNKJCv8lSHdUEW8jiVbC
lvYBajfuAPWsoPnbddyBaO+cdkCfyP3aXnC27CaZcp1+6wvxEWT1qOu8C26DwQIQ
ktSNtS+w57M/XZYCLpJJwgMI8SPZA8Nm8QnhI2AfZDPFSsEtkKLc5G45mzh0Fcoc
9iiyTOpCSGvVmcLFz/Cw4hm1cTxsWrWgsX6jU5mze8qksaFc0Ukl/iuS8jdzC5OM
3BuO4QRJqoUc49joefwcKgPzLl07TkFnPVyamX6M++65zXfL+aKwv98bQuTnRjUd
+VOSmtPCWonwxWfs+gqibSauEU+OJvnsrWtnukHhATryp2d7GrGsigegwDom3vnz
xDaO+E2X00JZY0JoUu/buL3PC70NN447vyxEt1QsBGhvIYZaJupKxX6JWnFrRrGQ
0e6sRlIDvwzE6tBQcLpYYLVrJuApLcU82pWFOQ8la2UIGpKr9e5gueHLuYM7URjZ
r/TKjgA/NfDJllBqRcdeY/g4JXJqQ+WflmiySRd4AqRB/2OCdw3h2yOGheItdAZF
QizLnILkaE/JI3UhYBTrEmN1Ch1rijPfg0TBoOsS1iHp5g94fGemm+jJtnVHH5x9
TC/Hx+vuC6DVC2fe2SAKp5iwvbgpNNCSGLPzggwP2R6CMyxSZFNHdqE/TbcJopmq
kgsdy2ui6rlFxxPGzKsnoRQwcaaN64iZRcD/kZjRtPTgB+h54jU96Z8x2CKpFrv5
VBQGuv1ezCzTGHXcZ687/ydlUxXYgGBxO/gfb8eSwzFHWwqPgEF+YZ5p8nzmpVXG
emISxnsUfCEwuu0uyfDm1H1ZtQn4gP4RX5ywBelcYbczfPq+lleP514CLLyuRNk4
GU0A6s0Jtrkoa1lIdB+8G0S2QDQBpJeDA+5c3AALPuOMe+hhd3QTG/s8v6a7ZFq/
Xxa/ZBd1F5XpKp6MLrtWIAeI9sjc7+i47AtF7VTkS/NDCtG88DGKIlNhtjiek4SB
6LpARqNwRxvdtqMWKxdvCVWEzGOAW0Q1BGnTQ+KwStdNzBCnxDEClhIMS3tieEPf
YFqB3L5uI8vyjmrkeP7FvLkDjOVHUfVWfXcJ4V0spn5KA7/ddD6jk7CupRJQK+y+
L+4/5hGvoC/TbYPa6Lhh9cl1FQitpnmlm7Me6PT4Ks0unOO8q7Rqy4C4xK97aLmH
FKhQaV7c29FBZbDTsPNxGTWD+Y2HkmorbLAolOz+aYhA+g2ZeAVle4fIDPLpLYkv
qMDWSuzYSAq6AqFlZYrvyRBeirMgU1qxXvcapeaM98jQulcTrchA5IGWpk43SF0F
OUcRUsUfQoY5oQUVqGvL2yD4t+8iB29aVyADT69D3NEzZNQHQ3rWDLhzcO25JDj8
Igv5+5LS/PaKhagQirT1MOfGROg4si4T9S+NhRWTZJLNARS+hylnaDN6qMi4jkGT
Gqgizu+LbJ5fTCy16y+ApCGkZg9oY+K8peru8Nxyek6f7PKGiHzD3mGmP+qrZurt
xlXWaTX63RqoaMIWuFKaW+05rHOuN5W6ofrgvh+iZS0zpWBEkrLKkFXLfWz/GB5x
yFztE1V/w4+f+MnMOxIYJt2xhFVdKqyrDHIuiDU9bpKZxDtrXQhHwitl4CAcLjjX
pPTQh8DJruv8S7O5lRPlrQPdUbo9xCsqkearMe+aCWd7iZgDdP3LeV+NbTRLP/Oq
fjyZCK7hxkfNB6h9XiJ1xvZEx5cSOsgNH4Dq3D3HMc0ezoGP4c4Dy9ICzLxgRvzY
Ermlyx10MNO/7D3WDBujlgYHEmXELaKK+X5HJpQvqLVQrsfaDbbQEy5RrShUbEKa
zvLoXOTe7SGqSeyzMNnW6MXsQYS5ipWHJRXjA0hLT2kbfoFBq0j+5fn9f026s4hc
NcDp8/CUV9IYhqlkKEu9zQ==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
H/p1VGuqPI8Jfl1zLBsMHIc37bWZCDgm+9HzB4l2sWBNHGPVJVpW7cyxFdL04XDb
2c6UJXouOkciQ1VQLVwR2TIinq2qOGHJIyKwwWMeiqUPWoCibpWBZqJEfWha9Stk
wOKH1sbls6u/SrHNc1uUOsJHvZcpfpa0AdEHSuo1n9Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 45200)
Y7p6thpkjmDgMaQtc04TV2R4djPVMshXGB/paUy3C3rza+HSRtYtCG6RIm9XGB8h
aL5bZI2ZeXPJ0C7iFlKZpaIRd1vFY7W0WjOinG0dCHp+UZ7ijHe2LQsbi7x7tYP5
ABBwP3HP/SR3gJkOOk0FDNPEclq1KGW2N4RxbtMPQBTome+KgUgqf20rzZCci1Yb
P592nzBEl8Kak0SvHWAUn56rhluPUGo+JrQt7+blUW6Zt99USeiiGv0UZoQLYFc5
OUATc5FBqWp8hapeAJIGYNQP4MCv/dRZLNPgOn7aOYmLMT4JznnmW1x/q0JSsWX8
uNR5Sd2te/rQ4jECG77t4Q2xO0z1Ohm33pZULGSjHtCyY1lwhsDeUmS6tyoppD0J
MluZcrdF8TpRWGatHjl7Yj3H9nLsp2EQLMTHMQgAtnTWEZFyV1NJW62YFz8rMDUx
3Vc8O6LG9QOwdntdcaGYpO1+OMWxWI23Yv5dj0k3cfbE/P5HTz5CnrjPMQNTLuUZ
wwwSOWK+FmjzUpHpRZw95i+j3HWNdqHE4LwKck4tQC8acMKUXCQeLr6WHTZX5+tX
o2xwCYTjU+s02XqhlZQRWJxLP30JkvfCpeE3FV1o0VJ/y/8mnQE71VAHmD24oJqh
Oe/GCqu0HY/mZF435+ZH+U/fU1hDbIFVKsQSMpA+4R2+41igaBsGj1s4bIhF90o0
RvJbQ8VUJTpixQnE77sRoyGKVr+5Bf0CQ3ZPUPIFCGX+Mx5jyQT4nVJgS2VeqtjU
6vhaT7OVnRbTWnx9yisyl55uDbyTRtw14966Qs+OClqu1lmY404w9iM2+pl/5qjz
Ult7Iu56ABOcd1sg6WreeUmAkCzgpqbC1JVHKqZhkyK7u3ZDnawDYU/vPZcaSLmN
i5AfNktLkn31tFUOEdVPUhH8AydOFfRLn/euZ8ScCPYFmezJ7BEp775B1l1PZ55M
Lhh0fHc8r0Ofa4nVhSjhmr+k0z68uyK1OnEqRYi9qFf9OM7R58Efb5WpE/5uKdi6
A0rJSS0QywSgAJn4OtyaCpbfWY1jl2cXZRlB4qTCWKkhfB861NrzgLvaUIv2Chcu
YRoVRd3hak4fbbb3MapxyPcMRR94lPujybu3NuHu/QMYXbW49JT44GpNS2/gJ5l6
BBOz7r84duXg6k8CoNo48NpkakWscOoVr68aZVhyU9cd0BGVJJ82NGkFpXKTjXuQ
lnllKblB1XZzl1oDMIp+KWInG8rI9UsLuyeX74dDDd/fwSdlGji1y9BScsXG8MBo
DkSNRVxqGz+oJAOJpyUieSuQ/Mob5r3N8gaVnk3EtEtTXiUnFyaRUx7O0DzLmKV4
eezLYGoYaEFeVjPuF58TWZ4y7zqhyGKA80iaWZ7PKwLkrZSXMLZaXDtBrjz7XUgA
AAJvSbj0tEOlVBTFJMUoqym3bSzogq6K3bIqAcLUlGKNsqeE44ylhwMsmffiNTZ0
G7RCqZ0r/KcJvIKm9p8KEGRpMPNej00BBEt/XO9IH0i7TnBkyXhThGPBh+3GQq9H
nJ+fAHZTADcm5TqyJNZH4qQbCaTP0EDojeCirn5bW9a51Qgd0wga6RoGv7OjSxL6
4voXectHbaUI/QkyuYS43ygy4PenpKCNhgj/5NDs1S3AGEVGOdBtJN/ShYVHZpt8
EYREJs6SGGel+hRo4fNTJyonZIA2zQSZ8MyMYnWI95k6eIE564wIA36LgwqxgJ2E
fduJHj7Aq7nQ/hX34EJ+j2HDdoF6Hmk+JEX+o6qyYru4Hsp1Q8K7mcgvbty/3aTb
J83Tn25qV+JkhFUCEBDDHosuNoDtKdB4rEV6vJTDwAtHZBNCNi6LPsaHClzbd5qG
3w5g5DLKFe3t9WHAXq2mdun4s9HFgr4RHc8I8xinBM8u6luG53hFJpQpl2B2ztSp
U+WI7MI9FfrzbzAI/i0tHsax4SYy2WUdyFVTp65g0Xz8vmasyq+vAVYvir30ESk1
blp71G0uI/QEfJxKRoPfZv5k/6eXH/YNmfoJGdnHNZOZRFwFVYWDm9AlEeroEZ8R
PjvZX22ZbhfkSBufZx9m7wwPm8gy2ZK0pbT0FoOGaGvuO0P1XymSYdgCbTEIUl6A
krgdXj2PJRJ9bD5y88ZK33LwdbAUN2ZSKLgjSdAtEe7QVzVEjxadiYyNjHYd/BLo
j01bJJ3g8vMuUKgiBkVnnzqFgMkmFz5iZA1HQmIlpXewJKGkzEAwFcNwDKz69YcS
AYsOEnYzwf28iX6Wod76Y1ISIPwiNmDx5E/QmmTS23Z3apbfdbyWvyUudR7db8mb
GNKVOZ5Ajo5n9ROouwWgC1M4iPZfpN5aZ5np+3CaKFzFtIH34bgYNqvrMd6nLmsa
rCeH2YtsRrxhkRu81bFgGk536IF+SpjF5/k3U8y80vVi/sjEey8+O7yi2TfqyzDt
5AUfv6KZyl1BdXlOZFRRZuf6o0tt4JdqcyWBcrJtwSQSbtX06Q9n1fDsXrGuoZC4
+Wm7ovRQtDbwylhkTcV7tPUqka4O/RbiurWP4ni+QX0QsS4VED7DQRZnENVHRgZf
+zZALh8tfPecFsF9Bq5q2ySJuMlWLEsNvYJG/cg4hCCdpo78Z1U+kkjerl/I5wew
Ov3RhbwJy1irQo/kFpICyeNA6awss/RwQMlry+s8LbbkU+08Cb7CvVxHQsAetKbw
zZ+52THR6M3UCQ1Qdlgqz92SZYqk1AzyE6PZSktxsSwW7PsAvF/ifYVtEAMq3l1k
7N07PqgohYIKqqe4xCS/10brgU2YYNiGOSofL+yegPr9W43IukaOmbs+f9iho7dj
pJ2EDDEYHq5LIwSC94jigtj2mTwE/arKxEUK3Lr0ejbGvU4hNikKeLONRtKA34uk
DMyl8GRPKEQV3P2bU1fvNlcgVvXiKtwkgdc+WLw12HSHMetjOrr0OlaouVU1jGYJ
Oc2t8Uh2B7sKqRFx9Z+/X6xHKSd005ue2pVQE314UDkMpH3yXv5RG9RNv0JTwfm5
pqc40nblueTkW0kBQ4uN4aqBNugYGJGRiHkxSMyAXG+kdAjJ1wE/TqNv1UFR9gys
rqI+MxDoMjK3P2hBxfgfxDojQvW/5BTzsQdrEyI9tTYsdYNUrFcVNI2D3btvpAhX
Uzp6ESj8Ftb7xL9i+LaEkWOvbKhnNpOyeUD/LzrASASj5Z/eTDTJFy9oWC8CeKhE
bOMG0oI/cLKBSUwyZqMZxG+vNbZ2ATe8edTg3YbtMnXrP49QNmPt4Rrg47Lgsujf
i9nCR2vgcPbXK0Y8E0YdoO8aWfF1pKxgHPv0ayRIlrwF7lLFrHL0fOAn/Knex+Nf
LL0yGYCKVec+h1Tc2ZugK2vFTmXLjb/xmpje2S6iF4upErLMCW5h5TT6Y59VUyLd
SsVJmTli9UxGVy9lnLhlqJueEBYXRsfnS8h/fR+ry4SvVAnVKJGVO2zYy4cEpkBv
eikuUrIbAieyKIc8p5TyATtEm02FA5Kzfio8LHbwoolj6TZg10VQxR8jUXRUwj9X
ZdvxpCRoVHVh0cRm/2IhewSM515EAgzml487xdnnnYbN88KEJsSH68HIMoDwsHID
5dk2xWSrdjg+ixAVkUbfrOwBl2d7oVoZp+iEh8+afOELKVdeDcBw6fPhXdgFprWf
y6aJCBX21xal5OkKfLkPN/+j86bW3xpX3vUIXGYeUyxH258NRoDKhssqKMRryglM
zr0cW1ynPGHDwH03/4F5L+oxccEp1+Zrn0I2vxhT+8JckV1ehQqs60q5oqrRMOOK
2Cy1EDVATZ9bwbLyUydNoJbAK0R5qrUTjqri3Rt4a0S2iYZSrlJNiZYSQbCLQunk
5xOzjhokygjth+BzcO2zDcwWd2NFc/SvCKM0SEu0VdWW3IgGnwFmy28zyS2SDZqJ
7g+m2dRrBc9mksz58Y9BKo53RWmb9phe0SirY5lKoPiNRjzmzFvaSOIQ876d2j+8
uygihgjXP6/6eYZ8kFXFXlSpETDEH00wPFDNa/GrqG6ezbz60UWpighkbEsYKxKM
BBF+j5cvYv3zVRDtHGMWWFgwMsADTcO4n3zN6c91qmKQf8Wy7TFfl1y1LCvgCCKQ
wldtNaYEnDF96baaws8Mx/Z7I13lBgrmmZHra33JX6eRX12Z2iv/w5uNlrkBaRnL
xQQyI7oKX+Vzknme1EnENZ/umWdUPXIxehjFc5JCvphu0e/p9s0v8o6vso0xSXbZ
llWnaqTJ7M7pWsS4+q0tGYiG/WZLtBH2lm2CycSp1YP/fJNTjEUaOsoUsNbytoGQ
9diXY00QPUntww3+LKoRHgIElAI9v03fMDM5GIjUznrG61st4EbW4ZCOODH2yGgo
w14Ru9ybNFkwUmXyMaAhsYx/BceVHaoZLk9t08hmX2yMOTwkQuUjN7/zOGqrw4QE
OE53Th+N+731yoNZpnXYMNBHh/ynYuAiseG2Nw15cvFTWs6SKVXmfoB6/pZfGYjm
DBJrAlbT/2TlvWEZS9jqWc7+1zdSQRxyGwehQ61a35kDYRBtY5TwjJhOcuXOtxKp
/Vji7PTlg4QwvY2pOKtFmwRcZRLcF5X1rp8EL0/oCHMx141MFBoWAiphWNh8lSK6
mElLs8wp4pM1PzO1saXYLcIOgdiD4ItGFMhpseI1EwLYoLLe3lWPiVa3X6prDe3D
dxpKkzIqAbnDYai5tmQu6S5rAqMo5bc2HwL0GKPFnAgEWmYlZlGV+QCWe/usCpHY
kW263H3LthXKN6QLTpPnDmPDWRFFDG6dDlGvSNJfttZDL502RRK0acrMQSmnGyJP
oYiVm57A9m4RMSC/qclbmw4J/1cxhbHj2/9vgEkZm9JPIRQM6HqFdI8RBBtMpCMY
G5XY0mwqb3P9w3ebLqFVCQqda/Q6X6Qkssb7LBuiOIeMCd5afPirnPm47qBv87+L
eQXynfQl0vhl41iMvVVcwbSZLMT7rAxuA+iV9rGx0iMIqApKrzp4b0k+ZwtkXOtc
s+U+RbdkDuUTSLQHzWT9ar/fEnP19y1jvVaMdlMFGRBx1xPX+vMkIqrsqQBRUDAa
XQmEK/b4RbrCCOk8bX8X9OUyLGon4Ilk6VDgKsZEJlaawhz7/EUWlSrPH+c9UQ/1
RxbiO9Ntu60Z+albt7Qk7/TSzcDBq3/9X15nLXSUVszgs7fMvbmjoYppez+jV4e3
Ju0qxXUokDtqR90Gnf3eRNLzrOibTyIdZzT776SGINVze7184qPN+Ej1LAqG8PEo
BiglXGPE759yG0uoreEyllhf9mttSCXtXfs5H8Bs4SQYy0w6qmzifzWlajun8crU
A5K4aC90/6ZwRJUVCIphlDCpXRAHsj6dL2LVX7WlD9Yt78slVCgEMBtVYF8R3avS
rqSAfLjXGsls3KqMToo4DygRVo0WzzTNEzKIQNsg1PMLkG0n0AE5lpMJFwaV3/WO
6p2qlSBADey3hIf96Rn/wun4woevn6Ui5ESwlm4YdqPXJ20UKa1njm1SyRv4X7XP
Tjqb0cf4KVM+6drL7BPawb7DDS4l8v+Soyj070iRAmGf/+F1VEwEQFPN05D6R8hT
flyS7qYL3rLfuK9HKIVYitC1mqX7dJGKhJ77zvLbRBS4lVT90KE0zlJ4adGSilEb
3hSZa53yK6Q1ODk8R+S/gC/fV1sWFaXo8Xglalz+/v+iOz0EgVDZD0zqXQZtOCMk
X9ng5OCGhwOdHajs9Tk+57K0poZ+wdAam43rrpfWWfVBNYyHZFYdUYFiev3X2gBt
bqeKhG/pJzvHyKSFlK+rkG7EKIkS8TqIYeYd+Ops8lO1YkfntVNHkdDzjCp6YRuk
aZ7v6f6Z0HzmjHbyNXsMBxtwSApjtMjMJxZ7SGMd4rLoyF1XUwUKUF7nq5q2FKUr
nnTbxe4U7AYpAvMKZhaD7cdicMXzseKkmOZ7vXF7YruNUr2QpsLWiJczFzERz6TF
tYJ7AvenjFKtgu6Q8UIDE4X7KhVOH8L2cSD5ltCcaKySbioVA/c5+tLB/e2qMiTg
XOVQxB6pCr0lYgpxbG4vORzqStz2h7DQuAjaXcb/VmqxIS4qS4TiufR7ONlkPCrE
TB0mcgSKhr8fVOEGWZXhiZl6wLB15QtwWB1owCdmL8/PSX7ZgKRwcqjbG2vCZ1BB
0wEvPrwyTPCZJbz0TO9cXdXT5/Rp4aukGc7OTM7kGKi0uhA8eSSZBnBD4nwgYE5g
ACEKwlrUw+CELgcM8XBxdKjVXgCAVKfFKQaryzVG0uiqs4c+BeS0ey4PPgDN3nIL
B5pt9GfGupEWFORWJFMqkJfee/STwpRNUEdUAC4uz0dgmr2rju0P9zUBCuSegIyJ
HQN/+CbJxcu28zgA+W26t34nlC1i2d+e6JADwYkuTuYTh7ab+x1pR96RzHs4Y20n
RRvtMxBHNRFBU5Zub7xlbpz2WUTgy3rjY9pG7K7A/o6851nJBJiIgMa3moEgmw81
2KwcNziIX2Dxeg9SPvy9T3qqFeXUz25++YN+IsCuHTBp0I0bFT1HF+YyYm/KTkjP
wBMGoD8kySzFPQMQF2mgdD/iBHSwkQxsm3N5EyfMqLPPyt4ZEsa3UR1R7Lhizn/K
JE+C8Ds1QxrbjKvdAJKpyzf2ycZu/k1A3Be58rDKoLVoyvqvV8OIeJ+SoTni2nuQ
GtC/6qjEM1cI+S/RjGBsFg3TRBj3cRvonqHG7B2L4vaIv5A3FyDOsQH1NgDcq0xQ
0H87bJBNCUauBInNeit88+I28DBY+5uMFzcbqs8uhFGNXD46gvdQFiRMgsnEeOjf
zRBMCJsnzv/E5ykHMX6aU7W/6U20rdruI5MUHS78qhBxyJEVA407grf5zaYwfZ8W
bsgESt5SLAHOtiZVn30K/07EqFe0aGFwHsqlqD+oO+4uRwwsYnlaqSFJk9toa4SP
he5aRahGTxqxWnIYvM3sEwH7HYJo5keCSFBN45YTclYcLlGLdaokMiuSRqLBYOHL
sumsqFQlcVAZqEGhwK2a0hzY4dQNn2vkHgha9ou+gSe/PS1Y8+WTVNcN40Q85hLM
k968T6ep7vfzYVvjFwfvmJ53LkBCpUCiRSlV+7h8it/6pDTYdXsd3HSx20+B0UOT
QlYvsNrP4jHnEUdTracDNx4zRFLN1GpbY8ZU6vj9akM46IM8QndmWJhkveooCkXj
Xh4/icWZqrSFPjAeUHfbU0vvj/YDZ2qndG0DjMrEI9jY6Di00H6O+TMThDLD6vVS
AZPziGG7pSG/IioN5Xra43ErvYXWOOoDSqEnLZpaou7Obaj7ruaLSy+JYexMHNSw
NZU1rnUesISLk1iHG0UhuqbRP/P2PFjPtguLw4u40KbKSNLu2DsG0u5mtB5pMT3N
A+HnchRnLj7b/5s2IBVQqvzW6e6TBe4RAplN/Y4DDZrYAPmBDBhaamzHFRaglTQQ
Om4sDfyQQOqwUdwSzxh8mggK5kWi6UduB568Skl8i6BxMIQUMWDqU1rf43oetbKV
tWXjC9fG1eyLDNwkBoNpaKLWd9FDMQEGdbpo0dWYnwJIBP34KjqnNhv90jhbpeO0
tuCIeaKWdlNyrO+6j1ekzhNHIaMoB9DOe6N1ZlGiTLA1QofCg58vjatGwWrjeiKM
yFHT3H8zj69Ws/pXT9R3zMselPeaQusl+SGD6vD2RiYU7+aGpknToGE6JGrLlOO7
N+tPo+5pULcP3dgXuOpfJpM6Qk2K3a+AbTNnnIcSzvZX7vuNz5iQd85RFv040yAo
gJcJoz0cOfxWcqKLPOW7pMAWNOMArl76EZrCMvfuO5IaessA1HbRmDXhdF1NSmiH
hYRM5AvrqPMHVc92mFS9imVET3fNmKVZ3LnEV/wJMbAF9BarAZEZ8hs/UnJu1rin
+3EzUdPSvteoIGrgI+M2sVEGvYEo+j1TsIiku4Ggczn7y8chbCtedCqxYBV5rCQQ
AdvP7HyQg4Rm526o/OJOSWZ3T/aWxhubknMilipa6mVjEESsnCWaHDNoF+nY7eh2
66thW2ZUp3se/Cl7PD6Y229ew6D/6/MYXAPfL3taR091MadNwiaNcWFqYMWNh+Ii
N9PEfYHkzm3yoISvsIAvuiDH5Z6m6IFNTU9RCs2RjNXg5cFKvJmd8OLmsEU8MQsf
onBwXyBkCaGI6vPgDa/wxItV4fYBmd5p9vyUNK8ODkxyNQz/x/APeNT35/3IUTqR
dOsbw84qqpgSo1ZVsnrEAVwj88ekmB72J9nv7Km8lrae1eneYBXS328cB6zsAe0e
50fdfazSKAG+myEhuO+D4//CCgUbY8t/VHUNUR9yeEIRUP9S1sHmDjFQ9YKk7A4P
Z29c/xK+HuJkoyRzcuBiDw81wy9gIiYj5o3by+qAoeysFa6JCZJhsXciLBL5vOot
3wqlFzzTeZU1V45eTzco3M/hzDaoCbi8ccSRXpKV1laIo7oaJGDdHqFlgK7z9F9l
Zugxli/26Z4q2xUQiKi3X/DrSVYa0lzUbV7IkLAL5ThlmJ6BXIVKHJuIE42GVPna
wWcPVqt/RxA0VUxYeBw+i9b5AlTVL5EYA8wzS3Sho3w9OrmusrXLEIl52wRQZIWW
j7viZum0VPmCTrOf8KPamt6MjZYt6jq0jBjTrXjucnoJ8vrJrGHpBBRRxW1CXkyZ
nCGfe/r9L+T0ZNyAYnwbiTf93jr1u9XjepCF73sj1wbacCu8f7KlzY6btpkEJhJo
dXnJ+Q75k2qNhhfXvCJaIk2ozsw1DE2RKJxeSLljcxZ/agFuQzvpzYBn7Qnv5fqr
wA+LeNZUPBepnsAhsS8xzDDd/dej61behWVL6hOWLWUB/6T11qQZZ7tOwTWeUbYK
Tk9I4M2rtWM2JChgNkx1Krlk4nwMl9zzwBb1RLGCiteVjT6Jv160yfwWj5ujeRmi
Ei3o0K9Mwv0zejFWCbuBua2TFJnGpXwglRwdkexazlINhquTY7HfxF+SM01rsRMA
9TLY8jaYkEKnOT1+/35CF5zksekzHu43atqVXtLWFCevKAqaZFG2VkmLKJzDt0xs
/yb+OavXFo00w1twMDi9g1E/ovj3rBschPLeBgEt3MtSXmCtffdVQy4PwNIa4/Wx
L4D4Ro7YuU7xMiKDk9/uJ4Qk4MQwNW2Yo6eEln0p5DxdZQDv6T7skqGhalc3vn1d
RLgf76R4+GS0GM5LxJSff8AiaxbTkQtlfDBMh9Wtx9sZr9WuP+EmTuzOcZ3tGCHM
KcrqR9B9R69E+v+AQUeA/Mnt5Yd417nycTeY+afe6ZV+z5iamq57moRsg7dNGtw1
bKaWFTz3fuCIlHdn9QSley/hCzxPCL/DkYsbnCdJpr+NMBqvljAUYFv5ND27adcO
in8MRjTzhfku711Is9bFyU5T5VbDzq3CxivP2+hsSF38TW+R9S9LbCJkrnRwdzWP
EACrf6wZGbFRFQfV0rRR3gN931SBEW/A+VAC3Kc4CnQ43nKbt8D7u2jLwnQGwYjJ
81Yqc4yK07VKphIKbroJtmgnfR+FFBdMOjcwpC/qqow2zlQNpGHzaP7tOIp/bUGV
UarpDCSLhl2UN20A5U7MBIFI+PXWdAr6EncbGbFLXrcmY94wljxpSgc8nPF/84g/
IxaJHXp5dGN4T+9zSMByvh+piY10Z3ktjt9Sv/9ir1sCzkd8IDBXfY1i8JzOwJEj
BpLfXunAzg1OLtMzy3RK1z7JWg7SC67kmBAotJflrI3UKoqib0TT6MHC9hUykKNM
A83G18XXbkKxMQ7r2ZIpZx7yewqUYMNE4wBWE08HbmdwoQvSd0NUWccH4mBpRCbG
9np+9rvZklrK2MIhl7TMJ47WUqkH/S6xfT1uRUGJLOih+Zei2xObiFm9mnJoNgei
B5klOfU7Xg3MDFQTM71jP/vAACqmnt4oL4j6PyYl3AO64YlacmwWZe2mDzvDhO2p
+BW62RRfTHdx0HevncdAhyg7lw+zgOe3sOe3CBwrGqQWLr7eo0xm7vy56xEstq77
3GapsBHprS3K+Dmg2ZL9cdjxtHgWJLzh2oZtNqtRsI4vatJ1TC52Md6F5pgYZ4Bi
rKntichhwmVgBnaZWSUmhBEeSvOKuOeUpzN4/G08QXKLO2NexUqxDjdlpGtb3J2Q
LuWLsBhQNzaBf6gwTw/LdPk1dx89dlF+Z37HTlzCc4hQecIreCj7qBEHnMSVFhMO
F/RLg5gmX/JKvNgWQqZAHDIeS4Mf/j3+TnChlBcHlHTdTRd/nKjkOeAVhjH25Nps
1LRtfSM6j0o8/6dok+kiv0LsJDIayFsqx2Ei9lCP2gDR/1lVpPqshRJzlrtnsGmp
/SB0hXgrOXdTn/Zr93Vxv3QUpqzCuGS6CI/oP+4+YgTr7qLrNKJb+HkNbuhtTZH3
Dzz9RNpzW5jgLzVrGVSDfOtavfpySWAz5c0AppIxTaChtwmFisI+6AVqPGzQzi+e
fiDeCIFuKJfBjrTNbBWcVeb75jKF0rSQHnTbAqdbuR1ErSNcsUOFjdqGx6mVCFUm
gV2GjfsDkdPttGA4uoTb1rkojQilJFjkJ6VmIeDm6S9IBwIQPKwhhp3M5sD7Bxct
QWJtLv4Rr3y1B+tnyBP218ViU6fKVFQoSDJ4EvGMFvk450QAQG1qYmQCgDCi1kVA
Xg4wdyb7jK14zU5zFDnf8H8gr7J4a3iPSKgUp5tMV4Un1ZiHOHbf5/3hYuyBiaGC
mRDB0xcahHRoBUneCAVLkODwnNb6HarwD62oWj+dbe6M6gsqb30ZyZlk26RF2hqB
tor8o4Qi37nU5aY5BwSOMbFNyYHH9jeRn2trFhVwfIuD/zxSk17koJuTrjtY9ofW
Cy6l00lE+BlhJEyN1b0ShdRVfaYnWn5FRSbZhc2r2jfHdcps7Yb/p4FvqLI355ye
iCYzf9359eYEgcYLcW5Sy+//MMf0dX3TSEdSJosJVdALg00PsXD/1vXJypCDpysi
70CVPYVBnjDi/2pj1YqojbbPYBbPv0u3TK29PnDycUL20vuNaINm99I7grjzpvnx
GGSgOTnjVFqKOC2pxZqMl8GbNeUyFWo8yHuQUioIfW5H3lnzcJ5qIufscjpw/3Ua
SFiB+JW930Td9p1S7kPczGfu6CeVVuRLNIhmMycgvX5NoU+xjjc10R2zIKHHbrUQ
Mx6TulCw54EvISLcSZJRX5u45KlbioGXDuGHTIqpUSWIZV2KfyPA49Cye8WmhZrk
yDu3+kloJbEslOtqHRWHBMwFTFBs1zUj2VIidpJW6LxBCUWUephVwM5E/0BujDfe
AkzQp9NyKvxXkkDq2obL1xK6EkB46+hXEqjSaLi99IF4PxBxuM1nNiQSW/gti2+M
tY428s8EziFpFmF1HRkFVNQ5T821Q77MLf0223kxfi0a85K1QJ/heE6w/7NRVsgb
Mq6mIxOAK9+DW5AGnBEvHlmAdnomGk+H+3uNYr3ACn0eIVI262ZLvhY8+OL5SVfJ
ly0L8dgwHWExo7bLxrqr/I0zoa3vga1wfAeWFIDix1B44+/pSxf8F8/+dPpeJYKV
uvZ6vhJoh6b3MVMpact0OASsqbYcSb1lXGnxftgN3V7598yJF6//MlFJCFpf1wXf
EQ52tW+I3shHR1YP505I34cIedmYkb4D99+78BWaqn0FPbhORuvegiuO8tHEv2xc
mwm5kupyeGg5MlSDYGSlgNQctGKv186nEr0Kef+dJkl7lNGyB6ADouKrP//r/BRb
0V1DrJocqX9FmfHF+UU//MIs5uBWRDwsfqUhj5oc+IpT51jozNYiWask1jLX9ONZ
Z7IBtvZDfhH4VKaKxho+IqmC06cueKVTSPVFRfhwA61s1U3f4yRbfFpuvcJvPlWI
+fOJGbvkZ/ShH00GQOB9UJcCdPs+JBsJx+clxlrGJAAyZuiSuxZuKhcJBOpmUgNa
9SuHJgH/SfQ7FIM2DRqrYd08qrRArwFuTO1tficnPdWr/1ITVpEtxL48qnQ2DrOj
KUJkVc9gIOSTRz80dF1Urx9DktY3oBM1bt2Tp2gv97pMLlY5xx2/xMIbTNOtwD1u
GmKnTC8viF41xMv9GqL/gO7IxX7DUNFQJOLs8noXlgjvIWpcY3Rt8/WIClP8bwT5
0VYBtR6ynwdHh+Km+NmNaj81e76IE3dCJA9rAdZBhntWXhkzvw47NHU2t4cWzwZ+
lgZEt/hjYZ7cR7y3EUH4JCJiHgYJdLXRq238zIGH0GzplqtsjM39uP2GpveC+gLi
4JP9M2Nx7FlLBDwQ5PIEf4ZGiPCa/dG5YdxXZpdrjd//peQiKgA4RR7tATveimtn
kLuGJMnimsluHvCF9Ah2oDbLwbC9M6qgT4j1WCeSnLmqdZohbWRny01IOOcbCn89
HcCpnwxvy93w9fFnBCCVlxDwXAfBoPrXJabTFD7SqcCcpt3mTtl8SHHZucev9zwc
Y18CFUpEscfK+hMWYiu+hPo2pigzemKbnMFPEgoTpA7n7xL1Kx3Tmu8CMRWyNK22
/o9aIdARxB5rXTeyk/1KIiLlJEPweqS5LTEEAlVI4AUAxquQIeeh6ZAAnfPGpsyS
Mg/hJuCbqbno8xwFpfW4a3q40Bii7jrrJ9y+8wvumiQL1BdiPM2g3JkczwEmNc0X
eSld3Rbt7729zaRhu0zK85GaDpzyNpswS0opGGINg4PCeWptFJgoVsT8vovtdHSv
upKwLHdmWqhyqPhmNRQ447Tx6T8YdX9nya3MLGfwKM4NYy2L/9CZZStYbHSeEmrl
t3u/mTWliS4kwZBy0BGJQRDocElKhb6cg8tirhEGy0Uc5KuyyJwvRDLJpSBjvBwe
bm6gaX4JVxuBs47GamcqvuILHemdiA2wbxzYnWjcJg4sz4t362WCoZVkl51wXdVW
Folmxh7gouM4gQymLscBAiOfDXT1hgEOQM8s/rjNSVEgIVOAPvHXSiiZifpW0VwA
Snd2YxnEnMvrdgIdEbQ4rIdBYzdobyhmHUv0u2y3/Iegnwhd6Vm2mEcQocrSqsvd
d8R48YzUbqc88YUSxqY7W1gy0VNJxjql7km9gkgIAXBX1tcMQQRiYTGbpqTWs0m6
mK6Wc/VDEAYxWoGATc9ypY52ylPzhqrYnOm/R4X0zwszDEOPp1eTyRJYxcOag4G+
4jxDy7CsNVCLyQz6yqxROaSxzI5G5HLGej3eY9zFatHUY8H+cUnuuTExc+Nu7UOu
srJGNk8FHom07uO3JoLa/IYUUAi0TDSbRsy4lBEXV4zvL7DsORSEbVMnPewHvvli
Ocqo1fsQxRIgR4U3lweN4UuH7tbdDtHbqqn1rcvLgruAXYEO4sGHcF42d/fP80cr
zjBVs+uoXznTDtYpCRbQHQMst0ytKytQ3U6YmgqlimhIBkts8C4TiFHaPG8fWzJD
SqhDdivSKSKTRzQ2Nr9ZdK9I2GQfdWGiAfCBXpiqmJF8M53emBG1NclYeQ9W4XZE
BIdLxk7ZkSGC9sSsN89iXAK1m8MYNyxneVIFpzGJ2fqANi1wpPcvtSKLJBS33xMn
1FYkR7jG6ZlPH5ATpYWT4phFh+XkuY5xZdgyZ00ZoFdqGaVlgSeHVp9lg+Be9lOU
VpTf6KQRxEagjmAwxtu7KctTsDu+tnNCebwIBrft1i4DkhhiySu8sRO8YPzJtPix
Th1/fW92RCYmZ1OjP7wVx0prQiUtUGr2geRsym8sa14j6oc6+1Xrij90AQN+3j/Y
0J4lDyQxjey4KJ/ej1ahtOQJmUvsQdKAlVt16FTcklLqZCRR7wMoPBv2bSRoQ9/6
Z0I0oAxiLcvVGYP/Pr1+DShxTaCK6U576qoVCu1LqhC05Qfg1uzPfKcGQW/EGzRc
OXDLzGBr4CJZiL6F0MH5TdfwEqvFaS3Yw0HG7EmdTFHhUqD0ExI3/PSpsftI7ESg
gaVx/rwpRODA9gtr4urrWsuc0Y+opxjE3teUPD86XNCpUR5sN3QsBdXw6EnBqzAg
dpmw3O5bgmo6vScMeTw8Ynb9TUuDv1JWn8Rofuyrw6wqxmAq/0VUwNWsxfjXGPKu
TNKgFRHv90EExzV4K5aJdRdlMxp8s5h7cyziTxhuY+fW3PjFBY2I4vnVWh3P/Uci
l7tSnm8p8JjS5zWGtCLcY/KCkptPzBXnpvUU/N8+x6KhjAVylh21ss4dttbrjBjt
PXSUumPu/v1NnNFKZV/ItlrFBKfvU4eC7bWRo/UmEYoaC1xvIJArqZ7Kz/yglovP
RQjWQYW4AQsLVi9OM8oBv2PsplU4jV6GI/gwJnJeB0thnppE1u3+zEuB27cvmKoi
WMrz3tcsyJEUWMO9ZqGeQO4767juCD3jL6IKktBY00hwNsS7y94ElNR6SP9ruURn
Wz48sVPnYO/vRytKNOmdq/01tkjKj/A6pI7UMWhMKJJUQS8Bo7UHTYZv+qAnxCqT
7s63EIGWUnuUAGlXJ9vjYkACDBg6VkoebQ+J2jKU1TXxlBWVtbOgGtrslOx4Wr8F
ehzGo8fNlWITGkzhXgf2EukuxSJ5IgUf0xMdMJAzp3gB3zJ2xaQaXsguPIqw+OLt
RR+aGFVE2TrQzbGbCFHAgZM/Wd/EGbz9IdgeDhhgPw1I96fyGD0d9RxPA0JZSlDP
zaSqItcbO3pv45e8aImsSDYNoY6LVOARiSeZhWVddemQxtSFNx5QsSulE95SO7W1
qJdc0PumDxKH+wILcZhNSzo6+DojtysKECkToJF6yjDySEFCglx7oLjehv2PLc6q
CgrxJF64Xw3XOEIinW2DmlHUztLwsONpA7TVFU+usLrZt0f/fXtWYPmO7AqRUbDh
ptSPK5e/k3fTs2oBmbbfEeJqO8LVAjCaJYTrdZ3XvDs6q4t8p9HUEyeDJNyLl4MU
U01nD7PTChNEVzHsvnuMOH1cEwXdJOdbF8Q1KqQUiM/eYxUm32WUqqE+5Z5ivABW
iEZeTX/U+KnXhayObtOFML1uVZ6i5CijkLibOmnSTrsnk+mcvY9nuCBqujIQu20+
toc517Z9kY7aAT8KC88tprxaGBV3NSK5NQK4QMKPQDeYsWfuo1xPyXL2GBqK/bvU
aY6q9CIdGTkQj/uKlBE5iup2ne6dak/EU9jvGdCd8mPR+sAC4LLQfzSqhT5JhC15
0P+yzYU3c3UVoA8yVM/IC/6xorOIZOninlDnlGV6A+CL6Wt5x/nlqyAUzF93+A0R
aM8QQA5fuQwTzYgHHG7eM0wbGrrkA0laxb6zqwaLccvPNII2IKImbH2pCiVjbD6t
f/HXoy1MpDbEHgC4es6Qs5eyeYekFA4yZJu/6XPxiME/sY2kOVNCq8W9YBwMP2og
sdVlAIuNXdqLITticIEw+8Bzo9tCQMm6jGAuXJZ9tHMfuPQJKUiHWDr4c1Bmyxp+
yZy3d32YmxSzgc0pyDqg772ZQYUBf3gWzg6qM2vGB5zdsAuWn+VzGqddJ1PZQ/iq
rZIBBA1fX5VeSusuLmN9c4TqRBLdHli4u2L+VNsiYhYAQGZEMMWoesQE2qXtw962
YOHz2kYoc8QSapbO79Ff5h39Lf991TBD2HXWo1VgvaZVkRs4DK8pwHv19RCuY4sW
uD+3MyR9eoBTK3dmzoIWdlaIQE4/HrGzza8C9NYXYSu1J+Fmi2+QjkYJuPsU40qn
FlI4dKcp+Yex0xMOIXfjjKlnSPD3Vg9Xhxz7XujpDtJJvje6DlDOsN4+KqcUwoJB
BF8YP7w42OOAPRPk5Cn9vihOAC+e60EkrVY1NFce/9sk7zkoii1KV2pXEtXkl6pI
rxrrkUORWpx50Ja7RUHr+/bHlM8NU9RpUkCC+WuY9JJthafdwSNCuXarjQR3pnPP
VTVpx5IuN33JwpWCcief8lookmrbgRULEIAUwsSmv7xnZC2HJ1dWogLjEIufsPtP
URky2ZxcAVjQP9BnforgfeHF+r7RzWgqdlQo5ow0MFZAFVD4/is3qKBgNoYWkuOU
VMC1krv8mpSTTPYKzJgv47I7WjGKg+ABNvVDX0aZoBP2xQQe5fhAf5cCjPX4HbH7
GxILvGZxwUTClBscKtd7wuMin3+8hkdoLLa4lsHSE3VoBj8F/E0BkmLYdaHexCKf
3Rn/XtSEfgMAhDIZXfehTs77+1JAHfAxFzOam5evepdlX8gqD6Bq8W+pcWa0utF2
y0TIRU73I9tGMv3jUemnwgt7Hm/QIhg7lprFcZ4X48fQuGjpCCyeuvWdDc6aLGor
6RGjMmdodMx7bK51gpmQ7NsrCLmqlWUuIXgCMKjttqxtTYSPMHlfWYsjDSYvks8k
6SBN2zp7B7XTvxUtvVwA+uLp7bPmVAjMaBTRAW/jWi8agMn0bUxJmufzuXY+m/Tc
+8TDAwC4YQ5tLekAaSbjPJnbGlzUJ2mRZfiGlaAr+zuQg67jyzWYaFZhU6+fQ+mj
0YhMC5eiV9ScrFlEbNE3P7pjjz0KZ0xz72rLOoi1nLH/nYJWvsWOPnQmkSXKRzgt
wrBAnoiXjC8jGzX7c1Xne8gyvzTMFMHHx2ylYbxruS83twvzVL3JWk4Y8tUQ2LMQ
5U29Uc74WjS1N2wErRuGpvbGmmH1TuD0ExubrLqDjTj+NlmhKvVjHGbtjElwTjpN
PM5x+CSBOz7RwvAD/XST91yu8Qb3eWocxybFT2GYobYI3IJGgju/FI9V3Tl6qpW9
7lo6+eSj2fX3gTcDMPGbRSUfkTgaFczs+GSp/DYF8IatZXTws8hwmfEf+GLVv2uq
ExBjtHR8H+L7jsN572FqtZRegc70YVfjAXFO1pM7ClnglDZqvlZHpG7zIvkajZPj
I857UKWXo7JLTJjGzAyzjFv9x+rVJ+4/Bu9UuUU/UOuVhu8mgl6Riz+d6QdFHFuc
NQFdVRpvi2lfE5D2wJhGw4aIVIxj+5F8Mmr72Kia8SBQdbNW0UIXIEkYR+3Qr08W
6H6L1QPdaOWkyg5ICKeKYz58zkfI22LOxc6CAKQLdp+vB5qg96/gbZ49X6mzrazP
dPTEd5zjrkx4RDD+nmKmmdyy81rjUY23LeAeisLuyhStoryTI4lSi81DNYrnAG6D
W6sO0Jns1G52Kz6+weVaq/Mq2x2kjdwNZFYYfhHhxjRArQoI8Cm8iA497yUr4C5F
u9sIFY+DYYsLZ11kFlCdWxeBZku8Oph+kdR37H6hbN/z4z3yVVpiSl1vNHv4Tc0k
9D/dl8gA+Xv0uo42VI45rtfEz7BVhw2XRS/VLQBmXKzbH+8my1ZKddcvIeQctPhH
VJbylNlLGdlMjUUzOVdaEzyE+XImwIrmAbwEUrIS2eb11jQlMtmF7J8HKrXFvlof
BLgOhqivpbr32/OFyt33WkxyxEeyuh+E50xkVmAtmf9RI/Ui4+VUEqgq4l4+fDK5
/dmXs6WjjhHchnRuug1147zwxrZtlgf7L4tYzs2IsdsA6kVulvYK/Y8lp0oQJy1n
B/cZBXPxsBziApz5kfBkGutRgW/TCYe/c3UYgMDdP1WyfmZnEdhgBSngejSLXur/
x0Abowo6jB0S1+v+hVSNUWUDnCtF/aOl4wAyTvnFzWdi6G4Ha81IZDTkGgNlaCNi
uKdFMSsA7S5bx8ciU4AEoQk50CAJb2JL7Q4TztWNc79zc6JpOiwbVnRG7Dm0Sig/
Tl+LLgJ+hB2t4wvYEbl4ojZ7wGDckx3AITUt32Hi1fQWga+/KHZxKEwqJaf8Yw76
eKXeUNf0KW+tGO7QMkWY7SpjVGFvVeGzT+FSLKxD84E7A+KqYI0Ttkfcdpx5Q0hv
06K+sXpzQFt8FOhMFu6SUC9+cW7J2tj2mE8nLmMwiJrWUSZMN5M6Vsa+pPs8jskC
9qk5I4E0zTaz/VG6PRlOfLbdVqUETcMO90i0GeAGOGKQ2nSggnEtchLrRggVsJmj
K2QvveCC687OleE6wEG/Oy3vvzdYkd4xt3Mu9AkWIQo1XYFDgOi2vlLRlpzhI+CA
6bQX2apNAPoB5AYeJ3nDlwrnCepKBny3PnVphZNF918+mj4q36CZ2u/RmU8SxZFK
fPwbR+7/YYKNThRz3718ou9/fDxLuQ9GudsdgCn0k7+eoqKrx4jmsQv6F6bZALoK
EWBbBtoYNtMFguADs+fXQSmXQTALvpt4fX1UgEUIZhvwVLvGDB6C7+jpxz2aOwLu
C449AlU4DOkRFO8Plx6CRlhgNxVDVnc7SRQQpARhb4frbhWod3IupArf+JxmNaOD
pDWx5Jo0/367jcS4pKJQj2aej04+hqgVj+LCuDN9eBJXWBtNKTNiXDLVYD3SO7X+
J6wCRQMXf+dLZDy6AHoTJOzEqvjU/uqr8BENmO1Hs8M9g4Wmq7Qr6XWImhAIDKmI
+xVD5aKyNNV/cOJoYzwsxDGvY+iaHQOed21b7mBpFd0OCbDGsJckZ551ip2Y2gqg
gTk6slIjUiJExIeL4bB+yWXlef6vDqZGYwZyutP1E+H6kuMXaYCiEQUP+SD0K2Jp
uN9Spmg0mJZ6yohX2MIWwGa6fRb7vHNsvmYJn78qmtdKfOpDeHnKhLjI6jMXRk4I
s5hM7D3dSIm2D8L8eKuU/6eUuW1grQkjVGKtExmBw6zIbzrkeMikbUiydLz5YpHZ
b2ISUyA6Kdquh5mgx6JwuMn37fgykWtJvQzM6w0O5KgvUD3LA6fM4UEpTa10Evmb
FvdDs1mhkJIr+hHuL3PBFxX/u8vdu2PPxCI3qYht1LeExsCMRuc5qAvvXz+tKZIn
Y1QwgOQshLNom5Z1wxTB+Qqf1L+nNyiEfeaFGkXvW/Lvat7AjOglgtmFAINd7soM
cNxTjE9T/YsUG++Q8slDCQnwPsETvIcQ7Pi2NmYXwD2F93ed8SiS3rUOvIsgrLjf
wX2qsHNUi/P2fHLw1scYleRghG/vRkXc/CUJ0xSdUf1VBN91q9ziJSCEGxdP6eH8
IgaHO2pmedtniVt5vjDREjPD3gD7VhTFoJUo+5hluvOpQardQ8wcC+Rcz1FeBivX
5DU1ZSQpXm4qEvwP34IjXRsH7HwyA6p1nK2lg2N43/1OhnY7k53q4OYIkYPDglJW
KxMr4axFiCnbx7RPpbVi5UhGOJ8Z1w2esPGk7fL+VsMxzskkwW0ad0KaTMyGfeRU
9PE2k703sj8LGx7MLa2ZTgwMbifcHCC+jYbpKkqvJskBsZnBzj4l9Mog5Rba1W8C
hCHoum0YlAlDPL8AjE6fz2Sy7JSUOxChRgCnc+gsJ0TismFYzUzKUNuFQpGV0WYz
pnSksxczGASb5BY3F6fwKNb9HPlYCg2+WYsWEW/7pi5655Vh1IqFUcLIG4WqtKkr
eUycN11Xr5BahwRmoE2IQc9rvUZkxoog3ZRNO6Oeah1jL5blYAcOXrNygbi3hfz9
TIGnmtBUQ/Lky3AQbIEiJ5AIvupiM999whrqw249ZKdUMAlq47EZ5V8sC8U6jsDp
Vn6+uHmbmp2sONqk/Ec+77VubJDE2qjJkZIZlqjJ3lKrg42uui1jR/08NP8+MaoD
jkJA5Qlkepz7dbmAn6zzfsCq53BTw6S0p0OW1VMd6WEQzE6YM/SpKSjjVfVNreiK
d0JwEyzX2kzQKapy1IxQKMLMmLMCgLFCvOpG1Urlq6FaYeG6oIqyvqFBDRDEnGtp
CYjh89WuRU9jAArXrDoAqeHqHH+tnKh1bx5IVwR9uOWkuspFltTDWH0bzlPv5mB0
3VtRSYpwB08itTaRZ8PxxkwtHXM52ds17aC/d0i1zPqRFWQTwrTauIJeHyqXSoF6
yDSZkRRlvak8c5auYCcOf7zVFaD3oyU0vcuC0Nj8Y04z7KNVI+Vv49QAS0rhYNU3
M1enriVwdKvNBkOgHhqMfgrql1TVEw/9Jc9MoKM+jdKyD44/W5WTU8VOBSChzYs4
ZSviMWcQhyI6LwVQx4KZzobYz0qLK0SCLf54u6l+CWn56qVlGJpQ2OHvCRCuyuPp
neNDxV0GJyuavpEggC/658hKM/+DQUXOZqskd7jX8uESrFxN8zU1VgoXDGQeoFYq
i2b2lJTxQVrr7yleMzhAbjBW1vuSik4i1kA3YCd7j8y+0QOzA/EbKgxJaveC7xMS
FvM77daGndlsXmCf/t2YvPxd0/geOBLClX2CENKCpmHtr0CgZO66CbR2OK4br21C
+gkYVE9+NsFJ767pHjJGvRhvNlgavI6MGlZkozNTaEbsDNLRycGUrkLFrHsKhMJ0
34HMXbIkSBdsAlyztBCaO6DfBSUWJoXk6jFjMNfiNLjHo0RgwJfflhsLceinRfjg
zj/j767qXSMPQ8nR0P2OnXdplFBX0M7yXCbtbGrWdA++RTifonLIhnM+IzACfo01
SSx67ZB08/7avfHtSbDEtrOk04P2OUANM1fGqyDls8B5myM8A2ydWPjr139E5YN9
bfjVLMjGIOgJFj8zf9rYiwC6FZPMSyslu8eM2in917HFZ5fhacvlUuunLgyQH29O
D9mi99CepBDK4zhYrHtXmwv6U2FIKjAV+mfOVMLnkXY16KOnR9vf7KGpF38rOobC
M5sDcEpxBR1j4nYNVaQyzOVggPn6v7iFaeUpaU7BZLUgg6huF5GYdOxlI0IRxcta
ygco44O6YaulWb6zARpAkvsZPGeJfQqisaXujXanLh8FAI+WeOGiYVGp74hr/98v
uh2P4MX3YsHqJBp1RhaTDIt3/XAXhlo+kOJeXsMku/USrvQmsnQ0ApfUNxcv/fpn
txGJxjZOGKdUtaxXTKLH1SGe8jIS2SgucVI3zbxXNYONZa2RAnbsbrGJS/T03kd9
YAiY6tNUoLAVxoQqMUNhhqWXptoAkuTys6IzMD02Cc6HfE8XNjCOuJiyr229tnj9
T1D1Qdf9XJT/p4CO7TA8pLhq9ELsTvJxhV9epEWO/7Nz1lNaBrl8bdMHzY0Xm9Xd
LrE0u9hUDSxboqreNN/IdU755AdrG6+jaCGhprsiqAEavkg3KXRyhAIymXa1sWB2
6eX2mC34qN6BuSQWpvi/C1yG12aiA6QSZO9Hj5bhpWPz9ebqooGeFOhwzOCU9Fkb
ULnuQMolJXCQgVd0E3UZDgHsQerkGxNr/b/DOVjk/5P0yhk0q+yMEgXWJmjamMB/
TtYPGDW0PxoEtnpAcpOkCwk6C7ubKMO8w1Wq+M9+pHzHR8heZRJJfuLylwBJPSiV
qepo9ZynQED5kD7yHx8y8nOO6Jh85vPl4yE5liCIRpTfQb3odGQI4DO3RqPGWCpc
XP547AvMex2RRonCZDMJn6ZciWyG1g36uBK3LY5hMQ+E8pYnCkQuJLdaueLPAHDV
g5hX8VmAvycie8xdjz+cZzxLZP/1JlpJ0n8Sv+EF5Kr95pwYmz7lu/wRe165UCMv
WPPIIp8mJQNFT8mxM6/Y47AWiDu0iO1eDb8Wy4PsCo3zqMeuL98oa3QLholO6tMA
4gTq+qPeX9OsYOOyjb2DgDIu/2e9tC2yo5oR01H4aVmqmdoJbWVVyHJBjV2vnWRK
CycHBe4JJqpr8Aj8B+qkJxCNmmg9XjiOYZuyp3YA7ukQ18SIhRi1Es8s7JCReg4D
ojMHVLrTqqj0kF34SDDV7oDZ65/+WWpfKjOChZWBD+tkgz7Gh7K4Z7TwGK9qn+jm
Bx3t8XhT0jvwoEx85rc/BuuBaPxlUvaaqqHsxiuZ4zYBP3U9SFjhNHklp2PGNRWE
J6voELqys6ZOtrc+w4UuUC1Xjb3aQVZz3OKqQIE8eqImcbZgi1bGLBYywnIM6qOn
Ep07SyhtUB3Vn3M2LAMDC1rwj/cjhRCqHe01CJ49dVOUxat9l/6pH3H96bis0Oht
Im2Tdd7ht5LQDPcU6IodVqGmlLZSFK8Jwn9v61Qe3Zqdcb/TlNlW+zkjzZrSaziv
k+89BjVir5V6O5O/d5qoxrgZaw+3CLyJ4v6Mzo0ZYrBnMiqhxzcp0z8dnC9XOJZM
XG/S/bzeYK0ihBhNHnuemFY9b1uo9D+sU/2Zxwr9nvfcdmlcMBMjITvUSrWTNnRO
SvEYhzod98fXmwsHBg15aUbNE+wPQ+rwmk6dusc6WIZVBoJ50mykvZDCBuQ5ut0I
iqW/aKPReIB77yQmfwIJ0cFtsBHa8nc0tyQh/6e7fbtMoAM4M8hg8S5IMN1DNCMA
SrbSNcmvfdgD+KS1sSWcIShlbgCCEOK8PFGDFzE0klwx/CaVJ2Pe2ZiPfZhBpgH4
SZaSY4eMdkHfro0BU6H5NSVxj2ODMOOZrJE1y0BD6/UHQX+v7TwqFUGpD7DJmShu
9+mDh7w7NFhdelKOLvEOrHV2lUHmXsiKbEKOaj+3x8Qh3IebP3qCkH2AjaQuthr4
aaT0Zpzw1cMTIpONMa6vrGvyLB1aK6Qs0bNzp+6F+WKDSGNrmZi1L1OulgWX49Yd
76pmetHsdQVrmi5TJDuIPsjPhWo4ZTvy0BYTyHiM/Hhj3anupHqgZh37gog4D5KS
w+lD6jnuLzIPElel051ACwfuC2MUVlHo0MIm7Wfcoz0ql01iP1vV/qVlWcvqN9wy
EBUs6XxNHEgVbjcVA9Un8jllbPlUXyMsmmSMF6NGC91WSozfrFGq4XE1KL4Upe6s
UaYaNsRD3OiRarhiMhZZYk4dL9bbTSpMuUjwoy9LtEf1jbun8s/Tv3BENWfQbG6J
3Jd6I3eQloO/7cu3YQY4F2QECCgThRwd4IsbznWHW5DH5V3EaBVxI8KPfkHIM8Ez
GbSlwpSUuH9VCOG8G/5S8nZ6H0RiEqsrXxRPhamtFhe85I0a7px75NkpvR++3syG
6Cux3CPN9Ai8LGuCS6msrD912EeEGCBb4B2j59WR57Bk+iu5tyR212fAO4rLmJ6y
0fBZJtCN5oNsoftVavz5EkPsu4UmwOQLq7A3pZ0xHi9x4yR2Rcz92skAuu5SVinz
hVjStAlggu5fP20yOcHCy4L6dtTg1bby4/VkqC6NXSuztoLO7LvbKerZAOirgMxy
LK1LMmMglHvbURn/+TcFZHHDS7Fh4YsY+XVCyFriiTAEijiiZ/F0lrGKvwFIUQfQ
WZxE2FY56IlZ9LUaDjNVsKukfqo1H+KoMyM6v1TKh0+zFH14QbEfc6XueGL5wuGg
qN6EkOiYSvVs/06sJeXe9BPwAND8a5xlC+001L2ne20OfuNhLOTNaV8FFcED8aHe
0XMTtfwYKf2OFkiY/I7o5IC5zuHA6ftQqi4EiS/UimDvjHi6q9NKZ5D5Qfl8VSz0
3merzJTAbuE+ujj/ZJjqZgdYapLZZvgY2ceuEylLh5FXuPhQtsJMbGSRx1boXDxK
7Kgr0c2IWztv7C9DLhoA/sQ0GNB/zgIMzWEDVKcHVhmRuXgjVUEQDlob8nN1gtZD
+wK3zFTZiVT100vPThBnrJxcl08+MD6C3snJ+y+6RanVWKPFlPejdBC/9iw3nHRd
I6Od+mn0TY49tEGba/1iP6TWt6si/RBI/HgUYkDGcWXgM9QWcqd2GYZARe1rK00g
46fPA4vg8qEvzqRmHseXfdNAZfKfpR8TO0X5m2YiSJKvYpOQIdd5aeZFvpsi+u6o
ihOf0HtuBsUnZJZezlYlj4j5RpCctZp+Eh8AF1IDKXLsvcYS1Jo5BY9iNNq2ftnj
60O0V6fd6hpaDXXl0qL9LRDCwn5bWypnwbul1mLXxQQW2sQuIMUmpLQVTy7Lpmgl
Xt0lvhdAgNzpJwsCzhPHdG+BoV+dAoiemkNrELeM81XReXAU2QpbjF5w+7/8ODP4
Y+7O1YKfbUuipPwMqFkzMTfZ4Yfp81DrPWUo2G786h+/FfwFMT3O8JmT+NUIy6ZD
nfVYqaBcjFBCUyUrNeq5uyTZO88ppOaEfD7UAMP38A7cNamnh/XmvIM5f0XkT8GL
9dGSH8bporOSuho/wIQL8brnDuGSKa0Wvv9iCXl2rxQ0y3TusmMu/JKYQWAoS88h
20LqpJD7pMQ8UwXBLFctiHc5DPs/o+zQfnSz+4Q56pxzTl6nWTN1x8fwDLvhNEjY
Ks05uqTFMm91EmxHS1J2YZu+qTHChWckWGqppq9szGGUMMlBqCxKpx2PuSDIISdF
mGoLcro9B2q+Z0vG5oDFzbdawTgYGzQOksxUugqKo254lUS/lBbO0ooqOTWfXP9C
NJjD0XUw+BCrXUjS312EOYq1pOOu1kgl7eKEBo0u2PRprvBk7x7StBzb88d9ydJA
ztpnUrL3wurou92+uppwstAuSU8O+qyU3Q6iB9V6ZK7FmZLO4tEI3i8ajK2L+HYd
iX3O5hHQBxTGqCFq/kH1DSbOjl7szqsyrlw/e3/SXCL3+0RXQkPIDwXJ6TKPwZEz
QRuf/BtnU1nMa3WGxCObWK2Y++ThxV7YvG+9kmUdwayvXcwRDZVZFTU9SyhKSeyJ
fnea9IJP7ekMYFXBZm8H0cwZF0bLHl/uCvSj/dyR62VjiKEEJZhnPY1wlaOMWjun
pDhLzKoqPreUkLtjco15ltCmCNGPgQX5fVgO4De+RDzojyMVSaduNzzASUFRQzGE
73oizyxU6/fTnMPEfEFZqHvo+DzidhXl/bE2AhS5XAFzVsewX+FTLpSi1T8o/RFy
ATb4XuIZYoJBkHH+FHSXFmU1/uisMtQRC/o3HRW7O3Ezn0srMWRDD947EaaL/532
xByIEcnANOGiN74WELudWUYJrP2Z7kqGaZxZJdB7+UnoM3yhJ1/u7TsOb6DZWK5h
vDnSVRqPsJ5fUoLJ7/hVrrIfqoPAket1cwEuwGWo1k4wRTLSyKxLXRKuqjXTf6En
5CbwTXCGKdFtYS3b2bgVAtZz04Kjly5GKWw71TWFf9B0liuGv3aNw8hO+8ADUaiF
cfNu2aBGaPw0LCkZtTVAGJMGDpR2ZbA5sQXhy6Oo5EWdnnbE/BzLCicmSEt2SPKj
AoccjmhVZV/7d6iFRsoaDdo7nm+HPHdjxdDDaV9eA4lZaed/4fLPPfBoUtwDZcNj
Jlyo+DjPjpdxschd36XM5MIdFDwRpTzh56ubaFKV93HnBUxAntissKYBImzofjty
VbVCNZNNx8FCx9wUePK0KIPc/DGm+jNL8JkffgD5DOE52gZIgQS/NPUnfbsFcDj1
cnqpKcIte7/HBVeDFiMAzFbZc4O0F2GBWbgQ3pV2f80eV3Lka1ySAgfhphkUKeXl
xGEUeGxrObg5L5bqJSLu4yBjf/jrTU8aq/lu58GyRPFV1uQFkAAXk3b9STvktxFG
lBk769d7grAHe4wUmEbQkH7IZeFOU7zcmwUjpyorTlpKJt1zqgQeBkVP6MwYOBIO
Hx8I/T6Z9QjTI9PGl2GXA8tGPAibVDH73JhC7N5atPjgSEtOWzs7ezEumhCBAWh6
WM2q5z4rK8j4VvySeJDPKaQQxieMABk9IKBwLkY5feou5OKOZmRTiz8heXzSXpbS
3NrF8Pt91x8VTH4PZ5p/yHpuD47kTyPpSRNUXqA8kA2zTvNfdZShDvGiYVBgVwB0
jv0nTeeD4UAW5HQSDELGIq6GWqpNXJs/5QEbdO7GkQKYdF+eyq4PeUhG8e2G8Nch
T/GERpUO0myhVRdKd468ZqfZjY1NYHyi75CLEQLx6gYFPiGSAQN4UX7nWh6T+4lz
9fB9NtrEN5fOi1Pje1Kc6ZYHLrwbzx7z3emv3+suXmPy4189S5Ad5A9ZG5hZeM6r
EfXNP8I6WxEN6D5VJh2IY9Ua1MMIZ4JcKBHHmCaBHIpM1sODgXnG8x/yGdXNi+Wg
UUSfiAn9s+RUine6BkiV37UdgUNDmcvLpwin9DRyZ+AIHzegJ5LfLeQ7Unncc7Kb
f/VgL/c1cEMG2s8CN6gXb1RQM1FbA2jARP4ILLzhlIE4v6QTVtMf46F/cHpIfXAV
9IgyvxNFlU4y32Ahox6NsDAH/wJL/VCBm9X8t9TUNd2BeVU4JHr3kLe3uIaHPPAj
2TzZLmG4bppQgG2Dx1kb4HSoODVSHua12TAxlBskCZkG9/MxlQXyNIM+jgjdjrTP
qoUVUdqLc2H2vzKmIswlxygZyxodY9oXf0AwIrgnhjFTyrWAC7rH9p7Zl/MS2qzy
lUMnkHPtmCCSDUXDX3MIptAFGHpp4MGrn7123iXab8VV2JqL1jTY7Rdg+z31kB3q
1PTXbWBaTtgzNOehNSf/pli4WiGC/frfKIPUMLcy+dpGy9tBGYwRbSs98vAVmY7t
cEQiPj+QOcvXRknaVe8kIY/5JotlP9bqfXMQS+2r5gXd5tKjOUMJyyn6NDpKwiYx
ycKNRJuijGh5V3dD/lGzmxvBDtOWyMiitsCxn0E77UzGsNsj5UDUxrtR5ix+HzfL
m0Z/Yiw6+LXarZpKKPGCVNWr0dd3MOnBk4bWY8bS0+r2rjIlDgACLGvZqNqnr3cZ
H7PNFmH3Bn4aRF1wVtTdOP90OZV90L7fYzQxUwEksSSxxP72OI28VVpHDQ7SicSf
Rt0EX2d/NuOsZVnjFS3gDAd9wKrIAJ2UU3Vx5YvH+qJQWPiZFPrgWwo1QDzKc34B
BqqifXA43AsKyKzTSpstdBobA2drIcAZhoQedBedNCvsVWvmw9skCYismWdkFv7y
uWsYJ7L/9k+ADwAIec5vMKaUzvkVy5B87kDltKc/icj5FmAOqa8MBSPshDkGSnPW
1ZY4njzxEe3rgHFYYUGkl8iHOHIbsV9Z9bgDFRut+IXHGO1Bi3t0d25HEAZ0Dk/6
y94rjCrqDX10613gxQduqlduKu/8M1DY3LCX3/oMCcxuyhckzvC36ryngXzCnneC
xaou4FpfU5IrrZu+bR94fYwOPbH48QLzbsmsWcRLgTHtc247Dwkw+Zi9PX1lIeBF
BqADzmUeMJDqzG227xUlvaUL1Mp/8KBdsAoxPMjbTowAjI89XBLO+rySeWoD+VG8
csFN9TzXnZBIokQNC+UeyrDu27G+lFxNZTzcMgCCBxxrF2c4hYbFjAzgKVq7QJNY
8RRSOJN9+zSNnpcz36LgksvpGsAlukbn/vV1AGQWI6slVQW8lcttFUdJJVdseDWO
7jWWaoaRZe84T24VTGgGwjy/dIk7Z42SF2Bn5Wa0VM3/KyLwjcJU7V2PuwplNhEs
LzElFk4AHjhv17+AMIvxiaVF4CuOlInzfeTFbos7Mxz5V10jUG4W2St1ZQDtqh7V
516t2/LslR4AI/XM+sJoIT18lyz2Lyl/373KE3D1zsUnn/TDaoFDuSksHWGSBS9b
U5psEpZQlCzSRmYH/dCs4HdPi2UtFybOMNh/Il9ErYz7lN6VWNay/XlOqDaihFen
zmFrZ/e5LzHhyOTFKukuDuXvTQugmMEp9if9zzRYcwERJvomhijY1EfA6BKV6TuF
tLezMmWZZY5c8TaWxDIWOvyUEypBDUQRHvTnFCU7z081rNLn1OjJtA3OvOijP+M4
psRKp9MGDM52TGPxeT+aeIyVychGARZ8xvx6WaEUr0htt6o7ebn0zvLpVKiKy8Ad
TDXYvHv0/88b0Frw3lDMPF7p2kggQWfMgYlTuakUCD6EHcL7IWcNLvRk08DhJoPR
PfTOvG9B4zMPQgOb6Ws67foZBt5vIZwIgCSI9htne867LF7nTdCapOnonBCqrDV7
G2Urg3sCpumfs3AoTH/p5baOMR959GShiPYiafCEiT8qs31K8nkFXv5/nKqabCTh
gN8Fukqee+Y4MnHPkP+gCYC6aFZlXAJn8rRmPf6v/fLkMQjpyTojACysC7Hy6xp+
P2vwbH2PUNUlaS0qCAJO6Go7Bl2ueaQ1RFLrx316RlgoDaoPSYMY7e2AXoOT6pxR
BF4MrtiK6OAQXL9LyC/suepTmnPrS2Ep6MTUwbUQf81+jarzxJGqDHwwdypK0Yb6
2+ycnh7V26yoEziaKw5pq0yDu528reABkn02e9r+YtHagSvgjOVTf3HAaTghPy7q
NESYK2ocF2lXwOQ7/qL52uyoE07K/S2VJg+jTcdpJWHXsnmSaOLmuoszxCd3CjvG
SXU2Sj2DreUCI6VYljMeC8ccc/GhYamTbes+po/Fxdw+cyk7lC847Ux84GhFg7wh
NwAa0lOZ6s5caGYby7mpA87N7xfn5aFM53jSuOvMqK5ZsedLgFrKaLlnQdct7xcM
tRUtnxfxF8WDEdFlrmjwcPQSCu7qiSwzflR+Q0xxy3bZV+/ibEsVTMDhSOAbD4nS
2nTAxnC30vsEmKoFrkKquwYfTBiyWlc+SQUxe0KPaNVwXZnMwGHwF6yWqh2z3ySc
8FK0NZYsqKzXQ2sdIMHMsyvPhRFW0NxPLFNRk18VaPPw7cjW+yyLnIeECu4OQ7lX
FBjZ/07PnG/9MyEQqUT3vb/5ZQhIevSoJuOf51jIanNP4foT+mVDdQqeXBHu8JqL
8pzMZAXPSv6Vryj1amMkkTqv2eAqt/poiQs7qfZ3iQBP6+NJP77k0t0/e0VuwW5p
9MkjfeuYw07JBTxt9a0J/sy26ZmsUze9IYArADn+NBzj5yhm57E2SiUFKZRUiqi6
T7AK81hIILpvD5Bk+9w6fh0sK5s1sO9UC+0y7LiGkJsXUv7mUprGaTfCATfs9pjR
/r+dXLXXl+eH+Ef4EYWS7UTJdhzfL1JHgATW32J8iEy0eGGj6Nl7xCJakK0cDr45
VWoFZx1fmzqFyNX8whEYuHpKLpgi3pxWExZiARKosyoaMfDmG5BewmnCJYwaJs1o
K9eCIEtnxh/WtYRTXE0EvJEq+h2YUdClxKhsmA8uv8XY2CNtRLNpt7JZigD28Ney
QptQrbcWB8ykWMUCoh16UCPSFNWTSNqaRUiXR5WrHpD3ifPNd4AnundvZEyWOVD/
6LIIFcpewZgo7nI4NHZH8F8QUd5Rz4F/QuBGSQuatu5N8yOYbamE1wvWccuiumfQ
tgMGzlD6RJBHAwzXyz2P5itnEuQYbjgZ4k7F88+QQ/JXF8aQgxhHfyY1gzSA1S45
jolY6STmBeRtROQ8prZ2Zo38dDu9fTR5RFWklflLK8bKvh/OmrVp9MnhkCNxyvtQ
envI450ulqnCnMWl6KuI/g9RkKMqh5DulovKHQmRvSTQTX7Hp+LPNWJAWYQAs8OD
kP6nCWsbH8oiOwmqG+JjFL+WpW6X5XjS7rSUOPOdrppAsGNQvpyxIBTXqlolxShE
wMlagRF1Dnu2SOqKWFJUc5XYx4H/EyvBxEOFdk8Mw+K1v7LvS1GvkNlTt+OQDAUb
7qi+THSp61+NJDjmdATLPymwnoiKDhmuewFWhGZcEXYM4zTkfUgoSUe1lNF3NO3B
G3iJtS7K2SkBiLDErsJoL7GwXVVaqbXf7qGyElb3i+y6L5kkCUrW9VPMlZuODCxu
avtgHyM90RT27VYZBHNd3sQZWY5COseFT5qEbsnw961J1khD8OP99XWB59+S05G2
LBHtggMEhR7n6pYKUsD1yhx8nKVq+99jx8t49TTnO0zb9YUawIDrteGsA2+Cg4jV
Ya1BT5oubUPOiYi0ToGBlwdjEssD0ZDpLs6cX/ZM+sMsJiz9MzjBtTijxGoENr3A
E/XjuYDRzoFkNUT/e46N2eYXeBmkoDtDHV/SHEFdxuL1LTaij8vai18PccCDegfO
5mpbAgoXA2+RMZix7gXgCaHa9Pf0i/QKE6U+W4MXfksbpCzfPhGCiIe24fELqg0L
qGKiJhXuQwmaZ8sp5hlH6nqNT/Z8X1V9jqpzcY8so7hkhv04rFsvhu3iVEYzw+AQ
zziqIC8CclBb2eEE+SP/5137AJaVM591ZIluq3AfrSZWGgUsu+s2TCefGyB70k4w
pbNupdG+2d73OEIi2vX9lsr8pEdHLDofudBU4SuE2DR+nFOiW25cPHuHhn78Wd/w
rVGQacWrML+7HsnKCO4Q0dcprSv16ZhK5nmkqXSu/lEhFCL8MisRteH1PHU48qpB
G4JrmrnmfgwZRhWZKns+4b19eBXtyGMPhofqgz7uB+oEsB0/s/xqxbUJ/LiBEGdy
euY7lYgVFuFPEtvm0dBfWE6n2iMZep6wXNw++nicIXZU0M+/EcImnxQUL/avN6Bc
k7KY7RekEr/7NRraXF0lCo5tMOCnoDmOSOGXc0spYuOrO8mvKfxAjmJVwBgywqpL
tF8ueCTjNeGAl8ylcQJaSQX/cE6GB7rELAHj02wCxAHuTgGB4QGgaOYh4cFqh/ZJ
EoGaz3FWJeTXCoLidRmtbdAdZKXjuM23/bz/YBSiGMrj5oH/CgpBYyEsergjmisd
Vnl2/8V8GXjSkzq8f+I7/iHO+CO7loAloQDJCo7+4w4ETqRrs4CUpKATaSCjQ2WX
cdEPZXsJaDUB6jQWbblx8pZ+tEV0nn8Wzfc578CKkvAEwwLo8RQZo8HjH/51sgLa
QV7pQvbKqQ17GxY2WrEkiEpilitDh49x0X4rJwriuJqbjdwwHGrv4KkJJ0zRvNVH
6NSX1GtsmK6YUUcvkYkXb+iBewyP1UMIsoikHB/hyYuHH0BEYcL7XtoXQ+9/j2C6
BCInoz+7lIqKXgE8ruE3dK7x0lxahpDpuw/UTUdudBTD0zdDDeGJy1wGF0JipaVX
TBv8e71CJc00vrIirMIW8eXMaSyEn1UNea6akS9wCufB13nnbloCikGae/TlNEen
SDRi5BtAXFHPLJfqNgaU1h9YjH58L4z6rnDLj6fYFSqYYBeIEg/Uo1RsiKNiplCg
hNBdEJUU2FfgGaN8pFBb17M9dZYj6/8m1eAuuost5q2IHfa9YsfVYFoa205RJ9rh
ODo9pm0fecYun2ygDJXNouDoNid+ojPkTTanHXJB9lufS6Z3o3CvkG/Vc/fHL3Em
0zlGwP4MvcJUCtsklR6AY3SpJYMz+U42gbOczwq4dIp1SBPZiwZFI5smH6+7qnbr
+Mgn8AMENe3ffyltouoZGjJsIPvdXL3SzcrpzQAq8c6reGNzm7pbI1Hp47qT41C8
s6WabTsW18D5iXbgBt7lPG8xR0wHOIMmNBZ3XIzEYNXaAncH1ZDjlhdnUGFn4xkW
Wbb+gzv+eoQt3TsOpQrUxfybybsX0hILLPO5gpUG7LtAp92dXK3jd8qsuojHnsY4
9L217NlFpJk0Ld3/IOPyNcfk9pHCtKscP3A9CWghSwB58BPwr2e7Uw50PIoiHYCg
NiFd3DoJRdxzym+PfX2vE8A0Cpqx76Uwob1Tjb2JUKaXWWRxLs/UcjXE7UzJ60M3
blTaupVl9co99eLDJnxr8UyIfZLYgACHy+14kCmDpbyC8IFWv0RPplStcZgVVRiy
ZjQnDj9J/1Nl/7NbDUn93iAXW5Qw5w1j2VNSLE/+YomMlFqqySpExSI8nGkbbQVV
ye1CFG0a1ctQ+TfQ+08E5putR7/O8p1SJ09dPOqMPe4Fmf7wHerZkaFYbhLYXY0A
W8icCaKXNCGFBatNWVo+EJCgUqZtg83WwulhJRmEcJlOtnthxthMJgj9xu5kudh/
tWpeeD7RIjvqVbR8VxWm5TjA5QFhVXfF2H+9As/dEzM++L/FWEz0LLM236SiJTU1
REfsVtM7Fjw2P0ISnfTiOoTvo/ItwtB9lf9hE20bsLSS+tbwbQhUkNJl6O6RKqrE
XjxxipxF3rYgWElQG21D0Pr7bxvb0pux3ltlK/weGlEuhrgNIGUbpVMOIG8zdv2e
FAJfMZ0A80e9/36qrehOxEODA7HLpvpr9bjb7SbWeMXCCAXI6QH+A1ufEpwSRHg0
jXghuO46mFQFBkwXUGRSlE7uLeRhwIpzjyHvEqiox1QKgzvzoPuPMdk3s5znBDOz
QvG6QmBffYADaYofOBff8XlT8y3r28ILKReJhr53epqCB7aDu9Hfn8nWx8/pUMX9
JKaBRSUDmKBHR2i0IFQZHBXT/RzSAsf8mgoW9e82SOgC80+69sYJlnwbF8JKlQHj
EwtBw/u5SReh+fQ2R+FqeWNXQwi+Qp/ZyVHDO1v75vpAt27fYhka8F/UlpwmLbSu
u7/lspDTT3P1fhxMKvQ0WDtxo7/+spa3Yr6buLVRQWV27myU+fY00p5qSTfNzfPs
HibPgZ22Oe0y+9TKG/GcmzRznEgf7PgZHioTZ8hzUTlFOGDOjA9IKGBxztR9XoGp
LzG9gHnH651ZvjjC7ueNVhrI1mXEu01K7iM0KAWO7w+iOEe90ZfsmWmAvH7oE/vu
t9fKUzw1+iZMhJ7s82v3Y0MyPODIWC5Yw3wOG2ByoyIvjlalUR4raHi49NZAOmi8
0GR/7RS2aIN4BVamZ4JF3GyiNuPC6mk2s7pMiujor95wCV4H7RaKpMvP7SUKl/Eo
PFmyy5pnYiBsiD6gPOdARbrCp5q6EUer/SD1mMhKUAvQNT7ovxEFCWODSKRR1VI1
CGyZRuup29MCK5Mgh671F6BUPQsphJkx/Dka3rHBVzNJmQBb0WdS1O+x7Lp+VnjP
Mg6zSkAq8aS0sfBCf624ZRK/7kRk/goRnbinNuczHREIyCc98HrmCs7RRIvVmdcj
oqdt8j+TNvSiCwzMSHL4h5euVEXupuKuJhjTqEedjN9rEDhP3Uz28q55a/SwyO41
AkWNHHpX34Ypz4VHWB0JZIKQH35GgYKNCPq65E6B/q43LYT5H20EQEi+qesXNkmD
78wfU8jUKuv3n0sHkYYtBcEWdegmi+aPvp9yJ91T6+dE/T2OLclkZPPjio+5TQsv
huknfncUlDA9ugajWfgfqW6gL8mxFr9SuvD6N4tdoJGl8YNePZEipldyL+roqDXK
UUlppmDuU6UpAItMt1vRBQc7hmnrjlgMSwCrLgJdTYmUJXMbaaLzKSm/PGGWRhwv
ucyRiPtmkrQxkuaB/VqYCkAB0ZS91ZEdL3Xll5AWQ4wmgd4VP2UtSnlkNW9nfJUE
HDcsL230XBF55z4hlK/3WYvW2M5HApNUgl45kDPwabESVqfRkIYL8n5HaoePmKnI
XDfds6Ifj7+C9fmhbA0ydlXgRDxfkI4NKndjnzmpCnZzL+nDPJESoHp4LG/T4Eqh
dgb6OjNZCZ09whTRDEAlP1CuOrLJA3MlNxd8wkqRjzoO4RaK4v5SAn23vEPshAhT
VWBv92VNyPl+54QejIzwGPelalcM9y4NAEaU71EZsAzWW6mRJnPpv2JhtaV5U/kP
DnZ7gwOFV+U881HGGDHnG7r0aVjf9BnLholXY+5Ile2FJ7dJAZGJ5Wfqx4EjVOGa
nuB+3RKe3TjnyGJfNz0lVHIEswKv5FcJXkW6ItOO5de8H1XvoclMEKo4bxxupBDN
bpuaNZFJYF5fVvRc//DE9TLXFdQ0J6K9F4Zg7nysNZDbM9qE3eAZGCXMEQG+W5xA
1DK/9I39hzVP7k0xWWNkKZB04EpFdjYc6anWl44YYocKbAlEP+ea8OEjARuQgyp3
XDvZmfrjwqRe1L6BtaP/Q9hj+NuHwBaVd4gXK2FPVHtQLms1UnR9+2InydWY9JIG
GUZKER0kGMVKPTBMWHnsA0LMeW/oAEJTcd6nWtXeSBQfKLjoNbylB5avdbo5vrJ3
H6zkk6uMd8kpZ39QUAQEIdEIkxguI3Cr+H4LPWDpp0+6OJklFc0CImwS1c+StUAv
zcDiluEZuWjp7n9kCOzkm5jljworxLP9th9tS82PxAbBEtwU/XnoO36vQJt3NmTH
koDBlgo9gA+jLdVoDrRyzPjpH68GG4OKTD35CiVxn1+WJZRp0u38H5eESgFtDa4E
PlDlSuEWjih2j17ktC2qSXvCyvlZWzJlI8l0UZI42jjmykjkLd28kySOTv48MaqE
EyVFlkaE5JiV6FuAVACVBQrBC0D+q6bgyty7/5Iz/P0qgIwnXhOf8z8HXTEtO2Hx
fccrY0KYUBu57CJut4p8rjP9y5qA5YLANyhW5y+cD3R8otDEMwORNu1kEzKZGz3b
szjOa5MmKC835TkDpczCa+x9j9Cdz+Y7P5OS/8aEUXjmDIHPafTSmBvo8PankxwL
7rXX6qIm+01w6aLz0Z7DMUJ25F6sS6u57y8W/RFp8uLawDwFbH/uA0VNMLbKX1LO
1MGpP7S1MMJdYaBSZ/lsqQsAi1URBy9ByC3FkaM670hH+ueJgrThtTkip/F4mkY3
DK01Efv1QuJxA/GD6VrNFsz/BJoeB0L6+MxZNzZ9JcNg9hz4QtwKIHdeWwQWdH3K
YGvbqls1QCnQFHGJvV8Blxj5SON8ZmdHECFVt8JsL0eG/8/MMpuyOl/OiTRBYwNE
kMRGkuyUq2vo83ETXEaXQDN+HKXVzknTtmZsLfyBWvEmKEPTwiF+QOnzWJBFWVYw
MQ4dItpYlZNlDoJIw96hs4VKPmVug/45Jid6WAUTZUNORZ/1s/wHI9Ati1I7FUWg
XSuxrZ+4YA1KGdDsXtd5FapIKJm9dbHQosZUrP5p+tHaJhpMnLioQA8m4DLxER6F
UME9zIfZrzwXxNPQbGrSzgfzC/vuPLJQgXe3lC8Kdrtx+c+lu9Mz7p0oEwqohxZ+
dwDGlGKVhu1Vy31eB/mb3tFC4RsPJjSYOsFGGdSKlrKJbonx4LmgLz01iTvwkei0
Dwhu7Q84bNgUAj/Gz25XRvPsDtgAy70wRnQc3tmq01NR6xVrdjX2nEdgaVIy5w58
8yXBRhiZ4CALE8aWF99ysSgYBd4XWAbZbbaQepkJp/2fry6sfnf/rOQykvr1263Q
EuSow3uNGZe/l7RKKbSfNFVgpIRFc8gjWkHhqk6T+WKr/TWXMEM/jYIJpx7I20eN
5SaC47G1jI8BgYOWT+5fTyqI4+KYYb+AYTQvf0OWdHA9ao8pld5dAK3qA6ryUdPN
IM1TF5LsRdC35MntI7yWvAYJ9FzUhI1z9brHCj16gx7+HABEvgC0ztkq+NKyhIY/
bIpolYybfKWIYNQ7UmfewnqOGKLzGg+OpN3ut6FXxpcaK0FMx+Wvs+WDkeKeTCWp
e/I1dnerT2S9BBH4oxK0OLgVP00TnSOpi+Uw1XddX6OaU75giDS0k5cEKz88sx45
CyyZEbtxU43Ejdf5kxG7QPCI94u0/fW6Dhb39g34MjvAyhAzEJIfHRn39md//7Z7
dvvPSGEGJs0Gpg9Za3MYjP2j/F4XqJuxyZI9oFums8q86VWIZW61CN8KcIjpzcvJ
XUU/nb/Lcft0pq1reSXG1fhm31IoSJHnkSLcFBtbVPCSdKwMrM+eAPSnFJsW9tsP
s29IxXOWFlEAyZjtgsmSpOhRkJHsJv/2XOElfo8eKMCrE+ZqW6DTyyA6IgM8vJjp
SBkv+Wx7bAoWLBWC0YF89V3QDAEAT/YRBPMsOXFULsiT73mj3BIeU+SsjZezmTct
vvF36+PuHCl9+Zm79un/QWjfC/9jhbm9LPr5pHeIwNhv+uTvGsLlGhd0xsYbNWDH
UtmzVlPInPh2pq1/2roxanCilvDyoACUL/hkEt98p0EZ+YMm/+BrIIRkA6JqZnlv
bAKroYErcUrv3QVaYVcj3DML6m4r31Pp+FzRF64UHiZUQwycxGEP5smirdj7L4A5
ymvWANbzkptLiyNnPjjzVWxc2XuQ6F47hEIqXSGUtXcNeC4mGl76nWqQa3XGQ2D9
GWbzhc+t/kZsVXdmKbeEA/YUyILP+V3JQyPQaEaDzi3vJmx5Vm9JiBV6My+xUBsJ
DiOaZRm/5Oy79ZTPNWBlLjRPOgawRrwuTRuMfDhwti2UjUCdt4wQRhUiHeE6ooLT
ANg4ySlsgwH41X8jQwnEjWRB3890hdIxkHWK7FziTLACh4dew4hRy9Wynkdgqs2O
vwAZA6/xkPqj0/dw+qWppbpzhO69lpwjU6ocoobo+FbcQzmYrD12WbPDC1azocLb
wULlqKLjCjww0hGoGV1N2lMM2yy1b3vILAW5WhX+GbzHFu/CSckceEtN8Qg+RoeY
Bm+H8CrGApFMV+2a14jh6i5frYahMbmvj246GmeNTAlXZkx74Eu7oOM8RrvUhLYL
+q2+qB0zmyrLkdYZDV1ANBhjNeNzl5GumnVloiBCccZrF+dPtMU6NTjZXPwokfLx
uujuYb5PTw96T6inHUuXemxsI+ndMARukzqlBvTo8EVrYSMU0gKnklUHKOipb44x
TgiZEuFR9iiQcaA0Mgmv0gy0V+I7Jd50Vj+7Lp1eldCfnRT/2oeGMetSPlKy45Wk
H8las93OTH80gcvqKJpmrL5faeGg6CwekWndUwLSR+CLXJk1OfwLZVOegNeo7oFk
0isgzW/uEkAj/kEH+1CAB1S8MUELVZ/AHFM8ItWNGTcqHdZsGRx+INwsWQcRgdYE
NUY5jd6PiNBwGlO9Tw9tTBYDrqEXvHyY/5/KiTQzRLKo+FOrYw6X/MIEB7o72LoZ
Bu9qv6GZbJX6uPVPONtdrXTwS7HwBhOhzG+XcoRexbGjTuceJ6n22SrEei7oNw/k
pWGllfIPwNHiHy7P7omBI0VJufumLfRtl32NjogeaVTPX1F9Yz108Sn/mct89V89
TTXdXfLgF4LAwRIh2zSrQNcQCP6YVOQFP9fEJE0UQdnHpUWUN/uB4lRniGIc9PB9
9OK3iy6HobQVeNzdCGnzOylt6pnC6hb/3O0ntc+1Jm4YLrZ2qBR/O2IPvY2ybT9j
vilX1kuBjUnh0BfG4aJ2U9OPrNGKLoSrCoERG7ymcbc95T+7BgrAsitD026Y/yz0
+PDlHvW5QrmKs//AeoKD1hDtqeM7TvLYaJxbFGafgnEBdAJWOnYPPIoSHy2Kkwkw
1kXg6nX9zsgjZJqtQ8sfo/p0UcHZGTklhFIMOCjZmskaw+Rlj/1DpY1WYyk/tiJ+
CyE6erao+iBoJ4ccZJZZYWNb3965vQumuh1aASg+jw0Ot/y75djltzFu7ntpcDu/
nDQ2hmOohv/Q0BI3v1CsZAHVpRdZQlvx6m9rihyltH+Lun8F6xVYUXMywf6DBzU8
FSKYnvGczPMTEc5/rk+G3IqCXSGV7ivpE0zVhmrMA8Rlp8SfWbvalqjEjM6yus6u
v01pKnqOxJKa5bypaX6p38nRXlu0h8zLydWBC4ovMYcItcXRPIuF9BPQpG/SnI6H
jDaZ5iAYTx5bVctCmNZysYipAE6avyNJusntpAKu47ZrhEyJhEVtiaGrk6lChqJ5
Tmytg3LmZSM7e8giYL6GoUV16s+avoqnw1vgHCJr/C5INxqfmfcgihiJiu/S2D5I
kFS35V4Vo9TD5VDR873boCMj5F2u+SxLDMmH6HOBsXp+CX82vXTcT1XxqTlzPypA
SLD6ln1SdqvShqTkDbFSlG1VKJ5eL86qw65+GeqZ09+W/OMZAjR23xUnMXvn+nyf
ikkBhavFD3Ta+k3XZJXqJj6Tr863yQflDUuAkcSbleVAAtjKEMI+IOF8Ycc6tzTK
q3hI7v9nUsuhOrU79oPi4tXtLYu8RSdMY+GgvmILh8PdUaXNxwwJOnb7kDnQqVe3
yb+kYMVPs/mxfC5VBFVbf1thThqas3wF9sOBPgzWgwRtVFmFMMfY4OqPCc8LiJe4
cTE2ZgcJE8Mlwq5uMLawoR/tpxvqx5I1iqEnbjcfX3Br0U15HgT3WXw0MKABUFQm
zPUbmpgh0+iPTnjZ2Gcu7PWnIKRiY1cZTD7wvJ3AHwVmXVifBUIrXECGWySGsTSp
XEoOfCcN5htfx/juP6T5rEvebV9XiB2hfmipEXttwkom1CGvbHh+8zR7CYXOdz0E
M5W4wDSZrbDCFhieEyefG3ejm3Di6t8NtFKYB9xtdfjxJJsYFf2sVcM+aXoCjFWu
h8ti0rj2UQdtMN/NYciybLx+5r4EED83LBmJylbAoFr4Mnx0d9jwQHWsTTZ91zG5
Aub+4BZl+518zgvYYnQm7sxGbnM+3wkv1rEyJodrSitKwmp+Jq02GS89JvVVdZ5Q
Z3e0Q1w5914C9Dx6MBor8ZnXSGzqjII35x4OzALt2zvRZ9LMYDoHfvIr2mU3CCh5
b8GIFB0Hozg8NYJiWKy4bIuqOGp/Jjwh6nquc9Zro3qRAPg96dVTti1R5ZqaBicu
lNMguPpabJUIp4C7kF0xYezfW/jQ9TM39khd/yA9EkLu0UlYCbV5wsGCA+VLEJC6
NxzeCI1+lnXrQTqbwEIIb3ifMmhUofZJU8ycXbl749cZ3w/XJ1OlhT50srXS5Tmr
K11VJzWJZlfmVet6D+ygRI3BU4X0NFhOW3BiQqOlGRFDHsC5hNAHxxnxX2TOgQRW
kJMmdDGhEUCIC5JJlDUOhYbxSjUdj4I8bul0qclWR6OkK0cBk+VRy0zCWZgBs4Ro
AWN2CBMPt6r5dnIFF4QRxSMDa90jnPdxJYsrNejCPgJHM8dKrk5NgDwgPu+CeKUG
CaBi0eJ7qtSw/MhYWYlTEi4IOVjYwxFORzaI/bbEIRMrCNAROx72ewyxMIDJy2GY
JvD+kYmxfI4c6fnh/gIQ7h6j6h55taGdNghAUd/ysWHvbWH1s4Xrs+KAqowpAUMu
xsHkT3igoK9HnOqP/T3djTVejmRlv9M+5SQCflEfzvykw4kDrU19H1tSIomS7KO1
OydPOhebYvvgziEYkHByJZfovof+w1f46UTu4S8KrfZs4Dim2HIv5nAhOuXASSJ6
BgnBwaWPBC5mF6tEpzzWz50xyAHJR6insCWLpLt2XUMGZijGrXssgow8yLRtp+qT
uz3wK2y02e+Ud5yUS/ooi5bo7+tXO2RxgFfY01LCfx03IBASS6plMn/TQXjr98FR
ANivvmg354omHGLlbVU+hOGeW9GbiXk7cmXW5xNQNIegd8E5UUkN+UaIeAAN+Yko
hPNVvj6LI1hZ9ERjSKytIxdvDGsoQIy2cVKMO0AFOXV0xMdh8GOnwymwI8HeCOUa
Ahqohx1LYF00bxw8m5lWduT5RaFUAoDI8EtWA8iMWJycKi9ONh9uNaqPxS8wnB6t
o/b0F3zDZ3Lqz3vKGWzOW6s9Nd8ndjf6lwSJArPX4B59ASu2bi1UgCH1s81ZfJwC
HBCyMRSZRbeEk1llnEWGuCW4krNBN9VAUcT8HkZ3/Lmx6DC+VxEFZzmI/Z1mum5k
C4PnJvCjdTc4jTcUeUK8DxQC0lmiwxdE3IM/4lgbDoRoo6xePJOJyyTaXC2EMTvX
D5XyEMiKGVnHoFxmXoGVfb3JIMyiANaNrwt5AoqO41E1GUSdy/XIvXlv8C24iegQ
w5nALq86c2MbXw+aZ99yQHKPAPMManpi53cv14qh+p4Ul7rDTaW1+xir6aS5Etr0
DtIfAfIGjNgHP+XoZlnPM1BWg7ElJ6ac2FXEEWvp9g4DvK7ACCDzxdqry/ePr/yF
hiTcLp+SzEnlf1kg95g+YC2yBK/592IO6W6tE+jAeG8FUEJSx0fUlGTVva/SMUTk
bR8i6Y/93J9GpQtjhV1hm7nLKalV9NLh+BIliVaU8MdfLt0ERFGMKzm1JfbvclhM
5QZbp+bIo3dHzeOk7SQnrlC+kxd6KYws8VEvIK6BrOXEHF/C6Y8SGEatRBug0srH
Ea2TX+I0UUhpCVTosUJSqg/oZQEsOZWEbjpDfH58JMdF+LbYoGDiE5KXcMZv7sVR
6Mtarm/0ztm8LFqugqxOhJXwnQERZw8GjAoIpx+MsXTcR+GhXIqkTMjtYmRTxAvi
Z+n0EYprFqJjdo+siLxnASyjfr2aWXpoYXBpcJKHtiMa21F3A8Fk7wJSAem83nUI
0/qSZ5dIPWo4ovR+zdrr1tsFR5rhrklQYepFiXHkF5MiBgPAIW8OVrvlXbVx76LS
j82HBjLUZoXNWkbQmB11EqT5/FXb+2kJQrsrFQjcM/T0vtVVZrs1rgux1N2pOfJN
0SJaCz7RBHeT/f3yfeU1wQAH8DkxT7znRSbeDak3rAfabd86lsGWWbR5ZS30Up27
q/YPkjjHmvbiVEVcn8sA9FZ8uQyvYOlsEpKXEml+fPNGrrMh09uJA7zSIDh87B1g
Z2wpb5EGx5ovP+dH5WOOWBRj9BuCjw0Z7yuHRUDuOnTxoStUIieBkTiIvaVPGDF5
gjSlthkG4nDwVRAI0l+mHICk3EKReN6s3TZYrKqg4rpo+j/avQVN/ammSrB5qgfw
vGQCfIclzoPzflI8h7zmsBf9uqCpqEwyPNmNaMZFMrgbg/looejga8pjMAkNLleh
NyBNbJam5a9F4MHbru/JBr3qVYtab/iRGdQ1vAa5IXKqARjsJvB4Zlr2EMZqNKOH
usmPjhn2nVLxTDPHplmtjL6Hu+WvyCb4m6+aQxcnyCjWQHGeOSJb8c8tzcYyHICb
rDzBqIKVTVVzxa+xt5A5iuoLrR6D/QcUVcLkMW67L4MOnwSVxA67eyGFEnISoPJ7
fGmZwSWKR4x1WlIM5ebZ9vimAWt7SRgFTheZaSdkYz9XK/rSqLTLhs3R2g3CfV2o
ty40w+dzHX9ErEsfHu3S+0368hiFWc6JLq4yLzmPi8llviiI6pzJ3Ei0MvOVOyH7
aEPOQooBUzg42dqlKoa5g83IVu0hnZrMN15sDIS00dZrEDqdQMnAygEyIffkxdJc
GzbFVly3POK2pKodVXiwdMI9gu28ECjyS54VFbnJueX9xZpuvgDaNCHlikfSazMN
GAe7Y/qnhUWe1u3PDvh++CoCSDebxSIptakqMgEHMzF/bZQZ4fUwAnqHH4Vy2/vQ
plDnqrLxI/PavwsuGq9rSiONK/VwhtvQn8h86TO3inEWxaUpSyYRVuL/7HE7y1jH
s5GToaKL7FEEnE6fuHOuQ67LqjoXF9ol6mKZ/kZA5VCMuxnck9xhC95k3ysBGT+Y
tuASg9dKWtecU9xNSc5uQnwl6Kns6Kh6OvVKi7wOYEVvZTjzb7PtE1YoZJGZ5iZJ
nzyMWRcL6244gsS7Wg93Bp8E+o4m+3HvI7BQbkBtgsCnngvJ8EEjfniJhIbENmft
XmmRzktW1bzWKeh8n9KqDWtkrYWRvMjeycmH02upYbGMvqNhJjxlw7a75DH84HCQ
JPuCvO0A9rNtIWt4RWotd0czHtxkKZlugEh3rvVuGyXLgzUmTtVL7o/kcgv4BvHV
i/A63ELZ1TfiT/dQ6dq2IB6zNDWH86zf9i8i1wyg/9dRsJawslkO9Ac276RZdON1
Z363wMhwdbQnwh4yY0BRPfEqz5d2Jz69uWwRZ7h+/NvEteoQ1Y4LlVETZqDF/D1R
6qon2wqDiQ7ie+J+JWEM1VLncLeRQzbRT6OCPWxyAV19oJiyjqisL3HTzZ3MJbUE
e3ZkWJwSBokKHlSeX2OAF9DegfwS1OX6klb1fV7c8K2uUq9Cn2XP1C/Qh6c/ynNU
blXOfABc9YsA+B2YbZ8v+3f5acO8GLcKdFmqZ5MryfdiSWFt9DdGAXcZWQnyYuNo
cYU1JHRMlApfFXBjkDLeJ9OCLURFJlyuUS4x3Pk7uuLUQP3fFs5hFfMYjBiIeY4S
VIRHRbuyQQ4y0Iguk7l1iwpBH8mL+V1mJvri90NLMtUlFp39UOOMlHckrGYm2MiJ
GhhM+VvHjI7P2WSkpodw9lMGJY7BXV12g3wljCDqCB4VskXSIF0Oa8AyqKazfnwX
2iXj/VaVzBStyTx61FdXgACeRGRZhOwbNBngOoq2AMrPVsgXW1+EBCCwYGXsSKSt
64a08mDYYmIzO3f10E0FlUFJ9bXyxhE31XmAyFj0/KwX9NVsIvk6uMNSqKtupkiu
Ael3Q934lcmIEONBPQ2qBKvZ4NakJVv3zaJi1nzMZr36gqIjGyRmfurcHbxiyPxp
RcVDpA3pNd+drwlsrOGkNk1B11fQtI32m03pS8ZVbPI6ZHJDqh+Xiv3vH7XKws/j
RkIOmVmCc60g3RPes59CBZCDIEYj/CmnosxCBdcPNrupItVhcnIHWOPPlv8wTf6s
jNUBk0nQ2+noxac3fTjKnC8gbBF7QHZUw1ad6ANV4JpFUbARHPqmgh1Zvn8Ti5KE
6LDOVZLSdcaWlxGukIkJTr2VJ+EMkOsA9tZq+VovujQhOYnS6Z8yQ4kwC07eXx5N
ImQhdlgdJa9MUPDyUygbCJHXjxUU7VzXCRRxSRHOq3MZawKSNOzKPHLUoyc2gugV
7B0Wfr6by4YvukNoHrj9yq3vu7zImTdYD08LA7TAsitO2SiWGyViIqQCVbfpUGrn
ih651q9nZGEGd02HTyL9FwWkTVzgWq3QzsohpHB9UQsu0Vd6shHcHs5A/SFpNiN7
YNkXLWI4Q+5ulmvMe/T4bPsCC47qPyG+//M4KPSXnzbihUOnmtfiNF19GDZgfECg
PTPs+MB027KV0+3UeGAANDkMSkHYwj5LP1AqtxveRPGXVBseVit1ME+xnvTOOa1r
sIrPe5Yvxnpx6U9IPKCHnZPyBDFsZJ5fBaVxnKmKe3LjDyDnxhvCWuTitDQuCx3f
kjKi8ic7EEkp1wSLhgohZV45l962/p1ZK/30dNvtGdR1dFyHUn7bZrsKQ2Hlh7r7
YxnJDVd6yoBl+aItcyFKNfhJJr5rbplVJ244yd1obnxzsNfdNy5IPesNIneXsANh
ZwPFaH3oGlaFMHG1pUnNJnyf9YSN0gBSSUa5DtptiuqPqJCkvcpaJmh40Vyz66h5
lPwpMvIzH2ShVqOfcM2DE/S36mAnNS96ziIaUsJ5cjk3qFH451Rt3ddEHe8RmHFR
qjJ+tfKoi+KEiHxKMInR+RoSgmcCaqzruYaAqDr6k0CVxL3l6y5zTwFw9490t6xA
OBb3WHaF48lFNkow1CNYBl1ZP/LB/iTSjXnZtL+CnL/BdZQ1Etvbi2z8w7oMv8kl
RMkrhi8oOL7mqMOdwoqLVFhLjpTEu9gZYOfnJCXZ3WQCP23WGVKNSa41gLlMMx28
pbALosDKnW0G9VBmr9ogH0zYSdEae6hsq/eAar1CBhU98iGdgGAJsEaBvMppquoQ
w/tz+vi1TIMgj/Q7erE2jZt6myZgHERyzuRtcU9U6OO+BP3gAyCPotmV9D1BNFzQ
LdtZbUbBVyy3P/jwCaGxAbfKWC2w/CQVnPGzusWgyMzkK2vxSdemsVwp7JKGnJY7
fUio4iFpbXC6itHN4Sz2sGbyZTo/rGraOQsQYHiVYjArvL9/g5GsseJCwbW6JY70
CSj8o+GBi8tbz5RQt1owtpX818sRnwNmbHX5oc22Om1fS/Ccgkfjam7gd20YVu7N
HbISjIyEtA5FppRKE2Y3x7OkT+dgfE7i7rbq4cuRTJY8WnIZGj9Yq2kZjY4pnmDf
V3yprqc4Yk7TReQmqgYq9cta31rAFhZS73q+KaF5nA5Or0ehv+R1u35x/UojngbJ
O7G8X6iQxhqbPOmYi5HWryzwlOf8VWUWs0a8GB1RSqMvJM8zr9vte3nBMYphk2dH
PAV0FxphBjCdeG3MkDm0vlJrL3HrRB+6itT6XjGxkRB4iOMm26UrAEyNEWH495ol
CSboswg2e/ZmPzNR8g3fTo9g8v3Y1SCmBi7pEP8LBy8V9PGchzrahHRn7w1IXkjn
RapcoxVl1F4Lo67ItaXAgUTISeobl40OE0R4dUoWnQmakcjFeuW7l6aXVAPtZ1NH
PYz1dBMhtWuLqxQf3VXs2oISj5WLLGZNYL+pkQz7xzDXxhJqgDlY3sj8hE/PC4S0
/IXYLpzwBv5K8oS5zJny5gIZcgepM/PcLOL+Qhul+XpnYTGlImsIwXvKr8jqAT7Q
WnaGEqgK6aVlJkzD+lznHzOM0wZlhkK9KPX9xobebbMTW7R+wWdVpdcR8Qz/uWOQ
DvuggI6K2PrdNpTzGldkpjmN0JdI0p5Kei9s7OxeHJvtYmMq8m201JMZRXD0oDBa
zq8N3lwu0haKkH69Xg7vjJrgUTypGLOJbVxBaeDZI4JY8rK2gHHGC/Bt1Jf1AXkm
vXeemM5g+Zr+euxF42Q6NdFIPTAWqvddA5jiW24th0QeTvmeUPuXEbQb3+2L5Xyt
/0bQx8HrIczq3SLVTKny3ritNu492pogXZFkCGVVsYpvIerN7ATt6+dpgXmAKeDk
mMkRnD+fw9tNsif1/e5ymIWUKX1mKhNuRgJ5Kv62olD9UWJC+oiSxnm6EDVqr191
d8VBRzcZq25khzDxpH/mT5+hB9lCpe8h++6+pmZ1iHc5TTGpD0B6tMSsoYf0GVv2
kyf1YT62vqzzpXZBUaHZiF7VYAvlvoZ+vS0TsNKcGNVI1wWLRjiXQJdYCMg7v6u0
oSzOk3VfndVgAAZnWSs/cowL3Q9ASlIQGXy3DXicaGfLqPxiQflg6T+UZFmMWEI/
QpUGlV8S0+As2QH65+QiOhxZORnxe5YZwQmkztV4DJ94k0iGGtRWl6tajA8dZmk5
6CGPKAXqfRBZFeu8RNEBQNGfn1uZlqvJZmJrBwA2qtDE/P3sJywKcjdl84dH57Cm
fotwhRwO/dQzp8RXHXRIt6GbBv0drh3XjvTaLVkXvst5mTjqYh81JGkamhp0mHtV
Fw/MLfv374Q4r3EKd+g2fOElF0jV1weqW+fAYIVeRgM3gBPHh3nIRxK51FjB9gqr
IKObctSEHh9LRO3TkOoKF/fcWN87PzMUc2UAqtYl1FN5MHDKIK1jE5MMS5IARYaC
oEFzFqcds4VFO9Ldtgyw9aRz6u21/HhhumFpbdW+wp74KKFhvpQgUSKyJUxPb8kf
tqzeKYIHH50DncHYD4EOGJ+BFJV7XHLUQbs3VnH4rSgMBE77bQ0Io/y38rw2gutV
UXHl/A9NedocB3o8D1VH78AWzlDSa5THRascLAGDReMf6th+s8ibEJLlinFdM4Kb
jU3+fVtzAmsgHrBZC+qVom4ftqkyVTI4xPLR/Q3WPWjSjL6Ahi0LfZz4u81qZ1lC
MwD9pxhw4ewCKj95FYkxTpJ2Sk2l5dsd0eTLmW6qBT8s928WiQw6aJfT/AZeUuxj
YaYK71L91rv1HD52ihhQ1YArhH+R3zi0FXrybpnecHDnqxVD+0mPhlSESfBcyqjZ
SpZZ3zn+CCMo/AHyb7vC91e65y3fq7FBTzdN64QBD3TiZdMXnM++XTmdR1vMGVOC
m28N85R/oz8zzC7oagUCPNUi4xCPpdEIcc6IXfgDHbpG58ecWQSY7B+Mka9bzOJ4
59wHLq/lshZYB1ZXN+mYMjyfCm9nEkWnxu/nGihLWLPL1e/NJga2jO+DsSl2sU1T
StVBw5fXCzIuDzPKVuJ8jb6w56nSj7kRZei1ZXq2vExnY2IKYYqjc1OL1rZig1GQ
x+NO9+SjXVHxAc2Ttc5yJB4kc1KexkR4v3YYSoHOukoMqSlH7lFG5YVbsrFivLmc
UiuQ3coznoxJT3a9cbHeVEXhxwQDY13I4dTSMJovPgbaWh22CmiEhMYSuwXuqkbO
BH82+NFYb+Iwu0Nz/ICh2QJxtTZ1EW2TLctrLS9Ha2TrRHM65OCE8fWaOad7c/tj
DSjjiQqm2xI/z38aUPWaqnq/E+yuG0xNC7UY5FBgnlTSksz5yupcHoVI4LehbiIA
l09y51dP1Q3SbAneyDsGNtRak1toGEOjGMnX7bY3Qk9PMxLVBpKL1tq6JWOOn8iW
ugJVrMGRhsJDPE17t6xguSxc+YlaPdyM4Xep769g2VecO+63jGFjvCVuR92ELPSQ
0yL0bXpbFWXZAfxtmd2bo9glDaS1y/wF2G1Su3E8440EegZJqqS+V+C0+3t7RPvB
sRm1vd1qJHwwfmZnphDTUuzyogTRJbNEfXY5lUNl9XUgcW18R10M6gaGelCsYDm0
aCfuBddXgP+p3i60EXNt3FeAtieO+PBcEYnEC1U7v63OlnRlNKVMgRPNTrDqSYOd
rs6P7TUFs8nuf1Akush2uNk5izQ4TYamNDkNS2vlgCI4uuOketOBikjPv41Toko6
X5byMOpgaGsYKS3AiifeXjqTgmPCmFb1PHTFlJxHxBNarNeRgxCQjfe6eaNkmnCA
WO+8ylutfFWz4vXHSDW9O8f12Ie6opLDLuBSlP/TadfXxZXMg5TyKjafNe1jz+SB
Yw5M/NAAkocoGlTcKWn/ncMwsFvPfq7ZpQY7Wpm55pb2F72wPrbSFYKI73skAnhn
+gfb8BvqsOxIpGdyOTgEd0CXQr2PGy8pqK7tLrsJnjIe+it2sEVN+HtQqOb12M0/
moJhU/NBMWneVkKXdBV0b2Qu35dDffqjJzfDhzMZ+tUipwdyobS2iHZ1/7ZyO7Dp
s/oTFoOOevhQiQYDqBjAqS8vQYrZeAGHxCBYhhsYrCwkAEhGXVm2wGsehDkDzwUc
b/QsN0bfAPWte0dYakpGCk/mSRVBQk9EeuYMBfWkyOHFXwpji4k9EdoYBb5WOl2q
4x8CWMOzXxaCO/iLa/dOUUhAcE5S86LBxIOfvb2qMPCsFXQQdFl81zHvlEwvt25j
VTz4WIMtlhyzhjihm4oVhXx8MnW/B9YsAIwgMrKGffu/PW3ZNvBA1NI4jFbVsYbd
hNqn7V7gsHEJdRKMRSsPnSHE1jNcv6WauOPK9fIoUdFfcDD3hKE9ylkQTlqVTsIp
NnfqAR2fesAs9Su6Qui/V2b7TO3A0wmUt0VDjX3LKWe2R7hyeynyuvuYnwfwVkZJ
rbaX06WEiAmFKqUfRhZzZoLM/rHMQBkE+BxTuJ5iOlFBBNrGEZfU5fd7C+rqirXt
3glgfElqzraEMKMH4PPc356QlkzUfMbhTtu5EYeclZmM5OC7s+jx2RlUgkpu3Gy2
7WmEZ0K4q9ldLDDpluruMRvbbyXQoO+MvZ9lQUQJ1jh02z3MKrc9CMHIWdLwlpBf
wiiP8XhxAHHGhYi1S8Juyog0u26QoURdKPIDIHTx2aIK5ekeOLAWT4KQq9XPkTnQ
EyXFmGGRyeqEnmVTJubw4ro0S3Ug3vGhbYIaHBZWYJ2/ce/4MbZmDBK7tZ1R6+wE
+p4SPab2o9LCVKOh6fYK7howyMoFOsePn7eCQKVsmikxp7WfGsvpVEFdRK2ehD9D
yg0Kmsk65u9NIY8pueczDYFJkIpVK/nVE2HQFLmuO/eHcByyV2EXVYC0stHB2/6Q
ZDXgQWZAtBeHjTF/1S+G8CYyrsgP3l34j+9fJg2kCxKlV7hFmkQ7YALPekr97+bC
4UKaPuWtrnLJCuKaj04dGtPoawaioxYqiJByFJwvvD2+PdITjbplhgwX+ZQ9kp+y
nuDiwhFKgcOkxqDHitn6hzf3emshKZE6zYiOpHGV7/kYhq4dHa6TqaY610INyBrS
hvD6t3AD+Gg2ix94xbzfJl5zOWImoiLuUofVp0woNm2McMSh0EN5Yqbr6deFukyk
aOuJW1K4/xOPQlHsJrrXRgN0fdfY+xayssj7t1xqoqhJzjmipwmIVFCLTPQbdn+x
51Pz0iFgNvBcoiSy6wVQXmvFgahP0k7e13kR+aHcI/tHRKxLbHMOHwnKR3zl+cv2
kRUCXB7VEUb7mf7xOgGAydE6fjGTOaD16p7YFm0u/Efk5Ymru7TXz6+peD3zgMnE
MmojRxOdL7RCeE3ZA3AFNmj+VJn9xPGmq41kZezU3RWemWJnUk6F0Y7ZcmtHihap
/zCg1jKdiT5tNgOn66KL8kQzXoYkseoVruHUSmf/HT//Aof49Qlwz1Fbk6Mbrhfm
ymZSXC2lDAsHv7DFDNCVMcbwCdGN7NhAgJCglSKeSGyJrkjZdRB4GYpdK8Ss2xVq
llsn+USEp/OHsazsQdblX0A5P92uWC7e6tc8MR17vBuy5l5VcmXx8cbwBGN5iFLd
Q6hdnMARATiF2G578U+3jUt42msl7Q1ypad9zznyDt4PvYcQ6ok85pJKJ2gsTbU5
Na4JQpmW3gqnkKgmk/nCRRKcE1EhTFcfCigwehu580YjHRIZslKnYOAwRkhlWt5s
qLCra7FcDoWzI2Jm51ES0fg96RAbIZMvWetSUt9iAelCyeZOTEZ8eba6hwPHKPlp
NGBOXXpbNIuESvhcVfx3rZhwzSgnsweEIvCKNdkYjPTjGci/xT1SiMHsbdFYNMqe
fAIzne4s0/g8dntZIBngNAD5u7oAjNypQ7sPnqVM81vcEts3dFpvC4sXgaa072Dt
x95WcHxwvBjAieHCvZKSRfB3ButUbqHkdcoJ7M/snZawV5ZKKZgHycrI2eTADrM2
mW+p4QxxsB1FcJs/43wb2WAld1AHCPiUEdRFOL06safJYuFHW5Gns2q64l9g3nZM
4HKQSZsw4I6MoHCdpdN7Ar3GwCbxV9E1GyOYDi8PVqeFDU5GiIu5Y+I9gxgDD0KN
n4l1j6PbHWWH8sf/heC1GTkrCWnGkQNPGg6BtlGXr3buvSfC7eqN/fQzjOBWqfbh
b6hYX1n6BKyHlx8qQtPTgG/Xd/FBogA28tjqkRwNYpMUEm+RWDxV7whpxhKrPIHV
7SgC1CAfxKHl269QUSmYulNMfQf0XykCmaScfJMnHcdNtI26eKONQOaGPWcfsR5P
xqqj8n6R9RcICQeYw7Wx5r6KHL64dKmh3VoYZ6jGm0Mmwm0SJypsp+6pphYA90do
PoT+gRPZ9S4V6PHcHu46CEI5K25QlosgqS7u3rpBaa6IJtPVuhgVeS8bgZ6t7VL6
Ikdyzbnrz0PV1YgjpekcYSE5FllyzG1omy8U7tEqeJG03CgQ7GwuPxQogudCnzaM
tU7W5kynWF573TSQnrtmvVAVv8zm3DQS7pnf5pUk1Fb1p6HJ+b5rYXAGGWJqbWCH
KYKIAaCdnqJQx3h0we3TnzRefJ475pwUSQWGFrUlzh3dvziFGGLT/OoM1YMCHPHA
d1QIVdy8mJAnfRDerFTsebRojYuc3YgnkjMhZQH5d0gdSKuppZgzMHlybE8kG4Ep
UFyDqcwOGR8ebfAAs7BDRxkARzXeQj2ANu3j6ClvkgYlMZhurMx4CbVPFlzoBWtM
zSp+ARRFCTPu0OPdc1nxk/MtJ0TgUbEeeQLCnjsRtbI3k8U/80oXcXp5ly0wbqgV
wBP9Dn3CgKhv7nSyQkFU1jufBbciEzkZH12cdkzcNnxS4kSVwAauP6OOLPHuuAOy
dtnqN/QTi3SZmqwfXNKupQiAc50phGKSFquUu6tdIlZ7ys8eNAQLSfKjLP+sIE1m
njx+CFhVmfHKoF2AvR/a6LZKu/HmkqReLotBssgVhN7jjcHnGr72eOGhTXlx5nqp
+uWRc/FN110qnXNRy6Wkq/dRyvV+hJSgk+/XqxNt/JyoyPBb4MTpKUPevk9udJz0
Yikb/4OEhuJ3jXZMZuNf9ZxZAzXPQ6wIO0nzbbR1TKOsbDoC2FYnEPze4fIlxm+6
H3cgTyDscWRc5yoRy05tiDRRa/38lo6PA/XTa+L6H141eaez/PatP+7+qiDqc+Hp
OQmdMwcWwJlPcEUc4qFYF32dJoqtT6ydKH2POig2DJH/55we78CoU71Puysi6ERU
oC9K/7SwnYX5Df1673oxaQkkBTna/uqzxN/oUOjmnEDnK33h+nQmnFjOrcpLV9vv
+FWMPJ5wZv5slXdodqf2ocOPPywRhNybM3/V53ZS5VPD8V5z9VT04HDdSfzluvqB
XMdu6aOVTGqITtUrRWtAe5FJ9MfuVhK/kIpXU14cBuEyoLVgjXhnzXhHL+GPTyPV
Wh+yeioBOmLtB6me5ETqqo4mMHQqNypC0YgBWZhFGQh4aihEqUhwSWhGONX7v6pE
rmmBm4rW8rL+GuUyPx/Z8W5rKLG4F/AHb9D3ZFjqK8ADqWRdWQu/vKsPB8jE69dC
SJaDhgg3qmcsySLYIjDZn5llrRwz7YYL12fzpwqw8JLb25E3hnr7sx5lBGmHptdw
OvFOKAA5Nqba/UenVvofhnZB12kENxsO9p9A3rJx3NiVXRE22pl2VTxhv4wc8ad1
TdDstTz763HPF8vI4vPREnWWkYmi2HQsMNCucmdeh2XS1Jr0nzxnFM+TzzEHjsGw
5JGwtuQhFhRaY8gE7wxej9FHtss3Jrla3iMn2T17zk2HGooylyHmHt2NAaZ5jGPt
0cwE7wxvfEO1w5DD1oy5YtH/lyMgZb1vJHyvQxh2ezSPpB5kvzOsyQkzM9/Zyf9U
I6yVRxpgfQcLnfUs+2ldig02roFgWZlgl0O8HyjHucdlBX6+Pg7RydlJCG40gLXX
LtskEm+ylxFChyICUD7nfQN+EeE0nzDd8nW07VeMl/x4u7RqcrViMP2RSnBDaaEO
WiKGD7nJrJuJJll22QtjWvqAnPg0As2lJj1AreJLrcYSmAPe9lX9+ZWVYRFpsnCG
FoHYpJJalvH9NFf+NGvTImBTvQQgvt5tCuGGOW0iEVTK77jTCvnsAPjle7MRpRFs
xAzJ6ujqYtV8zmO9YW8svNR8G2o8IFtl2NzFCrbZEw54ASC7DSowvWIx6ERoLLYR
C0VKJo87PxPOkK/CDXjkx8E9PbRdI7AO+aPKJsXjNQK917UuEPG16xTamnK5YzPc
jJHyhkOgySNyueiQXYEYwVt9xAbpRLYundchsSpZ7nd5zykPW/mOfjh9T+036l7k
P+ykQZYqOQviT5af5pbK/4SWIjKk0GsPZipF7K6/5wqw2uZgLC5SMSURchcaaIlG
/8IlVHnJqx4ADzim5uYmIJh3eBZtXhmoToBBedeWJ18ky9+zm2wU4wVExPKmVjXJ
j4jI8vAs+jppq7EvS+fPRwXumPMsZViI1TNKgRzHHTjg27jcr8mVzmcHJULQnDh5
L6Ck1UTU7iDpHtXZq4h3G4hsQDW84RBA21VoOoxMu8xpJDA511vNg9loDFepTVv4
Np6hx9Zd3JBAUFkfr2bC5FHd6NnsrNS9uL192kGXkivktaTJ55Db1BSo+kCeuNYr
ZTs577bsxtIHwBVaZMO5SsLTGq0DTF/QQDqXNML7VWKz/n728EUU9VCOhgKTORHk
UC6Ce3/invd7E5bWK0k/cf55vwjgVKlMJs9MWiJlp7GgB2mGO6aOXfUifYGmKrbI
i+9JvZwWN9aD/ymvzEs9nPkvU2QEpI+yxW+wAuxCPDgGdJZaQRyQtPr+06DuufHf
AgjF1jA9TXVZUfzvkVg+U9yPX1N6oX+fmBST3VnItwJsxNsUqwV6Zp83R5eV1LT2
sVwfvKnyRRbvp5IHL+YGOSejsags+wgKHC8yYm6b0qX94is8tU0iTVUw8jUXDxBg
rmrJak47FsW77H0BTOqNT+8edHYT5qlQj6x9DixjO+yLefdOQLx3q2njPtMw07cI
b3YefkZXZAIX9p/mJEtitBqB9j+PemcAQFGSjILoiPpAa7GZdUDSsCnlEkeWcmQd
+5bGFp7hs+vq9Ow+MYZHnOplPVNs31rsFsAVjnNVTLgZ/ag/SWhxmprvTwc83h6r
al01KHLK6erVQ4vsk5gtPNRpvsg6kq620zZk6Kqsf3kRBbp0k0EMPsT1PtcqxJQy
BJdGK8ZDXXc7iZiiV/zKyCCKs9m4MiQ00RiE0/0euNzEDmF0Jh9CaYdvTBJKeqBx
vitdeabF3ytbaywnGazBL4WYJLDzs9zhbdk9NjwWBDynmAgEl1Ezn/CZC/wknOzA
kaq7F/UvwN7iGzYIwLzCWNnGxxRQw6lJ9yEdD1lS6rLFBFHHi5xOd2BjwcV1R0Ca
XYF/jwI4fKvi1j0b/EU9Cr4JF3jomiB53OfhtNbJkHNTD5vu9qiAaWpwpUiVqOsr
lAC35uDImM7B4uB+ufk+L6A0ZdqMXln0pqSLUiy2p8G5j1EEJSVgxEk/yAaBjkPi
Un/Ua5zniD26jIKWLWlWlonvKFvhdHxm/FUshunTS+ygcJp62dfd2QeT0FZLcbNV
F2EPGygR24CqLlq1ylFN+gwJvlCpvA5F/iQuNoaSUCUjDF3YZ6vDCTyzAImbv3zj
DRtbK8SvwhQHCNrHa9bdDTljsXL7sd5uVLM11+p1DWuIONCbd8l/RjJ9fQs7CJHZ
jf9wNCzS7spid1ZF4cn6ytUYMzSA9OFSCQnCKsC6dtJNnlDvfmekurU8Ydr6RB24
tUpzC9Ry72kho7K6qYcfen22W5JXzek451uKbAg19hSlelrzmW2J6hzktLnZnp4i
r5XhzwQb2mt+BEsFljBTWREsSGEuS+IFrPgpJ7ZILMRuJsJ1cBR6R0PaY7qSrXmc
4qIYpaBxgvGYhUUvEZsq0IX4bzqm/8v95Jvyt4Y2P5xM6xSCAUTGi4Pe8f7xZ/Rx
qZdwdua0ypM6XCx80pdxEIz6YH0JiL4n5wQ/ln6DIkYCBawhZWwiM9o4EohuE9sU
CW2Ok4mI5Bc9WdcFcPzB+fuviVU7MKE+6NtCZqgcs2M+cpyTgsRFDr9AQb20Mjh0
9QBIn9MAkJN4Ri4ul2dckvTUi1wl7ZTXPJkBwnd86RisKpEjs8FfhGebSNTq/APL
5GZJwnmtk5dJDbmaNnpO8xzpLBxyzITubMU6m3sePXwf9Ttpf/1Cevm70+TxPuKL
0Hlx5DHFCbu6IaC5SY4XONz+51vMIUnQMSWlvAAUm3MJwMvk0A6DShKXQn3cGMUx
XZPwxAqO/NUl0X5UNyfjEoPrFyLgie+9PNoGMI/2WOiAm4UW8x/Ww09o8TDkKf2b
6mbvDb2ank2co/TFDhTbzOjw9fl/AYQxXGfuo0mZ77xFpK4S0lf4uDALMO0lbFIi
nave8Nq1ILztSsQcPN0iKRF1maasHctH6DUjCqPO88VRuq+V3MwB7fKhpcCoEH52
8+ArDB+Xrk8lWeSqDLgOCNu+h0vFIHDCAW6f9QWRpIZMlYMVpqVE4UDhnyrnOsFw
rMI8MjcPoTUKHXBSiK+jYlai3z0Vnm3l4icM/ilYEo0ctMPU91EJwADXmqT4qljZ
7wykkQSBUitBAERfCX5Jce/fdhQTL741AXoW0ClNK77NGDtAX0mg+vTjH/ml0/9S
ZA7L1yagnlY2sCHP15Z3A9mYPURqSdY+n0HxGfZzLQNyJt/4xDoDZN+IrGygzzP/
CbnfxZdGEOjLe3u18nHX/1NOh9wRFigTuwz4SGkipvdN+ms95/1XwC5iTUIJRCvK
5n5i1zqmOSHl4RVjBXz1lWL3d6yq3ntmAaC+PzGHKImDkn4P2zz4Uufj129oiOFD
pzvD3QRBKlO5zyurD8aqNUWSFEeynUkdzk9b01kmy01mxmWmvqvqfW6jwf4ek/07
2XM7bwEX+lXx1s6kisU4wBEgu0JbEDoPCIPVgRiAfONA0zuC11xj9os/1fFC46pK
Eaissl1+kdgHdvmZl4PZ5mzI+CV1dJLxEsSQTREg9EZoS4MbqOvJcrIV28MuTPZK
wIoNpohI6f052/GQPZdH6g2av/d9UtIqKSlI/KI9iT3MBHd5PD6KhM/12LOk0ghf
d8If50bKLCCsuWNA53l96477TM4mi4aeLBLAfhYdbLPQvIRNaPRbOXCpjGuu/+tq
+XrT/UmdWYcNR8w7Pz6+QWmyG0X8UpwF3FvXaeivmbczBTy5xeiGNNCbAn7oGbbe
v59AyYe5h+qwe9ZIqfs/ZuEJkWcMCux+VMlAucPWj7wX3sWXM1wByws2S2Vxuvab
2FR9YxXLbvqtJgHcUisg69wPvB2zfmxOu7VgCfuyMYj+VNcZDb1Gho4T1pekERh0
f7MHKvFwQK2uzTWyvtBGk0A9qkqY1olji9HyuQDOBDadeL0bM6YJJmepBirqqLuE
7T14y3AKIgA1hnjlNgTirUQFmRKO5oycPO3lYGZGwya9xG2oW1OrWbywqzSSCHbr
/EnFWKu5NUQdgRNbdcVlZiZtVdQ+lPsgSXOvKkJt3n7H6wu8Nfl90vonBrXW7+Bq
vCquxwMtE2b4EnQH0adfujNwqJBWtRMXxgl37WA13vSLD/4ptJlbk++JIT/OSfQP
+HDNon24c3q//piLW7pxLgkRZb2HTTBCVlBp8TyUF+ycTaM8Zwr04btL2ac6MbW6
XqLxfzG8JoKiVTVfsXClZJ1MVZFHBVppe9g20XAWbq9fRu7GdDRjSQq/FsTiYzd8
khVTWSa8akXiUG7kE3K8hxBMOUcwk3fO1avOiZkICUfr9UsteOANKPIPiqkvXFO5
FY78SAnHZQn93yySBHALewxOUHAxWS8Wvwmr9WH9bO/U1TS6t2eOJLFtbq+vpGtu
W72h9vEGu7sllNckqWp61arHbU4vVsTHtijpdQNyVIJspbdeK1mHAVcxvvC/XDEC
qSzb8rAab5Hs3pokPzL2mGT20llHomG+kZcGlOaHUuxmdu5FtTQPvHLYD6s+m8qq
MgmJY7ziR9iteQCxE7MIy3HdCYShlhSbiR/wLV3qs1iRjyVpCaQhys+ey4pPQKoA
C12wDB0rzOqJp1YbQxf//1M1UrUjGzmOuODDRj8LSo6guu6J+3cdei0A2d1cpFwA
bYWwuPIjAxoOHwJiPjIYqlKzDbP2R7wz9telwTPbl0UnrNjt05R+EZS9IeFfZqiN
xDL3MNNe8nTO4jSm5JDUFUZbcLFeWTDGwBjeJTDNrN0SAHRHbwv35sEhPkyXu+SZ
YDZeV/YdzPyVLS+0+SDDLA5K0Hn6qhj0RoGxj7Zh9n7e1+Jg6jKqdMp6mASQOk/2
TAzoWcuXytjDbwu6qotrA/6rHswIJ1INSPTw6sP/UnlfyWA0mOp9KlKx1JdfZh3E
JFafuVk6vRo98RCoezxPjY2ycuvxVAPzdXw/6eTXludMsbhx8t9zX0g3R44VfxIC
jg1m9lvESyU2huyDibztJlZ3wE3axymHYFb5wrIaUSfZz50Cns/ypzpYlxOHYK7l
YpXa4JoKgAlQNDHMfsBl/zjjkLwX6f5Et8UH/LupqZccBITnxV6wAbX7BMVbl+iE
O6RImaxa+fK2dYSi9I80MjYWsT7hgyC28s0UGm48LDMl/bIEIW4qVI+WzUeVV76Q
dbaX0ydepXLGiiHdT2fgDpmQpsZu5usmwoub4HZ3fF1zQHh0RgEGv5DkWtXdc3UU
iMu/D2Txv+umS3IcbB0rJ/P/sT+EpqGJhIpLaIEavlku4+6z/5n3dovsILIPHvE7
NUuk8Jjl2MTbZiBTjwmHjIIfdy7IdFpDdUnJuoXKnybIXlF7eqc44RQmPZCI+IbM
NohyCIYvWqhD4+wR/nxqn/N11y2dbHo59+12tpdoP9UFnw2glxe7n+b+eQ3lTOg/
jHztRnPAXMaW3B6nozsuoi325dlpy6lvk5LNp3nfOGP+RYuFvWB6r0qRNvNJZflz
Hg7q9yA7qSdbHxlDiiHLn2l9N9SJzhaVGtlpr19/l7/23pxUjAiy9K505p3iLFt7
fCA8Ob80YrPC2Qvqx0oRgDI2ssCPnENiboTTwHi8GC3C2zs5JJXiSqx0bKzOORMY
61ozlsmxwOOp3XP9Hxfc8FC4Mdyu1w1uLXBds2rtkqTuYcoBPe9a44U+JwO5KhU0
zmh7lvH9ydFZ49R6BKG6fPK3snQAaOGC7KQAwfEvxvZNCXzg2bJB3Q8fgDu+k8XY
eTskksHrgMr/UnZ//Mhcy/w9JwDHyMJ/NTuRDBm7DGH66S6RJuaG4tj/pKDH7uBg
L5TI1Dmid5WnTfzERzAwBuYdcpZR556Mr+X21BI2rI0KHl1413A8fFtq6lLkRVsf
miriul0KSZwn8ePRqOUquMrUjUHKG39y4oMJcTqkeRS0nSKcGf+1DpnK7/j4pngX
yM/Z2waAtMklmdvgEAzE9+g6lQ1uBZCG5+w/ZCCo2DoE+kIm70Gme+PyVtmgchce
Wdi6hCvsezPNEwYxUttZ1kdSb7r5nc+8zvbkihBtJXzXrwLahjgQ4uOHF+snTIHL
cPo3x5Lq+EtO5V5varNddwzJ1ZsJvkTOO9Qeppp5XSFgxHxWFUP1YREy9YhBN0Lf
SnWZ4TqUVUR69UQQ92XptQGwxwLd5xg9Kni3aEXMV8HUfsrs9N6PGwpIg1KjAI15
S8D1jOQw5TCp/eQ0g8Tj+veqWSu2m6rdpRFtYKisK4BTrb7jVOFJhqb13Wxha41h
aguIMK2PLF5IFgSVAu/+X3vjIsfFEaWR4DV14IdUzNgioQJ5Bup+4y0L4R5w1A5U
Ao155R9YgSJPromM0caJoviPPFegwoB5gXX+ciurUG4Fwmg+urgvEnoZ9Fv2E6+x
wtBz4mCcNyTubl3MVg95SM6JwGP22WDdx4Pn11LeJdGue/XcGEA1H/LOYF+MRArc
RVjzB7L+kddpwtj8Yqvl9sILeS1wtl7kxwjKNEJblXXroVNQEWKNdXYcuNpYsssS
ywrB6NmT8GM3tFq2OpjQ5U7NJneVY9ovwpocnKppVqB1Ryv+EtD1zdfS3CrUzWAz
aisloD9YIpkDcFVHzlYsdWGtmdxdHsP6WYGMpsgTlRw9SyQVHrqisUNkgJuJVsO6
DpWJrfflM9bl8svDxNfH8MiaqAsdDEytmDZI6d4xQ3quc6YR73tAFdq5FpzE+Tyk
En9hsU0onJ3w9KVEFpwA/7fIQRF4/os1QU/7r2B2XS1K6TS6/6DVM9V0LqZXKFsD
PU8S9T/s87RhkL27Zdl/BAXI1FsLdBHFguh8CGxFZ6755JLIw9YCfMthLcRSRGpM
uhg6hwHRtMEAoQv8/iibPljF1VcNVPsCn7kcGVOSw0aYECS9gwSQS+HtS/65Dxu8
EcXZ0XNjmITDRaif6vGySIjeBbycx6WzpXBPhZFs6K/Rf+PXXoK+GefXZ7U2J7no
aYMyd+3lcyrZ3QJeJls83e01/5ZXlvJr3SYoqeW6/W//kUz5qMbq3CjH+NYGgoZx
b6w+5wfJivtflBfIQJupnonEJD2+DHRYNK/X3ZEsWVO48ZMJD+7iivLONjjFI35o
E+x/C2Hwxd/msUczJBlyK7DtsZdiwYGZaNxyjkm2DWXpJwwsUJl7DTy2rkAb7BTc
ClkIocmU6IovhJjvJS1csmpA30z6cIcwtMM4wx2Y3kgGf/yKu6TXsWnI6NzMji/e
cpwu+U4Y0qlznZoAU01c100MQ3Irm+3/jxGc5t0s3gV4R0Tb5NCSNlBMD9rD4/nb
aj6k0fB60qzEOziiVS4wOU88nA58RI9HC6gl6LHkFCHse0/JYlRFxyGWeRSD32h8
yMGXvbWISaNqStEyDVzgZIwt2inPg4XUeyNKHlooe0WydnU8fr6HyjSt2h+aoT0Z
3pc3qX8i4Lbwb18d+GkHHGADkQ0mPVnVgsIXf0TrR7cdXZaKNbh0JB4DP71L8ZP3
OzUCus3JGMAbNEIPDAno9EsQrx98gFPk3sTiZjh+mn5RqU92MyldT/x+vu3UOtUy
MVCUYgVzHdEELPQsLxo8hjCYdp53qY+a/4XCK59DE+wr3m0ERzhzm2j0xgLs92sw
kNWPWRuH6ZTemmjGCXatA91Req7JcJyixyGrBj8AE7DoIfQhx5AvJQCxKsvcroMw
jNZlAt/rUlssprQJeVtR+ENGC4oYnRNKXqh2eMkHOnzVWdzdX26NN9CjiALhOFNX
V2DVOfVorV9Qt+x4OhQ4ykHoyfvz6rYRmbN21Z2wV6GTiVqXMeYGULiZFxgSnSXf
cu1ZQ4GU6fyR4+QRExnPiYEagk42RMF7o1jca43+CKYrI/AcRPsL1SJ5aZck9xbZ
nw4OTQmJMdQDhCTSDEsoqwnms7B6rTKZgnR8P5o8gwg5wD3y/K3wvTbyAvxoU3T6
fUtTkg/09i6UYCWhJtNn3RiSX62HJRJUiw0JnKPhbf5PGkKSHGNjFzAMQmXkDIbI
3kHXX9OwlKJdesLC/znJhA8uZwczU8Ywidz16vvOoYmOFNqipZ4Ne/tvE9/DEZlk
4U/ij0STjeUPLmKQErPDbNxTjEioMYVQbRllQgwo0LxXLe4fhbyJZqovSA5c8UKa
1xWfv0eFu+pAnwFB0PkJInhitpFl7R7h07apmZKvMjBGgzP4zaSWlN1wQb8T8jAe
KslhsMTVmJ7AZa8bjGFh2hQN3wU1jyyOHJcoSY7w1F74JoIEr4Exhc0cLL03sE+5
LLkSN2Gz3Fm84z0MOp6otumxLrhT/21jalXvvq4yc+m8Jk+rxZhwjgcm4oTkaLBb
3MidCG/ey6w9Ji/BLa3IBSmAJmVf332W4dCVlAkWPKSX90xHtAgXl85TfvHoX+QY
TuhVeNus7sV9JKy9v5HPn3MmotcBwepgiYkKTsFPF0reiC6n0xSmVkS5kS+PipHF
mdVaGYD77nEa3qGxbO/vSP7+Ni1Kegi0A+CKZxy/kg67cYcDEkgsbTPVFKAjr5US
FQEGaekQKsX/RL2Wtpwz/lY3ArB5EIfhGbrkyPQ2hT/Tz6S+3uIC8RzBGcKe6mPH
8Cv918/I0AeV+r79tAiPfzVeT2Ha74bR//v5TBEGY5+OFcsieIq3dnjzhuZhKB15
k3DX15NMGrxxj3SEq/UKenlOV+mDShZMIlEofWs4c/LTWsN85y5QJrQQPIqRVbET
wIIAFYr2oBNCjvNMz9mgeYv9f8X24iw/ysVOvxQZDXRajCKio7Pjwrzuy1LZlldU
PvTXfgWJYPK54aW8Uv1xuPHEraKOU6MDcSwL5rhaDkD19ROOaQiJNKEcQWsiY8Hd
36heE1oEdr/dq5tgwO3PilkFHISiWSLQ6PatpiIUAd3oaZUpz5kGholwBD3WpKco
2OveU2Szs3cLzMsX0uIP8ZJRvE5WedYaiMZWjj6yTEGW2MhpMb7ffzIjjETTJ28q
RCv2G83DGeYQSQWiIDPackYprFXLPsYY6fONK0OWs2wopwa7LenbE7i4+PmdMMsZ
Q+yiozc26nQXuulHP4B+AZpmr3Wbh1ahQhZFTy3O+WI//ICX74DmhkFO5VuXz+D6
JylNhusIUmE2VDQuA6d7gwKInp+bmiOTpB4ho0dXGWEFmDhNhuMqq8caAZybDc6Z
k1mPaXxRruWhj8kJNeq6Mo3p12XUCIHA3VTbCV7myEcJLoWXYvQgPhRRftVkq4Dp
RuTFCIrEloK2eOyXA+FDXy9Jo8Ke/HFiVZx6/OyRpq1zLVMAc1xf/k16eA2g2fn+
/NwDO0pLd6gQioNXDkXhh/yYNq6m13cxLG3hNptCNY5M9KoxKiY0B2ga5cd0Z6bq
Crv502xb7jH13Asv5sPeq3nfKX0YfngtnyQloThCE2KCgoJOEjIZALPYqbcckoM1
NftvhNxdcbdj7jW8oDAkXzda7Mig5HBTuVsYknTBHbrPBQgvUeWIU76liQGSCeui
J0dqVrlqoSdE8c2YBPoXvF/As36BXF0Va+AkwBAWc4BUOhWdyKbdGJPgBuJvsTD5
PEbkURz+kVqsQk7v0IVXcpfUjCVhV107mEFYdNeougJJcimaZ86a8lrXxvl/L4ZI
2i+Y8ErukW1QkNq+9QZxDVcDLMZSLVxodDzea8kvHSpZ8yIHgQR5Mv0Rzg8iubv0
OQopzuMICz8UsfzFlpc6Zum8pQmAYf6BLUu40ZElEt444L2UnuuUeh2iXGr2v91L
UGKkF+8hIxtlPwLHcsgz/JN976hJmtjuMcSnQBj6GaOawm9fDRJiK0TLPWoPBRPi
xU1cXyUZPujN3Cq9vLTsi0e7wZudJf85p2m5u5CWMqnVEBof28WTXSKGzHxtUqms
+YvO0w80mU8+VwdqOt7rbnwsQAHDxRLFa/y/D15iYBp3prIte1rGWhTKeEyMtZaK
JNnES+30sLGxA/O6PxtSUjY0KBnPWEQ1sUgYVpqPFSjB89XtBB8W87U9t+8+FIIu
8I98j9xQQx8oKGFvCZ3UgR2Zjbnj8xzuIs+WBEwYcC3HID1OKzB9yS3BhU2iWHiv
eQVCeEj8dL4oMuXwo9I9ZhnemL8V+7yAMRqbVwx0+dho6dx0wmxYGCD7dhuQaBS0
L6yVLI410GgUc4uAg55tfzxNY7BbP0imT/GohZsCXZ0f6GJSDenpgTwmRFn3o/Jw
VfqjMkwXnWOELv1NqO6kCiXqOA4TL2yeTWpD6vNenzKdu3hD58MWnt0coQGTnt5u
D7+59KOtsDR21zNgM1MJYcw0W+I/5r6QMyK1vmVbcM5z5orulh2FvXvbJxd8iCQx
3leOXsPKmmOxh4/crz4hVJg++fEb0gd5paeFCmE3uHRtnntbSiUruJbR117cvo6D
AiY37o2Oz4N/klraMBh9tZewkRlXt/9NECQgWo3oP8/w1RaZwNr9HHT5L+5/oRML
coOw5Am82ctX6u2taPX5bf7d7/u4/6rOzKgvKJvODj01J/04RowBfgzalGl01pdl
enMbvxw0ePQVIp6A7GiR7lBxRR7FkGvHtWirv2Dy8P4InDq/0tl6apppT3I+7j8e
lt2dGmJnxwU72Hs/wkuECRH9BTEDH7gZtUK3+Dkm31p+ZZAtf9jm5ZrKd5Y15j3z
dyaIBnAVkHp6aHlqnBNW9juhpfhz0+HPjI2Wf7vWx+N08yj6tBDHbzT9EWkkqVbA
k7EGbdhIchx+CNPHIkW6pHFE/7f4aP9V6Semg+TRjdEx+LsToSJ1+ezqVre/feL3
/hddXM4lGLFRMXX9ijcOkgYVvUMtVCn0GC6StdsOEqY=
`pragma protect end_protected

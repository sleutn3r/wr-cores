// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cf8ITUnp3WSY/eDwjBk5mFX9kG4RnLVqXxti5Tt63UQP1QW+EEGoPAOvtTuO3T9T
xnxLxosBRpFq3pKzez26TiPWN4dST3RW2ZLzvtRl04Y5uuvQSpArDuqj7NPK5DAg
g3kkXLia518gq3aGs+WouDTkMuZekwenL9qaVI+wtAQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22160)
JRrNYqKzkAfEUqopGJ7dPovNTnQ84cInhnhO3LZakDYn29wZPYXW2svG993Au/7p
IDqwBaWq5AubCgSM1MSwrEB2TI9kxe5tIcrRgGO7tnezA3qRk2P/tZ6grS0rLnie
ZMNOf3mkCMxOkhcV8GtYOlz+ayrL9CHBcMgjn/DBUPABt600X+WCmLEcD1V2yfuA
8kRc3bWCr8OGjpnM5TcYGgm6BRVCIv00Xv5jxTOkWNIGMns1zWxf/84iGpftycBs
LvjXGzKbojEsBLiZ2WpoilIsBD7lLdhbcKCgBjRgJnG3in/7ZSUkIIkzStZTQLOV
8OuDaIVTBX2nQ8/ilPoSLYnj8LHMprUUnNpK35ppf77xqjcTDr3Z2NiUYFJmfQ9p
XL8ZDd2jPoZOQTmcUb4y3myh2thCgCHauNWL6BBdPr0k0Tpv+EwPjqqxzk/TSa1K
qikwkU+RCLNjFyD0lM6nLOm/gM9EW+8HJVnX37J4USmnKprF3h98Vgn0SG+kdp41
xHV/+ozACXzmJsPl54EMUbFiQql2eseLvvPI5pZXVpU55gBCXBijTm5EnPmXVNPE
Qmday8UCRS0x4pktKUnBjRTP8DqiAPU1b6gU8HNfMJuQapJuN85a7EYBeVaXXYb/
q/Iv13Zw8bPPDFadf2GJ8GKRg7ubvYvTTFP8ZvDRz8nZiqppE0IcwqZQUr6BhNUB
w/e2uAojYib97F9+BmRFVgVjXvRj7AU/kk1xUmL6d1GJzmkXH1GKPQzfK/kR5Vnj
+3szeXNZeHNZ3pOzIzkdJiOpxMofS3tAEqxaEV2Ba1t4fMuGxJ805ejb4hQjWDyP
JWOLXJfydrfcjpVsRnlqson4W/CcBdlYUJLMC2aQhnmHcYZZAvgOGnaVaYP86GR+
WtehgCOUSWwmry+O2fQB9jxHuOwcbhQlyIDyV24qfeo+e4sMBRTLWwJ7rgYyG8jq
ZvAKL3IpZA1o1NclOaggufSzBJKYerXN6t6doFvzTNeO65YJ9WDa3lJD8cC8DlYf
/Su3wewIrC6Qu9w8ODR2FPRfm7IP7Aiy+8RDvy+SOy94+pU/XwmLIKA5VrMvoGvT
HwtLk3wRzDRgRUM12x89q/nrHb0HXcEjoUdIT3SIMWm307uEO9utM3IPrpW3Mhs3
MZjHnj4K8brpIh780ehUN4DWqaFGqVJ1JgAA+FTnjPU+VPVkVHTny30/fhfts1y/
NHzSr/Azjfl0w/MSzckHAWysNAD3232sroxX5ucGEkHLhUd4UMN3lMuqZystEjyX
CPc3nCqfDwxfOXuc7XKUvn1h+28+kwgoVhLvYAn9wuhYZYU+oIHMv/0PDBxhs6rj
r5dT3/F3+lHUp1E9dOfpUveXkx5eB/RJ4tEnNHQtI2d2lvGEUUgHQBU29ym03QqW
9yyal3yrUKeQhOpGBGS6b2ThRC6iDi8VrPYmBQh5PLnR2IZd2DLYBS74/2pcW+OV
3DELNpCECQQvkCA0Uhi1wSjGvMiul2l/ABTEnWTPNWJFUUZO412QKVGgeVcmoQXC
1gViyTfwFaU2SZoIWwqJyKlPXJzHEXhsQbOJQdZowuH1pbUJI3/uMqoyyETuQZ9p
cPnJM163Yj/fgKmatx9mHzjnkeuMuXdUpykt4CFYSNLsWNrUX2/JIegvz/OhdgC9
3MNbfweueUmjY8E5yeBGEU+N0Ns0JCtvOt7QRHQqokNCSbTaoiJ4t+KA422E4loJ
j38KDROa5Ieblv9/PYDo24xi2CHBipkifFpIOPXptwWi2dcVpdOXUmtlCDqHj3QC
W+cU3CQvlo7mdozwDFboRRBaJC3H7CDRSf9Q0846y6FxiHPHb4jSjuZcoXEvCWUM
cEd09Uu6kGc0e9tBGOkUFGqLjozEgYLGjSaQkJaDqe95zN4wcuSc96bImT5M1myh
URGhVUNImYe00GMybiyHU38XW1Lleu3ID4O3ds58E4HhWqQxE0Ah47Q3OG5mmqCq
lwf4WFyP+cnJECv10ZIOMR5RWvDR/PQLp6QXWcVlQ21NJWCd2wY96Gr1Tbo8IG7Z
YLZMc04pvmETGQs/T0zRWZ3XYH0VAQYFYvz3YtmeQ6oZxgT8dZ1vcIYm0C6VeSaP
F6go7hQ4FxoG1LdtysvGQFJSsFID+4ToSkaPIg+eVq0ty5mOcaXMJNSAFsGxeRlY
whNM5WHXx14PANDmPa/AqsVnZTdvAoca40y699oNhaNtQC6vUbAxmK1AAxoKAWGr
6pRHV4KMgREYER4Hpei1d4gqyc04I52dHEeL1W1dYwm9TmQk7ppeIxz9gXxK9eSi
/5fAgXV1L2bnGVMcyIwcZkXKP6W3orjfyeO2t8fKN+7k+J7v5Kx0I1iHPkjq7vR8
WCbpVkhb3WX6aDCHeQipG/005ui2Sj5qd0VrAUy1jgYV+ECbJPQcIfJVKcYY2Hp0
iVavUb3PZk7ZkPN3R3bdl0b8VaAbv+Ub7JLjwAvxKUuKDEMf9JWbyVC3ssNa2Vlo
E9JQNQB1k/3tyLaoKEaF+E3PeIKDFyZn6qjG70IkghENpf7P9avrqUTe9g1+7WLY
N97kF1tqjU26naL5peHd0gbZNa7blPRDnlkF1UCbbnSZD+bFARAG9gVukmG6BOEz
X4wZXsNBGxLRAkUiVTORBc7jjwKI2AZg7QuW2rj8TYO87vL5lwB6K3R8CuNHkWyg
Y++jGzg+geYt2mYBH9CCQUpznf8MF3wlpLThAE7/FeCYjdhLFmbKVL3joeNIGjfG
KR4avdNEHaU0LWuwRIWPqsAOR4rSyxW1X4cioorHVERWX6xbPUkZRvTHTUdV86uA
Fi/w1fcgMOUAQ62yn4BHsKcBG5xCDNDFeNcuSqDqDdCrGZzM1OuTac2ztG7D9N9d
/Ez0Kyq4qZH6XQME/4egU0gaPYqNhAv88OfBwIrh8cPXR7Ne38lDloM7VSihtelh
ldvKR2x8qI3N5e5U3rIbh+ZKkmpsIVO/Lo6P3n4aB3aJCtOY6qYo+Zc48i9DhZ16
HttGGv3wTkTuuUghxuQfNa/yjlJm1fyBi8/bGYvYaH79/1iom/SIQ3H/GKfJAgx2
rUxeqgXZfBjAPS4K31tDvQtmiYH/ovt7H/HJNCdseAVd8H+BMpAjYyMnFpl9NzMA
SNYzT3rf/vy0ib9ekOo8XdaO1kLBZyscqPtexkvEesDpP/QzwrHpoDcOTKRjxznV
ra3qb3e/TSydYzrecmf5sPu32YpeLgJ3V6iEcL3f+LoaDMRAH1JT4WJktXaeVIdQ
Ql6g03xpT49PlPorj8+PCTs18bp5YML+/A0P0dxZaRvBqu6ILlK3+iiKtdTCBcWl
fbuYbpBZWoGGTQigTKx1pvP/0AqQxhwgW9oUwbZoD7C/ZniiJ+vltOxGvIAebN1o
e1sN5J6e4e+z0hW049YiJvdR+Q0RnLbbxo0B62SwE1TwxaGgkPHx3cqq+E3wls5J
4aXe44ZpUw02yIgWgB6f+A9bGx18zJnepBXgknUqzJ8QW6wMzK9lsRn8L3l1ZRW6
X7IWVCINj+mH+vOtNWegIK6jGpmvBJohzZ5Z0hOS5hpM4MY13SqFUYM9G0vB3KED
UkaUSMhuf5JGY9K/Nh59IdhZhFngbgWdIdEZP5BkcX4cIBcZ4KP5uELvV44zxwX/
Uh/g4f2hoRBo9pQEmMSIKX8n5ExrmYm20CLGXolaU8iVXrDTtBmUZILadkd14Qt/
U3HfgoGpNs/hQQkaMRF2jxT+4dnurrAqTuaHlLRQSA0rD1X8Cz9s582YH2iU3/HK
Yl7jQrvtOP6yOTEbqOKoB4l94CdEHfbsfaI63RAxJsybHIYp9f4Z+vl3KvcQL7zs
8GzXvsg2YS6bchg8eHeCP+dWW657zH3TgF2oy+Z6KZdgQfgDl1J6RsnW5VMMxCDn
/AGBAAI6FCJSAv3oDsKz+rSnnhe+dKwokwXkL1Mc/v1jc0DUQqW/htSNOwpTyjLF
URj5aQO1WsYbjehOR49Et5ng86Ha6mm8u/0rqum+ExS1EdtvMQFc1MaC68F6yzVV
Ye3MsIgRdVD87L0jAQW+fMKzZwbdQFnlIht6TlpdLLV/BP7kgWjkafayXyMFHAmt
Gq5jRdiPneiQTYNSqpBq9XTH/L750L9zu1H1Km+4QSyJXTegX391Lb0U4DW+rwY/
8Jki0H2nQW4oqrNsCn+PAKHR5U+xEk2tdqTkfTpArT0MMj+abybArfjCmZOn6ide
pDnNRXCuICZmszIEymQ4EknujxhvqPLGcFJaGTtz68+KqQ94hItH0TB0A9YVcveh
8zRJKlIOmbpnwmV3R6G5fcrtoYpYZSniodkDpSR9psHYuspfGh1BaQOP4WcujyjG
6OZeD3KpGFOOLmGrytAfGWXaFJg9DYYmKpbNKZDefYsKt7B/Rp6WEad2Rm7FCASe
gbMxhvzKdff8Qbtv2wvZ2kXeO+Es2Qn2bPA70y5rVAIVIWtqqnV3Kz1AxnoIDuUs
bvyciSD55wcKDUa52JshI1on2JHttjAYYkf0u42HP9TWPYNbZo3Iyd/i3L7qrzqi
RAMjLtfJOwCAghk9BI6N2qVyEV8ZTel9/3vqpfHNSmrnISsoM0ZoAEbKZmM4u2/j
/bNfRDm8NNKXpfNLQ6oBt1LkEr6QBr9qURVXGaSVVKTNNIsIaX3Jqhy7taDuMZRM
CDFhiVCyIyG6cfwhk7FPJuGTUBE+dmlqxdD/eya2Qyv7Bh4rhjo2yg9UBv/BYlWT
I4UjRMzcpH2kkMXykeUn2dtJqUM5DvLm9slTsM9bS62k1du80JZMIspj+vqr1W/X
NusPRCtwXUHo7Dh5x4W5w/ikLcLlzuA/ilUZObU8+Nz4610majz6zFssDKiv1neZ
bwIL3Scs3tInDX0cplPc5boUsxwf/reBqhcqcUr230n+tYfy0YETMnwvC4PAOj8j
oAfLwVkq8jvJTILorBDjQqHKJzSgDzWKSICf9QrEImlk91tQqmg9YnCgDLPVAD7w
j/yqVTYFmG10p9Xkja7YXltIISTRWri+NCAUNiwUh/M/7YFaSI2Q1tt1opXHPD18
vxTWk5q/KjllZ6whWonjnKaChOJQ5wa3984LTN+UBV5zLMgTfdavlAhX3y626/dD
AYquu5udExfZlN81q24+CyD6RoFmI2aaODzsGH8Qt2te0pcODkYBCeALj6cbWyuD
R+j5etp5CbFZU2mN2nr5NF0u2jjEGiXqsBO39Zf2xSK0Mq80aujytD4KvCDoudl/
YPQn4QwqlSkeAwiNn1i6q0jAWrQsXKyYJWU2PGq6UVD0VhnRYDLhl3rwueGyNl1g
CXr0HNzoh1QRB2w7LdJ27nG20C1H7Gwf+YRfpEbQiljM3DnyI+tbfwgLrc8/z2lQ
pNXnAOKKYRFw4JSOOWywk69SQMVJ5syXHZrK/HUQRvSbx8ONrny2kc3ucOvdBiSE
WrsbB+4wcFFgixn2u6TnAbftU0I/0O6s3/NYqS1gI81AuVsi7Omi0OgBjeYILkp8
1tkk5keAS6bp5l/yAkN+NrjX3TQUcxb5dGN390UZ19uRPVhb2gtkqIwD9MnMX2Dz
cXlEF6G+ALnpCIbasJeJxX0XUmTPAlCb+2dOmQIGKvMDnWagbhNeZscxFdvOCQIL
8S3LIHXbK3H8jCvijyMURz9DE//NY8ixxW9WfRY2B0g6exgcE1FEpf7girxRbGPC
VNYg01guUJUnHtnJF5Yrs28BnQ9CsgWNXvQPzQzgVlJqqyBzk3+yyBRhp7dpCjKC
RXkVVMQRMxnu+LoL+ZDVNtMjU36O9AN2WZTnMC6DgIlfWHxUEvVKU8JzoAOq6skP
uxQLF1+4F9gKma+SAQm7SaD3hUnmp2pLyjW99penig+cUhL2aJcMUMKRkWUu4bHh
HQFmB0rBO5FwLTaDk35XLgKoJMBPCm/z1CTn6i3wEPEiHunzwkUUZjZNX8oHKhlJ
itcBoj2QB7DZRXPz60VmiWAZICU7xbEfeqypmciJ+XZxmX0u8Wc8K8ZG+sGvpwUM
Vn3jU5QggDQkPFY97wGKKPw6zev8Lp2VckzIIXqBODvHB8QPZeOifDaryKukyT3H
w3t2fzk07yp87Wz/t5MAVgFmt97uR9fD15l8NX0tIg16u8x/hjeudvi2cHMDzl14
0FjvwytHPzf/6KyXKGP3S6T1oYhC6JbC+g1E8mDrpRSxy5nlLvGohvM21QDxhQbi
2CZ5f8O4h4pevEkSpgrLwyVvd7Hnpz8lem6EX1PIfZkfBZP4VMb74gjSgJMXn8HP
r/DvBrWZWBnxqW6O8e0025814vhN9YDzA9GQBEgMHLqAuUC8u0u9Nf84nfOU9oCr
1B26PgAyQmNHYGBm5XFGtg2usoUUjILQdU0TEvZofSf0EqwCK1HQKb9GkrvdY5AX
qP7qJ4xI8bXuKR5plGrgueYHK++LSvyPnK4KaxEhcnPUkg2r3uqnARnVHwijdgqI
u4pEQiRH3drqsjkqRvSbg9HfLbUCrd9z1d4s7MqHXrt3UUi5I6BwZAv7icTwQxcG
jWc3XiYFcfaud/xN7uyYiHa7qPMAGmRUJiIshdEJzVZkoUA9UklevcCZxL1Ln+f1
pnn7mspBcXVusPBf8rqfddkqeOldm2axLF0vBTQAKTQ5U59Bu1zjJkGnI/mZBs8a
UYHV/37xAmuffAon5p++lOs6LKfpnlhyyhWq671ke2j8YLa/UuONZQVfV6YW4/3R
njv2W6zlEOn4JMm3ghQNjQ1nFR/sLEe4HnRTb/o4qjLkdtOTFG6SQv/lRRY8hq6g
4EyHfqI56K3iMrDFiIw7J6YDevIjYCd0q2CEnVR4TMXDZwjEyXfIsIxEKCaE3hsn
NGwdTdlN96lxIw1BzZr8xC4vxOLVn/4QGyEs2vB5A6o9TWo89XBW2eqxAtxgWuSD
o1/mwCwVnulKCarL+XG/BDzyO4f1SBn3r6hsa0gttRj/s85XoFby886HaXo7NZvd
8KG7Nb/64uz6aMdY/kJyAYBhesAOk9DQASpCm99A0tqVu2rJjJVcb3g2OOktFIwe
WaefJ+KpH0WLeUY0LU+SwQ+1gR+iWSHhJN/UBjmz5/l52d2EIzdtYc+tFJip+m9M
ZtM/H3KcaAgz3aQdlXK/0Wlq0UUsp/OKoJp7Gk4WJ9JrN2V4HPPd5g/Cg6c/maaj
yGlT02B0USzy7c4EiOp3qXyLWMg+W3HwT2EzuA/VIMNqsRx10/z2gH6Ds82o/XHl
9RBn9rYL2bUfOrfuXd2vOKYY+hJk4zkYKegp/3d2p5U3b5nQa/wU99AHhNjIgidh
ia168m1gAkNcmBlYSPYJopo10RVkMpMGHNKLiScVHWygRmvrn+n1AGTLgLf7mbwu
4buIl9yeOUG4V3CdqBEDJNGhibohKjc3Z98j+MP32Waq4tmCPUYD26if+yzE109A
Cj4UPfQX7hocR+CbmvMtdA08qwgwp0BFpt1lEYyiDBRGtSYp9PKAhB5QuLASgQnq
TUKLPirPeCMgfqAouo7zO/aoJU5SQQLt48GKQCmiTW0SX41SVgIZVgi8DbKtjIrk
4Kr235M2Yd/0cs2+Hr6/3dX9u+MevcrEUXFFUBG2QOdeciFVaeYItGesJCVKJgS6
gz6I/oxGWq03yAyx3vfl1ASiGFX+urhQsMeauWviK0o4cwqhcfl3gtsLBfUECZKI
GPQ14tttYE9HvdoZV8qTwxnmb37jkJHE52C6+OCIEWQqmLUDmHAkavQx0ib2VIgw
nGN86s/HSyqPMkUP2MhiSLZMn0nj6lJqswI55gi5DNVpMaw3QlMqFQKPA95Z0aof
oDNG/9W3y8ZwwbuSv1iwFvCM1VxRx8tHt20D9xI8bDOcndn9qU+65VT7CK9Sb0Tu
bG5BQ3X1kQnYFj+XKvjvONPVhoiV6QkFg5oSebeMuqmpfSAkht3jFvijlw2FAJRw
+7VoEBg0fZabMQ/leecR1/+HSO/ORavos4AFxfhzJFwLPqqJ67s/eqXLyWnlw7/E
hiZWxgHiIfU1LOn6AcoEAnPcP2GbWUXwv6/lw72gBIIm7yu7gUsRKdX2qDK/75zd
8EGOTpVEp9fmllwaCJaR6AlAZOen47qxf93urVm0+Q12NK+r2d76EIv47MumElFn
1XdJ6dEmtVHVlh75tthfXMnHTDOnsn9yk8jQeLAiz+/wmlRnVAgkUm6jibDvUjVP
bVLHF8GH23FBFUHakeIegn9VbCSEZYpjp1ktWPbQtXyA3QTy8nS61TGpIJeBbx3X
a/BqbwPzvEq/pkAQDv6irKhOUMPRfhaoubf13d/eAwp7NXssDa1nT3ikhby+nrSk
c5a7D1TDwZEsljZwtru5Xe3lqJBkW5JrO5jsefPFdtImNtQq+OPLHCld7agKsnsT
YnqNOWDL/qt9/Yjfq5osSQXY/lXSQKMxS75h/BUzJdnexvTuqzOaNrAd6xhhrP4N
q2jnWcHBTKb8nFxPIH9vMNEgmuWLsHcws2w3weGTn+vA90MGnsCQ7LHi3xch+1rj
VziNciXI2cT4ITc3f3Wu5sDWflzgsX7q9CRW75IxyT+1PMSU/8wuIe4M6s3+4Fvg
KM5AL0xGWGjkLWOo+L20YesgK9KP7AWGPTYlGLcST7nUvgxKPyP/rDLXt4+X68gh
kBgokhkbi3tvXvNvcrlD5nQekv/dnor4iJVF5S1WgOPAuGiigyiU1XOuv623HU6P
Z2oALHmWZa09vU6oze53iyOcBkakqRSXcgGcbvETjqwPGNikgkiTtYWu3xNsXwR1
NjqXXbWeugG9DF4sLA9Y3OoP5WLhIBvGR/sicOvPNGEbx5MUoliR8T8d4HPHEhcf
k82VwSiAD8uW+mnzTXy+CqcxpAtxbI4RVHQvIJv1iDZrDyfMyWU4ySBzX4RDOQyt
Rjord9fYjgy7PdNqikgwuITFlI46zi32V9Hl9rOL89cfiEMNf//ELqPntsgU726p
Z3zblqob40vJEyV0dSfg4XiP59DmYAC6limZtOw61lOf9GkPHyr6y350EKsWCM+t
r9a0Dn6m7RZwqP588Odswq1i5Tr/oFR9KXvfbpCx5w0APr1CWo18c1MsqYI5s05M
TZmb+8BsAy3lnnnh72u5PEcCD+Mq2O3hr3prBdBKrFlAn+z86QGWlcr3SaGDy6zw
Rqx7lhT4kt1s4hEOfH9SAUWQvkQSY0H8zLfRk8uQmjuMh+UIwY5UmRDte+Q2wrPe
Zgn5B98KWRWZ05jfnGt5AQwBBlWsn9cRS+4HPM7N7eEvYqo1p38LXQthYeRXZnxi
tfxqisa+h1k0K6S6nzTbOz5fbw1D3N5DTzgCOSUIrE+bXf8V8D3R86pWkqMmYpoH
sn/bgzfwQs0dqS5+rXgAGlU0rG224oNLoj67ATiR+UnjZyajz3c8LbtT35e5PDcb
Iw0fLimy8y+u3tEnpr86kzZmv1i4LsliaaJy8skXPnA3rZ7F9sk9ku0hNqNYtABb
7WZCY8NrWiXvlfZAZIHxk3Nky28VcANwUy4/dMz+cbGf0qxXUP9/l5yGaCBIbCQx
v08NvcQuw+/vN3atUT5GnCkuJD6k30W2wKlWOE7TgKck2Op3RQENsF4zoyB7e2TD
WfndD5e+bv/zibuyunMbYTLY+NGhqUKvwrQS4PcQua3GeDsMq7p4I3rY8ISX1S34
/Jl0idjXcLeoLZn8OXzPble3sCo6HHHapIe0x1pcO6oakLC3jfhuMcWFhpe0dHrv
KYV8iJ0osF2ekwqnH2n5/IWD/JhwXmq5VN1qk821p6/E5BtBLInbvKKK1XRzTgg5
XLrjKhG/9vLOj0bzRHRxNEulmvLvIhPAeKPtsmd7Y5sY4oSfQvgmZxO8Rmn4TrPQ
Cc2jjTaVj09hr3V9NZVEaoFuS/ckYNy8Lf5fuenlotfFsBioixmUujcNv4M/zUao
0FOzmE8PmgYNMi3lWY29YMiNu+0eLFnfOzNzdJ0nRx/F8D//F+GpaGCFG4sq3NBj
WeCpa0SimNKAbVq1IZfhu36AvbYyrRdA3SmL+v0n56Fr+jS3gH/wn6rJkvErJSI6
9llcdKCYSFQMsa3ePTKdqWQEG/HOyLNPZSi+hljC9bIJS6TpATcIxspofVDvP6Gc
tyrgIuHyWLypRaRtaMZueAJb+t7Q8x/nsMVGGsWDsXnBigkMvcw9FA+OKGEj1hjJ
/jtcDNR4pl+ZxWKXIIHMkdiXCVJuxsspGNXpScYizgUDC5CUxvsOTiyW+G/0RYZb
bhsz24bnh+WOhpTLcZ4lNJj58LkNVK+P/zQ/uhRWh4RuOS1SZB7y9YleYMyMRbS0
Ffa+oe3+PJaiwg3flj4wtcknP9ZWqOFth0+aJR5Op8oDJnx3DrTh8NM27UfueMER
6jIfaF47zV7oge6wmptFd75FZzQAYlkp5I1uXTHg+aCR329bnMJV89CBorRVmqFN
g3I/BXDLV9E0gpMzaLUY52+TjDiTb2NM3SMgfT9K2aSmWxcYOJd1IE79RMAiBTTx
93nDnrSYAQZT84iM+laPsdxvQaITpxBHNw9oGeF8ThxUHVGdvdE8rJ+KE7lPUrkV
a/2ACiTS/KkHaaFAMB13lNcxyP9g4aR7roI44qZquqUXltf+RvFjZPfSNDO85pc+
0xAzuLGUsLEz+txxZg+4cuFWDrceiCaQGrNbD+B8TYjGAuFCX8KI06LOlom9mRd3
1pHYnpcPwfKcoDC8ryatztSxDtnZUCv87pc9SUpaJGCrnLs5AoY/+g0mLXi51HYw
MFiL+O3cjUyQRmACbsbVd6l/lNQOpQfWwNRCZ+veSnCymitSZO7y65tskGNiCZqa
gGtlyrm+pl/9peGZ06p5ltXVeTAJiIU/Y9GnIWv/qCvii/0FlpaRbTOWf63Feeof
GzDjSs2Smw23zoNXQXjY2P/es0pSo9MbjSQK95Ox/CdPd6vvezwL4sT6tRP54uDJ
YSuOUVm9bgJcwtMA18sDyYgZxzggVrzw93zbZEySjV7oog/uZTc3SufKvdXK+ZZb
YyzDbYF+yb6vJot36GI45BGS9Qu98d3tK+wDo4cGMpubK4SrgdLoz1gqb7XBtbFP
BzJhEECm/j+hgm+bsraI3pHardOMTxJYRhlYxoP3IHsEQ6a4xk3Wp6v3opz6ySYh
VqNIzzkGDkY0CULwtzqmY+ajOBzESB8l0r3daXCtx2NESvWBXE9SgAX8ZGnGnPB+
wWgY45F5waxoIe6/9LHSmHHMrHNFHmap7UWvFkM9lnp8FNBqVdZUSQc68UFmQaCa
htDzFZ6MXyEv9/+KJe3McBKOfbVCTCarr8lMAyrtS+c5w6uVTb8x667QVaXybIki
fZXJ04DeZ5Hba7FRIJGUN+ffA18Qehemracy11zOOJV6ij8uS5NDZdY/d3EXOJP3
0E8kTYXC2s4asHwGx5vo+pqoYhrHfsvfvIYOabUSzOk12ZvH/uZZt4LTC+M7Y9Hd
2QY8K5pBlZdJI7NtB/69nfjpw1mod4aYqDaJf+CxSCrRoGlM705RTu+kcJjmUNlX
ls35RbbQCU/6Fa4bOM6sDh5yBT50Y0IjvuUuLbKOAb35i71VB1biAzyCAkg7nAli
SIz7fpzNcIDI3AW4uYpaIj46IO1EY4SPHoJrqxRtGvla3nQUB+wcnDetJFN68+a5
2BzSMMOGHNBEcIA6XHuUinAoSvnx11p1mfTTsvL/xLoNU6TBG3MvLQ6B1XgHYX+g
wVytC+XapahU3fXHl7XpBB0YVzMIjnHzz/W3/vYFR1VH42fvjOHfLbx8yNRoDPn7
F0xv2qWI3s2R3i2UCTrAEmAnuFX62yLyv6zcXckWwezPqVB2Ufv1w/jr0+NDgwHv
iIXQqXGv3nWD/tShU6aN8ZD2DjNwptyZsRa74l1D53s4/zvEHoslFTsfl3urfmJT
a5GXKLDMGPWIgtQoOqYq4ikLK9186NfUYNkeekBbfEyTLup+PZNIXRIzWi7p3rsY
SuwCj+mOl31IHaZyjLk81w+v+nrTKPbrRwmeBqq0J5pvUVOVPwClU4W6PklMgqQK
JVW/mmjJuxNupj/Ki2LVDT8OwwFeLOzrBLpiUgjU5N/L2QreKgl4Nttkx2hG5F7W
9cu9NBXMJjNc3TWTDMzd05gvCQgLJjXdVcNh4firqI6ftN04gE4+WoC1CXF6tk6b
yu1WKMeuYnammKWoJ2k0LfX9zDR3KB//5iKpRoXr4SeIc7fUYg/8uIL8jdHWwKDG
Glc+YM/xtlEYSyC2XFcoP/tJVBnGj6dX/byfT+HClymZwpglSiFH4FGlkHLZguUJ
6OZYILZFJqWrdhX7GfMb7SYchKV8d0wMoX5bsYvMFSeUOdVs0foM5qLXkZT08I8w
xm9cCjREpzwem2s34l5YMTYopllJlByx2vyZnWs6jXYqN2am6ejZpjjPHBEo/Zca
5wFAFCNpL7GMR9itSkzfrGvnC/PU+xHeZmcMMXJ5LgbIRKi+upcM/KGciJHL+6z7
BKoqnx0k34uwaBL5Zjj2oDjXROTpdHthhcbbrwVHOHYdl5K5tMpUpzUidSTxhvlO
Vm8Z/2VdgwcNHa0mzWE7lupTm76I6l7vER+WtKN9PBi8IBO9fjm7edMEsysNKxua
MRwN1sjz7dQlKuX+oH+l5D42X+FJvXOZu7MoKmy3yWdqqlXtU99LlXUdKBYCfYPG
EZkDI49WNWDycV0FdkTgf+VC2ZqwegaVl2Z03uLrwQiKR9D6Z96itwKYvzHJkcyC
mIfZ5BGsNzH0h/sKPXe/aaQdWoFFnHGgsbf6ye9XD9uYTwP+wqggotvafQ+iclyF
3nwwgtfB4NqVX0sz1JZvEDEPmvu1GdJ/yNTS+PaFbvq9dv+qvITfRDEuF8qTNtlE
BW0+2Y7Yknt8MxIbLbLzKuIN1E7vSQNejNCxJo/Fx3B/H2yUezTv8ZInLSlFAXOZ
1UtwQYeXle1JSIJTylXL7COQrnfQazduSbyQAIW2BbFzMecIa8vkpYi8eVY9oXUg
ANQ8ZGKcr0UWiXW+QPdEQJjtPYWLOirS9sRvhyNtRrAu17l10SGqfd4Futp0KEiH
Hz+F77Jbp5Z8G786Pfb3yeQ6gWMdFpcFCQGMQVhFzikuFLQW7MiLx9H6IPhdcaPb
T2UlhU8JfEc6fagVobEr0+hca/pVHgcSMplLSjcH/vadFK89CWVBk+v15XUV2VBC
W02K4/IqiwGpqz+iH3gmZNon5ZJPJyx/8+yhvNK/n5+BK6irBwAsoPVQAbgdDU9C
e8WRDAW8hjWODybk4DIRJ7vl2sZ3+ZKBRVzqea7QtfwxCL6W/WBEwlho4yxOs45/
rV75nmmQQvnDL0U4VqWpHWTw2rS9iwWilik/M3nKY9bpod/GxEDzP13+Po2X09vR
4zypFUN0kasmxHDbwMVgvOTPXInSiZY7a7WZ1qNaxawN80Lh7EHgcvX66wVmZTuf
gV3l7IoZm1/+V/qic3SEsBdU0nBDNrRccqW93c1jFnLvI+/my7pbWjJCH0o+HzJd
6xL1HI+bMATtmoDEj5ZOgTshbAqgKjYk1IUpMqHR4lBny1t7JZhCL8BBj8Qxr5BO
F+P/Rz56+6SzyYzcML90Isb0nlktbywk3TXemfa0tQL+jCGEIrNav1JhbYIcIrr6
Lcxa7cN3rCxtkwrNpOXs+u9lT/qGDR6OKIf/77xk4g+L5WFJSe8wIBkngxc9hGjG
Cw7GJIHPOQsaymEHtAoliuYrDgpU10xb4OrLhfRUKGUZcyBD6q1nJN/QD5lRnTXB
RqyCqr+DE+Gp2ICS5STJzgqJPH/J3/1FL46B99jH86vaD74xrp3hebNWWOakGUnZ
IWy8tUUHlg02l+fZJg1LPEJWqWU/q97ZM9nT/sxmuMfInq6eb7+OQKbzxLvY+G8B
nD4OmfC6GhihcydJSI282MCb8P8mofdO1eGIrtIsdMTsv4hpviLMW8sXBrr7Byau
LjZJhCgcj6/e0cTdz4AVQeB7HP6+TivZjyqB3UaFuZuXDjx97e7Y1kFd6Ga7KuDq
nYbPwAjkwZdhB039XZjlWAuG1beJmMpV6OyrY+oeYtNKXZYwxrA5fQZD5nNtEMb7
P+OLMNvydQSzAfLOfWGdrNT3wqLTtOfwL4y7iwj0g2RRqaSgpf5Gg6FCUeHbv3hW
qFXADLPLpSlhUfhuEZv9wcthjLZ6uuN8nIvUVqC8zw8s4I19hLpZpUoddixLVLBy
yWKyJLCY1mGsklXBk47A1gDzcAZZQkM6f0Rwsc9NnjEMX5wfzaanyJlZz6pVHd3x
+oBS7YWaePttwX9wlSI+pJWd0feHRkiKhStjSoY8trAGplmH6/wlaocOG3ha2jT6
25qMXgqfl+MxnuWyH28pYrECvvN74jPIyQMAzoPd1TcnFIXo/Lro5g4aMMXjYKKw
jGzGTX73rW/362x5O/haoavAbsrXZBWcg18HkORDITGLY4iX7jkXkHI6Wtg07PpP
VIzRflFI0c5xNoxYBA9fstjqGSLTS+jkjQRdlv6qpAPh4HxrawXZPPD1t8eaDFMA
F4C6bugTIIEDHGjS1SRNiXk1GlIruOqMNjVAYU5imtzIoZ3ZUYOkXwERV+dZbbWf
ZM2rg/EckwFUWRutW301OaONpRCRUduGWTdxjMjI/l5IaiUp6uIbzxPgjXTAQuOC
orBq9KYdxzT0Z3SkWz09F1dHsiQAF4HBTfMFnHyVhEn2ZiLxzoabRrbrdqfyJUFw
IvSOnE6XqFZ/PwfOQp0MIF5zW3FVwVi55EA3ky+v4bKObi7MTesIqQMqEOnu3O5X
IG2yDXv33Ez1McyBjinO3SpRS45+sVn46jNVrbHSQqiAm3iRackKj9JCTwRGm1HB
efQqsLCefQYPUh1FxmQd3OQvO5VUhR4YrsFxgxBbwO3e/a1I6mVVVeS6Y0el0JfT
czm+T3CiCRxvowIxs8zxK/MsmxacbKlLj65KOvta1sbgOexJQo8j+JXxkIRTkVuY
lG1eJPZMSStynpwtV8MpJKBvGEIw4SIbIulj5y9IDpMkSsH1IFrlSqpQJ0BLqGBm
neame13zCsYjcfOXEYcvWnFXc209G4iXObGyhlTsqB31DZvOWMSgVAZDzbHUeJwu
SakmCsf6DJkOewTPuHotl635BZhc168rhaBDcq8b2boNu3SukfknC7Qv2wwWvm85
Os23w+g8esjDVAjPOQ1OxQozcl8Omqno1zAfKFeXZMP8l/6/v9cImz4NpRURnjPI
Wirzvc6XCM9jn5RzctZ8Y5XiAF9RuewaGDwOYIpGraBidPd1jpGTXJfSIGfd/RMZ
GDJB2p/sAHwsj+oWwosLatY+01VXhxjnldQda7h/BEL/5MdCZE8uYnvinPVKV9Dd
lsdeJ04mFM8TzPFfRisWWJnVcZE7in4BLGYh7M09WvpgSgJrYBSKL4eFN+oppNfs
cjUjJUA1I7Kfwf/TFsHFi/k9e4f8eCyx6GxgzF40E8X3lfebZuM5YMLBQwOwwO78
8Tkp1Dw0awe4SgDMt3GZn4BsvM9+gXOPfuIuU7dNjPZwh5LL6bS6hN9tzbg2W+hR
bUNhyv7H6maRwniQa319ILHHH3UyEuADAFbsRsnwhdcf5z0DxyFkNQEkQRW36q/J
8bMWbCxpClWZAdz2hUvX2+U+kb1FcsTfjMtln5xksoCocc5tLoA3k+X6W/FdfjW1
7TaWaDRhlPBXuFPWOWobFBxUweLCqI7nwnsmnUtcu36Uk8WqU8FifUQYXyIJNbih
2NcqcEVjXgpBuLNWosRLi5CjNlEseld3NwRPsJ+cAGIsAXBZGXEkjc0Twukm5CMt
6fRCEMQA+k/hquMKrwZ1ltA+7pPvRqpYtii7U3BK2nxIDZ4HJn1TMUS19ViQhkjW
s4AU5MufaVpmYydImtC4RMTJobu/vDyI46V9UcBic/g9X6aAQZkpUuoGTJvcXrx9
86anCYnQdkQU6d+3sSfd2qQY3Qlx9MPeaM5vb3AbkBZWDkbgk7EuGNnUAjq1LIVh
1u5GuUGuPZHdI9a7heU17WFFEcyNsaVwv5Qv/9LJJcaL+MkK4HitY6d0QnoOluIc
AOCISwXfpcTu/TmsNNOkQL9iiRMIbvI2a9SWNY0zrgHWxkOkv07GjrNTG5BwTwYz
3KZlUcmTbs7mTVGSuyJbYLsNqWZ74/s824TPyxREWbt0bv3Vo11/KgFq5MoeJkdO
q/TldMP+RtJcEVceFBm7jGhwW8vsdG0CjwPurGTTf4qFoeLYoyKX7aEHNTxsYX5O
kBRLOffnnLVB+r8wuNIUtyxtH5nIo5aHTtBfIfV4e6tACIUJEI1Aw7NrJd9AV8m7
yFf50/eBdzXh0jtIqd/fraleV5uVuoz88FweZXehgpa35Wie/Vq/gsW1Brwt1fNg
iIMZLzexHytof59pyHbga4jDHFRzu4vIvlK4nSkBDc8dH5MAGRJHFAlz8gsh4KJ8
57egHGC65EiZEJCaPCOufawzxypXPN5KGeKb9iZxYfWVe0CfDRFyMU9mmdvOXX8t
Uz0scyu+u0oOsm6jFdShtD4Yxp6wTe6m+eZeOiq26PaDA50QGcrIiG4+FTo21+3b
fHJUO7wvt8pIWd1Pyzeori1xSEXpySJsdnjjqvBxVrMuc8LzARDRckXkBqkfNGbx
s2yeAu/A++mwgtrU8cn/YX4VuIMFKuBY3CZtO+0wqvgqeYQcsgO42rKh5bOqqEUF
HR4GhihRDbcgHcm9jmBhdIFZ/yRnqbOrGHu5fhGcznXuMAGk29jvgY8raMmTAWnn
IYwUfOaews4u99hXm9ILgKiMRMzLJ4/7dbVW2X54V0SVw6pwzCyZs+euF3VCRTqA
0DAvw29TZoTTjtfR9MUezblABBqV93ZLOZ7apHbqVLJG3j5RTxhgZ5ZtJNgubNaQ
TDXWfQfKiV3CcZyro3uSkO0g+PxxFz3t4K0yjgP7QhJLzy8igMdW8j3e1mxQF8UE
dXcCnqRtlHbsqMCgO1EoOIpEGVvYv8g84KKiftl6sfJFItaM/aN7DKh9+PPJp1ro
8sPC2TWmWLHla4IN1D4EIc/hicyjhVVWJ6fzQrTcB7RP6uwxEVJHxkP3t8zV0e/m
Vu4wyM03exifcQIMyLWH0Im14ZHJKU7jmTiu7EHWKm2AVCHOg6yE7VhJAMTeJoFl
ABzuHDSnqMaqqarbI5yMOCS0FSIkC+PUsfSrf85Nc6o1JzdNshxZtguW/skuF+5s
/2AWdBnGdUXwWo6lZZKejAhpLkOOBvCItpoX5XdgSA6H+FzVa/XU2T88p4ZIt2l3
4A8bCD70BSfUNATIn//Ro2QLKCc8ASjxrGuVKoahXP1WUPq5vrnvlffeiZeKw0lP
BJL9cnA02G7bvv0NKbQW1hw3PxYueh2LuVxeo18V/MCIgQRCZbcrJ3qGchFJmh4G
tDkVzZAPSjRXPqHcKG+/HKcMePxvJAaiBUcZ15UVLrErwDbizCbe7ObwtUmjXCTG
5mZRi9i0asT/7h1jP/xOrC0L38Rm7BFsA4H1NVRPrqhdT7OGzh1lsxihZbAR8Vfe
gvgsD2FAeDjrmyTN3fkkOBhei5EHDy1vYJIC2sVlPn05uZ+oJNACrLA50+Yo1myk
AZmFdMOUbkije36w5utnsAxMefMT28bVpbqasPbp5Eb14pqgAPk065afc2OZubWo
OVoo9T0i5cbRV+zg7ydMBmlhOTI4C7HElkqnJqJXOvUhklvBJF7OnF/z1PIqR3KZ
WG0e8WGPkyNcgogRArOG5V299vBBfdrK+qvzrYMcOJIzebDX2nh5pURBwCqJIcB+
7QTihMIvRDUm58W5fX7sI122GKTXKRFOrRyJmUrqA8LA+4N6GiZZh6J9nIQsDo5T
A1Hsbl2VS6UqASSaqLitSrWEm12DR55GIDA6kdwB9iuamPqXuotRgA9ghPyNAqMq
DQIl4CTgZUWj27tQnQfWf69c5enJW9yhYlFp/LHVMWAkYdlIt9bTf0sVpwZUm/cY
03Ar0CijLFoP5YfmFFPJo+6shqOfbIBR8jkcOI+P5UQ44wCujmQMNo5BNpNh7O/M
OQZ6pTDEq7j0w47fSBKaRXu0nmr1ingiZzfnhChRUKh9Ikl9y8FH/ZeCgyL82n+d
8rdypOKld5zBqfa8yIxOMdsI2AQajKBcFBLV0f9LMJMHGsJMlIp8JOkr82nDJAjO
6spvI18VD4Muckc3za8dD6enayK+fKu+TZOoeR954NmRMHd+RwX2aEbbdoLqgoaY
7Fa0vuEKJXV+FmfWYUmRmEpa4ZJ463hu3mjtsyO0dmjVT7k3Jt1FQYKLnvEiXdDV
0JhSUmRaYLZI+PVsX9oHMYWOz+lU91zhMFN+vcwoy9SKfG4pv8R9gBc4qhn4COla
twtPFIG4yaisiSwg0sdCVPQ3mWThaoq4gSIwqoa6iPntiZkERCQWpAZ9YGIxeHiJ
r//AnXqjyDnxZLRCHQzuBV8HJplMXQgm2WtgJUd3UTXZZ50pv4/inJNHdqNCCNCj
vpqhCV1CNPKTf0rZxQkOT6teZu2kynZT5qt4HsnJEDwokIi7mlOgqstY3VXA5zSG
RkgkBcnSnnRSf91bHNzxdqk8WVUa21ujFEY6VWkfv/rnjLRox5vjLcXf3LlpyHc6
ofzn2BmJMm4FzYt1EqiJUS8qGRoGAwkoWZoMGNZjArM0SIcDNxUqBai5lw0qp+tf
6FfSPUwubM7pB7rvwHh0Wgl5RpfrkRWByCzlJA8JcI+aELova4Ek1JaGh8QDMuMR
ZoVazrrYY7gsc/0a+yHoGSDEmLvBsOvxUb5430s43kjTwqwzhmrRLe0tcxjDCEJv
iZ06Er6C5adZMEqxKjfznDuvVqMjAFkUWy+MMb5Zpor2LO3IzCjNhocIHeOkiR95
gqT5zegp/ko/BIEVd3aG6+5zKldwxrSLB8I/kfEL0lIWEwIw5P3AyMLfzHdWEXDY
rGuC3VkKvI7Wj/Ns/ZYxeU8e20vtYQvEBtHNSrX8cUg0xQ1C2HYPS48Ig1T+dyOg
YfonlXCQevhEKUe/G/1mnYlyaGKFqYTIz2iOdw2UpIdJHmw56DibqF2YjB8W9bBC
FaoJnK/m8n70969A1DOnrdJgqLlzz/7Ox3mgBzBwaHELylD+dQVNvIJxJ3D0P+P2
e1iTC7kuaUhnM+GxWqJd/jyGVT7wKFHCRCMBc33n/nqVCCCRjkiLfOiURlh6OGaY
KIxnoVQo3zcfqUQ2Tyw1aMw2fKgMvEEvZiqdxpnhSyZe33/gPf8DJH/i8xlDd++O
1yCU+Xs3YEsLzX2+TeIWGOYyd2tmmAX2DhuxJ8jonubjP+9Z28LL2rMXC6wgGi1z
jFhw9LWhtL/M8gqXz/lxRxvyPj7Ih1onTFiCCl/UPeo6RKCceUO7LDPwXEPUjird
G+kHSK7/KgwRumsX1U10uoCC2/xf/qPgVsR6eL/HK+2Ee084e6ZUqGcd1zO6ZjN1
Mjzw2uCI1VfuPoiAvxtaFY/mh8tAvhklmnp+LCzRUYnFf2O/2ipc0o1NkseJLFBj
xdSasaKkcDvAZMFy+pTbSu36iISVWAh6V0ULDb1ZAAaag7zOS5J7rE9QKlfEr30L
5x4SMLn9HcD51xpQ/MTmnbZD5ZpcWwFY1UpgHnon4lZPNCSTAblft1Sus0UNUC3Z
ErU3Ioh/flMaYK9zH0X3LrUDnqpqqPC8P/1BPHjNYzzVlXZvrsa3kalbRJzocLiC
YvwdO21GnOt9xHlqngFjovqLQ2D8pN9Nhu0x+WMpiBfuemjVxh7OM9dAABySrYTD
xqC/ctktOT756SZ0sf+iBnu+lRacqdmB11OakgWnlHR+3vgKhQrngsxvdagDEhwu
8xdYztTfEjJ48L7C4Khj/R3qfPno+gd6+CnCkrIN1oPh9TAmuclK0Oy4hdALFd5j
TkaJD3s0y5M1smaPpAP9EOPHCjahvkD4Ch5BB/dnvDfNHjU55kCKT7hvVtFbAJ7l
fxrQG5SL1GlJUZRmCrkz/el+2fKjOtC7eJU0cTVcgZt4+LhlHdre5r0MT47XjUhe
uDqOpGU4lbTSJlE3yPgkU8PP+p6vnRW3oGiF6pOTQzyq4/MBr9clF/6xvpet00tW
TWaaMBaR8KUvxdSQO5r6Bn7wZT+wMFLyBmJKvTzwnPdhUY+O57ftqHhwMVe6Vfri
lqT9ME10AoAjvyb56HXomx/LYagskP0acGAL8mqez4wYQ0L3Dnc296WtajqYDPGk
ethuUSmnQAhyQv+E3LRzzEZ0IyiYMZHTn8GYRiW4gvBMGoVII5HszMkYJO90NOZI
lXtt0FukeUXAChuWZjsAw/GQpCNvejOtu+UmEqfnEyngQLGY9vs7X7vSBxPU17ic
6sXhgqnCjER9m3gDHEKINdVRWHtk2mdVoSDZ+o5hkAsFbQqU45REPDyIGAIvfBxI
aYbUC7c8xBXxFTCd44ioBgTB3/+uOZQcaiYHPO91mBW9efokNksg2xAJo/RPv41f
CejCnMVz4YdA/WV/AEuXP0OgJxW8CjlgZFDRYpTwd9GMNHHRVXt90pM9vsho+8sk
zbCidWDLZQz6YtM4ERDvHW35iRpjo1HbvUORawYAc5ow0k1KyH/veyaJR4ZPeWhj
uYmJ8pBgmFDNK1Ch+/ikb+MWDwPxDepmIY1h2qZixEKZHOveruTZkKPyVCQnmxD/
jpa5hUv8tscgPWZ27bh+h9zuimN6Kr4/AK92JkRD1oVOZj9vbPru1ErX0616AyXe
ZX+qtcaozDvsGgI8mbix7W60YUW4M2ZyNQkcctv7gyiv5W/x9Ge+y8GI40zICw+M
hByO30M4qRNEyqPQoHgCPtMLapbJsq+7bOimXe/JV0pVC9iKZIcjlbF2Ejtub/Ys
5b5PX5JZLJb6Of5DQtVxEo4TC61uwcgef22e/f4sn9MPSu8uMBr/9JAa46oSjkC2
Yd7Ni3OrDCrJQOLQPZjFTz/eRn80pI/gKWu+p/et1SMPUqP23wYMPFlKb9o7if4U
zAkO7rBrkWVRFnauPzOI8MtUkOezVvZAJFNP+yI/MoSeW8oSEVgcWuIhT6KeufqH
Mmqk7WvWZ0Rcj9bwsjoguzZ7mSoyDRbuDGhMWegmSTafm/fYwdQf/arFk4CkZEYL
bXs4f3oLXOTWgrHWTHIkUeYjVTKHqoR9UAe/ZfJJOZwUW4+YhFwwO4biDCqphgBw
VsrZ3OjNOmMiSDiOopBPRtx+FMBtNNqeBEVrOuKIH34IMtQc3VLnDXlOBT3NAuMB
YsYINvCZ8OYxZY9K6CAugChcJ3hwvTFzgkJ1EQ7oMOCNlqnaqwZ42OK5Ihzx3jUR
uxcrS1ZYbLHKdm9kQmmtE6I8VbO0jmcl8PAoH9sYcmNM+RAsd+BXdZPUOjYIpoIk
wwb2z8h49QuR8l0dClxZprhx5v5NzYB1NpOBL8AOIAC3qk28VSjiOsZe9xxfxme5
3frY8Q3UbhFosRC+ndXu9/qZSV3QuFASCj7HMeKZtfQgB1NAh+iIE45zSD+Shy8K
K8CvDwEEYQCjeP1VN/k03QtPIhDiugPNYITv4CZoCRJuhgi5mxQCf5ZMHsBKPdQ2
wPK+s9CWWUZWUvVG+DQ9n+mOKOkag0pYSLAXTXED/lt9eQ6q4uY6Rg19sIUpX7s+
WmV25zpFv4e4Q0fJxyxaWpHfPPmhFQp9FS0Ab2X+IlFBBSBOmzrByqDlfhM46vq7
AEQbj9HM6tJaDo/TKx9dBoPpDJ1hlbkiZVieTSRor/3RQ4tn8j4FBw7xk6Ru2g3p
kG6h0nOAWofmRy9qB0Sc+Xax16W/Fw1y7qE1ezA3xe5ixHin5qCnif1UegapFhPp
8UELxj82kFRpqJchFeQ0q36eIJeum3pQAlfnOfmiI1Hr7TI+6gMjyjQ/Bro0LUR1
FzTeyGdpEIX//UG9qqjpssfL6a5GluTxvxHDtWsJO21wjZHZY71HiMchZKWFBSfh
w6g7dFjVvuvLP8Jg0UGEIKZiJBmKqXJssvX9CWyfn1uadpVcpKDcHzF8lzyfIX22
fUflcGNovvQUI5ND2L0E2V3lLM30EeGw8O726WE7BYHrP9ZJmL+dti8EpGM3lrQ8
/veJL2uAXcxKhrWTSb78zh//sR+PB61fcTr34BKcTHZ5Zk2u2ecLdBVVY8xlarab
McTwLsMmEJtSnAvGcMhiMn3b/CR5dZgTrRRRIUmy0bkzDesDzE0DquARcMBPpQXE
DB3O1tmY5lsJ2Z4fnb2ykcixT4K2Pm4vkhDCeMcLeBreAX9erbhZOUqSPWD11slf
oKdeSrCjAt4uirPEbWHeHhXNpUDLmi/lV9glgbe79FRQSD6+1z45DJufBOf8b/jV
AqvBp7HUxPbP4vMMSbM6GSdfdhSnsk/TcL1YHqBL1DeUsaCnnXwfJC1NF+4ucQrw
yR+EIP98Vvhnmi0H1Z1YKPhMrhvuUE7r5U4zNUN4OTwjGbr92cU29kOGiATzX890
B9gaXYRYb8qEtPoLh39t0gzbr7Ng3XAKC86nOOYA/3xfDD93QH8GgX96qEBF7yk9
4VlC3VkZiA6mQLpTSfzC7580WoXev5rBxnDeCzygHl7SvmPv/5NARjcV6XaRDvUJ
+GWdLbctQj621KP14gxbofFMNN83Xq8TQdtAdxEOBLgqrpXRagsO41x5XTS830is
BEQAbps8AZZomJR3hTBErb+DtF7HwsvaCFUd/VhOlNHNz2bcBYORQNquNsVfYKzH
rjO8hLnGTuyWC7y8SOYln0rPtiLUZK0JnIUWBs4bduuLTQwjkkRHgBdR7VIrS1tL
i2UlrU6Jf4sjlNh+StN+cVAbNUFHgAMhnXujc7phx0weXFzV5CXDzWRk04AmNcW4
gJDcocRgJcLIslN4+VeJEreWMgXn65iMm3RgL2tSQOxslOBxG77+xviQRgiBrtUy
1uj3R/tn67mMwze6ZDQE8d82Q8q/6M2FcK//+2P9PDN0vOpK2yWq570StzZfIdka
5xVVpilJSSTVDmrFUpfQ1vOQJloW2Xlf4F+U5Z3ppOsRno/mY/hH2yR+xQFejHzc
+sTZq1qq8i8bZq7dTcUAmuoADXcw8/3mC3/6h4MUX7gtzaoOMdw56rk8sfuNLjAt
INdFRTPbwlB5ifSJ4PJLl4Mr8ZoGx3YK8d779KnBkBPYJovLurE0Y3tgt6Y9w7mM
es+MHDnHH2AuXwCvUDxBCXnV7W2diuwvCI4wHIMlPkST4ApJajdhQhJVAA4MmjyY
7xXm3/CLDNoM/9m1/3BaXyF4mHR+xbBnlutYDyYI4VAHwAawf3bw9heIq/o9/+wQ
HBTOF/2diTGPmrGImqkgPjddjFCu/9EzsPxI/rAV56As4JGmGkqZf+JDPxm40TMd
aMEZQHRSlHBzG0/p/MnSNGNfdu1yT22JjkaYb28B1UYuQc1zX74xOiBGZJLf5WIJ
Wnj+0BanjQpibYa48CPF3oNi0OdNhu+i8i1e2bTPGK1eZkSHU3Jn0Gpm1WXdh7qx
LFN9Teso073e/UCfpOJwp0N6MhVCg2juF9Ab/Nvm03wTrhQfmk4ek2evdZEjviZQ
PMhOks6TSRroe3SWQ87sp2wcF/1A6gpG7YZJRY4KrYxaDh1zAEPFIiElOOZwQO/6
EzrTLwDBLr3/v2GZPal9XvUkNf1t66Af3tMeob0wDiMCyx+4BM16t7A7nv3cVK8q
4QkFWM8Yf+jZENdXLPf5LoTw13WGzYH1YRJNg8DFA9LaSthrE0lAwmBKvBy77s61
xD5dn4zUHBORi19w8yzSuVhsCvh5PK+abUsv4pRMFtVvoEmr+fmYePPMshykyctt
nL5DH76PijkUDuKeGIOTJjIrZRGrQNrIw1WZtAnC8r0IqmrnZGgxoMi9d+8mFYph
gz0+7v1fiPzSupqGbWgi+RaKOk1SUBG9uAmqnq4GP10CLkvgg/59Gec8xWInyQPA
Lqi7Cn+0OlWX3sfpYy3FWX2pj9TRabCZLJ/yc24gq5wY+jHp94lON9m5EHpq3FPA
umgfshOI7vu70vGIOEWDG/yUUQGqPNjfI7riBQRjuyr6GuymRL8gp5OXyQlJHryq
nRGaU2VNpi+SovPQvY5nkqWVTurS+usREmqTRyM0jlNEjotXGnhxvwVc0C1eZrF4
42DP8cx/qkyy56+aSbVo9i8LD/cIWXr4TLqJAPo+gLOsRVBSSor7gsvgafwFPpx/
bGzgA+25xOYuisH/tv/ieacowoJ+mO3YF+gnDg8lS4UM6onwq9UOWFGPnqP5gcI6
wsUFoXZralaMzGPQyUwLbuo3S5JGqyo2g9zFO+dq+bAq6glAfI4Ao8PrcXpab4Ai
IrAgbVeLiBtnCJyLHocOVJgbi3bwWyi7jJXHClusX0MLsF0VRhvYnsLvtAjVinsh
R4fEtiypCYQO9eLQqXMJK05VMdvqxs2szDHhQTmuvpxK3qa4kr+RAUhrnB1WBSBt
4FJTaqciNeN46jKwYcrHkvpjST6Hn9k/gXkGwA1guS7hIH0SL8psjWT4+9gw5Dd6
QmMS5MWdGO8yi5IBTalcgfmWwAGZiRiW4ldTJR6w0oMWq7npdjpgROj0uWTvjRue
PEjbU6XVvzPr79uh5jJZLqxsNXnvFCM4S2X/uv9J+j+Jm+wnhM2gPT2I2fT2r4Px
usZmeNnIKv5oNqs7aF0gbvVdngRze075VP+jcN8KezPh0QKwoQsHZ/eba31i3+tQ
NOeS4R9vMkwMFk5gH2Xy/nlPA3u00NQMXcdvDCg6u0Tdaoqe84h3TsfLh5oG0gXV
Jyafz4vl9rW9NK1qhztA7A/hT/6dfEBrF3tj3RvVa3ZDgnrgn9Vuggn0s/nZia7B
IxOHNS/0f+iHW43SH+8ADtaXh4+yAN7RbtnuwhXKwJWeI2J0/8TjEpmBCXNDbb1J
yBSTdhYQ7ymz/+RvAaK41Ja8wQ7PT/hnwaQ3+rb/xsYdHYCd6t4pZaFruExj4GB7
JI+uLyqfpEZ3QL6U+SmR7+X44p5CPPZO6W1BCKm6p8scO//hBp5G4roJxeedzd0f
fbNolxHXpItDkQanP+t+GOxSmjx2Tu5MyaqmlPAdSBXhd8C6PIZv9l/146/LATgt
F60BXXGRwxmdJO6hs6x+lWB25ZAycXLqoKPxKYpi4r7hYSMhPwmIt2NPl7Sco0go
U8Oe3MK+wN5oi37XWP8wVdBxHX6Qax1Xn9fPcJ0b2/A7Bda9AFa2HLy7+U234+XF
yCSGM8P9Dj9TImQjynZHVTfMgXIjrxpidCZ0f4DP4Bo+1Fbjh12Y88zrfEpCGFgj
N0bvotbcx44GQTB4y5fxeViovf7G3w+yyiufMi3qpI0qyL3yE+na6/zvSkU6vDlD
xl4qZs7CzD+2lnuJ300CIg1pP9ut08aHAeUPrV7tC8fTmfD/ro/Hooxl8P2aq2ik
QbN/VfbrW68xuF+ugot0G+GZKXlnTCU6wc1f4FGKN+FXNHJksG8An2QI/CnrX80w
7JbU8j4OG8EuBjBKSDrQne3Oz1KhAxQumxTabvUIE2mfgM3Y51bqNUL34lUexzY1
XEeKiHZBEXKyjyQ6H21lsBVMeVMq+4m2PvVMxNzr4+488+PQwunXUwqCd82hvQwK
4AfTrGW5OWh2wsWKKCiIYrAU6LLDYqF7lOZAC0MdbKlMAZA4rEJWqdwajQ2pHwna
arRmG6EvNfydt84PzS8ZeOtZVJvXiPngBPjRhkXzYHbQORZQnLb0Ykv4vHSCG1Q3
OVq+IKXCsZ/Xp7gzlNumExp79fUt+XPNxg+5dUJ4qofIDxBdqZqMfobkRntXFvO7
TWO2MSbGg4r4dkBb9T+9LKEO/jydx5H/io9vsaaZC5f7fBRmO05Zs4inXadM8Dli
F1Ql3eBrJojHdxPIfkI0j8ziNtthG65Xw/LqH+ozGwo0hCKiTp/yGQT0WFxGB6nh
MMuwh+HRDLEfVQvVElcC8p7HAfamIBDfhuPrd+L6kJF4XDZQUv6A6EWUkAt49ElK
2K9kcjiiQ3L08C0w+Kr6nErsozyyFzTxlf0NaDOZmEnwKkt9YLojovs3rBZ4rwbT
4KWuknDtYNBdAOpqOcKDjhV9XCNdM2yYGherHsxmvCla17XtMvMq8ZvPYhyG8kAO
v5No18Mto6Wb32/sk9kAFy7onErxfuiPtsfSx1bZuYRM0oL0z0lWYrVcbMG7oxFn
vPRO1ZRNb9Hpt/kOX06UZsC1dbaMCzU61eO3378CuUpixfIiP+zN7Rat/shtKkBF
qno3M75P47mdSsDmeph5Rxv2yyJER8ThWeY8wZXaYoQVdNN7yb+K4kWBJcWRR0Ne
pSS6ACQwdGn01bENN3BkWTMlwCmYyxk1OOab8wUJIVkuvV4Y5rmT21OEOaaiyIv4
hbiHQxSS/s2rQRuDXMJAcaHxoVtWGFRcA575BnhEPdiX3EP4NNjC9x1wQ4vi9L/T
s26LznBJu0G8M7IfWc4CnxCPpNud2yrInCXxIDwaKqPd7J6r3BQkopaeucbWd5us
Y0mn/HHKqdzKGrby4ed8B3kNRc7bx0yK41LN629BuIQHLYjJPhftigx/ptbgnaWk
2cW+P6i60R0+fUqkQ8yrNLbYhvNA2wU+XsvdXXIOCY+OTtbvdInCBokVAJdFU8C8
26jCNcgTzFFtZLG4upsTpTiRhHF+RfcQ3bCoxDE5XxlYdIy0d+7LLxKzvsJFFux4
YPjfa3kkyLg6NdUjC2Wdj0uPs+iklR2SwrUEi0fIpocr/VLR41uIVxVw4Ca2nHJz
M+vvUKoecJ9Iu4+fy483doaAhc6lBhg4dQ+OK8pjSb4LETBHgeP3sgNlsHIaCGYT
TQCYEKP9gAzRZpx0jgR/zh19miq14ERiGrwEWxamO5Mbd6JugrToMhZOLlAd9eVz
sOIOci3G/rqNT458VB7EC/v7blKYEcH/0SR/lOEk0WIKoF9dK3XiqRChL87S7bur
Xqr/fdZ15EUpaW9ZSbtFc9RYegNN8/91LGyQcQKn6N7Z42wSGiKgG1twkTeLzSee
5355C7FWCKNAQYgPSyyIg7StEsP8kLeCB6QHnBECJ7lztwN6qerI2TCWbMB3Hzfc
hhX8oZRMZyvwWhCdKNHDKRNBnSH6r3vLDZaxljQGi3dWCG0NK3FWyxhRr/26QtxM
fphgMIpsGOc00VZwQgPBukFzwtbgcb2EZ0+DdiYO6Alcak/JkEuEODyh4oMXF9CF
8ME9lbNRJOGoI57/e8L7WBWXWhG7KZevnEOSS+Uq1GaUMpXWpypT2QbaFoUI1vxw
08HTAsCuJ0OaB1hU3tcXLeypTaBPMujBkUqMg+DIKzZNbZ+GLZi0CFn/XpeKXGz4
mWgavBik+9DP9Y1PgRhfjfhFQmHwuinZ3mo4mUDuKxdXlPbEpIbEeScJ5x1RvS6H
8IqeyttRrWefEV7dW9HzAD9lVhsBKde0vmNRjWSDgpPzY/XSwSJMkCDQ+fnLkjen
hQy7o/7HWF6T6rXK2WCE+UHCLNT3bb0/yEGgdBSQ5F+fSHIKUzfYBmD0pTFUcMME
2+LrnJUnFt6WpDPCW5y4M/WJVj4f1+I8IKk3Xcg7YfYO7TMy5ExXUwutqJ/agzjD
qX80txrTuVw0Lp+d3r7ebdK9Y6EknNj+s7BzH6Ys8uYNolltm73/61VACOmB45YT
OJdkjiMn3TTQjWfyIpR0sB5AcNlWSJ9e2NDyYKTKdFQjmBgXRvfC85uCQVNWqlMc
jSj6dvx5oHl6AlwHtvBAj7XfI1333txWlBUm/6VTOKI3qfSv1kklSrmsmFnAoLaU
+JFdtHlqbpLP9aieCatbSLrwrIFxRSEe4ewkktqCiG41DWCD5dRW5/n/LOIwtTTF
ps2gaDz+8zsyDIdFMoS0zrTPyw6hY09BRYcu3bCXwCwDYFsTCexIjOhSZqQy+g3q
ZkVqOeCQviG9Z0etWSrlRCS6ZLGXPGYn8b1oYVYHM79szprMfV6U1LwiLuT/F46o
/amfW15zi2cmnllGz5W5n7KUECo9c++u2iomcUuTH8pZ5j+zmQaDItIzuF7ZTQSb
n2rsKvqP3xTzzyYLyx/tSGf7NvNPgMyk/FVuSH4WAkzbD0AFXLxy/iMJTg6wavN+
khgtRROfwgyOfTW0iSYVAou8Suxz5G1pLLOpVzCHaAyVSzPcnjpGZrX7MpvLJWDz
vJAuvL0FyAZ0gWg6Aw4Ns3vLs13dei+g7wYgPreVNo9XXaXrYz9ywd8J7F+i97uS
lY4mYv0/qMjScOvbxHbn6+g4T7YaDoV6TGKe9uuChf+qknyDfq3xMCNb6p1dy+9l
jXDTjKz+18S7qyECiENDYtxzzzUT1D9CS4WRduSgkn+vV0DW0Rud1fYF5UQlJ5dC
2O2vttj4LVMO5jgOiF5hR//YMdsIjoycZkg3V+HhTlg13dojDfcuYFs5s+W2VSNC
79BrejwC6Ase7Wv3MqgLOp4F3vXqiKhwy1M6h1hXmjsZDzuc1DYu7hUgYLmzr3X4
2WH/BkoGSdNe+xsN68eCMgxbKhuapNYmtKTHwdZ0llpunGH9DmWp5+WAYvAM6y/+
enO9I19MowxQRCEHJWnDt9rpXBhI6VoGjha+uNgZxxUC3Dq46AZ6st6N7vErZ6eT
Pgs18cEUuiLyt1TvKByQVk7kSjErGM9WiSkde42ZW5i7QgsUhiYmVFBIIW2GGj1G
v6xrnn4FO5A8bkoowpkZMQedOGQPhQgRAtAJ1pqS5FpX4zRX3kQImeyfe5Hd5quF
BNJla4VvtoRY6gX+wHqxy6vawYWZD31nEt8wsl9Bz9gqGFGjINYyUDn1XPwwV0g1
mKwEjU+EmRMp9s3I2a5YftsqwGCXTw81AsNAQl4IruAwqNL/0CiqOyaO6Y8NNIwM
Gg3lFoNHHpS4ldKh9oji/qXaf0BoXdMlxElSKlo4O/ea8pgfkco79DjIDImXCbr7
9OSdQ7SmGv0sAR+JqsE647zi9RK0tWLxTHfmGTiSxNMibMS4Wiu2K4PtdUn0/+MM
Opjq/kvbKb1N9g0FhAjeQJBeoQEavDmfZ3AUbyH02jb8tAkYfaa9vvvlKmsGT0Gp
kFGzDiIXgZzVDEmFN20WllSKX3f1yRr6Fux0esBBYGhx14qPzTnwvnd9f1SD0jvR
E9uAYGefUcN2ziNshs79v0WDVMWZYHdAmE7s9r50rw3kkeWs5r68JDRW6P0rLEKa
NWR+ktDJZPCLbP8vjQ+1LsECB+KpvfT8hNDLsDNNUTQL/zwWrWb9gaDocYrW5jVQ
n512bbVijpB21tdEMh/8HH2tJv8P32TaE7HRbQJYmq/bqZuoMe36LdDdZTWxVbkb
QJsM7BU5/uZyBCD8AiCwX8Fjf/Dzj1vJYRSLC0iItMiH9subxo2zZNpSgxI39AmU
TioW3q//hY3+dYZwIx0z60Q9iPqOPPZsyRz5e/MiCh0FmGGwIihCvSJg/v7oho/V
J8tWmC0uX0Oh/T+fL5Zswie0kCJwah6hpHkKq6utziclPIz3QfwU2GTxJCsjjhqI
Op3D+YN1az4mEdUCwCZZ3RyDwaWqkF6YRS7fRcqafmM=
`pragma protect end_protected

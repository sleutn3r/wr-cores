`define ADDR_SYSCDP_RSTR               5'h0
`define SYSCDP_RSTR_TRIG_OFFSET 0
`define SYSCDP_RSTR_TRIG 32'h0fffffff
`define SYSCDP_RSTR_RST_OFFSET 28
`define SYSCDP_RSTR_RST 32'h10000000
`define ADDR_SYSCDP_GPSR               5'h4
`define SYSCDP_GPSR_LED_STAT_OFFSET 0
`define SYSCDP_GPSR_LED_STAT 32'h00000001
`define SYSCDP_GPSR_LED_LINK_OFFSET 1
`define SYSCDP_GPSR_LED_LINK 32'h00000002
`define SYSCDP_GPSR_FMC_SCL_OFFSET 2
`define SYSCDP_GPSR_FMC_SCL 32'h00000004
`define SYSCDP_GPSR_FMC_SDA_OFFSET 3
`define SYSCDP_GPSR_FMC_SDA 32'h00000008
`define SYSCDP_GPSR_NET_RST_OFFSET 4
`define SYSCDP_GPSR_NET_RST 32'h00000010
`define SYSCDP_GPSR_SFP0_DET_OFFSET 7
`define SYSCDP_GPSR_SFP0_DET 32'h00000080
`define SYSCDP_GPSR_SFP0_SCL_OFFSET 8
`define SYSCDP_GPSR_SFP0_SCL 32'h00000100
`define SYSCDP_GPSR_SFP0_SDA_OFFSET 9
`define SYSCDP_GPSR_SFP0_SDA 32'h00000200
`define SYSCDP_GPSR_SPI_SCLK_OFFSET 10
`define SYSCDP_GPSR_SPI_SCLK 32'h00000400
`define SYSCDP_GPSR_SPI_NCS_OFFSET 11
`define SYSCDP_GPSR_SPI_NCS 32'h00000800
`define SYSCDP_GPSR_SPI_MOSI_OFFSET 12
`define SYSCDP_GPSR_SPI_MOSI 32'h00001000
`define SYSCDP_GPSR_SPI_MISO_OFFSET 13
`define SYSCDP_GPSR_SPI_MISO 32'h00002000
`define SYSCDP_GPSR_SFP1_DET_OFFSET 14
`define SYSCDP_GPSR_SFP1_DET 32'h00004000
`define SYSCDP_GPSR_SFP1_SCL_OFFSET 15
`define SYSCDP_GPSR_SFP1_SCL 32'h00008000
`define SYSCDP_GPSR_SFP1_SDA_OFFSET 16
`define SYSCDP_GPSR_SFP1_SDA 32'h00010000
`define ADDR_SYSCDP_GPCR               5'h8
`define SYSCDP_GPCR_LED_STAT_OFFSET 0
`define SYSCDP_GPCR_LED_STAT 32'h00000001
`define SYSCDP_GPCR_LED_LINK_OFFSET 1
`define SYSCDP_GPCR_LED_LINK 32'h00000002
`define SYSCDP_GPCR_FMC_SCL_OFFSET 2
`define SYSCDP_GPCR_FMC_SCL 32'h00000004
`define SYSCDP_GPCR_FMC_SDA_OFFSET 3
`define SYSCDP_GPCR_FMC_SDA 32'h00000008
`define SYSCDP_GPCR_SFP0_SCL_OFFSET 8
`define SYSCDP_GPCR_SFP0_SCL 32'h00000100
`define SYSCDP_GPCR_SFP0_SDA_OFFSET 9
`define SYSCDP_GPCR_SFP0_SDA 32'h00000200
`define SYSCDP_GPCR_SPI_SCLK_OFFSET 10
`define SYSCDP_GPCR_SPI_SCLK 32'h00000400
`define SYSCDP_GPCR_SPI_CS_OFFSET 11
`define SYSCDP_GPCR_SPI_CS 32'h00000800
`define SYSCDP_GPCR_SPI_MOSI_OFFSET 12
`define SYSCDP_GPCR_SPI_MOSI 32'h00001000
`define SYSCDP_GPCR_SFP1_SCL_OFFSET 14
`define SYSCDP_GPCR_SFP1_SCL 32'h00004000
`define SYSCDP_GPCR_SFP1_SDA_OFFSET 15
`define SYSCDP_GPCR_SFP1_SDA 32'h00008000
`define ADDR_SYSCDP_HWFR               5'hc
`define SYSCDP_HWFR_MEMSIZE_OFFSET 0
`define SYSCDP_HWFR_MEMSIZE 32'h0000000f
`define ADDR_SYSCDP_TCR                5'h10
`define SYSCDP_TCR_TDIV_OFFSET 0
`define SYSCDP_TCR_TDIV 32'h00000fff
`define SYSCDP_TCR_ENABLE_OFFSET 31
`define SYSCDP_TCR_ENABLE 32'h80000000
`define ADDR_SYSCDP_TVR                5'h14

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OvK1IU5Sq6f6JDh3JZHnSC8dm5lUcMLPQsjkLh7IteckBmceaRa8w2nCRlKne+gA
cfXhMJ9QhHzdPmWrTofpHVLpS5s2l21qePSe6RiiYE4WQBTPcD92/XqorZcEYCZv
s3HNeib+NGKg3D3V85EeNykDdVpGtcqJqTuYHHtTJjE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17984)
B6VovUKvZdjrJKxgcDmHhQfIDp5nVxRkf4bW6O8p5Kq74XxFgLTPdIBhfKYuvDXV
xsg/sGOH9LMoU06Q0jbTQaEZpYgBVAoRQL3SofvzHCoKS9t+2pHXYheqFV0U2/H4
bpg+bzrg+2+sp0T7XarmCXhbKvWI6nza5QoCKCxgmRB/7iVc+IN28OifuAayxkvl
M2cHsmvDLgia4VY3GqgilxVlWNfa5uHgb5Jujr3YAI/GJsNe4C2yeX7kpmxbp9Wc
we7yK0dC05ul8NLHSsFjyqyFekPfQ5f5tbTEMoY8HjznJX6XA/SA8ZDIqVnTmGnJ
rZU52mCUg3eV2dtVbMFNdK4wKoyiA8gZTxuUf8+zdC0yGPFcuwr2QrroTo4U3CzP
T18oaxbnhS3YsDA1Gg50APR0CySZzT5raTSfPETjl1rGx8w8BLXFL/spoeAsQ0vn
ZZFJIPky8VEDk4j9jovDYOVBt3ND1vHI5dEadGVjtYgi3FgE5cf4khAPeB12sOB6
oj4GFnLYw/5gatZT/cb6DFfYtaeBjYERiHRtROwilmYJNzqmaj7Z8+oySzS+nNmC
TOKoUw/EcTn13OhXKI0Qyi3X5RZdzSADseJtUAI/vRJpXOTcjeMAVgnpQfm9bNX2
l57M1Nt5r+OexcAdU6RcysjhdhtdQ9wyzh/MR02WKlsMQkpcL0jY8RjpzI17w6hs
WuZFqI2s04B95kkZ4DNpsCCAs8wPEJ6e1wPoEhkdZuz7cUkAe52Ri1VqIv7Lj0sW
syr9VXgfvyj2/mU185Ibm8XHWbSWUww1yOhJdSB6YhnVaCo9XElHU8EfGmtYvHHU
wVPPrFt5BsO1qzoQnRfEHVjsrl00tfxfNY5Bjs/XKUAseQ9/DeCllozjqq4NqVa+
Mc7B7ReD6QpVQ7qTlpT0X8Nr3GHPK+oac3GYX3DOVM9DrjXbMUKvgjMIK86i07Af
0uKg7AdPyFsmHPQzkJuj2eX3qF6C65WQpEyiqDk7Tz1oIbGsQA6U7NXXTQFdMHNM
t4hTBUgpuD23UrcJTBfJEzMkxFGEHZFyGfrVBsvkxLZ9wjysb0aAps1q5EncYsMX
/mpWMzRqvcJT4CpVGMVqBhi11zqWwPgV+KoDwGK0j5v/XO04MPCPseUYB96oPwng
P+WQrEXz1it7XLfsSuRD1Z4ZDshkHMahyGZRgsLPspbhZTNfNjQZEvKHc7ghs5ui
d8eb+gEyWTh5br8FdNFhdQfFDaSCwN/ZpwNO/cq1sFDURiK16g4wH1hP0na+R+5n
lkHBKCWuKqqYKKspiRgrG3zIPqHzi/FwIGkSvaIQAQo2wBLzOQOa+wFlzNvHiu7k
pbZwbZfyuxvtviU9v3gIMR+FBCRxdlBk7j2nLP1IjaSQfXu7lK8J9ITbEG8LEHZM
LLs3xqqb7Gnt5NLREdNcJl27qkXZOT1ixhkKhcmIAK8/kT3U6zYXQ6SUkyTLHa/H
81K6ML+EPxP5J5FB90F94dzinvZxAsycju4Gy1Oq5nDrJo0L7jBzFxLC4V2Toy7A
dLcWTXHFIUTN5zlOVuNHK4p2hL/6xpmIW1UAKBxQcgxEkV3Qjt550ALTpotQQ77Z
ZvIDK4T1uOhjszcRqT+UQTWJSzgs2/rtx38ZTcM55ApteHpgIQv/Px1Llhnyc4MU
wSksLoai/CTc5ntrVCZpnWPJ8Yp2JUKBAjh54GCUS2BfYqQ0pcM3X8zKhTP8XOzD
BheOSN56gYHV3K1/63/9G7tWnQkaBFyevdSlpSrZDoLbIHWVtplEcc5l1AtWTXAe
ekLRmDtVqoePIC6YK1efz1oxLZB1fONEnFtNf3JdfaDTUtQlUnK1AGA7AttqaPU8
ijvT1BbfnER5og7y3zTOFGbZc2hzRI57oQWpVROh36CL2neL1N5TeUmla5FJ58w8
9ESjh8B0H71mAv3Bbj5m5/6vFgp0A3RgtiQeri2gj6bI7Lz8DAprl80vQzTxoFOe
iiruXaYFSW1sBngSZg7zktvGzX7yjDU8z9uleHAqRHs4h/7Xyy7RSmOyKbwwJCtm
f2afUqo4fmTp4vjLzi2vxB5QMy04b5xDkWKZ1anm1RrQ0WZ4nST3a6D6hOxx9ac5
jMn8/SqSnTlIg8gE6nooO4H0iknUiVsXfXCdvi1EExWfnzw+EJnQp8atyPe9pvHL
+8kt03QPXH19XswE6hFQ/rxWBKv6J5GFVnDknJwQe5PqmBsAprWwa3iPiLQm3GEo
YS13VMqaiZX1wSz9jLlV8KdHiseVM6r+XcxjB/9Q0WfNJ0BZBSi4V83Q4kxn/+jZ
V6MkCmUdnT5JjJQmxixqUuglW1RJ9TzKtf6bSWyDgWtGqwsskRQ24y5hrCKRhmTe
4S5x4ef8FIJpHyYOYne2hV8tYxD6DEyDCzjC3UAbru8f9uaw1pvp5kysWFYEbbUz
cPzMs6qqiv7AmZweNXRk1rJonN2cfKmbg34uGivUBgIh0vkZA9sGaolyu95pANfZ
Tw03iVmKWXiWTPD4LWtLmLbJUyoKiSqEF9619f9cUuli7U/BgiqE5W5MKB8JYgEE
eiIpzlH2xvyJnh/1vRYz0Rl8o2XUgjtdsdz3ggmFhBo5y2+gEuXLfgW+h220letZ
BZfLyHhWNz2E3Z/87NsNJ3JFWElbaQQXmz37MuExCcOTft/zhLN0cUgImZb5/tj9
BVjGtG/IZvPq3xi3aHwm3DF58LlDMnkogiFYL99gFO+dvPNUFw+qqCwIS7OhbMPB
PLtsVfl1aTpGZ+VlT9RJM/qGTT3JHV1+u3as3ZPgCE5X/NXaeP5sXqF37ndFPXc4
o7lV8XfjWNP1xrTBK3PoTVklDIntvHPF5j1JIWGFCr/AMFnaAqGcNqu9tlEbYGSz
VGxRA4tWZ0OoBIbZs+qEbBPimREFWLtDtdPa6BS5zuTNSCkug/yYl+P5ZTHlYPn1
GRhmKTPmeIPxfcWGizvNvU1ppqAVZYmq7PkGExSYQYsCLn9GIovLRm9RrWsOdaPM
p1fs1ZwSVw0AXU3yoMGs3S5xXrGvFJF1VU+4yAxBd3P5jcvQ0z//PIgGIE7bp5zi
Xs27+Y2t7jOlP1WaHtlf+HP1Hc56saFgInahg78h0dR+nqw26R8aVA5G5R42S8rm
1E1wgBRgJYYPGPtaa6zgJrDmjm7N+3C2VCN8NSzJY8b6pVmvymrErHvuo5lvWv2Q
aQJ9DZu3ZroHLK/R+WaJKTIhgLUSI+obqTp1TmCHb4OjFp/2DokB9zSo2upbqof3
BF514eU4SyVIK4rC7Y54HumEMFwyQ+G3R1VLn+ves6+zyWJ/XVkMzdbQoyVZKMZA
zq5EJDabEBufu/kn2nIBMp1YXGIbacFJz+oukcNiMBeoDyHY1s2hvyAE54gVNZ4e
NI7W56vTNAifc3XjPXujs/ny1PZp53KbfKKh8PCJl9sPTf8JTzJt8QPC3OepghXj
fIc0SIeLizcBEfLxQrSOfErJCpODmHu5J0A8Z7gjZR3CpgECBl43wWBkKGSoOqva
Ac/sP7CVKEs+21JSg+YooVvQMAvJOJ6ehDGsAAmziTGOsf3bY+TjlmqL5W+7boSW
0Ictxjxmex6m5sovwAmlN+mqGuNU5z/Ko+qwWP6450AE57HtZFbqGSpgXuPGqCOT
bM1QjADq/P7nR7Z5WEMVj5NWSMGF4mCX7AslWpGR3QdEtfYB6laH18IXF3LwQtAW
IBA36gPaVcZqcfOLn2vM12SfiC0XHyHWddUPzWFgHU4+YCntIOMNITytmePE2bFT
dxhnwfInFsJPW+L3kCP9kqA1yO3EezNbV9e7x5+mVK3gQrcvAxRtTu1FrvsAr28v
FlRXDAZ1FzFFv/JXChujaArwSydCIikNcviIqqO6L2V5USrMRLxEzVqXiymwnuCo
I8X9+rMaUv66VbafMjWWHW1WCrlO3lu5HYk695CKjCSZRCJbdau9u10WvX3vItWh
FF/5YwHwgRpL1W2suSR8pLe4TyDVroY4W4C0emx5vmWTlfihYtU8gHnyDCDRPgKn
iRRlvRLfKfBisQiHvVep3k0Qb+ThqBd8pv7FqfR0gM5tswpTbVBy2tum8Sy64MSu
vh2/mdwlHPndf2Z1AusOAeqnRcm0wnu5TMpJ38qMAKawi9g3I992SivvbrUbYmlg
GqNn1FQrSqVHUyVgPCEwEUUJw0qGiIhXS+Ty3HHvgUxcKsqefaO+8ypmqyHwqOtb
eKWIh9mFbL9HRjbcXIrbCJAlglIPsfe3xGZvzTNFOj3S/kVFao2A6kNjdxeo8SfT
mKZzXBTNGeZoXui1DMW+p4AEIx/fPShrhS+MBu4SJ6pShpd0JruSqM32Ty026SII
9SUJPxx9ZooT34lAfouUS6x3BjRzYAyMNR4SUv7ya1yvsHzkB2JDsiLYlxXQPu7I
CY7CGJ6AhDCYUE6SVma/dgBxrHnxOKOAppCdeJVba5wLaTYTAvT2kn2v022C4M+v
HV5rCfjCcM+O/BMYigqFbUisnxEUWUzMjIhngJcCveDF7D3OsMAZHNSx3SSkAXue
jfulgPW6A/s/tZXLvruETr8mCLM+Mz2MhwjWr8uNADWzTQmIO+UQQ6du2Xc0YBQk
PM3s3Kk5KCBM35pWAp1MZROZ2Xt+sK+Xom4e2PLxxuIqZkHSLud5FtXpXh1+es6T
Hr4aqlLR46jBYBmzpYlndzAVTCB4nbHr3pn2F4HH2e3ONROQtO2Anl7NJ7rVCwwg
nA91F0pZmvS0JzkqoN/vE4x+EPBiaXknCi3qN7ywX2YnuOqF6eY8aDhGaKDNBHmM
jQYtOiFmxwT2QiClQrpjN46LOV9dSKsa6lZO4IoTDRcAxqFK7txhzutD2z7OwhRO
lt6dDif+MNYHWxfdZYW4UHoT3DzV6DZEt8dCxYvQmMweD7XdAoLCJ6ZJwXuzYXs/
N1PtfiN7mlgcfsUQEYE5DZx9x7+r20NKowxA4iabKm3JDzbyNITRVha+X2EsvO2J
af/WF5RLi2HuuPOBHZRGVx75Upyp+Jc8PT4S8BYJwmVxltHDokPaXWiVKARukM1P
3HcQMrAzQGH451eyxwJp+KdCxp3Wla4pvjTRrs/cS6uo+3VkQsCX1wu7qahBllEJ
uadmDGFbwQVyhcvUaAjxL9zpusxepIPLc5Ex6iVz02cd8EhDhsZAVD5BM9uyGfZU
LVCQEmsny6F+cmwLLYcElF+vPiG9iYwmNeS1pQWep55WTMGbAtUHJLR2aXTwvK2u
aWDJR7N2e4IGCYm9YTJUZDR3VpeKOJMRw0IkDsXis9D2D2RYjGKwJhQGGPnaN0B+
jWjNswYr6BQEg6QY0faAw/lmC8Xd4d24IlEua2hTrgMQQk0lHne7M/LMSCd/yb5f
wUsPkFa0X4l7fiLLqSFQUk2KrLkRzo0uSmwABLnJCDBwUmiY2XRswFQfJQKTcxeB
XK1i5Kj8Nvo/akNtPe2a7Z4cY+E31my+OecyBiWwk2RqW1X7J8tMEPiJSqQCcup4
5022yDmf010wYgne/3O1r7Tn0RwRKX+VNR72X49BpatJI1A41iLdz0TjTPzftjUf
YWofLQSQ9Lj7mGqS4ifmTSVmGAuz0zp8ev9AvVMlRfrIMJOcwAmiL0S6q+qqCH+q
B1Zp/lxHlSswEd3z+RJKenkvAr5tXxOw8SOX7VjCtHlBLMMoCiCCuPbHh9Nkhq61
B9HYjVGqrM4GlwdwBiC5h9JCCyoVpgqp0TiVRhGf7b9cen992QAGnnSAx49fIe3D
ubectfGr1W4ld/f4WIJBnLOq5XV5kYE2pdZeG1TdPh/Sghz1G85J8wrNLTHj8rF4
bZRGFeFdfVAWezPaimMEv0S+AG3CIbBBpr6USiBc8RA2Iii2wsWR8L5DX7su/LIn
yfQuLJUuAJGCLh0S991EzYEz+xRHSgBo5MSpADkKdROT4IkezVAQ4KRf9Un9gcWw
UyNBho0YcDqt1GZtwADi7XZOBjgyR6GHi2rkx+4sCSJCXG99hM8KvgHdXY6Xv2uu
yGDOEgRKWmEfBYqrt/V5VKnRGIgecDpF7gK4MPFSKEIpsDUnID1nNAZvogOqtiBT
JX8lS28mY4d1K8XKIJR6+IysEKjKN7crcyOsu/uZcJh4fBxWf9TtDv3tpbpechnW
Xb0p0VOUYwzw2Zc96RiraVRo1UI2H1n7c2HY/b6SV4IpgzzuaCo0Z5TYsy2TAdQQ
D1NWPbfMI4Ap+U39B1LMnl1ZI6q8FTjX54WCqstt2kR1QzudFBY5o9eSXIm0cIo2
T1qh01AP6F1XC+cOaRemPcMqQ1/B3aMTCcW9KHRLU6jXXWa9auQ6N7GGe4ScMk8e
DzZb/UpOt7dxFHXbt6DyHB5Yj/kiZQhIvQ3feP04Vp+hdwNXhOPZ59VRs/N96lN3
iM85lyHPEA6+diWbZSGOWhF9ZRh10hD9iF21lDn75eBVGZfk21TQ4E3Z7C6ZCNAj
9h1Xf3ko84Wexn52gtprCVvzIVQwJPTF+F/7kFAb7AEW4ht0A7WML+04kq47mY+8
3/tVl+moKJUVURsWTMQ1J5t8UrBTSj8mRMx/k+eRPuFZfqtzDKoY/6lgJKki8TGz
fCGgoH4lVj/3RF1UeZFSCbU9CxKUu0gO63wTGtcj2r9t9Sw8YFhgKHvz0k6jrALd
iBjmvqJDoxpjtYSJahhOpgbVFu4RKhQlF24JSu3HqZeRnmkpfsiNIN7+KCj9fhRv
nmkcCL203XiPFWaJSrl9Yf6umfYRPd+wxDHBACAGZIKEtGcoeB/5jJM68kkfOOIn
H1wLVVrRQsjjJ36RTmR2Xbo95lPimKiCqhROe3gqph9H7PYV1ywIk0eKXqY+fCux
GjynDhnEmM1ERsNezTB61bN2VZKTYKbgoqhmt1UV3djwG7SmRkRJ0K7C+Lsa583U
7bLsfG53GljCs9994d1MX3SIkLUGUDRr6Z35sVbi1w0THGxCtYgafgpq05nWoRLq
tE0xLkRSwvqNtFFYV5+IvmTj5A4WPd5xkOQNbalPKeWJwx9+7Zr3g2e1haQFw3+S
8ux3cmYGwP3hwr8yfA84vanmqhxoa6wgxulqG8xdCzp4IetJN4sf87ud6FpBmMup
TriXMNFzPKfGCc9Tg0gn5OirH7DC1xFwwgFcSQ7p5Ywrad8ukLj4zTejIR3PxcK8
KH95zKjCA3XeGo85o/2qpWiFa9i2yxOei4Da7yvkCUUMM2S8hNajiZhaL3459IbR
Wlc8LPoRnua8ZKVsL0FPme7Ggr6kZXiTmg6SzDKwM+lnSLx1eQN9ByUgjg6bNcmM
NgN18llRhqvlDBjD1eXDBOQ8iiP0nkzNpdtrqq/tK1xe9zxPc3AJnsUoYFLjTMq6
c4eRkNKSsO98cWsgfwVBeUBMbaZAnKUA1ZBX2J8UAYOtDe/A3ugXQaT0grKjdBl5
1N5YFYJGMt+Ei80SU0u8ba5QVXqCpH/MY507y06ce9g6fGzTpogWsEugT+LpKKSu
xVjC7JYeP88noPkxKPYpiFW3WKy4J7WVqtCokdf3uxg9Gm3/kuOEBB8yJNk1r8Ue
Ghi9DV6E/1CyT6uBUmzLlDv7ptzA+UsUyAuxkjiKQbzcnjbABP6r6pK+ce6Oy3IG
Ot7RaYnBM8eXcUpSC5/gOHbS1vmySG+2stqANah6K+jvLZKotFUUKjzM0jd2MIjG
9QrLbeXgvXz6VjdfnfCkRqr4qA3oERrm0twNwfJFsv3QH4AOQUEjk696+YfFGK5z
dGZRDLWxZ5k0G2hRrnq76qcytDdFJYEav7+7+Kp+ygNmaukkm4EzCb1GpFEcNzX4
xjftmdjJmN4sgSejeMdFHkEffBcfaZIP7mjAO0nBQTDy7+ZUu29I2fAIiSiuKL+6
MIe8QaoHdf4FQl8EAqCJ0fSSHJUV9kYAgnTgOK9LQYPEvJhiWKnq89N0o7Y+uyfM
Z6P/m+BQXqstl+kxjlOUzzNismlndPCpD5EfOc1BH906q6SGvSEVcCjijiKFhZx8
TT4yxN3AuodWadBoh39U+2q44Ad+nkFKB38F2vpZ7JdCV8Z/p+Wju3osorVhjURs
leCdR6DXti/hW+LXpw7EhJQyUcwxwZ4kOaQv7XgcNGIFO0rCmRlJI5dB3w8eIl+M
1DF10qjAntgYealr08qp7w/2Os1Ca3+1AyT3I45dHPCM5Dkljrgcc/j1ITnVWPCi
pH9+hhhz43zefXJ9JMl9rMKcqpJjqI5yaLmADinuFJrizZwcBCYy1NwRlBqFOlvo
2oEZ8SJ+Mg/Y7deokMeA/3GeF8sZnsC3oRx4bY27/oVU8FmKmStYuxM4mhEQdUGU
9hJmEuRzbH3iED+lI0DyV01WoZWi+5fD/EG3bA28dfZbRIeu2NE//Z7lDRP13FBT
sK2wPMI5ymz5Eh+glJ/HHbaPcxB7sVkN7N/7vnFibooeC/tCVwSDh4tJs9/tfMz2
E56+vmE3Jm94mHYibW9cC6r4yN1aLuA357A6QJ5RsY/f7iB4l4va2DwH7BoSjd5P
ziTSizcBfDvIL46UxALR2s6GFTikAcf+Taqp/71g6LJbI9YfW/yHK4qE4eeArFZk
wozL0rUJq328cMkjoyRFl9NDoMCOJtAD3xYWsnsTkmR/rJtQxlFUT7VeUsPGUS3E
xJPMFMvDR1znb7U4YqJDVSdPpJ+X/1oJN/mrf3t2pOhCBHM5cpFwwtXEFhhVCDt5
+gnr2kXiOZB4m9sqek5NEcX3zzrys6/VquGKV9TlslB/H1lY6mU/cfl6RjpOwyY/
g93HGSVUV6+Afi0mySg40NAfSoZVencsmJ7J/3ucqSS0+VWxrjLOrQyMSs2uQSGw
py0019zBENzxBUM8IKDCffkX+Q7G14gTqNx9TtwwlXYWUN8kEud6wZfU1cz3K1Tj
NoBxPguoW72rkEqcwVOG6gl2Ec6y3xFHqFy+8MGZ2o6eedjFvD9XYhwssPj51QxF
6lQCUmNP7iTQA/7EQzIflumXRNX8Y6T9adf07ekE6F5v38hiuI/Ja6LwSkS2lBVg
s44IO1gNEPp43Twaa6ePSlLGjKr7t27G+sczjvB3Wmysw6GAw1KLcoyvz0YWy0CN
1eERhh6vDQOlRE67Cqg8KDIUm5acEllaeDHrgwrSt23NtOoii+VY9DOnFIGDyNFV
oE9o9AYVUtFls1oPW8SCN3ZmuCsBLul8S019gsbGOjSeFXMQ6NfmnIi3DZGP9TbC
jnjCZiUQV1QfliCtXEW6QhVFICcwXCYJFJf4NhMXj46hVrJUlKnSLRfcvtQx0+73
V7I6S2m6IxIeKOI9r17uhc8eBMx5s+kORq6vKr4+l7dATTDJe5TqhzyTJ+aDl9lg
EW3b8r5E7YZET20U0t5WcDylEFwo9kwRh5RMCVH0cAqePrsPpvjjeY4kLcx1t/if
SzkzfEi8RGzDbCYbdbXMGBI0BzKQxOgupyebBnC7NVQJgPevRUr105/i/Hq6nX8B
1409wIhypGJTlUA9s4n1eYrR96PRdy9tDRy36lv1dmg5O8CYxKEOeQ2u7JLTO8v7
7YFbzbe1SAchhtGp7tek54wM6TUPYJZwDeyoymEsY8LpBNooa3okVVU6PSTZmwqc
pBypzmP2P5j5q0iCl4M44SCiUasgm69YOdfNQOegbJ1Qgd0sNI7CTPNoxuIVL3la
VdlMDHXBgJmSouDHnUOY70lzsdqTw/xZnmSa86RaCnPDVlKftbcP4dgZ/ieQzTmm
uO9FpbATCi4udfx9AU0sknu8ybTjQ40gE7Io45r90d5IG1oDok+vCE7mgLdw7XA1
sOWDNS97S4V9nkqFaKLYqUjlVyyun5LwOSPXW//dMETzqiBryMKQHOxYr2DMyCom
MBXYXTQ6nEymTzYkRFUW0HlBxJzqHso+ccguNrV8B7Yd8cu/+q2NyiPezCThtKHz
/wmXclgBz0z0DjicmSQyFgl39GDTyevd2o4AuEuJ+RsdvjdICho3i4cvdGa/h98e
OjQENRpaoRqpR1xZQHPh+Rujorg72iHdx3aXledLPsDLVdpXcpZP9taDA/D51CNm
P+r8eE87oGuTBEej3K1pejTGU9xCBRMG0haUZYjJs28T3mfGl/kAA2FPm2zFx9GK
sB2BjH4VbSUgsEkTpLqvUH0IElsqwZZkR9djLiOl1/W/W4+J7wiR+pBoCFqVXAjq
BkIsimrabjSDNpdmQ+IdjavvLQWsnEjJFLEiKsIwcdMEtWlkuTMtSULOYIGuyxe5
Z/MSUsGIJwiL+h6FBI+iLPdktcIPImmo1VfWRjlcaTrolRKfCpoRbOlQwkFDQIJ7
tgAaWWCcPbVAFXLAxtnhTqfNzwZKCTHMeHLOT2uHu8D3UItodfKifsJzdyOLDHUF
kNVXgAwE9ePy3p9+a+2aDE/yXEikMVIqqZ2nrLjAXCgjI5uaDzYyZ4mpgSWOPWNr
wvu23i3bn2hHNW4gNNkcpLlGBZDTWz7+j3Djth/1O3BKWNC9E1WT4/JKBHkRH7xW
hciljlj9NTBjFWmPl4oA0NhJPBh2nxYEz2JuuSJVqDNoqvw1UAUtnwWWqFW6oYAb
r7LvbFqcX2CNFPTtLOM12hONbPjDKkN8YHgUfyQLU461EUsEwJs0kYc/3P9EaEOB
D2nYocT5UABQiGGNiSVldJmtHiBACHPreUSWyFBidGvolRbDQ/elJlcaX0Hpu4GK
NxOFTOU6OskXP36CNsrABHsHNHrCfI2WZGQ2vIm40AMVenHBUTp4/nfak9oFO0+K
m5wqtGIxLO2jJHZWOSkePpUJqJvA+DvC6PF1Nqi45SSg14/q6R3NF0iarfaDM6nF
K1vc8KAbmLwnvhHlXYfBW1ufke1IqZrnDLj9+bgjD7c4cSy7vTaSLtBkB7chC9n9
yrze3kvxJYUmEVxh4wHNH2zyK1Hv8syw0GMK/11Uy5lscYGTYUpDRIOj86z6we3Y
bwVR9PCCuFftzCkiPsL7NPRqDMi8RlZO8ZcMFENmnP8KJEvIlOMfD56pMel5D4Zl
nZayYYpnh4fXoBpivyW0vcKz/wVGFHRfFfLp8qj9ZZdun5UN5cjoi3Wb3yZS5fG3
9OIihQtxA7lL6OQCUyu6YzxYH3Ga437wG1uezSsggrt9ybCEEEt44B5iO4+Nxens
YiB9OuNvQjGh5jrr/2N/HsWLxD0wRhC+/7nDdZ3359PKGeN7fmzXhC0hgghv+knV
cOWyRf1MIYnjy3VtFXMy45B8vg0tmfmuh5B5nWw84KhmizBLAl5qPxrIuPc/x6hJ
phYfLIzR9mQhYVe9ywu7AfyTzkPanFKaOnMNsqvWvArPHyLNz2q4h5dfc30kySqJ
PRJCpN796Kk6tx4knCq3ZTS+eDbdgpR18kpVCBx87E6f3Ej42EcHvaDFFHd1wLpZ
2vYo2OMh009JFga1cHpZIHkrybzQoTiYK6I43FMkdk3ffeVmw3iKfZkJHt/bm+HE
vzH9AwQ9ui0B0UTVeu/aTDfheUfWaR7AqYbCoGP7dJ361vYthNby16oTPmMS3yCY
iz6nwGbcUL3D6JAr0CZi9CKwSjru3YQhf0h83mZE4ZeqjRavEvnXin4CHFcQArYX
DulJaO2VE70Qt2fNl1WSjtgEKTkYvwiC6GKOGMaeP61af7AhJtw3qh/vUgV5ntyL
vcmCryZzJxfZHmKl6m9iEPTv/u3yqb2x5ynib7Qd+rQWMjFHgzl2EbhQpDEGHx1c
tlyuTmn0ZrhXffDa/v+sc/rY4Wp/9rMY5gglgtYIWjTTEdGgU5iVLp/QmE5IokHK
bcaa7YxRKq73T14Zsn2P4UCWUtD2tBmq4v9CvBb6GODxed7eIJY7O6VWd2WR4RSt
NFU52vqsIaLaTh5YM8cc3P4PX1cYKkcTBUYPelqqug7o9SKOyTmBgr8fubIc3ovV
P+tQBmvHViqvgRVv050Ph+RtIlnHjf5eJZGgTIi94Fidsf59Ha82APC+iDJK3HWj
EbBtEl17nW72y3PdI+BUBpGcpbxXUjnO3nY+Iy2WQI2elX/7sd3Nrz04pVWO9qi8
MMix9iv7WKJztioGDcFY1boO7BrOVZKsqt+dgTy3K0W6kL6/fZXhbDokf2pUrCt9
6Wla6MG6tsivoSGxTJOXTjs6NF9RjdETEUJMWlwfCoZRbKBjlCbisIU9PIxxdtf1
hVLArcF4eyheHguim1RKNl4SxHs+6lrvU5Lk91Jm0baCjaJmtDIMeO3ObBnezujw
6Upx/cgaVlHJqXFvnkSSJMbq9yJnaol5i7GfF7Z3/wNGGbizFDsjEvPJ2bMds88Z
ij+n8ROVlmV/bSKY+l8iR+nvrlGyw3m9JwS9SpRVX2nXmLxybEVK+gpI8hAF7sZS
myG/L6AC8s3es/SHM4rHlil3FRAQE1Td8dVv4yj/nhIU7KLV3kmwwR7QOUPn3aHc
OQIWMzNOY7xHp3eTPcNpilrSfRdWhPzaJ1CEXbqrfwjZqfU6H2KboFF7WzHP4NkU
Dayrenhq4VpYqFcOAJn0xEQ5W4HMpLp3d8OodoLNv/7rHPWwqr6Tcitc1bQE4zH4
/daptmJdSyRNXWVebtG6GdBnZjvCQG8YgphVg67Hxa7izmiDjEerZ3AI5d0GESBY
r3KCrAA1MkaobvotLQMbZWFxiMIn9sPtYZ1Uv3IE8uqcxT3FIB7B8dLaU0aL6858
/FPq7hB+WEMi7P3kfkHzNo6MWIRNxt9v8yTJUPht8zgFMCmwkTcZGPHrEIDd1KnJ
4CFeCr8QRav79a1561ZQd9xaG2QjlNpxENnTL4g/onxbzB8EwyHBpGfWJ38lM/V8
ON9gSxUi/PkH0T/aseTDkidXzyDVn4klZ1grRHEVoGyYXYyWe3JM+UPTM1cd6YBc
uXzevUDrJygN6eNfZu6RyhYU4vU0OxbMqMLpESlGKCjL0UzFwM9NX81m7Lu6Bw1/
h/A/X8cQ1MgePHpQx9Acnew+lfJ6Kd0fPyWQaJs+7oOFB9gxLQOZRRIL/fOOR3Iq
X0GnHzRLdyzv53HFMUKMZX1el0IWqas7HKRU3zhOudYnjOiYyzQxWsGk6k7CuIqg
cymojZ6O2tjVLd314gPrNlV37IOuVgOHI4upftrujVRgzRl9y4+2v+hmehS/fyZ6
S/JkXWtPzbh697PY7I5pcAYo/oZRJtonnpQJ5BtFXEPQXHbzD0cOyZM4MVimGcEU
CQ/F9ALfRVXccu4LqcQPvA4hMN8hyx6erjgL8vLwvpq3mczYRdtWTI7MW0rHoSe0
TXM/Luc2tHUWXpLrcyCVp5eaR3MXeBe9ubYTAzHxK3yM7c+gzBTpFdhKmoPbKAwB
+VaQx0O8TYmKvYOchCl+AeExZ+VcTW9Psl691xd/roSW1skYYV3knGN0rBk2AeYP
44LGg+/9BalT5tYrEekkRnfAB6s7+oxtgu/Y+vGtHekxoUAtjeqxdm0EJ+2c5gJT
I02SY2XdnyvYfvmTKxBvLCVpbQaRDY62YVSkhUlqjevIpUHZpUt1l3ZBW9v9runz
7UwgkEjSRkvuTZXT8DtwOeKTXfVxs7DIbHZFmL4+Ds7lmngELo6tJM4ZTUcQDGiQ
ypGnaoL5pu3B2ojF4mVnTBqSiB6Un6ryIIr6QNaztfqxR74k0sm4KbqPqXT0Vkf2
mo0crCWtR9Z5jPnr+etg0CYeGdkyNywr5qRLGV2r01VkKuN6OudjLg/8vNl1i3Rv
mEgVPNmfb/LEnNUoM7pItIwiu/svbDiH5bJg97SL/hf55uoS93lwxWRbbd5CIqn3
0QTmHLXBCOkbtEeMN2Yvpgd/dauJqe+F5ZYqe3Rf7VXulKZ/nqLF0+3BEUINNY5t
jH/o0eajSmVf9gJ9k5+ImVy9IpGXYAQ7CITfbTNfXsT9yRd5WwgNVQnhgjO5Xlzz
hg2aMPMzXi/NYdDy9npAqsUaiVSpvnt2mzaDlVV5doRnZNidB5Wgo4x4VxwTIBD0
rR92wCe1IHufE3WuGGB21wgjxRrlCErfG8bOUyp1Frp1xID9IRuhgl/2JjBPkLzH
lDs0RlnnpT7banzwaD1WlOd/pbvQThywXN3BQ4cW/j+JltteqNhpoCGXxiZXfcLj
bP45ulSbjECf0LQrc8S5005R6fiY97Q9jGCUt2D1E/7LOgZkgSgQSCs0FtjGhX/g
QUzqA1iwf5zriT12k32ePPaIN/MtVsd4oFL9MMYx259xfxNXGJQvLZQiDrtiaKFZ
/zopdfrPeYnO71wENg5LpAFxfd0K0CKzqJMLo1/W2Xe0tTPsarsE8poCKgI57yub
hTwXcge5iqaJ4liN0legwhm/bLhMwomehAecexgRZ48HWQ5mCd0HZeo7oOZzw4BW
rp/fcf6jhtv6Q7nkxvG/2bPFzBfeZ5kbwmxOnKAVX5H3Y/JWY2uMlTiuzQMydM8J
2mrqLIRVB5g+BhaA2gnSmICfTBsc+e5LPz/+td2QCiF9yqdl8PqF0bouFjT8jaV6
dNkG8z/xi8IWiz0f1kp1P6bhddIaAu7AxcC/5iYqOsZEbd5qqkdSpwHODGsMpf/k
lkUD5+1kJgvPwkiYox++Cf+OsYK1EylcsaRkX4LPb6jWpWemEvw6hJVt68J2ng2v
HVOkQWwfoybxVvVj5IGLW+boAnvxAmQxkwtpBtmIYb8Jm4er8vMoVEuCDSHgddIu
uYb8qHj8AlJi0hVa6JLyX/UXBXDQOd7x3Xjg36JMzBV3LDZo6tEK1Hk0fQrgVUcw
VucIcp7j4fonxq0pd9dCm0x10E7h9j+AZAHOzJ09r5iIpmmfZppKRAbRAEZgZYyW
7AO/+6iTRUGVm+Jh+WL0eTSqlHGpBta5ik8w8MPTvvkk+yaKEP6WvDdbTU4PP5nr
nqoPHuQi9LF1ib8VFisaD4JjXMty0oBzaTkc+UttAuoKZs9mPONVWCXPCzaywBu/
M0AvB15wzjydiraAXTDlduyJOhkxzP5TZgj65oInPdjdE42mb3sHvYGeblT3WwUW
5pFoGsOPUh+YTwhR8aVKXCBJJfIaZTdv6ewMwXZ97BqJ/UuiQ+rgv7KgdEi5m0Jm
B8/dqWz7RkIRDTeMKxoZGseehzadKIBKBELM0n69LMdOp9vx2IECWyghLp/XtdqY
lfYGFITgdZAU/3PgKI+nzmViUmnKFwMHBsSVxgwddiaSKoGAicpXdjPaYgxm8d0l
XtUIRryhZ2mahoP36XUcAobSCDuFFpk/svpPRSdNObHsjzpbsrvnXfRynzPdZbHL
j5PD2mYUEUHgZc5pgXJE4r3lFGDJmxtL+RdzDhK/t9UB87mxFornm7Sska/PWHFy
gkVNl4fzgQeJp5xHnRWJdP2wLgJ6fR+o/wxP2Rx6A2uZj/fiYa7dJspUBO2oEtgN
HKsNowg1I+bkFuOYZrRud8vEGfL24BsSyKRXdcmtPsT/9IUa/RYIx8tseqT74nVT
3Pv53+YkFX7X24FOpfiXJOzcqEeSg6V4ikg0TJaOLt8PTUasOlaWZsHUufUriL2J
gZEiXu07hyproDP5WRZnSSGYI8HEjIOn3Mv8qs1SoCY0mK3Av7DZvofWUDFpf6Sy
YjUx/IFzai1yikkBYgDpdflsesbKRzgbkEavI1YGf/fSy8P9ksY11TGXBVAIAVsY
9IQtH+cbRb1MQYXEkaE0FmLMXVtNfvBNvnmUA6pXk4hTbfrP9ql+3hCggjE1cLmJ
sOYY1BmSdd/s/BEc8UGAdk444eP9E/IXIj6sIyOXWwqbI4y4RlnQ1jmb/NNbXKCg
VW0JnpvQhqk3LOFuSZOtfpA8Lp+MXY5jUZ7bp5ZU1lazRzVZgzUFLeP+bHtTtrMd
UF9ncRy9qbkZ404OddpnXnDDOTFpR49h87LHXL1Srzr0SpOFvbBSNWzs2UyR4gm8
YoIphqWKZSLYLseq0Jm3p1Xfy0c5vuGIuEJJCzV3giEFgiF7kDXcWqu+JwHrlzYU
FCug+G489Sp5gjNCSYc+Kuuop5b6A9S59ANQ0udAzlUNgcaiT5WQ4+JOnOXqWxtZ
JkHCClZqKgQVULa8/HLGZHhPXcB2oSh9D4rQ/8nSEGkRyt1z0XEkfjw13RJ/NfO4
i2FGR88yoGp8yC4Ozy8/eVrHAI9e8Wzk2YTTChwM2+tE0y05QHE8gwouaa/iaRF2
fnNEJ5nh1jYm226SGk2+jv6kmI7H+9R6qTeyxU1mx3cUD4xOB6gKLYIJ8MWbf6Ia
YyDpphloNgB1M6ShA4ITwmHVeqyA6MAf6BpljqAP9QbX5617ODc5eFC/2+KWzRpm
esY5oprG0Vuf9ohMO739Xk4tGJp7NvvIc8I67xv5KCS03k8IWKY4nOe+xfPBC/g2
nhP8xBfKeiJR12gEeudJrB8i640Z/g89vS7ELcxJa9G83rV3157od/5hRR1KjopW
gN30ye++bkikxix7hO1JBufCMU6ZvN7Eu3UORbzQnWSDuF1iOkCCzatBBBBkr2m9
34ookJdAnUivfY84jJXvWgiwKl0fr83GL/KNB6r7WNDrR3sjI0qjR/cCFUikj32G
CstrJTqCakPvupoV286E1+81Pt5hkdTDTsEXns9Z1PdDggebrpcU53HOGoJOwEsu
tOLjqDwd50K31+DdTMJJZdRB64FcGOuJqZHKPg5frXyR0tFJrD1burlKtvLmJAe9
yKmVQZwp+lr2Uzfrv2nRpQ0Ff8jXsO3j0NlLTrA6lGOOvxt5DRuzqURPBlZU31Hc
EFhrmtj/EvKBcALnFSjfjtDr3N2a0CfUVfP66uPMaD7RWtfntauoVPGRrNl/R1Qi
Asda4yNskbrdwmRJUfH7SM212ZZHLQAfdc6/E+EEW+7sX6bTRhAR23TRE2DgWyj9
pevuIMi4Yt/mpTDAOtXhkU/COEzYLVXQtTpjqR9X/cmcTwiBhbynX8tN5HczwPqX
3+1dw6fTaQoOqEG+4klOPnNV0Bx1L/aFHL9rQ88vRwIglByyNE/xL4KBYbmuGMFK
RVyTU8JkfAPqFPu391z1ZD84aksV2OvfzY+ZuKf7Avk5tzuriOwJNQDB1QzKM1iY
cyeESYQiiLsR8BMoXV2O33U3kbRV+qsSpkUu4A7Ig82EWZ9D1iRzVqXFUpbHyYWL
usr8rGJa5TVAghZRHet4TyLWO+8gbAKnEm+zqpax8xzUEpwGocknCC5HQauzIVJZ
MV6TB3whGB+nLs2Z5GBF/VcRac177m134yy1KGnbZLF10VncCYOvEVWa2Q1AuSr2
zB0eYAgKaqcNYIrPQB1BCwIp2rpWHDhU64ba8rVoM1+1s1FpTyWbp0awAdLDoi+U
f5s1+oDdE4BpE79+1xjU+EHJFG3ECDFDtfajKhXuk9OH5Q6CF0aacIm4U/WQbmFb
4shG64tWmYjDs4xaBuXAqS99InKLVksdf0KwtBBM3d7Mlt9cBiLxApwfOtpNZq77
jz/8PgmKUQZ0uBC1sc9CMVvun4bMBVekK3gKlCLqsIujRkub0DB/o+7xt1+huBCJ
kULpXNCfKnTMmwtjoXFnd8fhXXf9WvIkbVSHxQOX4M9QqmTcODmELkBqN3i+DvUd
RwJUkqq6gcnAKECgi/p0r+qyZZkAgsMuBhLMbG3TS4lviP6BzFSttxK7ztCzYJt8
UDiy0Ebt7wC6snZ6tE/9EbtKfZSjsFikmv1O6oimACKNDywV5OxKbdHA0+RvVsh+
+Kjco7Qimpbe9eD+DCfIOYY04qhB8OsopILzko9zJnjhUfEdVk9UWBBlCYKgL5aT
2dmVYji56d89vmOv8i5nuqaBGrt70hjJ/NfruzBBwiH8G7TA9hx2HG4o+4zClY3a
G58F9JrUhY6SL/vNdw8/gSN0LnzQoYYaOBtPHwvn21wVwk3EcCmJkEb3a8tPlB1V
Kuf3veEI/dN3d7kNqQd9eBoscKwnW8S3dyBDm7szliGNz8Gw9laTSjYp/X0gGp4x
7JEzBPxJspDLdOm3oVmhZirXKKKbHpOMXCawgiB3J7+Lp06K0JQVWcIvrxmEFFJv
Zw8JtjRMw9XUSFgGbHpTJVFIINzn2v2/ubK0hFp58QRvSLZcTwkz8M5/xIe+6f3K
Y5uLP+2NKu2l37bRgZaBDvJkXNMSBD6hDJhZpVHQ9WF6TI4iW9ut4UtK71OSHTV+
9kZ0mgYvxlPXvhLPjJVjSn9GooHTE9bmJHxR0FdFgnXIzb58aBhjRyJRAi2oSdFy
C+ld/mn5aBnND/NyIAtJaQ/g9buZoj/toq2FW9YiVfYUqbSms6Gj2T4PcMg6vk0b
u5taxGrrnCaPBRPRQfgoY0w8QAHSIvx+r+1Ap1gjeXXswMrHN9CIPlFiFypS350d
jsjmv+GmlutcaUKOL7bv2rLlDB9Sc2EOjYdAWquOF6fiGjGNipLu4Ida/s/lrsRG
C8KekfobOKv7rtL6xQ0xTrHLY4uQf6sYah2p63tQZa3/isfn2GwtSr4f+15LYFTv
CcUAijRMPjsT33Ih6EcFB9/X+dBPyF4dJRfCXwOxFDal1NuEc+YsGf/ZVSjw47Lm
q+01Sta3S/Y9HfBOHcKvVtv+ufaBZ2zavNVSuRVidh4ggjmi/ARCgvJl+FHAA2IN
VG1qcRmywdGNn7PT39eUG1K8XM8VQoZ4hgnelhfmT4wbxlzacsei1Xp0PXZTQed0
dDv7wd5ZTJ26CAsnZcej7Wo5++IL19n6fRC8iNkrepcToH+LlkcBw2vZIsfGrM3t
02ZDv6HX68FKSafhIJ4FJsqHH+gWhEPAxI6NxNQYs0g4BNwA6YmQAow20OMWhCH4
lUsKCD6llgcCLPBDBtosWBs6CkEjuIgGWs/JCDi8WRhbmM+vrbVlIwCVeva2E3kd
WycGTm2OrJdQo32cpZvJ5F4KkpyS0lzZsb9vOhkcTiTAMbNuXpVYHuv1tBwQ803I
E+qUGJ0bwt//3qeZjmdb7CzpY0KBNViqe3kCgGRUB1CGPnadLOq1eswxo7H7IDkX
vC7C6ondQT2pyGteBTBfw++mh7IiPX3LWg7CsL6AC6qBSpVtaEHGqsIE29W1+0Lc
qeUz/AalKV0Zx2vUc8TwJ8YNaADgnSk8UHJrojGtGjXkMa4NwkjseJv6R/i91a71
xPhNBoXk0+mscLA3+cEbX9bRxeEyHxAcFH6Wp79jXxYord1Yu/jm/BCn6m3VN1LE
MPvQpWAJSf/K9juzjLMhjpGsTC5kZ7fvtb9Z5RP2Qp6GXW/RmIlPMWWQ3EE25aiz
XIyAEU3jOSYTNqsb5PlLPsY5mGEll81OqO/kJiC7lkBxLWxc6fMN5ZcJpWwNoN4P
FGFqGPlzwwaITjiz5qTPnwy1RQAEJtDBYEC4onj7M9uL+iBjRfo1Vd6UkOCrjjJq
SNn9bdM8jPmq6L4GzvVvMgqq2ifoH9oa3aU+C6Yfiq97BHGRCv3BcE93pV+Kl5Oy
p0k3MJ/S5JU3vrOJwcQjo1Km3+xJrUWnQZqFszfBG9XuXST3sA4muYKIFlwFOPGw
KDK2VKfHz7HPHxX22H7s/DpMBtE4H+JiYxcqTI2xqSNn4woNTRygqp3SvFAyNPgR
LVbYZrBISSwD/OJVUptHnVrEW9Emsrmg5U9cd86ll89uMG3YzziCUS0L1hYtZjx9
jOWW4fEJk9a/xqscuJ1yaAtGiAsBg9E5sN/lyJ4QdQXamhzKCBtCbHAtxP6k2739
KKs2Igk167dXn3v1UbkbmAUuHLa9mhMe3wenXxD72zk2JTY2GvnoAwTzZ/MGY+NO
aoovfjXkFYmmHJY83foNTYpWWL+EAtXmRagOGA6aQ3eVjvy3b5LJ5fIQKeTd6+Uv
rw5g5Z6YAjuzZHpXxH173VDF6nQGVWV/wb+BGePb6oFutkESWBBVmMg8TGETKyJF
736ZqXcBxTwPZYJwwIzBRK07XLAfmOYFVFyvNF6lye5F1Xvr76jL1/Po0Wn/kGUr
QmgWLQM3EZv9yyBOI/fnOFdC1iSYyOvddKeomulH4K2ERRT40SmaV/yjrgt7x0AJ
vrtUACdLQrlghptTFZ/U2iFBQmySNGTYBVwuDf6re/CxI95obj71LRt9SDEkob8D
REULvV0Sj7vNcJa0bSLcZbZU4qvpsEeE0K1VkViNFTWZfqRplJBLxTZ5WCfuMaZj
m6VJSrKUvl3qlw2WfC8AyJryi+TwV9N+kSCWV4z/uyZJbWNfWBdBVa6Lw/ZpH6eR
7GbKyUMY/kFaG+GSNL5uyYgYNVDQqWH6j2JK1m0VXBn3OVCUeSRoVhmzK9Q2GLJs
TtpeH7QJwUav2u508tJas939vAy3o2vBEd0+ilNIq+Bn9sAfjQ2n3u3tI0kbeLKt
8GUNfiCqxcsibUR3WXr7jb9LIjqy1CGk2tJ/m18GjHFFouRAXmkf/DVxi3Aee7or
bRKnAqR28T6hBqodHe+xXvfLfO0B8DK7Ov0joc1sknR+qkq08p6Gb04jdKJ3Qiu9
2b8auGtivXVi7/jGpd4jRvjY3q7IaD4wlmOEcagHX1UdX0ogEm9+lwcxXjvTP8OP
BThoi1nYAYovhcQvIJSZjnkKy03CT9mmbry4ZxF50OjuUVPENuVhdXwBVoyZFyXb
OLnZLQVImi9LjRIe2SGJa0EJ77vPNxXOj5kyzriEZ/yjBCzlFkyKgAbGM7aMf1tb
FhW1TkZgR0qjs6mHmE+Mob6s5kkU5/x3Sr06F1VHf0kzraaG0azBNrjJvH9Wm23s
qhg+aTM7ZuQZ/DS6SlkdCFwWrMtz7XYlZt8DgEUV1snpAJxNltj7jORoxcToSfQJ
AHV9ltFrohIz7yiEND2ohYTCZLCL9AwXPHGKdwPB9ZREzFACoC9R3lbR6JJINiOk
20D5sauGuoJ9eLjIpQ2pVsQAYP/sL9T34O/Q2CXdne5keaHNQiwAwjilPyaIFX7v
hmCyCbGLSSQILzDGEx4f+JfzXFn8hCbf1PNYMYFqrFZ0oZLrghh2s0Fw4BACt2xQ
JgsY6xz4J90ONf8+2qhouYH8LGPLM7EnF6vLY1lP5frTRboU/NGfmsn8uRIZ5YSk
MXMcWVMhoR0DhLtiWUcR6OZmxH0X578aLWD+sjs03C+ewgqmGSet5ULuMYBBuBfT
MAqIKvfadgUII0/qwSBN9xjvIHPqiP3RE21f1u4i61lpprgXzjOYESREa7AhFleJ
mu91AhNdNAD8cXTReEWWO0TNvRmyI4zeYuRhCtKt9sm1exCd9d2wzQjoLI2tPFNl
eaxMFsq3+0Y4w1By3oOgagztqLLQUU0w5wz1NT5NyapCq1OpYRSww5Z2bFbKTrQa
1wcK94Nuc6BJtl2Rw4jE9/CuE4jAkr4TGSZmClGwEoqjiWf53RVkQpiLfaF4dj8w
O65ZY/6KS4JrID+SOM8FGrW2cU33vSdAFa9kAEaxaKxkQkqIR8l/2wCTrQhiASbs
yuUbQJX6CXA/C87pMLSZ7xf/ne3zMTOEMPjpLo/KVTo6R7Q3vOLhXrMSFHLy6LTC
KjDRbIwaAPrcQ20XgHmKk4O77DuMt8scXgY5TGxzoKMXCToUGzQNloQmXkuk7nYh
zDzNIBooeCIDXoiQl9tleRFJOCVC+gxRJVNqUzvjzRzfx1/Ko4N5/FyfrVcJxdbj
rm+mo0t9TbGTMz98peA8/lJLiLd65xp5pN10UyDCzqbfPNSZ/7Y6YbdscJ5Hdr8p
VO9bPAO454e4fphwsSUM1mcHBvqSu/O8GI9HkwWXccC6gmM/Pr9iTpz4Ojxclefo
0mJFBA4Td0/OTFWeghUFg9hF3kBch5Cd2aZNQgODHsDFipvrIba/+P6WoOCde4gt
S1x9gj+rz65aRC96IhohZNibcYO5K6tIMcKqGkQAIsYKwN+XNgWSdlT7wf+YLZbr
eFZNhZ8mXIZqXS3xMPVxhEMSjoot/XqaQEDELq5ez9NSn+9UTrKzVLvmjQakJSSM
6OqL4wA4T3fnHFF5f+3iSUZzBI39ousbzyWY+2ONARbXWd+fxLM/C//fa8Cpwqq4
f3hWUbG3jMGat36CKVMospuUL5nwEx9pUeu32q6e5dv07MnvKd+06zA6CyT0Jal/
vnNKC2hTnXjYY2NGhNxrLR4Rf7jvXdNzvkVbfSrujRdw3Ftmv7LJz2bcM25FcuOS
7zBgoU2B9bPm9HZV+MmbNWAy5WxZzBi3G3BuS+MuTLaJEthO8LU+qaBqJAGkbjUN
dM1+pnwrKE/4fojfd8UQJ6FAESK+++xd0WR1GBxDulSQB8pzooJFuRPeCrsXxXXa
jvS+QvjremQp5esKOUMc1uXwEiZpOZJNVbQFEytwfl5tQWAfHVbzNsL+ILG8s0lU
AcYoszkkohCI+cKPovz1j1B6oSr18cSLbm8uzSQQuaG+/jzBA20RRKS4kqPWaWOK
VJfJUbE9iY8UmCnEHw/QkoMF9zJZgJUd0rO7OV60QR4EzcciFx3sh8j+w1APThXC
6iQqSRgfWseAGm/DEpXcOXJHgrqLaPjaUbrADGs3+LGyuhJgl24V7LHsxb680tFz
HKUfSubJmPt4ntCUwHooc80c9DggfhZeWENaOyMz7/2wgVduVGpprUucbkdNYaPp
0Vk/Ecxpaaxn/jLipjwApws/3tVlxIwnz43NpMjTyKdi6cxbg6ChY4EtdmVSUDYI
Ejy5gz2O0XOL59upby19SNOwt8o4DUxPUftiKkI+i0nfo8BMCbxjwt2xBO+PpngN
MUpANOj7tCgx1ijaQ6SWVY72ULHrqPIIdlkN79NWAe0WYa671N2qH2ovsl4PKbRN
aN6K8o2ujBubyGWYTS4qRcEs0fNvZZmlGAD73fffGkqP/35/Ep0YnRf2GARyt4IQ
dE2DYPvP94t+UWGp4nxt38ibpcQtsmB9prxkRW4wrsbP05cjn2VMja8Q/ElB3AgD
BTgBFy/rpfW99TwcK32zv5HosQhgembGb6OydgvtXWRRlPn+s5GR/+2eOOeUWMnk
pxz5BSSCC6brUI9JRdEsdzpEW3DJs28NSN5QyoEP7oHjBdSVYemS+QdyCi2cmKOw
XPbxZcwzmYaYTHbpdAnCKKqf8qYi8YHW8mmm/f9DFQ1YBOMo/PVxLRMXjhq7Gu4m
so2EDbaIVCO5jzTCosH5MZp19J8NvQCT7/9PJdBnD3rIgWZnz1J2tjf0+kKAWsur
c5bR0hyaD0DDy+qCN7QHbQpfQSi9kclqoKgjFzk50/AvBeyS2s3XvDkR+/NTHseg
4J6oavIFCYMtU7iYOQwi+xCBCjzKZokwY/EGKsl0x7Psr6zlAXWw+jPh1jHjaNJA
DcuQPHAUUJEDQWwHOXWOD79pkps3c/sPnTdAW6c19w9nAQz9ypiYGYYDSXVtwzhp
naCce3wREkSzevIZB3wR3Ip/zhPq5tCvnAEmFh1Dp7QXH8J9vRAWfBcaiGYWUDL7
6u9MX0F78ZNXPQgIwpmZ+PUuhcZl2W49GPOTcQ2btK1ygeJ+1OcGSadRlRAUWFix
3xsT0UoVPd9mShclFgr+BdVW6wIOJ4AT3KfLncdBUKnRDWLCXJuO2fNUr2wALbP0
lqMbOLJEhSy6WYleZsVrBnWGpe1qXHH2wLTKj+R0YmzB+aST6YAXqhZi1vvrc8p4
qLluiOtxOg1pInQDrlYyW4xWo+Yur+40gYiVWAZte/1I6ytlxNyZ8nLfQDml76Qi
m+kw+fRve7gTiyrbMLZyaUQKqlcVokEgp+r0DO3mLdasnrP4O7boMUA65jva/arc
ZdKyknsfy+ycuV1Nm1nBMH+6n9ya7nb4XCxclQeSBnZaQ/FT0Z/I/onnL99cHv2u
0hTyjViu1ZdW4tN7TCCIh7IUPUM50uTPhjyrb0yUTbm6LjjYgRdG24S2m3n9vCH+
wVbo2k1tvJ1h7aNQWPYGTXQdTQfmOH4U7+0Vu0CI8f5AjJSyrtRHdoRZaz1x/WXU
Yh5PhFKdUqUiirn0tNfL8ArQ19bSj6Z8rcKZP1pkkEQoIoNPo2/eFJOJOXjkWIjM
+jOUVvWYeaOIOYnCyvvQ2+cS8OCcHBkH46dOMPdw4kU=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
LboqPFU1oN1l80K17NSI0NY24LpheDDQHx3txXJmc38ZpJJ9UhXgM0VylDRnPbLH
qyzQeXoIhhEG1P/LmS0KvC2szAN9wPkzTJMX9zDYm4t9jVkENPj+ajwHlnzSg+26
Yh/+waxhBRD0t+J7TEMRJTwShkYhUtwR0ZXEyNwjg4Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5328)
DBxuhg8lWE2u/RnXslAv69hQBRdaWhCUtpnk9e0RTG4hRxPQ/ox6zywJyCfa2PUM
3i5y/hrQjoUZSWLLFgq3m96Mi9pUPn8Kr/r2SRnfeDxLb3fHEtTRKZNJRK1la8l6
y4uLz4cPmxJC8ZBeNd3Fm7DaNbswU/2mgYjEI6cjPvBwrDCq7fXv6IvPWMo4xvX4
iR4Ep6uxnEb1aiSVy/ao06cBbFua8+jAOERtMBcMj5GjhllPMKvenUeD1DKUXnAt
zk0M6Y/Nr6Y/egUPruatIGVRdDX/51aNQb2DPPpK0yOlBWdadovFyjnnqPMYPw7P
OMZ2J7IsVv20Vt+Im/0vV9pWeK/NvtYbw/1cNPHhOwokSftwIdJp/LvFgFnMXi3h
N3r2slQ7oANM2YZjstTiLqimBopsE56f+v/c8i2gwu3nbS0P6Dhz++VoKFHGglFC
wHsqZA6F6+LJhNzjAaj4zr21FzQrvqd1z7kTXwFC62zEW+h+BCPS3uKm/NjZv6Ex
i6S0Ye/5gNkwXdSjKWoMdNUtZ+dZnkGBFtZt+N7ad/XTsuMXsaqfUaTV2f12jMG/
WsANHQiZ6g96cUfYbUP8nLsFA3rk2n+F8Ant9Jz2ooLl2tzFEizYaVkw8OeVXDKh
6htYM0B0k9u2w65KZIpsVR5ZApuEHJ5ivKhDydsmtsnj0DlhByLYTbgPtJX+CncP
1ZAMZKabMVdfs3xxci0XLmASTIf0XlWCEZSR6gGq2wRLhy4jIIjCAwNu4+JE4Qe3
Gaz9Jw6HGgbcBvwryed9ygdy33VtE8FZTLSBo0qhUfJmpr3SICMVzFmQH6Wp1sRU
OppFZpXejkM5M90OeNFLF0apAUkGuPex9dthC4EppBAbb1Gel5VDurqb32XDQftA
IDAjnYSVlvWac7xDhR2VSyCJLUgYKSnEVHHj5O2iasvE7whdrpRlvOr2lnjDSTrJ
mTjY+8lMFlaPeiU9u22jORLbDN3grqa4/uqHtTAgJsmlo7B84YDbv2Lf1kP2iPxd
SeFwE4T3HgS8XMy0qMFhbz9qlrQvuWHzGK/So3qRE5DsVI3ls2mWMDPJ94SGzh6s
RyqI7Zd2l3mlDjAtTA3uePzPRQq31QDtbW664rnsmCNh++eMkxtlPoFo/LtBK7wm
5B9gWcKCgH0m7LAsKutnJN8VxCypzw6lzOOoOB234Ed/kF00fXydCopD4hL0nkA9
Pl13eii1cN8w63HUwGRafRAnAUYoH1Z2ciTPI0H62Sfw+MwZLAeAIjAg7a8iYo3H
fgdDrEYMND/UKYDupeR4LOyLKUs/O2KxbupL4trT3MZtSMQjYDCN6SNH8GSEb6lV
hIPbv/UKgTKqUkX6DThNJUfNSu7rwrES//0gLtElWLCCniAvRX7RU8Is01iG5Xha
+vv44FTiL2I5Az8SLKM7ibHcyNenPMLe7Aaif+wNiZZXGGKapwo5c0VEmJCVR8Fm
9AdnkHP2i6Hvw7/Bb6HspbSChxozyPSD/ZJyfmX0oFTiSWcxWBTjfz09WSP7wtHJ
Nwyt5STO2gdP+uDWi3tsl6mFphl1DES1+jmCtbhxN31oxNEXS9kOkTuypy2sVKqh
cUyWSUdkfVDPSzLfVk5g4DZgL978QB7p+pIPcYHu9K35edA1DGq12fHEzVsqZ18X
5HUBy8Z5EEg/eXWOquB/RM4GcGBIwdWJ5IsPedBUiajXwCyO2VKi2ph6WtqrKJLs
SbUEgLZCFFAKgDQ4SECGIbTWc8mFwrenhh8TJ2xSsDwQP1cYRiekBhKxTMEYHHWv
CpPe9+8bSBgvH+e5w/6abnFIB4nslo8voUVVIkWkXMMxlvpH+Ar63eA6mJEOP5Ir
1cYXPm3XgdbnJJEqyVnW2i1CQUy9Z0XZjMfUz8U4HVm3RLaeQOb2aUDBp18CNX5u
rQgBZNZ7DLQDXxusaQ4bTu4Ch1aGDn0IrxwIaHcE9s41jpa52a6TVF+zI1KABYVf
cuU3OZ+zNQOjsYYAsdfk2QuFSBxKwxXDN5la9rdyA1coe2GHgDejwtdPext7YNZ9
WdGx9Wej2mOUEj4aJZGSjlXU5KmAZykCdkcSPAg31U/BxtKdVKrK87UcfejMD2hx
bGZBWQnn0lhWGvM4BIB4D2StlciJGXjFTwEiMHPaNOqCa3tnrMWo8qmO4TP1tLXN
hFBsC1NtgWaBaCm8uPu4TS1orYB2POg8Rp2J1BYs7lzkjFebHGH27lgTRsNgtBXd
pB9WlKbnD6xxB7fQwqHwVe/5gP+vz/nHcc7hPcv9Y2281O5041g+6Q5jLO8XlbFi
TOpeyWz4Gz5wMBXnhGUMv/6X6prfOp/ZvlNcP9o6xmzqDnJ8WN/lWMVJl3Ko6/O8
csDpp5X7eqlYd31VM3hVpTnEzey4KizeEc4tDEUdKM8sl9jf/fy+kN0WNJ//+HTX
0M6GlH3QgBJtPfklXZHUhU3hUWytHI1Y3/v5xMCPt04jDg5FlTPcFn5MMbJFYcUg
qDiXv+9QnkV2rxKVbK3ZpKbWu9yF6g7rE+kkyBHrTACWzbFCZD4a2N7w4ZwX3cq5
6Nn9G3GtXqihDGygMpedRwXLCuT4qKprMF7k7OMeAfCPI+jq8fOgxXAwDfSTUEHg
8iWkBLWJjyxBrM7YROtRc2GUpMLFIATcBlNkgcqlhzSDAmitCopHioqxLrpHRjD6
G9BF/uaiYHa7HxmkH922EH2vJjrDvsI5jh8dj42qqjLNHzRREqKgcawNfDwwEgnd
bfTL4BF3+wialeNib0QhbSa55yltEK01FPr4pOYgDV33vLPLQpUN2CA8UC7tHE24
r3VxpUGHsXTa8c3ByCeUh0I8OzdPCzdptu/E+0GuWE+4kXtjC6I9S9ghmihMvh+8
odaWVoDT87p5tMiH3RupXg0a9W89N7HKSuZcVsUGAGvpKTSrRfUcnfDPdxm2YDRP
OhZmeDu/di4o7brgWbzkYRAXuhL66YxdejIUf2OlB4CYUC4nAKUJLOEJ9gGU8uD5
DAweZ0+ls1rhGjRARdawUBdy3uETFXp9JuMsUDw2wwNcNgJj9zjQtYwDxSWWAYEb
TlDS2zcuydwL8/IX4GL5fRPpoo/IyM/K537CHXQc/QU576goLKALRSybzm7bySma
kNTsig9SQS5E2TxXN240SIE5HlaUlXmDT6L5drIyXB9zd2LX1nNa/IfQd/9g+m5R
3IhEJ76VhXItLehh0kLG4G1Z7Tr2xGLriiCzzgbGEpwik/Hg8L2l8+lLFDkr/yW8
VpY8dZ7Q5KGjEOAP1/AMaIgwdOl6nSgbrBM7AbH5JoS2i3vVrW1df/PmZ3F562pp
E5nCfifzXTL8tHQ2bfgDrbdxt38tWru1YV8p66uwIhDHfBJC585QL8XfA+eWuxOy
JkhgdMNYEtJcl43w3cfJwzpChhucGwpBGylBNW/tIgrcaHdTVH1xkyCfVEEiGIoQ
qDAdFCPSNQWzhlXGLgZnVyzQfBF+IhOpo2ibFiQ9kzDmOUjroteXEfPDYMuK/p63
WSGl2xrbjXHMVXLpip+7WknwS7NmcpMDghyiukKYQyhFlWcC3Nwa9q+7PsrwQf7b
utZA85TdK1xC15dQZJAsUQJwAkO7mxmGnHvl6qRD5grffHmXnKRtav1wCleM6PHQ
Lhc8+twKmxV534+OBxC9NXyA4TEN+zyCM1FJITpgL/llKex8efubKiztMlc0n79B
lqa072D6jjnhJilc8GmS8Jj6lja1xdVzzxNOjCrAuWHVOXGuVDDSA9eTZ8JaHqVi
WQ+ld6hfwO5XAkGXFQsyk0ZmysrBNffmwt2hJYWXBl43Nu3lWLuxYkMw68MIFTT3
IFh60YCTddL5cE1nJrgCh+oCRQwzAJX9W5X7pXYQElQNjhOHSZrHCZaLyX/ewGqC
s574dl2WG1moL2KwpQ3TAC/8TMxNxUhzqLLSKBGiIt2ldId1XOQ3WF8qDPUQy1gR
6gYDtnR4iR0aEHHCwtdzlPvTazoGp68fCnVOI5IHOLdfF/p/kxSkc2AmBcsYMR67
2KbyfezMqdFLAxSbxmriZOW9gnoM1zL2WQYVhYfVB7b5zAVwnLFlTi70pxgty7hl
81Fvxi9jfYy8tdUjcQMRONSiTZ8Z0zMcIwNx4qDE897hizvw0RFLjNlHEcvBXV2C
ymi4Z6CZ61eHdCB3ELhkREq0Tv9CRPxKKOUI9eTbYkNbXOA1jbO/4yO2T/M3mtvP
R5udTpD1G5l8NpAqtQcAh6qUTO9nrm564FLReO6GHKNeOili4UktiROntLcVYrTq
PIuhhdjB0y4qqZgRLxe2z1gXiqHUmRlEmnf91RdsYlPsxDdJDwqBNm3MvDgXz3xD
BUKFcsqFA46BUKVZlO0doEUs12M4Fz3DRazAk062u8zpsUy9FAURXs92BBKZEaPs
bnD76QjltKh1xA/1ff3wWl7DZcIHsmEDwyBv9+2oCwAVg1R9t7yVWCFk8p3jFx85
O62in2iakLE8JSj2tlwaaaUgw69l445OadfFzlfaN1rv1p2JO+FDbkXANu8Hxfss
2xiNlJl/i+m3dcxboalRoiKDrUI2irdNH9z9v+qTdrwDo1Arrnr4V56OZgpBnSlH
QceZheLnU0hVPOYo2y8aeDwdz6DF3gfNLSTuwM7IZLD2ycl+0cUzmpBwV8qrsbM9
/un34ly8PRPz3CaALrTUVRwmGP4ae8D7au8G5DkB2Khx2K2Gn8zMWvWyZqWMVxJ4
iv4rhLUIfsld8R8eq6hQNWcm5iZPio2gAX7090vCl9BTQhyUFUT5wlLDAXcsjO6I
8hn3noAABrNDVafcA6CtQEEfmygwOi4e4X0pxLlxkqt/j0i33F3YFUneKktyoxeP
MC4locUpB42x3FmqH1wlyfkGXGdMmHso4HturokACDvT6ZbJJZiKfD13pNDYbS9T
oSQbWwHyvTYl7qwuqKJEbf+C1Cv4u5SJLROdSEx2UF3ew17jkG730es60vAUqIGi
3y69lrk6ygXK6VLFtg/9qNJxDYBLlhqcNSNEKEE4p2hJ6o6ZNar145FbhQurGRLt
lwtkeIdDsAGrMk+dD9MIc2fvoH42YDAls6QpvYuRpyifNi5nJFuqTFp5FvDRBemc
IO9MyNPyeomWyGCCep8HvSnBGI6i/rssiPtylwLJeZP/9aBn5twxvkahn+YcMhXG
p/zZ+HWhQtb36B0COOa4JEwUp+Lb9ZRibCBeY94ld59l8fzmm/g2WQ6Ni+nUFdDm
wXZZpKBuLCcyDcIGWwI4vvI801fdmGWCFq9pSmbV16Anet/h13gKIo2Lffahvg+y
llWYM3V3LACb0uDIbM4+Tn778ikspz5+0Pd9oFA6U3jA5WmIaY0wCZ4TpXO/ZZOx
m00zQFgIExea7s4B3MLO4V0mDtODO1XJ7tG3fAQQ27rEQ2Ymt3VbfOFn0G7gFOIJ
PSDYr/nH6SMYM7MRf3c7t3retEczurHmTvYVNtOfQ8DAGx3+wO34AVXkKRx9yhiF
QK165Kh5Fq3iSwmeyD+M7fzyD45F6XnTdxN8lJaNkppEXLrgj2bOaVTL4urztavA
gShgx6rz1hR9Li6iKxGyEiPlxgDe5DQl3jOJr66feRF9RSe9CmwTPGmGsbi7C2O2
XFZDNx11139/MiAHkRrwgxJFJtgo8B9jyHiNhhf5OOHHQ9nEkNQLi09vBTRPP4+T
jmy0A+ZdfYntxDd3wlFW1pB0bB4k/BVqBuL8gAQ/9FvmZ5OogdaZuUOkQ5gX8+8q
yThY6w0VPGPkrvV3zuQf/pcpyze/xAYG98vcruI2PGk8EOn972PI5gEN+O6FNh52
b+53r+0tdG72lcrsMGBkFJ8RqY9daa07Z2mdJYB1klZ4TgvXA1BAPMfq6kuuJv+i
+Y7RKcbGHu/202NdNdUOT8HKdjauiW6jisZn1eYAyY1MHF2uKmpofR/EV/ZyroYU
e0mJNvNTosa4zm6HrP6nin5qrtjf4odH4NtSCN7Ykxz99lWOHUIvSda0ktqlYX0s
1l4Y+WKzWAHPAebEO9ZWubCdS9k/9lOe2++Naoa+rB9tkqV/LQTWahLJtCiluBgh
Aijfq0V9jBPM7H8jCXdjVLBO0rwfgf1PYOb3gTbsEpvlD6XXJ8HJx9acHc71lhrw
kdS7N1JesxlnH72DYB5lbBr71ZpHEtaUlR1sJA6v2bqZzxTihNqmmyR+fcB6+t6n
/JYntDOsUl/ILEq1VYUVsoSOYX5GiVKEkjozKTorB4o4/uWVydDfXf/3xp4rhy6d
ZF8v4p+4menfqJTclhBZmESlCFGr8lYUYmdYpsXTc3pvflNyfANRPKOKeNzuoZPQ
EgYKZ5wZ6ztJtGr9mjTSKW/GuR6qC3Jx9+bTxiYSfIyeGSiJVfpJERNn2ZhyXMh3
UjCc7ikhUgyg7uKCMt74jcr7iNv/qrIUZXwk+6pZ6y2yn6FDJ2fLLYdpdidW/eQd
KzGkuUkT1nQa7uDNvfCCrKlzfDe6SjXm0LgIyPZ2d5fWCi28HRF5M3HeoGxbnmn3
kv/cB/Nt1CU6TYgc4jIkGvNDzG2keffqVhlbH6RHrLcoh6cH/Jtfzpxhj0aM1M5M
cYIdu6JHppVsXHpq6CHT9808OtzL+aJ6SKJm0cnzVJMC9VcHdH9cG3i9mD5uum5C
4PKc1f+ekHBu729gC6bl+8hsFHMtpQhtoZLBcPPdX/CX+YLt5qGZ9vFjYvSV4vd1
4DMS7BW/jAOsT+fX9mq4E6EBkmXWDNqcbllrzVmUA8Vre32sNkjUiQf6zis7ut9d
CbW91KEuqr3HlWjKmshjutKcV0l++uajsTvEGT3rC46gEclFj+7/T0VaWG87mHr6
4puciqJEPT/7oiY0PTbr6ioG5GkQ08S3/tWuHqK+9U+Ve9WqY2DSd8/FHO9jt6i7
+byLEggGq1rWSSA6M20iVOcTn29D4wOILqyf/+ZufyLVhRtEnvJRvIiTQRvF/LHl
toSiJXFHpiP3tpGiiEJmW8d7lp6WeRSEWDq0NxiYGeMKAz3mZYMHqI3K8b9drwwi
L8eNoMw2zrZ66HEWVxyahBpnvB4Y7e248WrvneF5ujkdlK/ab46XavdFZb+BqJPk
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
TDFMEUhL+jZ4uSkDFdLvg01EdMFfNonUl6P8PLjkxXAuK2uNbAumS4YBIiKvbWHu
Hbs0bgWonnkgfNjduskOSp9YdXS0lLSuNh6Y5UDLCcdpJb78Cb3TV5twlcn1aDu2
RmEbqmIk21hFovIJySC6Ta+/qd7o4GTz3DYj4J7Sz3s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6336)
5e9YYwnbOFFZK1vgOYBOkXNhBTePcahhAqPKTTN3Vz/uTUn13LIivhmIsn2etzRY
UIizJkGnlfVtpmXTr+hFg/c1k2RdTWn07BTSgM79iNIv4HrnaHqgG7atTUmVxBj0
2Y6Hi8HMGkM4YEPnEpmwmudFxWQZ23xh8y6H4328wb2jV9g00JaP0UPncaRk3MaX
2D8++06dRV0QqY/x6ixut74N5UbPvrgk7IEsS2y/x8Z6JrNrmoskB77F0ciTT0F+
CASAkuUYsiGqZd7PgTVAA4cXwqZsc2loIVLiK+3jKuLOWSlcs7/WBd8DpsGR0InA
JZyMJPCxa2hKFY1pm7QmGsLy59M4uTuTXaam1+ZXd4r9w2CIlB8E1dtjgd39F8xx
Az8gYTUGuRlh6MsDZOjZdUNzw/+V2NV6DDxCIF65Hbz5JDFaQ7waV1kZSryvIewD
gdYH039NRHG6ToGj/xoK2Wp8fYCPcQsFRtjPTdA2ghxrI6vXapw2LkZU6bLIg6Sa
JPs8kT7ESli20md2+4YiU3yiDna4h0hZdt3xniOEL8TNASoASlJ0kTRq4Dm97HU0
r/MYMrwjkp7RPM6dkmmRCsv/BuIsGpZJLzvEx0ZyEmhej2ivszPK+x3oRen4lwwu
xM02U7Iwn3XYk1m8yMtJwcYCmm3vlD9+DsH77fTWRkzETe/HNTF58spnBZfqnodm
5jS+ta3R7cXaCsE8YbBYB36iVNqLcKL9bSiYQIXCGXpRP5cV3Cfh7luCwJIIhUHe
cH8jpSHZ0aGa/FmHkuSGlqQSuWZajzuATXYhVdAD4aHGYQW62QQPPctrn6VpngNV
vWrg/OLBirluNIs5B/H6tXvX79hEYIhleht9pC2nLvj36ab0axMoDXIGU5qVYnvL
OAPWS0BEMpJkZkui4SPSVuM/6Jewv/BI7taimEKeypLzokZAUBd5337XvaS03Ri0
FoSer6RC9BKrQYoWLTHD2ILGnhkJNDNPS8qO4F9TqARky2JWyxBWeAw4Pk2Ats43
GdTXvGJOYfLCX2MFiJh1nyA4SYd+an//RHEcRCRtCJanamtT+op2bKL0ZZGQoshp
ccXENUuyvTCDx4y6OPAl6yHMMDJUasam0gLZGHkyiDHD7nsu1zNcSUaKhLt/BqlD
PiabFJUqnbiFQDmg1DDV8ylfdP9klPT9mJPB8JO+xIV9Zo4KFBjvAB+49f+Yl1fh
l6yBrmw9TJ3zaZX7d3mBoZYM2a6j7j0Mxhd+sVxqkhVkfmH7QkvhWNoSM28wAwez
DdNPgi2R02UsT+38KQ9lfdRUiGDIFtMrh9gxt2XcSxop9EWIaDztwwB4EAylTpt4
HsQIb2raAJExQUD/2y6U0HoB3gs0LibZWC+2ncnHr3HkiiUhBhGOh9OyGXKW/2KN
ZDA4hssqehaeqw4zdWqMOB8QQT0kRRnYchtoI5qVMSLFrt0B0WiHvDD7e8akmQUq
dLUDOCaDRBr6x07VRYqBLj8fe3hwfLfNfuknHbxA/mTIHd0sJndL0HkGnh/w5Mqr
IWCR1XgoNR61/Re43LciztkINOEx2/aBXyXdVbBRFIfzNLsRcMo921GFpiUHR7xO
1jDk+hJNVUeX59bENaFp6L9x/dgbWFxdXdPq8+/pdUTso9spfM557rUvruWvYqtv
wU0FFRaMUSuVL5KtXnc8fo4+KqLI6VKTNsr0Gfl8lR0RhX+kqFJtjsY2BcZqwfKW
KbLk8RugLVwFl/ERsxfe7iDHaWx17J+CEg0aUhZGrC7MqyRpxV2zepWOlKDbs82a
5rRlYUyiObBbK9UK4MtZP7S9JV1JsusMIhxEHeLgnf9BuFYxMXrvXuJ+i1feUGq4
exk4Y1WrXqX59+a9geI1HH2QZWfR59QmwpRdLn9q/3HSVLtaHoxjR2oCso+dtY/F
CYgfN3/QKZoC6++C8YUcECW2w3QIzfoG7vaVSg7N9LyprmyfhpaknJ8opgSDqrt7
EFKlF58CLiQ5hVTq42SiGPJgt5gSpOxoZOqnPOaO9wj74MeK3KY6VJJJhBEwMzrf
+FV3FD8O+E5Px0ei3t/d947aaWmJ2i2Q8/RvIprlxQMzx69p0YhgcHZLc9dbPBYQ
w3f49pwmtqiaqNGUYrBS4n5UcWsOmYrsOTyeUZ6nJJjIGp6tF0NB7pS4fSpUCtRL
ibMdU/oF8PFUT5IqGeugxZI3hb8uYZfPyAIs3rTbwEdFaE0coA+sh+qHoMlfYp2U
omo/b70WTTj/BHjTlglcKzPJfnTkXAKmgcTksCjhhHmZNWUk7TSqkyqnIYoKi1mq
wubNgk3OboBCotxRXSLIbovwa2uHOwPmTacAIDn2aynOBrAOhBWGZPafm+1t3jU7
BIoWptw7WgkLu5eKfaPbkXK1nP+43cg6CV5+IouWKE7SP9Zx+OjPgEFh2EzepEIG
ERHl3sojV7rgtbnd2O15OBpGBXUOlBbR5RuBsexThiBXDz9mNh9RdGGMv0MVguMb
L49VinLFgVOJINjn8x5qR08q327Zs+hGWXe3hTXbro/JqD4J45RhPUDcn2MTRSQ5
wjohYqrXl/GlREQPNgvuyXl7NL23Bk8mhMYslrbrikrYAYBJdSR6+L4wInjd0648
PeFVEcP3pkO+63a68Yhc4bN/QKj+SxNUc9mTUf9uy2G4eXjZMiy2ApZGGSiD75nl
9wspyehd8iO8uaimleFULsQmnFwyD6SaqvQVQ4+OMvCjUCkWQs6xURFQgrO2QGeQ
pL9HBI9no44BJnBoxOCMxher4DtAYXFK7lv0CCe6hkuiz6ybEcbqLKIGv7d6IFqi
Ca/gHl9MQDIElvNsBVdhBFw6yVrYu8ughn2AhUbWqtaUlbl/+qIi5pLJp6UaW07Y
wnUn2MMEhhzsMa+0epFtgzbAvQ5C7AAcbMik26+3V4IHHsKQ8/bFMUlbhi3wqjct
7vgayYdqLEBRMBBi6FVi1b3oeiH4Y5m8QlAlsqfeQyB55296praX9NcuZMIFIn0C
uql3dhye2hvqZ59K9z6QXHXUqnnd0FqqTdn5rWKvg1dtY9CvjpVB8KIo0/l6ToEg
8BO055n3BJzydb8uvT6L4rO5LCKmyDx9y3MwldPdk6oc0rDZyUmicul66oD/YLYZ
UT+Ea5vIqznFcjcPONqLlJXhGxfrYQHwzRU94Uk54AdQPLaCzB6msAnlqSnkvvhp
jhe3d4II2ZQoufzfRTIwOW41aiC5PjAYSVkjLKr+RkWFf67NeogcEqGTJvwnFtzO
PWbyY697d5PizbAD1yf6FgjSBHbRNTFa0mxfWtGhANUBND4h+wuw3etOsVd8CZnp
U4BzcZPcKKYK5i++bu9jvXVPZ5xE+5CvjQMQsQgc9t0fLzTV8VcnFbJC1PntvxwS
3z96bz4Xz67ETIFXSsSvIg7wlsDgAi4U2majXhS6jwIIU17M8oe5tmCtLJSoVhFZ
I8FLwuDH1U6CeZwrlGTqWjbHdWAcVg6lZNcFHGTFoNbf2v+Tg1l+7Acu0ZkP+q0a
jKNQU4Rw8DZF0M9EE+OmC1t/8+PeYw4qmqoCM4QeitEvofucfxsZd+EX9RUva2hl
dS+I2sgS8gsdkoAh3PsMIOqHrbL7rCoY4uAtySPq5w+dfsJVvJlEFfjoUFpq73sT
YiOpCgIWvADDSz7duFdvYtToWmykatGE+FlljcCaysdwZf8cojIgodYfhjBXXyou
uQVsaFoGdlfDIIcjC0fI3xYMy5kepKGIf0QRezice7PlsEyXh3SE13zgamT92/aH
JAsHyIeoLGqJPHLqKjg70W8aYpSu6Q52c4g9WsVGrxE6ZvtK09oNHhvRjbcPhsY0
2ZeOg7Y/O9qyBM4PCnIrSpZE+M5dhOm/HiVRbkacx7ixEqiDWlEww6H2fmtR1t4P
rjG1XgoxZGTMJtwre+Gqe2AGbTI0+Pg4RgYN0puju8qSFFzP1OwPYZtSqUVtJRZO
XHLws46TyRcof7r/vr5oU13fvS298t91XAfExeMCMFZs2zSKwkMkJ4Pk9PRe1FLi
xEsLoxBlx8uy6T5XFm6mmIAcq/ZUOCpwOkNcAZn6AgkhiGjlMEEs8tOISABKOqnK
jApCawgi/Fewcx2z/v/akWbOQvWYTQ0PdwmLXVzBEdu1a+6mhe3UUNIrKmmiMgwM
Pnek/IW4vjyX9shkgKS1OqMMo6eY7RJDzRgZvmhvRPqMvZSTZQFakE9Q1rzh9d/r
gIRjchg103za0jsyltxOC8RwzVxesVtMvsR2jMFh2Epn4BFMc0G/nUsdEijW80sQ
JoG1wOUtmfSqhhQkp0NAw9gg4VjscfmWelVRIAMoKeV3FjjH02efSTt7KjIEyhea
05IY4zhWeT0DPcVhFONKcVfNXrTtbXy3wuYIBLHlTHADDe/WEjeShiYvDBR9gXBD
WCFI1HolZdB0glC9QxJKpBik209z6n95OnAblgHit+6RLCtDGC2iibimVdCmstqz
XKgtXicjq59KK+++oRgMI+dhyGFOGtnR/sZctjL7998lph+TofkDMyIT6Zi4GGJJ
lx5GZfd+rj5CJ8XRZ9x2BQVcLJtq0Sh1E/GnsCrQpi5HJzXjVX1eQhJKLlVmdF1J
iko0FasgxR8oPNoPofj6aBguWjBG3f1c3fzyWiVYpoHxmsRV0FPsFaj+AgaM/rhT
2nYnJLDhoT+PyiqAWWXJHgGk7AXOnRPeB6dy5n1hiTMENXij2CEkzxVsjG9/Besk
99d6tOJWi4CSFRcqoMcS8UpsmclyxKCFlz59lVFews7d1YqnrPmXhgUAgndHkfwG
XwKJxfjhXqgaFYlI9WPinJVSuDAqBBR+YXEwqPcemrA1ShdB6FB+Srs+lZQUUtwV
2LTPSz8rFiWwXcHTyLyNzLAQVVxk8tuPFMw/fTWFTMR1w51u41HY6r8I0kOBPrwo
PdsoXsOl5QiqgFtVeUJP1RbTK4GRqkW/Cd5zw317R3ReBJkMPypas81+hrM5FVpq
xof5J8g/JI9eFoWrwIaO4gfd6ghFwrLaP7hKG5ZgfB9xLNY0c8EZ+U8yXHFl7Y05
RA7mtnzF8Th5A2MlDxV5ijE7TNxB82b20ygx0Of37D9cmt3HPzqDH77YgkPfJH96
cc9I697EVruuBbZ58T+nvqlqkqyuvlTmUHVT0ggZKIzkc0Z8J9LkfX2XGTwzf1LN
fSePARGt8r30SAj1VyFZZrxswnoeaj0pE+enIvsvDSnIkTrqDN0xrl1TX4KD2WY5
b+uH1FUrWF71JaUdwZLbnrXlAk5EYFn3ngT9D5dRi7xfA8R/fY12ic/SogQRiXK4
0REnut4hxbKaMudnHSmRIGxenvwoecZn+YuoB8ZSVB2mgRO4YaLKAlPuQtn111HK
PtWlU54Up19tn2MslhHrujKLhKiVV+ZjDEzUYXF1AFAopASIR7kRfk5kWn8qQHFU
gg7gf+kXP4Qog7uAiefIwxDDIg0k6MA0j+MMccNibd6MaQxf48P+pNNi8bgfhhjc
RXyqfY9yRK4o+gRpy4mV3MSBzktiBHlCk/TosnNZCW95DI1abHr/hqTNDGvDhYKu
ofh74Fp7rb2DlgfXF2UW1Hr4yybaT9znrtkN/ovFD3oLMwI2jnDtKJdCZfirqUf3
+dYJzBenEzkDH9X/DMJRl02jpYmzR5U7yws4ZFVMKY2U7PpK1xibyFbkm5s8hsoo
sg5Mm5PnNROX1lTLDOkNsvGH9U6l+hMW2ZOxrxZjag7tZha83da2U+2ygB56Y0Dv
F3PCUzLIKc1pERrzm/2Q8YZkkvBXpJXXDiRkJyOnCMRLhrsSHgJXygedhGpyWJej
WjiQPpvVoNn/50q9/cQt3QPp4dxWbaIpvaff8VZ8BejpAw/+PoLwgkluOP3tZKoE
983P5NzKznEhLgiJzAj1avkjRgj/FcjYmlSYjAiYwdrat9IleX7nM1zFNQi0OWiy
ggtVJyV77JfnMGRLaiBzBHje6x3MryyzEJ7AbRxUBXc81hoqX0rtczAs18BtIMoR
s9ZzSiHOoG/MgvRcVMzXTMcZh2/pM5JAROmftMg6Nlz72RiCwnhQMITQhbzcOgnt
YKf3keVmkScbVKkOjgDP92ugysJ4JRITEAgRfHSUUH5A/5bKTeQgyOrq0fSydVg4
3Tf+rH1++NQ+Y3OqYbnpHDjgRJEbvgmKOB9SOgfOw8Y68GLQXea8pJWlC1s3o2qN
OalcKXolOPn/AVIXr/SRRwmpGxovhXmJJ5Q3o+xhmAPxfagAqfSUqRc5kvoUwyT/
/OELw2nz+R2HP4K5lo9qpmfHGGfZ8DSfs+GXTDkW462ufHR8fSBXutriDyXmWUjV
6OnUVySN3S0cY9NvWIFp/1Ebfq7yqfZlhqK/dUds6fdWIgnM/ViusDNycusVlh8+
psDr4oqFe3sBEc08gFK18PsmfnZPOb+w0+dqSrCBCHz92g9AJo19YVwqV+Rgslfx
NHPg9nF8TAMAvpM41ZfVIFPJuFqsuBSgR33acc04jNp5HUJ96GVX0EJdFENUZwuY
sFFY5ltsi6GnZkyX/Tn8Vaw6vNd4I9YbWb+S5A3htjd5Y9ZDAGDsCRwelwbm9PwJ
1+xANSWx4OCEdGiMzUzpYTAVNad4Gme6GGgiH04c3CMmT/Se1iQqFCAt560Oywgm
wC+G5OBFJN9j4krKVh2XScwJXdofZOKXNcqNmb7c1s306EzJExzukTGvko3HynY+
5T5g9uyMrt75n9Y3rFVWyhbGEDBPlcdFEkvXqMx56zChBYxaBVXZjQE+QXZfw9mc
JjdBJ5ZStDxbctNv9TtZm35jIsV6SFvr/2CAh7Y4+izv2RscKpv7EAqSsoqMhQnU
88z7qiMfaAPkunnjMgEnaCB2gMFZoMJ/sLDIVukJk6/6UpOacUYQOIdLD5cDE4aV
1bvXlAahk3U7kGbqEPghJdO6WbCfkAg1KlHO798wNpyyiLWHSUu7vxrBppEblXaf
1BTV6C//9vpwmjhSD6wE+ybk3+wu5s32JxeKSSoke1Aqcwb9xDry+t1h8r8/zAPX
5pCG5vOZIRKAdx+KzX2BNQm+7zp5jgk3xJTmKN/qz2C9+8XyWj1u1zujXC7S831a
O9Yx/fYK2XaYfvGo6duD0Kr931ICoBxH/oZWHjcUjc+ZzNWfsStgm/++s+KxTiZ0
c+wcM44sDerzevCJBCNQBRdPzewjXVZzsZ/auPa4KGngI6vsTrmfWYvQGZivvzdb
jp+YFJpwSM155aJyUR3ZmohU6GlsqO/4JsH6ym21JCP11be50/gvCOeUMAvd2oSd
ld6EUGRs9x8J00g6cmNA9vo0Tk0Z1EEUAhXvPX7KYF4hDNrcNWYUdQotQw/SPP9S
lorVjct2q+zL+BMdsehMvIOhO8/nLgKVmqf0l7Q9IiTa0W+l8clk+OFs6K+yHZX3
Notkwm4NDed1F6tjORvywqcqY6aQnU2f6VkZQLgUEYx87GEDqXgoR16GA8LFS16i
9BfBH/vO9mtwdqGCW+x2PecVZZ5myKXYz9BG8D25w/kEyEztGcJtCWSqOblVaSf7
FO/hPjz4RbFzIAMtmmDX1p45DXo99lgNjvYHTWhNOrYSb/sdxohF2Nt2hs2HN7Wd
vdqNH76NPBcteJxEyeiQK3KYOnNDxsKOcWlboaRZ/ifQ4j/GZItLwed/qWts4M2g
bFYhjBJk+NvKlyvP4lhMH+H5n2m8y4Xw2Z2YFXTPN8OdJ0hDFanGhxLZo2ew7X60
S30sAQq4yPnLwOsCFXM4O/Uroy1qfmX7aqIjZG7nWpcLEfd6n5iFbVacbStEfF5d
qrqRoB5O6wq2ciknnl8+CXTZASMaSi1A3UD2KIvyoIeJwoCgG4e9Ru0BAmdY14ao
/mbZqLBELp+g5/EO2RRXCwN/gXmxjN+WuYSpFX37iZzVnxFRZbQLP9CD219fFDW+
00ylnZ5yRdzSZZbPdCmVyNzxLUbboRzBhjlMQIqTMgEjudFBNm9TZCc2iJfUy/1Z
Pg9Cf9rOW5NGpEcbUxh1vt/ThUkFiMY3TBIB+lDFyH+xG8CZqNOK3s4X30qW5qwd
uneVDIlnWODZN4oQazk5HCKk+4PFjoEn/h+fyOHR5FOQ87xGccV2zIfxrk4qvItW
uzzAsuffhU/JKGFytqtZplzacsZkAGl427eozjYuoFhlqkDeGGt0kGbSv7HVV/q7
rgVdzLQIH0qQuzhQNLA+HjFxUyGEQqkEVKk+KVoAOrh6S/uDbRdB5fQ64ehsFOtq
p4A8MWPsjOzGfycrymPoArO5mYpn6bj9dDOeHf9u11z+sddyjrH5WV0aOgir/kJo
eSeP3dJwl3pFB7sPskI/SScHg4tddA0xi3M8UWMkg7CrjfQd+NGq6xLgwRdi0xaY
B6d2O9UXX2XjJ2t7b9dN/hUiVbjAFGhPhRd5CtdKtBlSthLnBFA7KU7BMfqK6L5M
`pragma protect end_protected

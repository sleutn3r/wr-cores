// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ku+sYVBRBWXStUX1i6oMEptPpdI8C+GIP0AnosGNo2mGEmomrq4Otjd7XVhNuUak
K2lHAzJbTkagQxRohyf3hGf0PEKJN5kGkuzqHnk1GZMaWjCdoFAsz/hDUASovYcG
seBnEJ1OTtm7hVKod3nf+5saBryK72N60W4eN4XPnN4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 27696)
+YfZpf5W5vwTFeguaqeNV8/JvILt0THUfh3p78oQ0Rmqg9xdK/KNBkr3b7SogGc/
gZOMui6iDsidk0SLx6umMvOWWqL2ldpgT5V35RYx4rAM3yxOIuDBcQeWJhJJQpt6
Fs3LNPA4/4Iv8NaYV1HEAc1uniLNiKXideHZHvfbNSIbLrXs3MkcG6/E77EQ1QQ7
90v6+enHlyud0R4y1A6PEWQG/yGaOmC656BZ22F7bTjkBw9oyWeKUyFgvas0aE/X
/r7Ng1VuNx9irUc4cK5H4z8RRKplmm7Rk23r0vQWB1ONX2Zsig3Eo2UNGwu+L2gi
RAsI3r67scOrJ1nDovPhEfiERt0AplyoLiQlHE/eEJ9Kla3/tVUWxBIufsvDTpKi
KlAgai8vSZS9KcQLtLs7q+QGsjAMqczU4nsFngzpPnFJfTQNUwfxv1UDUMxyeqOa
blECtt2Dfjln+BLswRKceVhAjTWZIFX8lR3Ii58At2LKJ4T2cDGhAEUBuvmZoQgQ
fAk7OQFGnT4n3wcSqzsPoLlz09o76r6GHim2RFKdzB/FeQnzxMLDwCyYk0IWfGYL
KA0MGQsS3rkIavbgEag0YDoRfMyb2Ew67+VxXtEV+gbR7EUIo4O5y2fNXLHWr1jp
FKTNy3873ESACobFap+hZu56YTHUtmEJOSXdVj9uWqkN86NlpZYr+OBVmYGiIJTt
8LYRdXvBR10Du6BwRISyT+N3c20B5cKlYVEgD6hhDwtHw1RnolcQrsl+dLLcNU5x
R8zmMI7xrM+QLBqPQAIFlf6rYj+oS9fSlSI8yvbmti3+zAHVL+aGwpDuxmjOm5Ch
aNTuQVGOqPNlgynI9bfv4We6XO2CF5qn/c+C4+5TYKf5Skai7lXCMhfaIw5rgbXM
hZIEr27vBXXzdsQsd2ChwhMiHUSFoqcAwRYd2Bmm4GUdRZj/uhJWY/EUTIWoxErJ
4fh+7E4yhIIZvbVY6DmyDz3b7P/5yQSEAn83MH5heswICmwIu4cI3vSgNE/yUjwj
LX0AHqkOJ/bFaVR8Hqe4aFaj8RfmO6f7fjD7oPnbM/l/XMzAmAJViGRXrHNKARh0
s3i1205tj4dCITftUk7PwX3/sUMPMflYNRV3HCXy6ROZm0+kWe/YDvxMxZyV83Tk
H7bn1baWQNPmmTf3WXqF2qVYLH95GyQyF+Q5Qh4lnJdd327q+SfuNdpTiCwGB4a6
MPVVi67/GBfvcYgODOYI2scTdXceb1a9ZSC9BfC1dRg8afr4Y1u4co51/QK9ldhx
UIwpGqsS/DDE5OUyBqqrCPnvUdF5ynXLh1ZFE4TOibSgt4bQl6klcd0F0gviewxl
VIZIsmb9vtq4Ho9pT7mR3IOK+YTjQeHzRmilGQwmEtlC9C7WIfuddoYXWkqIqILt
6R6idSX7W2LtgCKTusIpZ/f5CjvoH4bW87SMknC/OUiipn21iZjy19Kt24pdYB/n
0uI/w8l1/glkurxax3BT04msXC9GJdhq3VN/2Gh0OgoHHeAuEiTSW9d7PsPtXRua
G4ilo3K1o9Blhp7KN78nnybVT4k5FkPA4l9WufAdzAhCmsFWWT+PRexOUX0lsqqN
JKOz1h7DvfcOiiZsvhg3Z5wRLgoh0r9ORSbkDLh6nwJaJMaCnvQx25N8vF6ulDO/
yDmrnoOxfPFMMmVpL4M6GrhzUDMrQddDBC8+TXtlnNLWeLNT78U//vWvmJoTaqEH
3sgx8XhRfKGOT5nP7YbT3BeQz93MmnMaCf1kmbw0vf+BSeqIsP9l3XuzlabSfoxo
iu3oQ51TXJ+y7fdN4b1uwa+LHbe4d6LaYynTadcFgQBLo1zGKJ2PzkjAs9KFcSjU
aHf6z3HTsQDa8h7CLrrvHS2Zcm5ElGkYuv/rlbxU8eYs8Be0g1SKwuJYuwx4fmOp
87L6vfnITroweSgZyN2KvB1TYZXneZXgz0cBWK0OOBujyqJ44B0bloRnq9/q/2EM
WhOl9iAUkd4oM5wlVBpgZxeo3R9Xp6vTYfVU8txHwTuKu8QnJon2meIA59XGAYuo
EYu5kmNm2TdAF4mkdwn1XtWJZd9hB1j7iP4ch1gO4DIoAaKfk7mPwT0HNP/Urm9O
7KiW1A4huBJZwgi4n+HPiPvhNc8N+Sj4SphgS74GD1a5aKyoOYkhMFRs+VreAZBT
/eGZgEJnI9hgm+N/R0nehj9IycDgdtDV5/AyCI1mKOvmYUL++WUL61xIhuuyuhwC
3XSw2ZtFhyAefXFmBvoO0p8kW949MSDtvVJwqJt1MJYNyg1QOfLWRBD60j7sa9LU
Rau4lwoDWjka0CzED0meT585/RL3cdvGGtjc/Oygf6D+Lp5au32pE6rJop0VqaEz
bny0UvsLi1BEv8onH7F+wKR9BZXfGPi6m5cH3hF8RS/qc/d7Tvsidz1jOm6+AfHu
SwdDuMCX2Jxl8oHvI+0hyForz+L1RolvINNJhfYdxOcE/CJHmoQZ4KYnhcD9sfjH
jPays7aErAAT2y81RK+/iAQ5l70YJD7X/MAWlClV0kXtVm6/pel+H1nmrwQTt/WR
diKHM00H5FNogfpvBxO7nWCClLCZBUGjcysvTprn/ksPFOzryU2C7T7U2AfeagNu
NUePFbfvhx6x8ArQ/VQCsJLz/3MsISCAZod0HUzt1m/RfzZmzBlCj0GtyipsBdLL
Vf+OyPVonqVjQ2xnZAmr/sR4SnQJQDD30gDtSwK6xY7TtJwSbVMH7evZPbuXASCW
MCde/1NGVWKw/6bH5Gg8tD8IBF1zSCq4jSe8xu/1octkJJjEzKZJ8EM+Xrs7Eezn
S8oYAfNVWYvfoE/6enKkWN9taDU1AODRs3KeazYnD8jlzm6IcGA/aELa5BTk7Xsb
HJhUfYasOzfF5wehPJbDCt7Ke0qmp5itrWLqFb4WS2OICdfV5LziKJLsOPG6qqDK
na7SwrFaIhpxEiawQMZDdjs6RtKvtuN8kkdmgb+SEbQ0NoKx5r7LnM9Y9W1MFJQJ
gHEJT5jmiuM80lp1m1g5ZTc+bDOq3YvjrL6+j3I+x/JLj1JMN9ZrpbRzYUrGay7t
wgVa2jYUNVCAoIWzUjhZwE/gI1TKynmd5vVoXHPdXjgb2cxjQYQr0Q5kAAQkbx2b
wlGm1jqFiOAGOh/cwrXDNc/OSLo0ZoLEaGMBS0CoHDqTBvcpAxQDIxfKnMxbsw5X
jQzyI0FvUY/6Xa9TcFRMWbbfuAXGbsAa0+euJo50AlTcaEf9pq5u/AN1A6vKLwZE
jBnPw1S0E5371AsSGoWEJ921pZ6EEnKeoqLmbm4swCb3zso5r9aCnqDGMfsWTKhJ
ZzpWfJP+DkQve5+ie9isHGqKvUb7wkM6+kCFfq2U6q1ZJ2iUTaKjlxLF7Ia4OogF
efMcOWvd6Ffq8TfYeKStvHWfBPGadE4WIub27L9qSKh+5U8dG+2YXeRSXHeOdA1p
5RrNA9D0sVIQYArhkyWRiUrfToIO+QieVj2o+bOyXxU+kNJJR2XKv0eKXVTBOGov
3I1qc5qysg2RDw4mDPSEOfW5tYs74KUBzJfyvPVAnkgs/yRDS7waJGe480ozMqwV
1k23GMEL4W6jUBV2EYvVAr/d7E75znl1ZMBk4zJtoHpArEFOMjo/drfeL75JSmVh
S0g8wEzprkBk771bhTY2nd6Y/3lQzmaffANebhh5x3s5PpknTx5wtkC+EEipCe8N
+NwtrFfEgl9qfwjYCk+OKQFP2QGgB9/N5rPfMBrYrgIQwiqQO5OgbYE8LYnqvOBS
5jGKTllAHgAPtdEda/WS7mjfiSicjPM2+1JmQ9mFr1WUjuebOAAJdCeNFhmBUpHc
PpzavgHPh2OH5zIPelASxMeKq75yrzRO8sqZ9uwI1mTBq48V0IRzAzJ0oHjmKKRm
eG4CsE3fz49pUC0KO9iKXtBgyHrVyc7mzIaJKjWW9GFUxYf/819uNBv1nqlwii4Q
BMYlkac6ZsFJ8f+ejCAg2wVcrh5aR/sH5afOD8HCHeFBGGxok4vtzAMt0PX6dbhF
Z4LeKSvtKXEbAAxTZl6SHeRRLoJpUWn8GwA49ZhgQoRvUC7j6ddq4UPuI4eKYSdk
cL1J/e1UqVf4o0KPtL4dsMjHB8mueKTalHOARX/29r5HpdjWL4pDjybwAwm46Ae8
2TF14IhFJA6bVwZVGRo8Qsw2mYU116+nJiUdZYj8epzCyzeDV3Q21c7csNyiVjJC
G8CK6XxvTaxCT22r3UtMiiHOYrPTn7sH3nZkU31X+jcEwVvLRuVZr8yns7waqPDd
M+8xsQWFsTO9C3SsCDKGtC8ZGt8YQ5QEFZjvZlHaGP526TmH9pVYIEeTULyofgvz
qejh85QICn+gpcVeDfAQ6bZR0UCqWkHZztGiLS2TqyRTsFdPnggOJmjKPmCx8bBz
gYXa9lwlk47pCWYVXevoGEquZ3dq+jEwR4ZtD2w45ySs8Fe3gRhRDPS5kVImLnKR
+B2dUX1hSzb5ejjKmkTv8pY3JR5f3SZAad81/X1UzkbWxfCPpe4wuIa81A/Q2LSF
Q/J6EVL/wU0bg9C+vZV8IFd37XpkG+fIfXv+M4rZjwRo+YypKpvVwEM5Q3+5tJ1b
3V//zfCQhdHW1VSiRuEFuG4bQCZb6aKiVSBtAHjaVlbqXSJcXKFOeiD0OkHTswDw
6dggZux04AEslF6JqEgCLdmOjkp15ArasAitcQwHmMhiyeRvGc7VOJYtyxXUTmN/
c3lmo7wayq47RUOM9h66kYi6dtzcofrEeeEhx1vqGj0eUKgSrrJC0b79Okbdvudk
qcMpYfiIZXddSmpC9/RbqVgcQ7dtVpHfbk7LNKYGDg/encrimjTsLj4RrNL0xvXF
l9GCu9FueieHxg799XYDJ9Fxk9BGKZyuzDl476sh8HZMWE5eZog3jH7Nx39ikCU/
GmpWew63m9DvdJSnAwIsi7zPay9ZxJQaGT5PB0YaPNzYlLtXmoysP+eM1qq5gvB/
OC7oCC0oTT5/3FGHGw1HggHQFDiCN8hZfRWsYTwhyz5jM8xi4BU0EpziVLaFX925
l+bOhhcUgbVHyH8fTbZnaYXHOU1uTKTlS4fsu1nc2sVJToZ4ZjuB9h8GaMnBfctH
HHYraBNKfIR9uR8kVzUw5CWn6bCte/spEssaYXJqEEpP1DkzMQUgFf2hnu+u/cWX
VMI8Q0E8OnagbqU/Mkm7cAnQkCiM2w4SDqg9751hhqDjpqDaAIaveo4Fergd1CqV
dEGfHVoUdtxeXSu6T3A+IZ1AsL0azJ/LaEXd3pBTBqsOqrSCslfeeWFSvDKwfARp
iv3AeUDf47A//6xpgL1fwA8e2AKgP7NU6cCXOxjfhNhJk/uzCa9KiLWD5XxlCB5p
uuXK4CkCfyECc9zi/Gf2KY6XwdJDo14Yb4K55W8Eks5wLUUiKGFcWUk5qQ/iFM04
PDOnLCzAxTmLD57hz35AKRqqo/Od3ku03irIAVU/PE5KVwN5vPzixHFn251PLEQY
VE3L8E4HkbVxTHyvTOrFMJjVN0r+IbqQVG300ycVHyhlzrnmCseJCVA2U5j2Egmj
G+VM/bLPcC21OO+ycN7NQdglWh4KzUh/RYSlblTUTBpM0Vr1aow9Qrxxdq+dryLZ
Q+uuzHrWkgYIBM8qUUIs9BH3KiwWyJpO16rFA60I+BcISKrGG8cfUUao+6/ijBhV
g66xcRLRBi0IvkxFuvg3kKQJ5/2th9iB8AV6XHFxhHVlBI8SwY3CYD1xEjmLaEsa
8AvFCXcuOOt3Dqj3BVAAiv2ZI8AMbcUtCD4z+NcZUwtG72RivoHWhlbKcgrWnYSc
yKzeO+8PQkbquFEwzqToBQPz5czo4OgVdTSPtbepqJAeI3XqvIKk2LIqcehrxaZZ
4awlz0e8MdYWhego7sPbRjHYSzItiOilQkCSWdjgpI7fVIIwzpP16lHGvX7L2BM0
dwfqgo9BETPeo/SallwAnJgUvo7YB0k+L4TDLYcqmPomsxDJyxz7M45dvziRwgVN
efeeMqVA73RGWOOTkSauk2BPjoQ3Ud73EGTAHnVIKGKop74uQR1Ote8FJlIUihPg
NFqz9iFVg45tdeAyxTXbqLO3XEijyFhH4dDFvpFiWGNI/NvV5iOM/PlgOy9TivgM
YxoPpIHgAIPmefHpc6lkSW3xPewz8m0CWYk6mz3LZ7TkBrz0ywuMkfQdr0PWL6UI
qNaORELzxzRYh65NCIl7igJfet3qDFRZ4vpKnAowe3EIIW4mT3adQ3sk87VzpKTT
wh9jkpW7C/Oie5MuSAzeB6Cq8C5pCQ7gX1MfTe5V8CgZeWTCC+0sN/mvXZceW8hF
Vf3PKk1lYZuQdHnFujmC51v0HgeuucI2DFWQQD2V9UVR3/p9LsQrmT2RwaB2cimv
OunQOSMVmGHbgJWC63GQT9aBCbvb0UWJctB2C220rHtS1eXqyCfORFJgT8Ckqk4U
QYCfYCz5sKMDEKCthvsSOA1ZQY6m1kYnR1enNuAszoeoJY+Obpq+qhcjCHbk6Je6
4VjlpDY7f/ee37V2Lk1xJK8QZjPvC8wBZMNz29j0fkLctTi1E8zmtBeWXt1A2n7r
b/Mtm+KBGz8KfmAmkQoOGuHX8IdZjwCH1DgUXfhxgZ5QcmwSKLQK1uSxfB8p2nb0
zmNZm8Nwr8ruLN00Xi6z8BkjLtCVmYsyLMU05/7OGGZD1HJes1lpvsK4P9j3Ilf3
5Dnoyo+H0yZXNe/LdsjfnbfP4eWUl8vR1Dn1m5UgiZEnPW60toQWxpyrjJx2b5BU
0X6fzv7PxmgGE3ODyrYv1VHjGgkFzDsvPiBIlUE7WN8icrW/YpwCyMW9GOp6qOKu
k5+lC6harKydmv2m9a86QiXhG0rDfpGSrtqoyaRzXqjB5yci0AdhLI5RGOyQB83v
LALc4761xr6430REDtXlAVUNQuErO3ESFYJvsqW9ea6mk7fq2hTjzwvy0xcqMIhG
4YFpLUGAFlMjYQetpjvqKOOA3tbs0tXeQuH8q+YxTQwKblNAmarkvWhhTt0qv9k0
QsJHMANiocruLua+vl+M3+ViDPkB00WFSMJ+pd22/TGoFUHwsuM04YYzAk9jb5fl
hbj+Na/ilDsjkjtx6Y2U8SmmAo3Q/9mUJ4IN9dCQaM5J7cYL54iagl0zxs6zF4IC
alqpH22ddhsPIBXSh25dEs495iD2BoPiwIIi1Ykvea8qhT65nTeXg/18f4kMbXvF
OCCwrUwTn8soNL/SKR1EmFhIWWGBdsbMj8nMNI1wcefrW7xu4ll8EL3jdZqWz5z7
tgKXq4waeAvbnEKCyQrL2rEX4pdilnEgCwGxfwAn2uDgqlaiZILEyfpTPOuY7jO7
B68Rsvaerxj3vjtJ3wwkivahbZQDQ2YVtTeUvXtJ5U+STpf4QZ2AjvkfXClqpg+X
xIBD7s3DnotNLKTslwNaK53hXNPGSf6rM5xZHG/eIXaTwU0BObfP8Nsby/KejNeH
yPhKRfP+WYNVqYrDtmCxrDbgYpQBXi6HbFc4ySuNRLebSv0nLmKzjZrwqTi1odVC
OA0/Q5Ug+S+H55yFUQN0vOCKTU1WswhptEms0DDkRKDPzcThKwdIAE9ZwtR+Di+L
JOE3qVxRIpWhvm4dXUYnCm4pB49s8ioakTt+r1Yru4YvMV3rJVXaTMV0bvJunpVk
fr+FBDOrwuYlyk3L4zc52LdpqrQrUw26RqO3t7KYYdYxKueTpVxmgglQOExd5Fbs
4cdSLKWWciB5fAgD3dVOuMMd7O1jU7uuEWM090SM3qbBR1eYeEOuKhKShqsi+oXA
15+8jjSYJPww3KyuwkXd7kg/Y2ScTNRDLGHHGZDQ1Gy99+Y9SNdjeWCxyEfdlMI3
OzncIr1Os0V0pQv50pWN8HrrQK5GImAvEN8QLptlmwEIg3Qh3W+SWUynMrZmzyyb
WKeGZz6j9ldkOGMolsCV+jegeMpUUPekK49AhnNJZkeBDTbN8mCpuPuh0Esuxd0x
BkSDYyo4WWPYUty9yXGWVq55CW0kqZxM0z84MHVAVB+PxRkXvAuWzp0oncdADDC8
kksKoA4kDEOa6gbRU2o4t2APsizgoKLwwMtBlmNmPglakUq+8nR+675/kaYrkLGr
yqwV9iDopNiWA3NN7ZQgaokFEJKNiTTG1AcBVGzdF2H6EFE0X7qybKbVM3B4MAJo
48hPVmsWyjSWF6eEMwWwShkHllvrB69iM/yNV27JrLemdw7B+Z/AZbI1G6HJL1AT
cRd1zcSv2jpwO2SZd63F/FW6yodE2fWatsO+FYxryFFQD+60o3pRDLHpAR9aeyfz
L9EyjTZasEm6wS0+dH9ZPpuZMSncxZd/4WnwcFtPZiGP34hnI1cqAW2K62u8AKvC
BNeqcsfkueWezg96wXL6gxj+9ey8JQJxqRkns+gpJ/MjJQlZk1dAcW2TsY2+hVS9
OteFv0nKNjxl7SYS2CRl6uUgD3cgVnKwN1DdUWjkmtrGj/FZoCKo1KrgmRvTWqba
FMJRWj7YQa5enEDLXvf/CZpNQfpFon+M+QA2/Mtwbb5W67BfDo2HiC+omOriugp8
jmVN8QQlAecAa0K9sIaI4AA6YSbBAiwNosh8kdTZ0TVEntQHturiGP351YyDvbGW
uLWWpHJPmgyGvqyDe78sbYJ029QBEg5dTavn/Ua56nGsH5HQuA+JpSAAibwOPI3p
AR5l+dQDtr+GyAiMGpyqAdFkAh8Q2U9o0n0lQjs8egwybQwu+Qu4xMssmfoPXzMd
AqlFCZcdy8nM4MbcmkMjhFDoj3GfCqQ1jS4QQF4VMGYjNoviuBOpjzL4amya7RJ/
TMrahmI3ANdlYGm2xXn2EkYjjxC06n/Dxwg58kSC+tkEyiveZ8ekZ0A4Qx4/kMAr
74ulDb48jYK06rdr8Xfj5vh90TX7eD4/tH3BMki/ldZjWeWBygevm+zrVsPXnVFO
4LQTTjuaUli8RfAIzds/k+6sGpiH+uIiptfJj62faqjCzhrKqlFGBfx8+o+1HJZA
sWlXvZe7Mf+tHURPkAMCOZJvfREwnk6C8YcqUzf5KQ6akx01TdScZNqYy0KD0OGb
PE4UZxuRfxUldqfPKdOBfj3N6BKoJskMpwcKhtC2G4+Jsi6sHtFQM4iy3t1ScyLh
LKKvyUVXPnvvZ20/VYvceCW+caUV3cRKsyk0bHYBf95c1ioZAqsWdsa66QFxK3zL
/kWcd9ZRNMhtglb3GyDPhUZ2KNcgVxglykx6ukPvv9668ce6aQKZ3G66bG1FetJt
n/d1qaE8nVViFElT1ddhA+t6YlXhl4dynRvbFjQMLJZUubVvQgTUnQeyfATGW9Pq
Zt4fHZdsGwWfwyeR0jn5JuPj+ZHQFXZiwrvYFUYqE2sd+KaPazeop1Hb5sYCwZQI
+wdWQT39yr4ywfmELgSJASNXtsKDCzbJXECJpG+pMHss/MhYqoMQDwqS+TDyIvAc
u0g80rzT4VbGUjpW2CjzQE/AjvAjhF2/dSy3CUgTdXlYLvgbAlgnDZlUZ8l0XOOO
UJkEx7ge79P4Knjbz+etfrMX3IzzUOhHqNN6pHsE1I4vPoszjXbLrn1j9WUnqHwd
PWQ8VRKJXnoU0vVRHeaUIsTVjU/3pwFeCMrnZ5Go1sOmvuq+18+25oWEcLd+Kitm
CZjeTmWYjAkCcXerexyI4e9YJjZrn4oBlaxWELN5kOLF/ox6xb0cvkDJLt9BxftP
lCQZmZr5jKVjllobGrXwLCJCUTjijEuI5pm/LmaggXobuzlGNgISUZMVG/ygUbkZ
tvwDP6uBWOLdr7GPpliM5bhgY/zpyUiKV8lthVeeJ76HTW892jeDFWEYO7VPuYF1
VXWx6SGrHQZpkDPlATZZesoRdJ6A4JQAMRK196zqLtgAorHBK9TvtnWFJWy7l66D
0MxJ6PhlrN0tOOZypwIf5jCE11eWwVWXmpZcTsVS+RMiYqTxDYehK1j+cnzOpWPG
WUdu2dLF9U4cL59SLgor3Pdb74/oJhYVN7C3fU9YN2qngFr2YiJbJvq2uQLw6hXX
hwQMiyOMAzasu+2xFd69atZZji9MHVuZ73kN0aWFPW5BhRP0QM5N6WDyARgBR5Qa
mwKU0fS9+5U1no1QuoExCA3s8yFiF8iTpuFvGN2ajqteU0jFdQuyFIsIekACyhDK
FMrCzHzQ02JyzS3sQ2b62NUnxjfAkBRvz3QOFNjXdEcexGmuQhPXDPAMscTBGGhY
pMOlRAtKIJGNFyYh5aDY8QUrQHiDpC2Pko4LGNzJMJW6s4PIEZ8qOsaN2AumCdd+
YNF/acj0vr01hrgI1VOiCA5Eos7sJs5L3ZPLkEXEdHkTkesKaMwIUJcmqPjT0GtV
5Lpi2rhT5TNHlOUkNTWk54xr9pg3A74sLkz36i6To2iMaO+0iFW+vIJGQXBT+POq
+k+kJXofRWpYmPlSmynrDh7DPuwrcjMTToq30MiqsHk2LDajlj4HQFWJYoYoRKXX
gJzWGxvbXb8NwWwALL8CQi16MUHzVdswR9fWkisv3SrL1ytKYYsX/3qNZvjXH5gb
DgYScR6mldpgm/MvuE8jgXYxgb1ACwnWcEqaOO6lHjSxp8fzXBbihQWMPsl+Hrz9
r//ONj1UWIAN2efjDbQBJ98gzUrmhFUVsrQs1Tc3BapERjlT7HHgVdU43OjbsAmE
OdzZYs41B8JexZTLz8Ei2ERc9Ig4Ofi0mcd89QHi7iKePUo2sVOKmlEkSW0ZK6+G
nDCLV1e/MOSKEYyqZdPq8OPwiyfwim49ARzZGBvfTeQB6dU2iUmq4GRRmLSFa7E+
Tsscc0yc1XO4SDhLyAlD4gJbQsLdXuH9YQFNnRPP0Q4kWOU1XNipMpt84F56tjqj
LvC2jfHauv3K0PXKgTRdrnicJkNCjOO+sHiCVOsiBp4zebeHc+Wk3fwBSwTBPbYD
5tdNYoIyFhO7iB1nV80W6uDuZmZu91GC1SYgJcgozNdGshmKUKewALb0Oz6mRyzL
y9G0Xuj7ayvsrWGuWDAsZNZqFzMWxgsALIuE0aFhV22tEhcBBLboIxX4h6l7sGtf
w5hzKP914CQYkI85smoH6YMshGAKtO2Jq6thDH1ljSiRh6kbsC2lTg4ICJc97ZJO
FCdm0GF9BjawILcO5oqf+R7rBdSuQcWbOImfNcg5RsYctuxZSdwZkHShgsUkSPE+
2UonCb7qtkfiQTtEC8DavvIzCrAWPApcoDN88YhvQkYy0IHlqIilIZsKTduGJDDM
e2X1ajVY/+h19jeFVaMSWlPemivXQwVbB5FvvRQupnWQTjpiOPz79FLPaoFH9nsd
sqohH6GpU1FHZT/h+1YCw3OeIF87IjKiqX4VNPgDd00IqNhBKIvjOLa8XGJBURhu
mUxg1XAA9iKOSGqDgL/f7gwXk1XTwBQ7BwQW6qT7350Tgep7wWSNqXaDe1rXa2cj
GzGf+ypvBuGd4Y5M54ul4hIsgM7eCGeHUmFzeWApmxIQAY7A6H7sg9QCDEXf2bzi
NbUQVnZH5czdklkNAUcmaBt1ELvVeQNA/5Ql2aQtY+83+HjH2uhZoxBwvTsUcZ5D
/uuyOZW+PxZF6NYldibeAv2B8r/8TrIzQDni2zpKhLwvBaPe/ZGyD5j+DZiQol8s
pct6d8O4TMgfjK9mmT7Fo/yGZXMICtXo/owRxKS03mIqorcD/9bvZ2tM3l/sJG+P
upD06+madjSaNAxXvzSelV9m8TaURYvZhnVst8e08VWItvHb7rMyyWMjW6ifn6Va
GbzeanQ8T6rzId3Wyab1RLkKOUFJyGjQWn0CjBuI5Kd6xyE5bTPvomAESQXE47Rs
55AaDcTlTL9oTFHSLf12K+yryMwYa2tDWh2P5/ivn/ZZWvdC2mb+eGLRqKKBNuA5
hX4UnR1rwlC0T0XaZcCjMXEc2oSopBI5v13IiJS+LiRuevP8a500aRdnkDSBlkT+
oHSDCJVDpHMt2qqgEmDaWGbndXI4YBVxEfYaACX2Oh3RZDVVmJRlTgwfdyNhKjsI
DuuWF+G5F4l7aAjkD/aFdLRBm0TtbEMBjEYTCG6zCxzMRUUG+yqX6UcbPE50CV95
dU4/LI6q/mGxK2mEuxf+m2h8qnntwavDDnhzkP4Rcotb8TEqnwQ5x0HklqYMTcoX
owl7Dco56nPFMXqwiSsm/dmGxqfJLQqBsEYbyKlsICRdw54OCy+4kdcCLg4jPUzU
Rr6Gwqh2aDjUYdpos6Aux4vbCwQDq/PrvE9kIpeknIcCZLYDIhGZouHmsZmIrjFq
hguklE/LBPwPPfU2DryXp0wHl6b+QmUao0lZCKi3AftStsxI4hbRX+uDMbPDmEKJ
xZK2NoVLo90Wjie4SnrIwACEhO8TKffPeVZj81N3jOwqPvK3qJ8S9Bxide4KI+gH
+2f8Gnz9Rlwff81RFbLv0dW5ckNabouhUqz5uNySEAV0bKR80whtIeSnVeMAoQSv
hrtsiJat+dYipOkDiKLKx8wSZUu0+JtY96pQdRfpXM7c5axd4DYgFm+Z1YiGS2/+
7ss7eMPBRDI8dNECt4dfiv6nxjDv8eX8w0OS1duGNwLJ22OgvLo1/K0Eyz1nSp6Y
Aj+hDOHCbgEQ6paOj1kL5AAVTPGBEeDUwgkTIpJmVXWIlIIvn0VqWK+ZqrMJFVvD
0XldM6YZTq/N0bmuKNWtyzChETHZuGnf9gkDlGsHw/GCrpOju1H3fPuWTPLrT6xU
cZbyn6wxVg+O10tF76kZ9AMBDolnBCJAAJ1WNALVlck+pDL+wzHEOt5tAX4QmGf6
Tvv2HtFjAUlVAac1zu92au2POQ78LR7HmRGv8LxwtXAv4N7HKej2rGVnRp5caNgH
v4njdsiQG5uAgmC58WOHTaX0W3QqRxAMYT0Vlf8A8i/fPzwpZdXEp6sWVzgtOq3c
pPFeXh2S7gQpfUOoTH0yH5Fs43qdDrSe/75YfSOwnmhgiHs3mJfCv2BmQAx0PboH
c+aW0Zngy+Ak4xiug7qVmwhrlnTN50dJ7lGEVy6w6jzNkcrGY3B8xU67nmcrZOwu
P1mJxzFLiJddWYO43olv0cRgTSDaXuEUwQJFEmWPNK/oRoYWLsmOKWn3xkh569VB
sMJTZKw+OQcQkTjtwXcAh2kn0C9tzp6vOQvAGNsOpuX9okSx0HdmRRHDA+yY8PWx
wlWHUJnXFOu/qE8VUuIugcGWdUdEhmP8bvrtKsA3frahBi8iKazc+YMbq/dvkviv
bIggl+ngJZHHGvdRDHKjBCcvuoAOj9j6194rSJfnzyqvbDDFv/8kVp2jsrOkWBiC
PxsK8dfwCptl961Ubw0nK5QRNXtO1LzQX290d4OgE5hIsS7DS9acqS2Ew3Mb/EuT
jxlYO2bOOIq19R5OIv9cXHxU010n4B8/06+Us7gj6LqzkWUenMOErvxuGq0/I5YG
o02xMd0tSFASjOErjOjN/K1FKXuIA39/GbXXMpnN1rFjx2iUce1uTj+IR3XU6coy
c7V3Ydd1aAlmb1K9ZoZYcpjTa6RxDr0Kt/hPkZuf9Lew7M9gJNiQgm6v2Tu2uREr
R397/WROsC75odm9MOPHIU7TpiumFRwwWB5Kw08GRtUmqo03Qiwv0dY9J0UQXnEb
RGO+8A9rDV7iOH6OcxiuQ68s73w6ZPG0vwOPX1qgMkgVZDAOCkAxmSmvrMnX6Kgm
AjwWsNL0But06NZEiXtj55ZOJFDXLVZxDtcDgA0o1rxu8TmL2g3X1NsdEntAVpaU
hOYoNEwAcmA0x2rSomty6fycdav3nZlskdp4FQShGyfLK3oJ7NHhY/QP3PsxsoMI
IytJL8vTCC0Zwf/TNGpYH9lFO7wwXRrWSOfCLonRkV2wABht9FxsSM+EnEFbW+kP
OC+IXuuR8Zag6oF19hOejF5jKGSFP6HdcIbnqD45Nt3A9UgEsv+nPYVLqHyJ5rrK
BKy9lUSUzHxo2gZ9VL4nLCHRp6SaaDrGWFfuRhKtCCW00o9H2o3TLJHJxn7z7slq
2NW5ZmEW7RXCVPYMWzS6FwcLcF6R9lQCeuyNAWmNNelMkIcS/uFX16scGmdxk9Nv
iHBMjRVAH7f1BiqfxYw3aAlmhLHltlaRG8cdhFcwco9cH7EbyN4SrAZ0XphOyZDN
G5m1NPHN7/RvymFkekxMx1UFHBrv2o2eL08Yf7cwRfcIB8Dj/UAyleDGn2bZsYTD
zZm00KwvQu3h2SOaQGCl2/vq1lkn3Vyvt/WP+shx1eQ8DzDb3epado6JSzIiOWS/
TszVttBI+nwpNwruCAuIMjQqiNxHqsnawgPKyfkGZtJmbYagDLtK4Sbw44I7DNuk
UeNdFu9B18lkXwYiWeGyN4z7l9x39Jbi5NTHUX1/JAzx2YfPYE6CJf+6lhafBtWz
r5+c8pW+hci2+Ks42KjQ3iksbDgA4xAR2BCg/Em59fdS1CPJmg/9444Q1RNE3kXj
ltmAxL7Hx2cUgM3rUCwaDYl5NAMQAm26P9cXHC0NGVAxjzcQsS59KUszP/f1gggH
Or14QjYa076FGj8JrueVW3bF9aVstGRVCaD+dwvZEGk2EXOiTO6WVmHips1RAxVc
2uyMTG5Szc2qo9/AAWeLzTmOKRaq+e2CghHUDiVRS9mL0dZt65JFOK60Njm2kgbY
F0M9mLlhqH2XytRGAJC8W4Vh1JSqpi796AutsuibyQG6MNxNUtzT8dNTPGiMSfNE
lAKcFZrMveA2tffVr498J4ZMIAkximn9gYvacD5gxn5T/RZzK7vggJopx6cPBeq9
T+yoPUFv3qWr3aqqx5V/H5EVMdqa5hlGp/c3y8HejUPYHqjaZ5hnejSasOW7M2fl
0WdckSD+ShBbJmzV7HPkBPmfcWTOhTETUrbG+5yPC1yflIIubTik2uXDnuf93bji
8fsHcLl8TM+9+0GXBIgSqzY1/BG/LyUbuvjRJVOOjfLiq4iunDLXNLi6fRdxCbKc
IiEbQcDCHn50iXiTBJLZaW/VYPouB0ZuIsWm++uA8rPs32mRwdAlxQ8riFFH92+f
wxtoOmApjJK62goeq6hD7WXK8nWpv4ZdCLcsV5W2qDiQqMARQ7cMI41de8e1ptBk
MdPMCNdcBSle/3aJtFc27zZyR8lRTECaHwNsyE2Y/oxFZy952MOaVu5tIzkBl7xX
msiTc+q9qyG3mfIDGtDzNblmNuDcmiCpdLyvIGte9fFsvGhztPfB2U2z1PYjZX1f
mcQAAyTCMl0ZlDhC4DfMmgCyL/Hw0FPiKTGFZuyr4LyVm6BoQWtb4hU9QN+vblzV
AohW5ND/baVWOIbS8dzSmsnNFqOfJyFLwI7z5eBtaYjlXS8tmpI3Y7J/dsx569LL
xaN/FW53kXof0tE8EmMh2t/RjZsce9zAkegKSDhmsqbVZgQ4IwMGIFkTeR6fsfZa
tWZQgoCF90wc/by2mwBv/yg84ul00D7zcjhONmk37/O+itAMDb6dKdeBlp2LRje+
D0X/12mpWpKJW3ZANetTd2VcIC/J1Vo3RqVpSD9ARfPjDJJN7fPM9Mv4ZziqktqS
FcDvZmaHLF/vC5A80uEHcqLvruvHJaBaoIehyO/L19sk91ZOejMXDLyh69evTGLp
xcDQO0zPIuveWgkc9h+zssE5C00oupPozwDdmX0s6vDeACbxu+H6JNIlnBnEa2s3
K1I6OfNKh+BGotMZHeFSWRv44Wt7QbkmwBvX0eS5BLMY9PbCHRQ0tXQbmZYp8oDo
9ChUK3MWgGWGZHIZFlB1B6ckrzVg6rIcgZFNNKf/ThPrhuShwNcZtBmLcoBait+d
Xr/R73q4+PePEgTy7hyy1Uqp20E+YVOJYdTK5Cvhuf2z6Uj4eBga74eoLYL5Ng4N
QrGrCCal4xSGVYIqIpOPnar3ywqxspjLzyZRJA29xA9CO0Ktm85b0hlDji2BhLLc
KFALj0Qx1f2Vs5rOndVAp6kUHc5iKfHIH24J8/xSYvCnWm2pcMYONBH05V1edavW
tutHRxQxBZhL5hf5m3hdoZkb3xvY1SdK6vyypYRzmU972PXZsjbQ9JXysTpHJdor
qyw2c9iE6kZLez820hukZvf4mauridgUu+5D4yUv32oBpKIlsArvwrBIzZTqpgOX
Kq14Ql30hGEwNzsF/yM7yjrGpLDtvn5T924yHxhq508d5f/ZdbGask3SEWItAxH7
cUF9wifJSk3I/Cj/Dvbxu6OMc3eMiLmU9uP8arWcfKGpW5TXUH7clsn+ADkdMmP1
7yD7DFJgNyMjgyDNVoyRxcsJxYkIMsq+tUJNjEplDrIzDTQ34r43boy6TJEUxQbD
paAjHr6bbim7zwTlrhwGUVUCpbN6yUF8CoEFELtHMyW9hRlhBnkeAwHB8ge4vuGj
KGG8PIHu1zP9uEfCjCXazMmtN9tFWwOO+hZoTQeGTUY/riA1H4uN9U3q7ow8avDZ
Vg7uLZI3pXKPiyHzLj4ueip4ZLLUt5GsoBCKsQfeliq5baWn5wAVUO0Qx766pbou
5GjOEQusLuCYfciAUYSZ3iHvsgAVl1LYJ/wJUoK9CokylGSduO3zD7YsOS5M66eS
bXQU+NGD/3W2w9yckYrdHl5fKL42cmQnszgeeNhLFBa30ziswBjfLlo8Pac5P1um
bHP3tct8XuWyGrTelkAI9xMkQcJ7RzgRx5I3OO68R8i/Jz2kDzN3nqQjAkBIO//2
pByi9vOLtS1VDnlFnt6P1m1wm1saoCXhZWF8CNm1p3xV+fg0rpP5OrzZBeLNTIKO
wfSJjd72taMMasdRTP7D4XC7vh/qPAVLusrWgfov+313wh+Yf4seqkqRR5QpF8sK
ZWwPHjdCyF+4BnIAULwQlORrKLUIJ5vq1Hnlhx6DYUUIYdFCM2O3OipU8BiK2thg
8i7wJimRxDzrxHX2Nf06ZCqvcGgzoaT8OL4tFa0sBQYymdPpPJFXKtc0rwaZWz17
SOhiM4FqlUxoIAAkNZzNUarlxHWz6ualfgNxZl7C6PWJxPO0we2fvux5DngxzGXX
gLYGVMM556DL6U71/mIPQFT4HXrzabHoZlYhh3ZKaFBxGIG10XaKDjPdM++kkiOU
SkvYwTeymAfX22I5ogu7Vj9RPQV5iSDSaWzKrfNCo2HgEHbqK5jhmGa5zmNFBec+
D1DjGIzUrRF/Eg87dSOdVO+62nvFVf+xqiNizJnWuRnTFTlhKM6g5zF0KJu9z1B0
nmmHx2r+7tOtm8YVjbJbaqDuZznVAFHQhjpcZdklHWN47KD1oZ0/32tKTfjRVrDZ
fDcm4Lsyd+y7o19VGsrhY97BAS2a0bMylbdkhbdaD9dwx9g2RYZfdsZX8zgfI4to
dXvFaavzoWMV2ANAdNWPkEs9uYuBsoChFOpohCXh3De9XMFNc4AM9jH4wPAih0Z6
mI0ScPuInckbep9f/OMoIo6SUBUiYvt/nzWeSQ+iMDv7R2shEsNdk3lDOeVD/daX
DQVpdyJ9RS3yfuDyMj68F5OyUyLioOZB4b45JqNxy3TD7nLWM8hdXe486oqpVbD3
iKkgYia0YvCiR7XFrewXwtlZ3nYJZlO9I6zGblYWNOVZlZQfQnHiFHZHWO7191uH
hiy/LstpArgDeQ4szQeHHZwF/XNJtcF9123pJ+A0MjIt6/wZ/Ys8IPWu4/W12BsP
N5AywAZ6/EgWCTQrTchjAFZzIbFzqazL4jixNzXEzp5Jod9jejLX0RQghatE6hv2
VrVFa5KLruXFvmzZ8kGeYJqfQ7dM+jDFCSQ3dpcT3C7RjEDG5eElOBxnP2kPN093
fSMYLf0VgETbG2jWD/51XyWPexGs/+PLCLScQ2UEOTBuUaUjvoeMtTjVem0RUKWV
7/vGgyFBfoieW9CZCPEQFZtQXLrM/xXe0j/vFYOUiHIALD5+B5YNA6Svh43dr/z2
QWY46q6VmrL6G2TLNc3XO/sLuZQGT8NFt++Dh43nxE0SJYcRQLGYrlVVn2PhSqtI
6oLlDtwKhRoyLWTIZFlRdweFII5jWqASBfjMRALagwODFy5sCHhy2LLMq2an/y0W
e5hsj/o0JAJPnBVFGbvJafT9cv4Ue5zHFnA60Y5W5S0BLHKyg7lCXHMPp3Vb32nv
YCZqhcuBNoP7NDdcyrJMFkpZpmXsEnGGxn2OaxgwbEH9+Eu8aDv4adzeLv2eI59Z
GKiHG3rmLSob4zB01AbnQ6yBzetLDQ2EV9zaaSiR4ej7jJTPyOsVEVILgkKPx09x
+nX89P/bRc0Ow2m4+KeLbQYkkXZtwK92GmbuIoWAJfcoEnafH1OIqhp7Q/RPqXbq
g0FYcpLYDB2NNPh4WeSjraAMY0yDQRU1JSOBriRJdbMkFtz5aC46nG3AykuJ4hts
0RmlJy0EH7NvVMsVY14D4LKHZ3PgN5Ognx7aFwzjC+VzpdIocu+GduFEoNuviYS6
FTmYQ0NDi/z383uCI/JlabL8X7YCXwAkz2emwZ63JZdifyJ2azjuXnfbl77E2XMD
4Szj6gz6b22GQ8UbjS9bRuZwr4OgCDHpqEiLkhSsmn3vmSW0INELb2KYU83p9Ayc
Hv1Hpb0d2Im2Cd1+7dRJItAhWV/vwHfed79/2KzO8uK+yGsoD+XrCX7XJ0IRcFfq
RFP4TDfybz6EZWH9nrgffJJ5UMMR3QQPyZ0Ip2lV4GycNMRiKt0Y84zy9qj6Fch1
ky1cgT4WmvWv9uv0iS9ZQUfcf3U6PN0qWDtc/jQyPyE9wYs0sD5i78ng78TpzEwo
PDQ9g5Zr6AH/wp+juNYByJuLU+Lp0AMVMhVg49NqTHkopW/iT9TupgODxmQQi1p6
X5muFbqKNVjKRwHzzWkTBxrglDKelIz6EENV+c3sgH+wDo6h9qksAmjp0v3GZb8o
kw04DeofIWPw5dwzr3F4mOoeZVqOuqO32CSYQf7Qqbuxxl/4AQjq/a+V8qQPenbV
MSTTqYe3qhTCC4E5Zwv4qPMqcyH59zDQ83ATZxhuz/bn68Ho/BaXooh4ztUez86U
DPEyE0KKKGyqWULKaj7exekJROxqQPOnBjfAx+r3S/Qw0anKIuGdkBP8ewiVj/xT
wliiTh2TFyE3vyKJqp1pXbLLZOxfeL8KOGXeuCGzTOmKA+ZSXNDp+sGPuYW6Auhz
62I6hh31A7EsJF0dDxozkxAqm1RlVSivQQ1YE/dS/HXj4nGWCrY81cRHfkKeZkN5
i+fyib1CZS1Z2UOw00VJzLynd7fEUR3iBakm6+xITPPT37imlEKxHlDKJ2rSlKQH
Ssn8O2Xm56UkrEjjeH9E6NktZbFllADI5mWqZNt9H7jMHHFNe8MW9Gkl4VovOLGi
+g1lgQvOwJx5zKpPjChxBJWzShu8BgvQYQ5bAv+ajYS++XKF01GV0WGBM4pFUWMZ
Q7IwAR46zbRFlaRow0KD/pLCMGDWSwldsEb6Z9A/R8PXiq5qUsmy7fSJ0aPqhqc5
Wg7jp4VOKGoFIiKrzKBcrqrX4Mx3/wuYcpKicU+Stgh8Td8HjzA+GVcATsmrrHYL
/XXOG+FaOSr9THUh/IeQCpLqfbu0kK64bncLCle8E1C7I0zfdDn4sZQBMcFeRZ5S
JmaMh/wGjMyYsnzeImkWDB1OiIBibflUAt+yqnk+Q7YhJJ7L/PFF4hgC4Clch1qu
4QCvBHMHAwri6Zm2GLZxkLBC/DcC3oIAwGtc/w8USgWoE2O2LAN39WCWeWsQUmfy
UsgRbzaYx3XOU28nu1nTF25emXKaouLdKQ/KOZotWZHbhAUStMuAe+9u6Wb4lcV7
VfyUIsWa80kicX4IURsox8XnfKlGNDlo1xORuEqykzLk0gTe8Ubw1lWgnr1kJGlH
oY2XTfUIm0jplB7aguVvEICjx75enqpLAfIjfFaKfPDe3dekwQ30jJUbjYdxWiys
R1F9DphixB7Tu4vO4OVeM9/MGYTOFNgyzwVwJGB8fCO6KkibqlUxJPTDVWTSDXw2
1YIVsgcfb9Tih5WD/meXG/4hB3YThWs8hb2j1Bsxeh94OHBzzaaq/Ekj0Do091RX
UkcsUh0o75y86Ig3zpa5VVrh13Qx/HESLkk4gp9ISCw2JWATzfObUWT5mAOROgyb
SX0G5ZvpFZHLtai+MJQAGz6kQLGWpcPKsIS/p3F1X3sT/FbiL4zU5oR68fW9KJsg
MT+pGZ4LeACBLPOJYLNCs2BNMlf0MFMAfoFrh5gzqi+ypKwrEaYqQ7tWbaO6M0bu
u7CMUE0Dm/+gTHtIVtdEVOq+njTi+UCnnUmN95oC3T+AoJmAImiB1MW2w5xVSQ9B
GkD7tIn7ZHICrF9az8/2+vg+/vfPCaZyCXD8A61zWXo6FBdbND2NH+qlDHbCsGDg
p+3EvcVdP1JprkGmy9/dOp+uXh6UW4JBTXHzKSSvmBd8xkqFRyoSJbpCvu1ZhxHn
q9gHDQfQfK6y4nH1yhM4rQ9+ZCoL4RTGbccOfWoWdpUm+y00cUZPsu3ISIepBBuU
0s4H3OwaVhiY8tj/0bwM0uTv1E6iaBEnJEzLFnIieTZXMMX57JXf+SzG7z6tRryz
Nmlm7WYpPZ57cQaoxMcC0eZL522oKkz90wGMrEP8boVVGN75whfqZeoujgNPgMXY
hy8IFu0V6N7CBBxUUe+qop3KUIVo8OpYTEzOTMOd2JaHHmPtjxugrHb9bguXd6D5
ZzuSddTPkYJ00Wrnsl9bw9GomOE9ygkfZ/vWFJw1LKJGveCV4R17cG2YneApjRMq
U5mxqFb0hAz0mk5lmO1etSayHPu+RdXV8h/n3WjHM74oAvIxCu7er9mYAwBvcLBs
5V0VuVNQYShd81LNteD8aHcaGlfOTmTXqfcObfwytQjdeZitFwTd1kqMLDEpUh0i
3/NvOQqRehjovKnt37jUT/V65GdY9GEdp01Wjmo1GaxneDRLZmxKzidBnSIOF94A
uLt6M82DQqqWXTQtN0rZHdVVj8RdvG9fBdGplSJ6uS5rDo98PmD+mZtHGFkfPvJH
gJgljvWTikNGOhlDeYbBZ8qxuvq2Ff9AQqqzFt28H9c10/67hUk+7O9CQQKbwdFz
LniGMD9U/HuH4WtchpSEARH29IGnIoaIQwdIiEONi1J1jCUJePdmdSROMmw+d9qE
/fh6tc3iqmZHdpque/FVC/h1q2zsHcY2wrVRE3B72Rz9R202QoOSjw2uywc9yxgO
W62UTQdizvjk7cxDGyzJ2kk3Ybi6r5EjenvQi5j1sUp7qcglAQni7yqdJN6K2E2w
ovNbO60QWNyR+iVp066/0V3QkKA8IqJWmdh5tA/wb/fZ75+w9To7b/GdSJ2+R0Ta
/LDc5d+uDMnY8r/ivljTxz3LxdgqcnNTbD3CoB9I+no3CbAMVvA9Gdkqj1tkJzMk
ml0SUoNPe/BveVGKL695LnsPK+ZkQjix7jmR80Pk8LVJMtaE8uho5LOzPIW8YnHz
SsXxgCv19CqAbVL09AnYeDKKFu7kdG6uro06bMsERhdspYlBMNxAHsoLmmO/sMLK
+nBt4wwOSe4oOCTfBDVS1yuHnSmdYNtVAXWA6eDVKyEZoHwrwnEkJjtZpFp0htVO
KC7mkWDUx431pKAAm7Fl4SW9vCDnPffBddlP13bwvsnl3de9Y46xYviP038mltUS
nuAnqhbOzHmKK1dvkKQZGXopPB8nDpZKR90Bp8rzdXeqvy17hiVMconx0U1V+BDq
5Y7A1AxLBhtVRszFPTQMndveP7lPjzJ4HXTwgLip83tgdj4p9PP7T2rh56rxjiHL
2nPvI4qRX3UJC/dBLUjpmAQ+KsrIC3SgW7/MKATOMA+dE4NpjypR/2kkd9QouO6r
rIAVgqeobAs7xqJwlK6EHCxkNfRtkqQld7a7ilpOO2lRU0FNz6jRoMOI9kJJcaSY
HPE8yy2enZUF7LStzn3NxW7Q/WXAHjaFSa5M/wRdl+2P1tlQGmIWdFFkZt5B1Tas
L+LxgSFodL4mGxQEb4Z0XQ7X4pdeqH4Ip4IexPsdie+Cas3VfFMq0h7Twn3+GWna
m7fzOzz115HVOA8mcCjtvf9qRgqtmLqLBSHxAzPJMnRSGcmc1Ac3hfK3EWZT0mQl
n2ZB+ilXjN8qlaGA8sZJrT7jrcHru0O30WDCWsR3eYVdCdeXxIyT6t0I2Vg9wW/9
vdBeqn4tiTvQkL6vXxp0sEWagMZmUu/T9MK1bBDqqt9YrO/wSEGqPv7X4036nplA
WIk4OKCZt+HOSBs9bRETDTEIUeUpF3d0Erc2qCIR/IMCxvQYLlYn95r9YgLBZ245
kVJmUgY7dBftG3qkQZPe+xoX1K8sko6CfLNybn0gSXR8WE/BUVkwL3iMYJI7zSTv
xFFJK6u/G/kSHEbdjtgwUGcCy76qUFXQteb4hVo9kICXaOj7ItKuuOK5JCQnjtIq
KYTGIJZ/aUyL+nr8qoPu1iEpRTKV2d7Egbj5z3suEC/YuVsE6GKuhp38dz+DJtwO
2cXpWAT6ziUZm6CFaVJVh6GqKGbKcYZMChL4/+LhEJkgSYOVG/oRXixSKtUurlw2
fDnEq7MSTa1Ux3HX1kK86Oirr18Mec/tnWJf2Y7Ta9Fmk+8LIOeIUuChIjrt3j15
Wt2r7mhI3khOsTMEcssiBibO4hXJ37Rf7hk0eOGLJvXrKAjkT0skYr1CQgPFjgr4
pw3rYSUUxvhucnKedklUOH4QYnsBNOirMwTrm6EHtmLr6fZ2T65cxl1HTZTpb0ou
IVysBl1q9zfqAhZxSSvRuVfQ5YVbnDUFj/DCogHm0o3bWx+UIcUEz7JyK+4LYbw5
UrX41+Mx5gPMs572hi++XFRZJ8kgtpkHB10JM/sHKZMj9Cba0eTWZqobvV+9YZHr
0p0iRDU7qar/qZ0DfSTwR8P0369D0gKi77id1hEAPIdC9xzM94AoVpgkxsQaOxdo
YjYOwB/5qS30Qpn+oxCxNunIzUb1wLq5kPDe2qgVhLvNvW03/14g52NPmU0rW1LZ
ceo2OL0Dp86BCsxBGQ9a5NmaET8/klnbkDhScpBWixwseezE2FfozFFld/WbbJAu
+JZNbXGLgTtLQcBQo1CBdL9FAFHgNfE2eJ2DTVt4RWCkYme4HTJwVywXl6zE7ZyU
yXdVCRlQhzR82C4SNDUPxZaoLo22Wv0Zz1HntrorskjySPs+yNJp5ufcf3aMuhy+
vvtO5NOaBxckLii6Oq6vwsOwCyQn1ucMPXgmKbb5MeqgrMH/OwujOM8mZp7QOseI
dukqVc4Va+fcd/4j1L6EVRhkZ3VIM/MGKvL9CrAN+cNjw/Bc3XpIsqQrNErpzRdF
LRiw9mvyEfjTkCStrRLRlVavb/jn9ZwB6I+VQk9X6l2h8dKnHnzVfUb8pZ2VPYql
gCip3mqKxxaeIePk2NhHh88ROhdHmeK9BZEnQ+jMqDpOpOT5Ufz6oK7exafjvnOo
4HFiJ///wkpKC3ytN1kSjLF6iW/Z2WMpnyQbmMrgL39Ty/IowZ5x5iNd8DbLk4Db
eomBmkUQwj7BqUPJBXPZkDXZ53D79v95G0yJOgDIYm5ZGpC8a5dqGg2ge25RsSpp
REyxdmYpEDQehKdB4WI9EbXwTEQQnqGS4w9n8ieECQ84p5Qadnt86gaJkrbsB5fS
/uEdgF0MS5BbE+OW36qC1nHFWfAyJdpNCjrW3R+o1cg+80U+3tdaDV9ex5jJo9g4
t7Q4dCJs0KfNXxEWIprA+RHfZ/2gN/CWyYahTz1k9gofq1y4E/vb+wXIIJnfkFaE
RNuaP46DAzY9rC0Ouvv8+5cRK7Ha+39JVatZaE5ljhMcflHClkQ/7nZ1Q4axPqYL
YuGHrfu7b6Tt0ZWxITNSwZqvbggcsjiWpPuXL3p1KvMunFdRb6/tn3a0hcKtYVU6
buxvlJQ+ctatZwFK0GXOzFaVMUYlbmeApQQsQcck5zbNz8n4M7RAOliL4n3JAm6u
dGa8O4fonvzSCkcSkJm4WiXiIFl4ABCm5tYbLK79AtI2ioqR+BA3p5IWShwYtRD3
kHDMNjj0G+AQngmF7ob/4Bi6rpN+VkrEBUNMvpXSZ1uwuCsqZX23PsIfJ7RNWUSO
XGgKZSzcJ38Rd5zyffsW8tQcmt1hhjTnKHje2K3WVg2IJ4TuAwi3ne8WO4+7wCvE
tyKh5zTPdSi3MaK9z8nNdBCNskZObhD4Lbx1ptSA3xfoXvQrGowDm7kcOUwgAP3B
PpYKTIw5BR1TGkZiVyP74zf4K2jBMcEwdpgCD09NG7pIj/jNE8mVG4vRdkhMhtLL
fGJhPXZZcik6f8hGKcspfNoxADK37lJEPAsNgpwcdp2P6ToblgTQGac9sYBHPrb1
ZsBJ9evRDdGFPabMn49iIilMuySiF2NehSmABts3edWdSikkGcfZiqKL3cx0HyAK
5xvLMerEjw77+yEulECluWT3JsVjyJVzJpI+AuCc8riEMi7gY/E03m8u4ZcvK/I1
1B0BVnazcb9L1zYpiX97KREIiq4pt4cdhTUA0ZY85AmTkaypgkFHx+hEYLQGA2Y4
JdnVJT5bixdg1z7xyjCqmn7nfwq833gUdu/BRgo52BiSWLVVhXs8yDGfxscDPKZ9
wFxdIcZ8KOi/fkptKxK6hIxQdZ0T6zQyhGF+pBxW4DWImz/4iFMWv66IGkiHkLMi
bQtGqPDnCpn8OlpgkqoS2QxW149NVwQLYxNjfAxY0uteGaJOdgM6U+p6rzfWgH1a
6iuXcBbeBcfl7P7haRGcKjRgzY55jgYmmo/t6yuKGEOnuiz3gTYb6llo7tHK8BKk
hq770VsAVCn5ZQUt645iUO7fDeGrqzEWLNnskYzNGTzR/GJkwSYUDPSrmJDmfezt
C27OJPs5tQWDU904IrYz9Hw13Kolxa4DApiuN5DSjVfvUAci6mt7H8xmim2gStrk
cPUe30rR9G694g1KjcuXzs+Wto4+zMG5OUUyLNZUwV/uAeKDk+7GfeCBVMyY84nI
L3GBRvo8fAk0GytwvkEygEuBm4318N40/MnvChzmdmYXdCzl1CNXCi6fFl3Va1zH
dwBuTSY6W4fFJEQXsiz5ypkEdTphEaXl5y+lLatM87szt5G6nl3f6OpXwvhMY6Md
xvmvlN/kVYv5o/Q6VPxMR8o514jcJ7aKR97vr0Gnw5sFbP86+SuegnoeEeSGimSD
J2tFP5RDY3fpaguIdai+Q+KKo96+BRINScW40A9RyTwXDEIKUBfD+b/7/pmLrAK9
0+LDwcmYDPXE9CxfqSLQS/zfGpkNJqgY6qcW5XHFlifG0Pt0bzUk5pqhUTpQDpTB
ltBsoTygV1k9TuzUb3saSgmt+9j4SE3mR0vwHCbzIz0cEa9wp884cqRmrScJnBx+
bmeMWK0/VWu0QX3fKpWTVTbae9scNrs/enEd3dlWiwGBXVTQztgWcxwV/hfFagBc
TCy9Z3JiZgkuh+5UAgIF0CTqWwLMOKHhkOQxgkxd3R2UqY6Y+lQuPguH8yzothOM
bRk1MP+mmldpoS3JqzUi7kWTNB1yyi6iUIKLMvdftrwQYkMjWAfzLVXiPyQIttU6
hVK9pfIC7PfMTZdnGBTGAX4kq4XG3a41GgxivMO0+IiuFlVANVlD1hYxvaFpBiqu
LXErIaBJhJa7X11Fa9rnA5Zuv36L1ScYGQVt5qZYQ9Q7wKkTfM9W+g/MRwgOtvmO
FUdt+xdmGJHb7pU4sX6Uzjcz7JSjppVgAHGDNafJgUOUuYGMOfCIHBZeT+UcYUQi
QeqSYJigGHxW+gDDVFxE5/VgjZepAW5bXe2VYLx8/3CfUEEPCvExzAqzGSsGFQp4
47fiRBfQeXBohcF+HWT37gCKip9hjoy28ZSkDaBll9/+dwqePCHPVaePa7nvvkUm
ZiwrkRiROcJlFsxEBv0UhotSi1X013bKY7Hv729kZgJ1DX1hEGMbSCEhwrUfjZjf
nZazr+Flr8VX9CLaFMYEdsjsj3ZW0Lal/QckJfrRZMFYup6yFXQZCuAJrOdWiWpp
7+EHPyr7kCrmRCCrNU2Mr865/rjNY6hwdio23aBI4vti4VPHjeWf5xNDpL4qLmTn
6QCtmNL3asCVYU4e/XGInUu+M5O8a0BjMT+BJLJ0Oo8BOREunQKkAIgx9L1MASfA
ei8M2JWPucWvqdJgBgvmnx2SKVNej3kv84EMdcSACQwRQYx0evEuIDudL/3+0G8v
XoWiq+5LlNwUXsFfT77eHAtehwy82Hvb6CrSuxmoYp7FV3u2mRPG4RJr7eGL8bqw
0lNlSTJkudNBSOgafhUHWIJfTrhqG05GznUpRsTTSnIJNugDjO+w5EdlHVRb60m5
lznZI2dIQrBoaIZNebSji9Sqkdw0vsyFZIltQMsfGEwabb5bugaxiuSD1vQF/+sc
4zaPcPyTocyl/1V80Xf6xawTU4kZx27c3tAcdDC0zoRiacYqHUvcyOf2LgxbnADb
OE10SvM71NiAokGuGRSzSYFStWZPYoelBYNnMVLkrey2XIBO1XrbCkvTbs7MozU1
Jn1BEAWCTJ7/DA1n48W6rUNe1Q1SgxiVptxJvGX/dNXgCZgezBDBXePh2uvMb6gs
SXzjH8Btz8NK/V7KGRF0Yr/Ac2PO9POFvoVPbN9EJCjJ2YJiF54uPZF6k+gF+sCf
OSIT955RfVYD4pCqtO072agK+fIScnkEgHbzwsf+gEoUy+J6XX7KLRtZr2ZESzrk
L/veFF+WKKhNGILMIujz1hyRURjjv/0JZ/O86NRMuMBVDhdAsbWMl2B80m4zCT8A
1C1Mkglh13Jg/DaygvnCVHWPprz4DzxZNj1nSUkwiOHM3I39gT6k0RPJitCjaRIA
/zXtb06rwZX4/7rEgYbKeJeQxRpyWubv3nz7EfekAiBmU4xN6wUCiU/f4/mS4r/t
ReLXq6pKh2BbED8flKC3629EPkJ4nHCwIEgLZsf0zxNZUjeM3FiZXm+l+X9q4bHp
JkoAOb8J841HhWktMOvwtswPfk2DxSK4Oyl9iYZYzhfBJf96ShEdoItqJf2PFd+o
2ARj15BIBFB01BlHPPUA8wNBSqGGj6xiApShqYJBdNfd6xCDXWXs5eTmj2oTtJe6
Ouz7UqkOCquf5O1sWC1jDxp2KgImasbxjqUU5TwzO3hxkHCGRrAp1AoegGbMmdbx
CGbBiqyNfYj67MWA4PvnZgOPmhJ2JjJvMwZ01a+CVLhqDyqDV+kAfsattHEmnu3t
V9RMo1VYgpEi3rRIGxuBG0BzOFux7WUAutGqYTBzxw1r4/DcgZFk9lm2NPVwIYYk
9Y/VNwCodMcLJuYsNJ12RIUCqijNTCOWt6pUCFI4mz/i9NZR28EWfmp5PJ7GA27v
FbDkO5et+lW3qhLUZslu9zt7UR3RqmULMYpi2RqKsLOps+RK6xKask9VufArcAP0
Jzlj34UzVXpi4ZV7fZHvouYewEUnOASLRxwk724YsdkT+/1xcsBSwGTU1RKQzmly
5fY+Lv8n2Uyyr3I0hpx3Qj+GI0aMFamPAHpfMAt1rscKXTx6wIKxF2scQjzZoLJm
0aEq7MeYAsDsuGLnCZ3k3rBw1BJHYIwUieJ/a5sQ5Nrz7ABvq3GeUECBRGT5fBpf
zP8TJto/RufUNuaGk4e8jperIjPUPW+CglJYEU/u06i+KvLB/Z5SpphkQa1hpN5g
J+aMXn91YqnW7KsRAFDi82smqWpxYsghJukuz5p7aZMEqsFmeANsf96gsFF7BHgj
8MIH9nHA9TCnLbF3l6Toyjts0+3g+SW41qX1oXtH5pGeRtcfr7I7HTdcm2QhDgMk
WvVg/4u+RCkLs7bTg1yxNtKOsuH75XFu8iYmJaj69yf+FfAEOO0JLNcpgF3a8S9V
8uu9AaM0scGQ92unevyYfZ8MVqlzH+l0Qud/okSzRoWtmxlpeWkPjJ+nTNFD1pDT
fGCDxBskOLsm2oxBH2v2T6PkQwuo+eTN3STvR6vHN6QqSWBRChZ3lsV8K4QCx3/8
zoGvMEzEjG7qjJ2q75dXVk+FoGDv1gzPg6XktHZOOiMjyKl9j9tynSL4oQfoxH7W
zGpIzC91Iaqt3RZVdfLVaHe88s9nnPUtM/5A6WmD3WdJwA3VlQBmxdb6kH7LB3H/
WfgvBbuRasimEgRldbO98JjMzgqhK/rlCUERAhiygRhIRkksW4mPaydBfhsPmjH4
2syoO3R5502tYhPznGIpvIiVqn1+ANiwAtJajXXIik6q+Hc5NvDh3JnkWt5mx20H
qpdGdbdbR9kqWAtOcgW6w4y8QrEncq7CD1vGEdbxV3G4LscLLDr6NWQU/K1gkyfg
Mi/25mryJdcgqATbEv4RfngVQ2+EL26lrvyUyVdj4Xaevkeg5bJMyyaxMcHbvb3v
ImMD3PjyFZc216BSO4FhWWz43VB4S8kMU5wZnY3P3x2NfdjAK1/IsRVvnl4trM1h
6fP35Mjep6P5ExqOKS6K+BEJXKc3aMmQr6qauRp+346+6dvY2l779LfwSxoobC6q
iPXQhFtq6UmE+i2cYHsqRh6uPooM+/xVvw8wsVRlsskuRinHxmYhtWrWRRmFonEN
iDY1OjabstqQBBvmS3mifKVRcW9yaHLfcZE1RlFODVp0GaSFJD/KWdMVxBhE7BAS
Qz1mHPF8oGZ2XwR1GAsOI2byRRinmYFfTXZI8bbWBCl4QaxclcygHQZPveX31CLR
jz+xOD7qas8a7rN1bVUB93xDdbfQldPBrPv1gtxZgpIqpXb/0D30En4//k4TKU4R
/tZ/tl+3I34UxN+Om3Ris2AF81BFRMdB+LbNMsdQdYUT/kyBMAWsbHrh5ZZ4oX2u
5MTcdf8lgQLBtVR6c/QBfhzJWRguPcJC7+FqZ1d+cH5Lt0yM8VU+BPW2blkFxADy
5A/Y6QaIjOGpyKdPaeCr1GvR2cP7YKLEmTNt4XpJEDg/LXWIuIVMdF/MRQaj+brw
lkMqVkDxdOHASKVW5QxmWhfiVaQjeiV63FJ1EPoenKDJ+AmEuPqJ5mUjaB7VS1qU
rtN7qazYMiLM4ONuKtXexZxsuqLe/xtKeheHphywMbGz3dAhMv9viLZ8xauUKtq0
fmRgmEYsXMWqi5i8aTflqeZXMfocZjBafukC0lYmLKVwy/7uRR+vo4Zu72x3fvGr
QHrDPC1Dvk1Dw4wp1L5WFSYBh7KbH+ZreMqRuzRsLxMFejoliRC/6pWGx/ERgZQB
FuoPQ/m45ZAKwNiJysM16ViAnL3VtVP8iRqNOE8TJNo3RJxHXNBARJu5B7sV6Amy
LvOAO0KEcx+9C2mM9znr+6xAn1axSSp7fV5xXPayxaXZf4CebxzACCsm+yC5drb0
8w1VXMgxGKHM0+smKRkDte9Wjm8K0M09Wd5LlVwM6rqw+bhdkX6RM6PE2usiJPxS
3hYe8ywpZByyCvkR5Y7S9qHKFbvmicvYCTE5jYvcpqG6QgE870Pg8e9IULonEhds
tEMR1RHfKyYkQi0PyNn8u1MpowiV5TPCuLhIhhWMbImXmmF2WOaRjhNXuTVRlEzM
71U3Qrf6N5875wf7EXgaut91YNT6k3sX537ZymCfuUmQ7gWPMbk3iFOY0IMVNpBO
QG6JfXpSVwLAIUEJusu64I2M1z/WikPn1lLtwPm2hmZonCJ94wPgqrM0beyz0G6O
Sh/5KQkPAiWE0c5PDjNYUs2gd90JRaOgjDvfD7cfSzMUSXE7+0zU//XruZswkCk6
Pz5BNGREV82ulrxVbXnr777rsDsN4eL09B9Sn8neBnXLX+EuUqFQfN0Pf7zTGL4i
m5/EIFerwl8E0edkGdKprjBVT30XM3nVbVvUE+H+zaPNfua82jSsniO0druPCbpd
1FIo4enWkiF2LBHK3EWCgiNvg2lM8EuDCp0BNfwVp9FBYTyMcKv6HXdrtRbSsDEK
OToUpA0F/PVfcejfZpZxbVpTK89Nsk0r5OwCVQooJ/60QlyVGEITVMcx95ehKU1P
WQtdzie2ohaRbRxIaaTK+lgDJYZmT8852PG26Yd+pRPHQ6Ak27TyHyDVqYYv10z4
Tn8kSSfkFqzOG5B+LonbxjcEoCqDAdTH7U2yEL7Qq2wfA7UaxNa7axgGKEpNXQ+W
9JWcJst9CxcNWWCoe1M2V4pw0/opVwkdVbnKYvVzxz89+Eo64sSEDSMArX1u2Fnj
OHiCGpoWaBLsWbqthwzt0vsnDvMYIr9P6jtKRR4SFGyuVxvzYXjOEuU8w4AyHZV4
wqd9M3OvhdcIyPLDBb8w2V/OO+zrdc6fFigeDlxzo0lqLbOysZuiKZgdM3WAKLRG
81t+9UV+sXbINphR/N5gOCyR56abM5f79XEIeX4Af9iw3gxNm5salKVJUGO37IR2
UNkX3RDvZ++eW24bzLzQuyRJeo5yCjPA9Y0qvzUWXzXZ/Aq2SeD02S0KDKTeBUKS
YSyJSGUpAtm9Qlo908H4saouuChpzrXSrOl34fcyKUCg44tlR57Zq9qt2cwVYl+c
zPhcdM+QUNIko3p4qkpRwURYQMuuG6pmzhSxbSQUnuhvqQQTLEIo/p6w+hKfPoHT
RhldZft/YHFVRlovK22hWHR7xoMzkBCdSHdM3BfBNYNRZqm07XKuiNbyCo+Hd3yl
EIsOo8YdEFYCi4m5XPOKACkQA4+3WD6LIux/7rb+FWGjhXQL64yhE+9s5dK8DHLd
YSo3p6KAy3Pf9Zipz2Wsjchm6YaC+0YAE+Dh8rWfMTy9aNWm56QXZYXfX5rNJ6ck
Ba+XFS26p7VWBvgFr7tFha72QRxXt/EBXxl1MNaGSI6URwQIkfIs/SSxlIfH2lHM
+VBySbEaTFydbenI3ddK4LsKa6/mUtHkhhd3Scj8/2dH2AW6NZkyYH2tPMtRQQY5
LEtX32Qe+NqHcH1XOz7FYQj4H6U9KbJWMDYI1Eecbk9zytB93TITGMzEAxswG5l6
rxNETkslEmOgoVyFyuGpJRFB+3xoAHVkv4xbntKnZYdytA5c+fW+QvALE1vJIZXl
VEaK4Vj3GCKJm16UIaa/xmp/VId1JQTHVq2VYoMT1GtdUMtLmf81Zil80RpPkQRu
bosqKewLVpjKIKTozkOl0IKDJtG7/SOPQstNbMsxDm8JFquWmixofuAoug2yidOr
b6XePkmphz24ReVKiEVReifxMEmFlD/dGWOoXg0As3VQxOgVFnuS+laZzd30hMoZ
IpAs/3QpzuomnjLjNYNyHemDyIEaASTsp0e9ws65hCEeDV3BxfHki0TYGET0Btds
1jJC8CvSUrAy5vCizYtImx2gHNzCV+ZsBB/FquW4wXSQ2C2RIt4yJ+7X6DhOnjXY
GGz0gAs9rtpNwHxxQM0YkSo6inESBRSmVpdkedzdD8I4SfVzd/brGLjqKOtnDu7+
sjxdnSHbPaau5wOcxzkJeBq5RWt4/ooLsOjhVthlhPplrjRIqlS1rSRlerM0BCiy
bbetofcY6IJPn++9oyv0DDOpY10o+OVQnN5vZv3/R9Q53QknbzAqrhWqu30eRrj6
5WJQ+o45xye5OQy/SYAqs7hIfc1fAB6ktRPZUOPgYyTDpkpbUu+cqvP4/Z1zZdXn
i/l8CQDx2mIyaDWx/9Yo1QhifyIZrefJSV5b1Ck9Y0CAPAb4U4VEs6Lfwq+Y+G2K
CkG9Li3LtptEqZZPNT2k22lllxW3KbRYRNR5p3t4J0ZPlaChjxU4Mr/OmPtbGUiJ
73Y30oIz4OBWTdYa8GSxb1ypqYcw5hXCdHN5n4Y2Pc8YPPHrkspwfw2v3X1hHJ8g
8E15Gd9synlGlvmFszNCll7y9QuUyoRIedJndA0irCl1x+whSWJj9k+7M95Q3uaZ
fX8d/BNL0dnmJV9OE517uATJNe2jwv2yMSPcLWAhlMbyFp/e4c7tSIacTgue4oy2
dvHux8Zs7BDvVndOyL9+U7Ov6JK3+ojCRIK01pCcR+UxaM+3GvfgUteI8CXwIY8o
yy21CQ4qz5CSqrUYMTB8qhP56g7stlQz2dxHLyEID7pQ8YBcpsqyKgwFAQggIcJF
/Vr3kNczkR1hvnM8lR8F8bngTOYk66qX1c+YGJHA9r2gh9A7PwkXLHfsMbY0qE+o
LyG88fP/sGmi7sqhWitvnCFgm6K+CZ79Y5s9Uvfw/Uh6bSqF9wJJDjY+ao9/w5j9
NfSaIYo5kW7lVGX6gZwlFuANP6RuSuk0xRq8PrwXYNG6l/K62UWutHGy6nxT5apK
rRsxf2BugA2cm32dsVjhrxhguqm6cEYVU7fGpxImj63YsqgEeU/TMEWyd+1Df3g+
QqZ8LITsfXUZGHBz/BVnsUu3rHK6PUJhORdSvf8kn4Y5Ryd77ux5yCe250LEhxTW
5umJQwYhh0ecyq/tBqFf8qIak/YFTrR4s/tTvZuoyzK0m2XI3LILYL/zWqfWfVHL
DtrAUzHMfWLyN1rwFnviAzVCiaz2GXEbi3qvJiTyWdndy+IJl7lTRGtoNCWhnvW1
PHo0CqrqEAYkTem7Wk8VwTDmXQJcTlaQm2r4y4k/96JLNmn6qHL3kCO9VAfVb7Lp
34bkOJBhKXlyUYyZOFYnGCR8m31lbhQggD3K1PguSE+fyn58/xARmDuIHlr+7yPJ
PHh6Hxqa2uWelPPhwITRcrdKx+pfX5VC6/Go2i4SNzwi2UpvbCrlXhVJb6Mddcse
4mh5YhYqL9kO6mg3t9TR1UPZKk6xTS+OQ7aNDkW+RNBUCmssdU2T6g7on0lAdRUS
vITqzkhnN2LXIjmosN7xBMXOKwKMRRsgJ/96H7C1Mvj4NukscfgLpolIFcKFQs8d
Yehkkeb5u55cnhIDc6GBYUCZCmm1ijC642dsv4Q9f8LLwzCD6ilL7sypxAonc7Yj
qMiDNIk7EtDhIMAPW+C2yBrJkbGlF5HOZ1eMyuFInrUJq8ZACDEzkCEuLg89GtWo
aabozG9Afus7rEVQlUoYGrZgr57oFOEYEGdseDJOX4Ao7mhH3nRoF3DZyH3euN3A
PL/lbotnQsqNSJrDz71sWJJ4W5+9U6xOp37S0bhxUC/9sNSXhokXXsnBskLj7Uc+
V9/p5Yu1lZlNaH/7iBZA+u4rRxkNO7XQ6OG9oXoz6bk6Dlf0TaDE0EIRV3vhcIoI
wiGL4lw+SysE6ajmmNtIgvZWJzcb3T7g/nTX2sk0ZH13SXzXp/fWJa0ws2WDNU2F
wvsJLDjzgfM1EintNSySZCdxPqvyxiJsjaMCo/TqqO2StqLitxgENbkHyhMLEeAH
tfz9koVKAtb33uhs5gEzH7lRdeFrPAJXKdrMX5r6oUkHcSVdkJRGLfk3hzzHxIil
d5PICHnQy5ewn/yYKqXck2QOfDM/mgJBFmdBFjRQGUtgaERX7ei6YDiwK5vmmHk+
u2UuV/PcOIbBk61C9XD2mXF6WO+JzB3+dVmEnbv8HpQModmJ5jGkjpxCIbMhzugt
AWUbCinejKvf254wNGLhpxvel/eQOT97D8t2I3Zj2iIzx/9KRp73Rb2TvB61Zll6
G0zDtkkn8cXQ97Dm8HNdBSsuM8GeBGdrvM+WhgEq7E1pYANmRYKhxTT0ANUngWZJ
vDRHFQZ27hNR/tCxa6VBNWZsMGfg/kATz5NdLb8P4zEXT87srxupe00+oBL/UFZ2
5PhwMRTV2eufXVoOuxpJBfcOsooilR/v/jzEwVaEFh6/NO3h11iNqI0uSg4tQn2x
wcfMZZK3V3KhNyct9guQ4xroRNPu5PK7Cw/3y5L5Kk8Lms79YuZoJ/ZWfKSkeg06
FbOQukSaSw1DbzxyOzy7kIdtKYpbCprgu54axBAg5oreMnwCyH3So29+orOQcQ4E
Xjg7m1qoU/DEEFU2huibJBMai384iWWB9rVHaMo9NdYZO9rV+Yr8BSKqTynKnuX+
tfq3pCwGgi1BYrTRPKRGLa1rRhzhQFVmf31x8kiH//Vyv1Qo4sZr9EHT7dUJXBTF
bUPmxNZx2pfowXCunP1mKS4Y6gb0ShnaowEzcAmL7nG7xps7sn/MK8z665LlrBfN
XF17vdpBAqZsCd2gxpDNS0t5+wSknHK9uVq9hiFKKLyYHty4leurIjTELbSZ56kV
YP2GJ8OgRJGR3v95Ja6moehBBjr6LGiOrL48SbGDdc8Td7CiWoN6OsUrIU5DfYJ9
NSxyazIAlbXYkUAa7CLhVK1AhBPJGG0LB+hTM5SOIPdFfFSD8CI9YTdbJ+O0NE+/
CFj1fnpMxVBeLfsVv/yj06D/DgHbhbU1b1jvmS4FRb0eGE+64yJqj0tMSepCjpY8
BU8quqOQh5mkWGsTB+5IHKWE8mWt8Bkicvdg4J6oWo74gyaBrM5HArFrevg+p59E
MLVNNoe3ZLrvnKaNXjSXSPqrVKyiz7iPQlzbqgGHha0QIAbF/Q+AlUhJgOhE9NKu
0ZeEUT2XKt9ywxsxRSmiq2Tb9FmpkiJicroZJfvX38f+UbA7Yhb8QellqBWGmgip
TqUdYldLxyTdU8OnxcRhlZT4/3fquQMWlrDTDV/iV8JqETTRnbJPJ4Yed3/ij1hV
f8w4npaRZVoiyTe52D9Gv20wQ6FKl4SvKDV5hGZWFK6flS42TbzoU1abUyWS9lJJ
CMc0H/57LsXpAGVNvPhMptF9O8rrvRbAPfEdmPKAFeSdMXDYbFkdur1+EMsj9nQg
oRonF1NhinUv3YRNl40LikqTfKmk1oOz0Z7ajsSr8AFB4mhWgJRnkcHBJ3yUtq6l
SLlG9pDeucEGWDXS94ac2/ZrrqqC3YFfidj0oDyB0CVukARFeoK1jU+PcaO5aApC
4dl1oP6VwzDVShBUWhFJ3Pl1a3OipOdQ7767SsdkZyDqlUwO9LqRUyxPkp7NVJfV
QhV4Jt/JW0M3i2+2nenGTKq6aYPUVL75xJZHU5IqVwRbCrbJ+yoQFEVNRlKZ/qOZ
Am/EiXvPoFh3TDq1Sgp60cCYVZOQoHHdi3CI27zkZz1tH5JOgg2XsMgvdhPz01bQ
y/EOm72l0La8gGFoCE4hlagOwMrOkbeGGo0NKvUoVGrqgb4ZJNPhKzr9a/kyNf7o
aBBBaRThtGsVs6bAUA9i7KkdrxdbGEBcZiGjKNhqtQ2EdD+IrbHOudvRS5xhmBC+
WVizt890dv35oxjK2zg9uQE1PyOLiny05slGBEXMlhHbnrFnm3qLHoSypAO5FBho
D6bCW6YNY6CddDt3ZZvlPViGXAtw9YKqcl8CWkSRxeHjGOlWVhSxyGvt2HOljgnX
PPcNeXcCY40PneaJ1YRrwkVscLYFYmPRCfypz46xyyl11Bt19E2wcOZuTPyt688d
DkRFg3KgQYyKBtaIKhY9XZ2eMduNTssD4SWjG+8CieX6vqusqHf4jKL84tiQXjLu
jtuOjcjm2QKIZc1gn1rpSrlv3K8EsZ7rR6iiHaKtDjyFkw3jykONyi5qPpbtsRGz
xr26SoM9ww2BaWLtx3PLJSTvhrf8Q1+lTQYUuPlQ3/y8R24HueCo/pCSrS/PrNF4
ITq7lS5KB10ezs9536Ff0JbV7PKcNOfll9Qn5iQ6lScDFPOGwbsqfy5/moaLDkRp
04ksd7SF2zKmCDGt3plC7d5yFCmYFT8iwxZ0ro49Y+4J+q1X1iQQ/sywQlsnIgJg
8iCknw+pHu6I63oEQIQrh7iWydNMx7eelF4lc/geP35SABi31Z09Hon3QfsJCvnc
tT73dF2Pn0NbHW7DbwyRR+pU1TZnr0vfDiMRNIp5kGreRa4E6AFAczVYxyZwLAFt
jA5EyNlf6/PFhfusTehvu1IKswLaILlYdVBCuWQTB5grwwyUGZC/QpTAZzW310Kq
oA81snklbZCWhuvaHrT7Rbj/IHZ1XqIcqs10BfcpXVk+Pa/hyqv34REOTxL9VWx3
6CRKOgJwOjp3JJbgmq/yFGM0BkGxNAi6F6yeb2lWts8a25d8gmoWUHOlhACimH1S
Lez1K15a8srTJifwA5C26+7mcNNKO9IFczPCeFfDlogMBnssXsAxMgZrj9IXd5ob
s+O70VRinuBycZlEQS0RlqEeeQmlwC6xV8+jOh19invD+YUF3tAnB7wVOTRqIKUb
c7fZBgDoCahKsx0TGLu7l7bzokamjVWfK9DMG4K0tDjYpqn3+dvVg6oRWZMofQN+
LKgNTd8gq2ApnS6fdP43YSVZgutPc0645lVXclvcti769QTrOLFLIeeT8ijARyN8
bm3HbcAcuJ9so9UEDD+ZLccJSE14bkX8eiTBvATSLKr0YMFIgzvxFDVRW7tJqlEv
xPrjQVlPh+buUqTv2HGJFMmEpaehQsHZUyXP2jnltKT5Tm0tzi7xUWuRHDSPgrbu
6awEyMdKXrIpc2gRcKKchLRmZ8AyFv3yj032W7r3KeKss763BxpEq92dlyiDk1s9
9ynfJ3Jb5SIUbcKmllzwezOHXt/hFafXDAOOrwaUvXRNvBfNDCezQPYZ5hm8Px4s
H1E0/wHpcA+6H+SvYVXQSVQp1jSy+0g7qnhoxNgrqgzfzNxVzjs9OiVu8jZG7HoK
EuozE0IcTEOOccDR+JSFgiYDlWYR0e0zPGA66NbXL+FZfk3uKq/oMOokWFxWOdVF
WnPYz+4j07npISGs50hwNhSZFP3eOTXCHPRhq/ruATcgyz5JIcUTwLTHNUEZt/bn
Snnp1KATibCVLtkgdhvGta2Q0ty3mUt9WTchM2wLKa8mop5n6+hkROisX+ovM3VF
MrrkuADnnWeDl+XQDc/04R6w6rPPOf2N/ZTxzR6T7g0MOYxFyb1uRdDT50LV/tgF
sfTCe6b1M30ZM5kvoz3JdSOiuKTFpPQKuqh8IyD/pkQCgnQVxAEDqNFoD3WOf3f0
/0cMdZPvm2wFWzgG9u2Rj7kQR5dTCy3RSlNk5A7exPTb5uu1zIVFT0CZwbua/sqj
Vl69rFxu7FLhMQHahzJUyMCy974yqX1FSOjPbaUhKdis7DK/NyW0BL/tlae4ym80
`pragma protect end_protected

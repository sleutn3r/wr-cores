// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Kd4xZBGZAby/28SMyyYOAA75C60WTH4+PCB36Rg8jlhquQbr1zd4MHVRoJ4/Y2Kz
LZjYxWa1Ffi5kUTi1sR1m7AiRTxlgoIoJBoIpDzp/UdOPQRA+PIJ1ztrzNpZDACY
waNwx6nXjSpY41V2qj+JeFx9pcB163CRdg4/enx9oDA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 174144)
ImZoh5Pmq4O591h8BaUXv7kU9s4gN16EeKdWdAto97/PTusWoTtZ5K9AflTzPpQH
mczSvemZdWGuRp95DtJx4BBzVjW5aYUMBN46EdaTSqpf8bNcAt3SfTa623+AadP1
f2xnsKfv5UyfkY7hShG7DP6sjfx3YlWLRZjsDx/zbP//oEmzLzeJxFdB0I/+Gc2e
nLsMp4rz3PPgunGS9md+wK0/M8mwfbxmHs9XX5hgeJ8A+IxGutl4TenXUXxs55+R
hegDbs4ZUzO8CXq3THz6UKgAN+hLttJjK0oDkW5soDxofKP5FX0b737xL5nwWa5h
JOqOcil1d9GQOMGK0SPhoW65Sfwqux4M9CktkNXpElZ5o51dKIK9v06b2+YsSs90
H+xkaSD5H/bEspAR5BlV00Eslemllp2ry08t1752jQvgNgHLdyL+uqaRjvCEEJdg
kcGOXDlScbo4ldMUWqcY2SRM0J7k/BQn9osQTcb78c3IlSykRS/441cJanm855k2
0LDC4pWgHsvRDkJA0HuwpIF6MdA22sZdbe1vEXRoISXubLr5fw2zdaj92BPjrvLy
kU5G2iGncima8bQqRXwcvSdFe6GE5tWKjDHlJucH+d94i+1ihl15rhWWZTrXLS8z
krDJbrSmrJV+tyD0UQieMbYi7gPKw8iNDs2d35mj2ZesHRo5RTPYUL4xPqNRSQUP
3SF5z1mqnzT3vUkBY2Ut4UjUr9UBllUs6rPKe8MEJ7sT8bMgri+QLzft69ffUf2+
ZCnh8Q5W7qzA7v4SfR2+fKuJQDxGpE59VdoEOWUWE7oX45fRH3QKPVwJeDx3YnP7
TquHQIlzz1Nnc207ocha70KT+7874pjXUdP1jJdiQM4aRLzpEYZcX8jvtUl3iLkj
l9wMPBcVAdOrGs0SSG82gRgubkm21D8BeBCst/uvfRrn2k6CMR7o7jLxfnPOHUUw
1v8pKOpEFAj6O9t3S1TZXhvfAfp9fKAY1rkv5RyTakNmG/I5UPJbDzqQ9vO62ha7
7gYJTQ+p7E8a5+nD5o++SuSJCTADnwXQPuObN/4MLqJPvvGW9R/E/mCJL9Ber3/S
LCi1WfArbDh9ZsSEOy5fBndnQbUKP7wUmcQOUrxeIAmj0mp0g797GU9WJQxxZC8V
PNlmTNt4nOnhPr5AUaDX3xzFoy2TJ0JNuIcRU8J4Q24QCTlsfbKi3ryZ5iFWKRRT
XwAdtLffQvqc/zAel15NXyfw6LJRpFGqdBaEMCk/A5y3+SoD7oXCP6bkMpfrPUq7
6zCf9b5wfO0s56z2QgdexNB7L/4SF0wxesvedkP2beeqn4YlO0iXFDP0ip25Rmmw
sBjYhLzZeG3zAr/j1fU624hRZPy1mFVr0jY1pBihZvNxcfGd8PYcs3/M7QNA0TS/
BTGwSCrERjA1Hvn+dprGsSPWvT9gfd13JIbO4S8KrzWoDTuZWqYVfZCDmnr8ia4Q
lWfqERznh3EUGDjVBxJ2cIHrPuRNriE9JvzEV8g1PEkusLjavnculgEKZveARDbE
K3Ysc5UzK2dFDRC212qOQYt4bNS/vRoSrh/8uXSy4kmU+pAskAU+3IGUa1MXbmsA
UnhKDwjrcPZKDg/NEgskSeVgZyQsVWJCRgYf7gUMM1E2kgo+sUSmWNBwlBdNlKQQ
+q/O3KEA6EE/3OWDbDQpgrzKfUpNh7HIZZK1hA1+lx6cIzzJT2SLXZsV12c6mQuw
Fli58upusLqpadX5LGF6p09ESaVGLFxsfgclnllxUsVzgdorMSuPdWQmOKhVmNnC
qfSNeFx+1XCJPRmcunKeHBwJ8FTDzQBqL1LdLSU320sBrR4wYAamVScEEJsRRSk4
rfN+vtej8jC7kV4KpK1d/m0xUrklxVR8rBT94EJOP0Yap0FSVpTJMLppP9oQsC8l
QstBURpvYCDT+w6hU125F3DHnbnZ8dU5FNZ4kqrUA5SSTSuWJ5V+C0Ibv4Wx/p9p
fNlvZfWoDVCkrqZqJtvNh4cCEn+Z6pKfEzC2wTsjuFdZoh14HsKJG/Dja4qU2ZYo
Rl58fTPsaYIMteM76yLBvWfABJ6zr9vfBO1PpkEhPg2NB54T9CkZB5VolwiCFbT6
JZEElU2dZVkPV+baFjhxzQpvThxAATYLD8omwTip/KywTrXz2D8jS1O9lqnkrukJ
waCtQgJR7fAZ+JI/DRMGMgiCME5RRxigbgwkI1fb22/0Y7ow+4vCyaQiUbmFvqmt
P7iYLzKmRbAuPtBW0lmpGbQvvWxG88FxymlmUA+2UnIkkT9ih9iRaCZZeg7/5JW+
+Y71M42iHKu9OhIuJ9+X2fySDAYlFgxqG6FXdrKoPNpyYDcmvOSYCgZ0//wRqDUm
J8fPSeeMXYSY2UaH2orpndhVQrQx2DSPOlSKcGek+sYycPvEr+pjRVZYX1SoGSrO
EFNxHOvAyDyXQzISjbYZJyTQRIQxERaEieUpH+34OVlwcTREeYt4NgMLncrE5PxJ
xJiU+3qyNiFSoLkP6RsnyyF1vRgGJ9TT5u45qmd51qn+HttnM4CqKk/kAC4NFI32
vFJ209pw/nObWEnvq3vLUdrJObST4fftf/2/lNCCqVNbfRChlHSkHNnzuitzm08C
ZBa255Z6FQeF91m4DjF6Rs1KM3Pcs1J/ljeC71VYFcTwR4bs6X4jiQZDQ2q/Itfc
gYb/UECP0tCWWzT6rBA5x5HNXmzH0H94hnNMSdcvs2sNL/Pl6lhqfiGUvjuBmNcP
tG5stZT4kR1XzMGkUULYCJnjIgdOwJvm+r35SqYPvWIC+4p9l5pl0ZW60UGE3H1h
Az765TYP4C6RED8vmqSiFOERH2QPXJmXFr22ePTWKwbsnQXgzTxEG/9orZ2Uf5Ww
nvRUonKXw8RT0uUDraaEiJgjq/KqXwI6a7yKjNFyp3Uo16iaRrcDKTqtomz4PAIH
OYzb+AxiypABFzLyw3SzyFkIG+KMXQUA/7Y7ud18pxBRFd2/F6vaxDwP1Z2sRX5L
zADi5Ssl/MpHGL7F0JUwp9Eaou1vLLMakt+t/Z5I/LRcW5LkTwq/1OXviVSDLKnQ
A1w+1S4hfJxr7ndOiVc1BRM4VgiIbcj67frg34byuR7pGgNB7MV697x6ggX0e/A4
Se6H1Ji5qJXNDNLKyBTLHRSqzr/TkodcHSwj7+KSOIdW6p4cVr3obhvpXSd7F5wa
+5RmHQWgq5QVW/5A50ey5h5MUsmnYL5rJEeWtbCSjNuq4G6m2TMHMAXMaZFliJ6n
NySmC36SRUTf98kNrMo6gGXq5LTBUNGqgKRDvRUbCMOmWqAOakZCQ14Bh6KyLW8p
rHbZaSS5cI4ESDkDRVxUx6i2iLFhe9uC2JRt5XND6CsxPwYyTyFpB3I8x47jHhPN
/xKkLX/1VaOz4W1gZ1uZtzFYTxLkoc/wBqlTyAAt6MXMp17Wjmmyvk00NFjZMCge
LDP4FamVGKQcr+0SR/8G2n60pl0FPhbJD9L8xfmfyqaaPqtyEjatLeqjE4NeLGIM
BmllHVpex2r/B/UZg554IASN/nEKXcIrAgyCYes7R1H4WbjyeTNhccMUoNYVlcoz
HPyx38T0lCzheaEUKErpRBA5hGc/Pxq7zfw0P1cYz4vt0ePSue4+bNcO71BR2wtS
DJSxvlKp+qA/YKXfl8/oNNc9dFAuoXUVZqihT7aMVWsffbLvxFVhjTJ2BWXPmzkX
llOWc9/5ujI/jfEIa6W/ZIqq/blgR1NdIyQth0NazOhXZ+8PXpTcYBtYq0GSnTmf
2qZOHz2rawU+iDuVTtA5BTcT03JcCT+yBUrwfxDA1Qg++pvpvJ5FJw0MJR48S64l
jpnCxTAFPFqW1441tgQYKFSYvDLaJVLpRGedrjjYJSXecVj300NVBf15bjAQ4UbU
ALnqt9XD8w60+qT8Y0FctSn83AoqMD0wAL4/OFPIbFf53pW1UN86GInJSoQ7LVFn
Udxuhx4vq1QHMj1w14W4h0PUyEebWpOINHYEyo3Ad0X5+J1eBKlfJmCCMh2ptEMo
jPIXXVb2b9QoG4pzIMVSu76LFzTypIgAyvMQ6rqg1QAM3aO/5R+9z+tJAmlpcXr1
N0kYDA6McbkY0vIJdrxpPxknxCqt+6ViKhj9CUlHyXOXFiQcL0xute0lYWRI3o3w
agtcAxir0FaaZL6Ta/kG6yGDnQcjyqpJD8abWz3zO/DKBNqVe3kcUNKF4FQbxxHz
t8dlCxpXPcSU+J57pO+fOPKVYQzAKKUme6uXDvn3ht57vJ1lXJ+7SMzyvYRLBwsi
YjBnlNoD/tpWmvQ87Tq0efNTIJqyy1G30PqBDEk9LJ/Pl4CQ3mlI+Fx+W1r6uobx
iL4vd2Kiy4UDe3+xpUUSA6KUfWUg6YtwufEWWTQv8AOOEhwtP1DwYRa+65Gjbt//
Rkjw8YdHRfySCj2lNaEa80qNZy9BT+BW5sT2qvV/t/365TLldYm9APaiebHiriCZ
BtwYkfZtgcAr2NzD2kZvXF+4fIgdusNNPr+sj/o/LBCSS7m6h0201U8NmwO455Kd
zv6EPCbSAV8LTOflP4ZLU3lNM70zKfre1Kmbb+KPrfj9pi5AwTEhaGf9ykX36rad
eBhgJnUqZipgmaottROk4bQbQymiFoFTVDM2WPx8fEdqImbAS5SIGtTAEAHe+inf
aNpN1DaAEjzYaH3RcQ+SRilivT6TANtEA44UwPD+QCAaZgQcMuWiG/OqJOEsSIm0
mfxzsoIQTGa4JYtQoyAg0HdeOFrieZlqwvxFuTYpjIu39IYAND1w1EvmyuX2SiyV
KXx6zlQH6jEtjkHgmkKu0t7mhCGqGjOFGztwmG2ad+vTrkFB1RLuCONRu8/6D7WZ
SZkTLAV8U0iCw3pLtz/wIBXlyawV7T7lGynaa+eea0+6jhS8kfOnChVrj8+6MTHG
t3eScF9J1iSb6SkoVkz5Psw4iukstJHojUAS/0S4Kv/YHY1wAQnwWNPu3dOhCU0f
RhMGi6AEyMnwaOB0g77q5Quo81BP8mkDbfZF6zfTRwq9C7BN7HGtIINaKr6mPcp3
cz3Lx+wX8daKhVjuwfQ8KZHhW8DPDhL/W0rVpOHm6UGq/yTcp/r3N0Gm127fgroY
OFk+qEsZBX//8NV2iSZoLORp3sEPTc7/zCGoVr00GdaXYxjQ5WEwTkuXLIoWiJ7Q
SY+W/arrmmewB4UE5lQJC4x50aeV8xzMXuFZ3BYN12YtjOenrhLEY7SolBcgU8Af
v9eN8q+Z1ItJbD3awRuxtTJlgjBDP9Q1K40H5HnKtBEoesUd9JAY7QZjT7IH2ajD
GfcbpwkqHBhuAPSozKuO/ny2qEN6645RuEPUfFUbK9VS/1WT6tW4kckDMzt9AwWA
R1toffqNeGj8U19of+ZQfw8nPBcnz62BOQB6rthYU3LdLWhcy2+Ee5ZNErgGwqZh
zf9cHNGedTazuKzfL1P4q+Vl2dJv65GiH1d2h/aQbJWl11r6C2tmx5zUhpqYbX0+
1uU/KTyeo38SPSv9BI4YZ4Dc1aHVS6jWWsy+zPajoM5Bfg4fGngTJeV2zar0yVl+
0VdwBmxA9GGS9KZv8G/TwAFltiZrI2GOpkEMfKSM6ZDtZMigoDAXVCv/Uo8DOWDR
apg+5jNb/77KTVSPp3/sovaYb+pkPaSS1RXXWvD3M+TYVblE9vjXl6MCcJDYDMgK
WH7nFjEzsEMSliEy1eHAeQXvTMZzZ9sTYzc5+k74a4COiGV7X9++ryyx2muROOr3
KHSYPFfF1x3eYNbaMGrkcYx0qkzowmELL/6uxiswO1T9iRfyqyaSCGNEKaC0VXiB
IOL5tf4fG2ksOuwZCKwuB+yEFVu4RjLMzTxY9h5YzXKactNyO4Czhbu6NMlFC2wi
6/AExGvoUEWJUJtP+3KCdfzEu9fYPEW9fyVmKFyd6Uhubgq477NVJ0ialkw8rs41
eSseqBd8/ay4NU0Jl1qDh8JbAn/2jMGcMXLBnBSMxSm+KUbj9TLmD7ellqC1sWZY
Hi/Tq2c3HokHWcqBkzGQ9jNxatyZWrcj/3rHH64jvLfboAIzwnreJQPmB1ZnyDBM
kk8M5Bfk68foYq9TvTm6rOAnFaxvuvbbTzHwivkTq+KjBWeiGHpnj7Yw8hO+zvyI
k9QXUEfLkeP5UTiR0XXohXTOXImdOozP6mJ5v8ghp0GqMqoChLIBtb2wrTe/t3UX
AdSEgcCaBZkE+UmdukWE3sCnyOzThy9rmvbKTM2PYXEalwnw1o6NxLi0TvYBzfzj
8OO8T3SC1icDL4DjWIZy1xqui4l9gBoKccSAnzLVudLqx7zq1JXQnYlIw6aC0U0E
YkkvySRFCIpKXWFYyPQAsf4HlLK9HyHwtOXCDa4LZqYpW8O8M2wJWugUKVcNPdRy
aZZQdGjB4zwH6gvYm6uUj3M+nKf9tKlwkCsmFxAT5Oc3+xDUwf4EvJ5/TTsXbAeh
XiKo1AipngK7ummBnHLvoH767S/7Wsd2jSL05II+hso1fxxbvNt//Qq7O0WW70Kj
UI9jN3p50yEQK0ufkchWrZljQlxXO9Kav3TndJA3qN2Vi/KHmKlTEBCwB41bGICz
yjC6gDTMxKznfOpHJbJJeMjNl2yO1qf84iaHs4rchZMUqEMWbIUalBskR3NOu72Q
TJ0xDSFm1PlBoByaq2/cZmdsB4isTGvNBq9bs6tJMRoaIi3rwEsOwO+F0yD3RVs0
/0Y0p7WcoaPtrWv3BC2K2n5A/GP8YXSeH2kOWPVVWkkpX6l0Sy1FUYtoUyag3uWb
3g0MxAQtNE+acaK3iDpqKgZUZUevGnixggeCOE8kyBVzYNlLDav87FjmYfVBNrS2
K+FKLzawKDhyMi5zzC0J9gO1d+IG43bNt69m3TI1QmL7y0ua3TqhIKcGH/VbTn4f
yv2wimJ+YfAiHhYs2D4W+4J1t4rKcsbw8KvOYfYP3nlvqDuHmSGxVfvN+Lx/l6Ii
meo8tZvfwNma8/zvOzFgV2BK5CvoVlIgiSK0K8gftZnYxlkyLDRVNM41b8pCIHUE
xUmhdFpKrnAnKo2LvkOkOuYhvBWg//T0IjRHkDPF3y0/G4cCzQk4sUc8IcbKpz3u
Qh7KV5RPKoJ97NMZVPMUTY/XGnK2v0kJoCiqNTdeuZeTWHtbEJQonTlzpaGJqVmJ
9PKJ5GcQofJl1YIDa+iGoze1+NXUkufNJoHGfqrP6Tw5IZWvjqKW5vf7J7d6Fxrx
QFIlUYGRcTb+lXkWAj1zJFZHSbE1H/lSKbkDE8Ihbkh2fvponW+Kx6GcTFLGOFyW
PTJNwo/L8urBdrVgfRtw9QlJZoMzKTpkirnQ7nnzGtNiYmU6coez6DU1z363R0ua
G9BK0xrB2MoFrV4qorXGQUjfTqK89I+WpSI3uHWUJTKN2ktOsv18WLQeGgkpgu4U
SGgt25wrCbFrK1IXPyoueDxAHDuzMyAUBY3yU0GopLaTUHOwvoVbRw3h26mefShI
OrmekIUHFdB1RnkENWgUaS5B5S/lTTaqUgE17Eb1LgVupXKG5IatuevxY44lj2Zx
uSS+EWHXMmrfZE+lxUX7WSAcMKuu+J15YgpSrghlCjf8sgbhT3VeAyYn4kLPeWzq
vU5K/FUpzrWFvZL0Bn+mssguG1bPFblE0WwuBSX7Qnabh1I6pODu1nqHvMcpORqq
HJ3cIELzbbyfNwzK8jR0AM1kNakmdc0pGO9DBewWyqq8NQuP214Xgpu/XS6K0I57
TF1SIshj2ZGUVDnSUB7NwcV6I7Ch/MciHqNY81Vr05RZ5RDpQJapiIhhPBZYB47f
y0DpEHf+HRiA4In4n1z2YoRdm+ychqJ87XtmboA79LG0QogRJZoCdZs4bV/mtPia
pdHbEG38EOwTHej+GttRiqDWFQnlydXXC1M6PbPqCpNrMpV9xHViI39ZC8oC+gOz
YABGGVoR06QZJBQwGmC5bzeKe5Qtwl2aPqEG2dhTeH9dnys25MxLJuRchQGBeKuN
7U4fKTN40wBKEhxW1+0yHu4+2d59gRZbRayTF9ad1uJLH9lqtvLIxvRfWyLjKX1X
rWDWK3txVEnVEZLdXEhhAKmIcXui1pjdxRb/USvWiHYtyOnz23UFzwhprd1n7Ekf
Vz6PEwuEYpTaM+vkogFT670KrSwU/Z1wqL8Ium1PTqCqz0nMm6Ojr4wZuP/I9X7t
VPsrQc1O7f7xy1lh2B+tBpJ9fyE1nw5d2rmOL6hrzB5aisE7Xcbm7I60r0bMfXUG
SDi+hCfXoI3RvJ0vysjJ4hPO17PhcIGKFzi1LLzPIrrhaHsB4tt+8So1YrgIkQIt
RSnPLSxPBd4EbNyKaudgCxkSiPfDJYKFJByU27xgovYT1hUnN/lj6+4pogLl4wE2
jHJqc0Us84EsDSJqefVXYAu6Cl1M6a/nF3CNTri6bAMDtCqAXHSd81wy7y4DBxF/
kMJo/vqy1WbVXM3agytamsaxWKrSMSBY3SUULfYwNziTyiv9Z1ktwoAkokKhjBdx
We1sJZHMCyZKED7Kzp4sv5cxFoMZl/HzaQQxT75MynsTsZyUWXiewiyORty22e7y
Ye9NwBmY33YPGUwaQkCAfF8ThCD4owjNP4dx0R+hrFWy+2+yW0FkMURf/aDbcpJM
c63btp0i+LxyLLJGyOaInidNql8v8dTVkvSt05nbDWwwhvOhQY9OKcFswIB5YH6Z
s7MxRe2LqVLdojXo90EhyrkP3w5VZ6vTo1Cg7ZejlKzsZq5wzlsFmglw7NbzKZXt
tUelyABmHfRA60KOfAamSn3KSfYEr0drNzZTOAfuGWSE5WZzQ5apT6lc3p9mXVuF
uk7i+f2mZOIACPpErmlZLu2Lnh/Vp1rH22XT2mQvuOzjDYvKaetimC2fG+cIsZTo
UILM7pu9+oOMtpCD6SIJMxM19qONU6Efr4Lu2tvwiG8BWx3WyUIrpnYbka7yi7cH
Rc6PrzHtaMbxG2plSSy1pTtpULDnOSjVloAOLqBx6L7OeqtFjkCtzJD+aMunZAnP
+S4q1T/W1aK3GQl0fFlCBIB16ODIEJC6cJz0hUI2zI396gxP2FIG/vALcMnDz9K1
Cytl2/bRlpMmD0eTPeHl0a02utmRsr8i0UDRGrMBwoD4AT2CM2oEhEL2RVIt+sMF
U3CrGCtfGn2Vqpp+rrP7lFqQzj+P6plw4DD4vRT7BmW3REdJ4BtnrqG2jMbOs6Iz
GBGWwSgqRsRg1aZ9Z4Qcs1bJoA6aEVJK1BNKKFMk+Sxkv5+UcB+u1Kc4StZVtZOj
kcjQDhcaHzEtTOXEv9tQ0NrwO+f5lNKcM6NLVkgVKSlqQbuuGe6Q216bD/KiBP+t
d8F1J07F+x2dikuOUtHfKOC1Hnq78yGeEY04JRbtm899fhWsf6XmGjceT2virodw
n4tti5vmBKSWSQ0wHqxpnBKWAPbiyKEHdoTrOmdE3DVbdTBMvoDu8qYy2qYEdXoZ
vveki0XBsipQX/DcMXG/IFFFa1GQVy8iH4hxivQKsyxbdbf3o8qjg+w8TSbhxO+U
QraFQYCo7wJ8cEYsDXMFE7E1U94YDta6iV+4Q47Vj4xTSDZMP/SBOBfdAGxv5WYM
5fLSkhsA+UFZFYXWotUQUiLqvtaBjIz3Da39NzdD5IvG2tVOA6oKOIs67NSUJjzN
t/wutJv+SpjUfWaowQA0ZP56OwCwF6TTAmnO8g/J8HXD/S/2TcK71E4BWXvvaAfv
eMgf9PjFKcVtNy80o61qasNkvmEeA/ksmiAXRNz57cCCXUakg9POQHUQLckFEpXk
MjFA3UWg0EZnE8vvHx09I/hDhL7TVtZuQwupTy1mo1GyHXjzTfBzjcFF66SIDI1l
AideI4OrzB2fiA9G533nEyikwlRUdcpgBcDhj8rTx2/OmJRGabpUjWQi4C3Y7iFr
IGxesyhhO4I2PfLRsyFWsAsEUUdpRlHPd/mcAsTl5D8UUYS3qHJYDQMp+JyoXM0r
X7xtzMYos9dcfR14ZJCey3SSFyX3fxgWF881Zz1CTCi6XYqp72LPorCXxJe1xa06
1EP7YqOitiEfLeVu7xL1a1aDTKoA9Z+vSSPAUvgSDbV7ECTF0ifrxLbl6U8fWMro
zU+Wj5E2Llm5zUAD2Ei0kKp9s2UEetOtuqkHdWGIV2GLWHP9m2RWZcdPSGftd8m3
lny+v7FFPOxI2c03xZDpysO4adXDvy4s0+Y7/xh7ukAPb9kaUnPnIGWI2JW2ojMv
XSqjWOaVT7RRGyN+UXV2XETooJoMQ5GMoX3u33Uos5+AnkqHSBQsV7kaDUNEwdFT
R+Dfgrs0KWs58wommObfBsonQSun/bmisaIW/G6YneBHnCnxAOnPM0HFzG6tNPyL
82rlE6A/MdYSaLIrD/0KCmT7sIwBxz7plfMC+Dig7lvP5mEmQSZkwwnD404KO/jp
WmlMctVbXkDdjN7tZhbiAor3giIlyaerhqe9mrqyPnuZKxS/5yGmX6xqru0n+hau
JiEsSA38O2QHNewS7HsekUEVRjnXZZYpNGeBD4hrsxi3CAobHphf+zHI2fAbJ34x
MShgTgOnmWIrubXYs3CVNM+jJkkzJL3DyE+CIz090v8Bw6z3TMg7yL6yCE7QQKLt
EsPjk7rDpFx1RC2Nx4crzUVE4qs3v7sN3DB2r1HeYGr+e06vlpYy/y5tj0iiRR2F
kEFA5sfihCbGMqHIBhYMgb9tF5wJcBLs6CPpGh/toOjH7pVNEXSDR6d3366s51pu
1//XM7zXNqYdjTrcga5i6MggG7KZMhqmy1fijSxyv4QA+D+dXni9TynnUeoAcXhl
usRI0d+WxrgAmBEYKVmzrX9IIJd+zpV/v/XhZLI7uWcWyZWjsk6PxFjVl35FPVcB
z+nVHsRaSNw+unlAXIV4FwxSmA/Rv51W7VcohCA2zbyoXKioDlXPtfym6yutky+Y
y+USyurEwtVnKeAoej09+eEKQ+hwm5i2qmxi4KvjuRciIzMrhOW/GUWNy4sEleBl
kWC/LCqoxYbwkZPN7bjHL8rXGQIS2MlAeJszLh77VOglYaRU8Nxo4s1hfn++3IEi
6BOM+QmUu3uL4PmSvQdYH3GWRGxYeJkq3xIBYOa1DozuwDY/hd8J2OFRS46W7tva
9/od23ML8S8RVDRLLiwClHKuzhWf6lde5epkbRlyG1kiVahjeq4tBnkY0SoZu8ar
mwpOqwYTipTJHKR9dBQcQx97/B7EmDHONAvUktu95GLaPc8zPj5Tq/kTEr6JAF0a
+GnC2P2QkiPeh1ZYggUlfQp5PYDvgca93Jspcz6sqkZx2PbyowxXnGmvnx0PgxDJ
fAi7YM/JEG3EhInkjEYQoABoJuGj6pSRByaOuO5mr16YzFN08VwuoH8H8OZFm8Dd
S46GV4gQ1/ovnYjS6fpK4lUf6Ddt99uKHAVFvz1Pmn3E0SkHoES07EEbGm/ogOuR
yAbcCwfdvXXyUkNWyaH+CjhVOId1+jyAMpkq7p7BkmJAPJLEn/ONHRAbvzp4Q5e3
xFNhEJu+kjejusR2bYMGV+DSa4w9eQg93OzNjhFEN7BQ+xXoO1O0IN6jwRnF1FAg
TnA9KB3gOXhqAe0TMWdJbI8hsTpmNhastXKEconhuq7A0tzRY1pyz3Aii+WLNfml
ljsTkgykq2FYn71MAP+rhxqta/5R2jXW6PR8tb/bbQrAhvyALoz0TtYBt5yuHqRy
8GcBveDADftykmeKkfKR3YADtVYU9rtSt2TUts41+/d5mvAcyGaWlKISfipOUJqn
Mf4Q0YXGC7BNfo3tscLb2M5EdwwxxrUba7Y8+c/v6fMZSqOl95hPzD5OUTE75Imw
C7gelrlrxmFUoXD7YNKESjqbaVdshOL5zbw/s8svA1rx3JqBZJNexOxSk36BIY+Z
45/sk1lwLdDYKdcsGPnb5zWnrwM1Obzn032e6q7CBrTBdMH77XBGVL+ScxBohD4f
wI8hK5++EgBSh0yOJtFOKtmZwJl7y/6SLlNxXLe0RePoPgGWawAl4DQRjnnTMBbF
VwIWKWuOJr1crwskKfVsl3ie0kd+XsdeJhg9H76q9El3t0XglfrZW0bzbhbp5XHH
/46vAk9FoDehyMqN8HuT54EX/csh3cEO50rubSbzGkaUBhi/cm4SvWH3lwPDsiE/
rUU7oh5LP/aiNSfSG+KeFS6UiJ3b7rprq5RY/qserBB/OiTqB962UJjZFuid8j2w
PnE45cbVBaZSQUdBJpAYbTfOLNvV1aGkBENFtghZ6PNgoZrzvi9lBcOJIzEjiUCn
9bnkQTx8PdrEoqKIRnIOr5jvMFF1neV3XNiN9W+CG7pf6Ne71lH9bXcFJ0XODXJs
Qpy9s/XtFsd5csG1tvrGNUgvr+iFcwA72o3egGavUsCkXQEFOTx6cA00oMicf0F6
zU6MftEh48IRUv2I/rLdvCDV6i9V5j2bcVF+h6XcVEjJgvLTyRYX6oLX0TdzpvxF
7X0YTX48FF8gE0zluC8cJ7nLioFD1qz390ETccI3HsF4ajVcUotw5BLIgEAQiIEU
y03jhxWBKle/WYdsITLAZ3PjD8cgUY66UGG7Df+gSSB3DOhLdKeOYa5lCckDCfuf
FWfCHF7OBfr5+rzv9J9jp4pFhG+KQqt2mgROiCYQmVEch76ldIUlsJ3I5EBQK1dF
Dwxk/xTRklG8pXBnsX8p7YlU4nIiUKWcBrlAWEPFXRR20jy+v8+dxxS3eOBYlbH4
8lwAsc0np+k0QjTxYQAawm3tXs2ND2td/Krbmyd48134wmPc/yfsBFaM0u1eqFwt
uRVMqpI2XO74RqYGZVdbJI4rwbXZexsnDt1YDHASw3158KYrSihqfLzWbkTTixe7
DNP5dhh4wznrhjf7Y0gFxAmjwY13bd75Jh7iJNM9vrlASfepEf1GXX89Su55ZErx
nWGAtsqpI4zSTOO9z3OL6d/7CntZoBBbK4UnFBZPCA3hfgJ05zfvMgX2RMJKs3zr
Wb9LfSfV/bRlmOklKIa4p+bRL0CWrKrGll4iUkWfgvniQ1lTpvQUdIK7wS/1prQf
J5R9CcWqyqlDNKntBRaQiVqu/tVuc/AWKPm4y7yj7AIfGVgZP/l4SIMLKVRM0R10
kP58gSc4NxbmpDQKhCTgVXFAooxfMj1wtfeqbqBS0uQTD/0sJpPxFBianx/Flg5j
vlMIX+ci2o+wJ+wVTZ3KPKxxC+nQk+WHfhgUGCS60fiBo6H3aR894aEXwCDtknQj
UUAUgT6AQnB+3pP8qYN4VRrMiquasZ9iq+gyA8N1RVrh3VB/G+BL2DR22Dk7Me7Q
Fz7J8X8CrHIWYPU7qWtuVt+yXGa4JelG+We47vkQNyLMLgw+6q4cTlmATh5EMcZH
kMCNSJ8xKfQQCgnHC6SP4Jg0vTPrpJIVyRkf+0JsSbStEkkijnBlKwmfCIvtmMwX
nfJZP/bWzMfg8lYnw1J9ZlNrVk1WK9FAmsIVmniYbxBWWxDDgzpncNhm9s+jl5Cv
bpC34KgMWvMEyjd8t8z5dUrUwweHqhmSVIr0gaxALwx833yMhWDvgxv2C5A4yY2X
6pbc4b4cO56UwWFbt/Oc5e4IuhT7RhUheMcgTP3MopB3cTom5DksTB7qdDFjFutr
a/h3MnadeMBy20agUYTTz0ZAsZJkKo7/+o7o78x9rheOsar/UfxxI1PNWSxvp14m
uSE3bMyvxYful1XigTQORpQiALWWi7Yc8HWdoHlUS2Q3Sb28yyi/yvz5ZkQN7NDI
A0gGn5UTSXpDh+pbiTwHpBsAF2b0dpPs7tqdaLnGIXGYPOMkC+v0D1Ibnuu18sYQ
RQdUNxZ24QD5eROBWocZYAcBBOGD5bi+WLet3Bm5bE7f+kJo/HsMawzZLwjZY9IL
y1ZaiBjERMF4909wamZUPA1nNbfu8KOHhIQaEh8jJdJ/XIa9GD+l/6vunIpYzt3S
awV/pB5SCj5XkwH0jHnhEwl4sSwe+C3vA//sj5Vxwu6yLrFFm/x6n8kswBsNGmix
Eyfdq6I0hgWZe5/HUBlPkizuV4M+Sij21F3pTieMub10fTO6V2yIXCvcsqjPF30e
qskmUtKlcG1JrrqbYgCcfYmQtvo337Pm4tEveKuqZzqYgowEh5GIt4r0wp4eZZjJ
SdskvuU8piOuiPrx4ZrIbucX3fTYUe8aAjkUjscce7zFZozLR0lFYULf9cCaRfeI
kOrGNBbVTNCtWfOWXXrQn7rQqN0SMj1tss5LASKtrT1arXsNsmKyawF5QT3GwG5X
2ubFyE21DkfgZzAoUwGyxW60GmWiQ98K+Um2BPALqd8Xcs1kl6VxowKTYcmi61p6
hHPpHgsQOHHFqQMGRfaF+OcQMa3wTRX1pgSh+UR3SwItPm9aHBeyYtHG9+KT2ZC2
WA6zBH6gE/pFji0fN2MQzxRSK3t4zJEWrzmsebDb6/rOpCujmVBv8EsXsCkdA//4
GiOCuPOfEeVWiwIjTNROgdXJ/wENOpO/ySTxnG4li2qQ1mNrgYA7ubjXVtkgLSkq
NhnmgZ9088v9/44bc1erOTqfOCF8Uo1eg9036MIOcqWIFuWfSfB+6LVzGvappckd
16qu2kUNikbkLS+V418A4bFQowc7qYz9xVerhgtrcR0B4ay+DWJrhs6rxekxHaJ/
vGYPWY1UPtA5eWV1pWfoz0BO6ejPZAiG3o5jaTU3y7xKEpDsIxZHZggT3fkDlurG
oj3BCRv5p2Og6Vn9XMnpfNIpxI6YO4c6T/Wh5LGZuf0qTDDJVaRAzeVZO2jU9yR9
G2yFLIf6aryqyGJdoFn538tU9gRFtbvSJlaXjzDuq2gLh8bIhD8eEMzCA/wIZLP9
oWYJYn56ZVFEEkocXbsU+l4TSX7wcx3XfcGLEZH5ZFACMihL6dSTJ2qobDmVDBB0
VTvXPKb1BT+6UI0p/IuBmk9+qD8c6GF2gpnViC6Gw1NSK25vgyn1Yre5hTvekj8k
JWZBKn77xUtPLu5jXkjkWFgRCCH7O1aZwl8zZwvKw11oQwfCKmw6fQb80dZG6iqc
Z+/mvsuvT9TmI2W08er/GpJL4QC7p5tYgGfClqoALDawvm5Fl23uYpeqwwgBowHO
CjgI676CWUpKhdiCLJpfFwm2Pcm4bsLVqgf4MYgq3qg9XBLylZ42zvoEjGmNs8MO
SLRiH9ABuQF9H+rabo9Ha0Y1M6O1n0R+fP0XPw2/fQbv0+18A2KXQ7aH2tEvHT9J
7RLFiNy+0kVG2W8F/66qFf7Simr2OTX9Czn512hnvI/vlgbiaS8v9KrmMazXsyTX
97Q7b769gNCB+j+P4tdVJ4OVIU4W8NFC+Hyf/cpR2pMYD9NMpYK2BGrHNwiRoVum
7SP0Tj7mnTFVGK6l/7MQHeMGNmYvl20thB6+mFR/hH1GrIxsmd+oPg7ZAsxzC0LE
QgKW83Fbjn5rWSYxyotZfEhCP8tpYbjkTkrhwQtMZROSe+OpxrugSNRWBz1/wpQv
5FXX3aa24JFM0aRtjH9J/H/GhQs+nQLqdaOIxCNsbUyHG4p4skZD2fqN3Obu5hsZ
5IpiPZqFnzqYapyruyIrptStsEHSHhlKjwzpaviKLnslj0UCrYvzukzl/5xr+sBr
fi4bp+mzUmsERaVmM9burAKHw/pJsmDBPgw/fX1s8aQ2+/ZXwchIefXlp+wxbBeW
ocDME9z3DQq2keSzrosgQEZTjIGHaBKj66rKHsJMw13TZatgkY92dQQVDYvA3S9h
QNZ9LfpoxtoENAygMmRvpBn1piZdQ+AEPo54j4pXJgcnl15g2Z30e1NvCuRelxSz
pH4bCwy8TM8cU1IDArLeF8oO70pXJ3WBs7SZ1OQz8O1GtrtE5pMEHKCxqJa+P//C
xawwTh/WgJViU8EeEgA03hagUQWgleNPgenj+QPVgSbki1MQXSymhEbjGuPO3c2s
4y+ayqU2ZDL6lSPaIk88AcLl/Vq+8fksBY8qSYC/sjbW+dDOnKUpYdlTKLgKCIwp
h+8aD8AAp19AGiaIb0m8G3Z98zeiZTuYZFK6QkmSiq7LFvRmoxxoIyILKbAJ1M8V
aMj+9kYGpYmUseP93P/1TTFTMGE3Q4SoERb3pyhwRS8db5TnV4OuZK09oFPXbYp+
PJad+VZsSCENqc81iDnKw1oltQAy9CQxx772y5oILHOBcVYSOc18HC2g0uukRsXX
cCYG0m8RHdKimZsLgQS6Y7TTKF7ii/+KrE+F9NiQaotcRgHt6m3dUBztBCXoU4kx
hvb76bCVxxfckQUneKVFi3KVlTI65ED4p/PORkK/uFMiVWDpDelPfh8txZmNmsHS
RGHQnWOqmyvT55BMh3RXjg/UYlqpFXFls//PJC/tvQ1n83K/P1US0comI4F7h/eY
3GPnCuynXfDB+nbU3FyIeo+MG5eOy1zJIOod0OaVlnnC8Gvk3uut1AXyzR8fnrMY
fDP3X8NxqCKIFRNDpEat3EXOVfhLAXE8RT0DLZFjPNY5yoRwrVy6xsHQPozdBX4L
M0QlHJGGLKweaKIHZWlOBnjDo1FcOKQ0ae1bfEC97pc8XmeGNwpDNlhNgCLHMPrG
SNUpHiP7rJwv/N9JM31OGKpewtqI3L4xNIuDolc3E6XNJdEl7SH2eZq8hTrsl31k
NOxTQJdxsuXG1lI7CTdSNFkCpXO7B+HUs+C2Oh2PgUCFXAY6B29zEKad9eWoHwA1
QtKgJa7RLH3OHutLAp7fCaeYJWPTi7o+hs13ymZms6iHjS8ZXIUYrWN4iTj/fFwU
yvpJFVSL1lWXc28WI9fcGkpaniHIzElazMWKeR/6RDQlBIMqZ4WIgdmyFhyQFf7T
gqO9DwPCQ+ozblJTsT05yDv2203b2rvZ/Fu7En1NtZ3Tg0Dy94Rb+NJ8Y77NR+ct
ZTaAywEsu2/oFcpg7nfJA1NsVo1Re2PiSn0YRdRgJAYW7OgpwmM4cl/203V7xe/J
+OYn7de/LJBGZhBRshCrcERa4pmMyN3aqgM2MYfqjn1mnVtRzk+QQn7NXcZ2sngu
6bYiV23bj73DDSeJg3jbL5Uk3M/zK3h/mFx/Edo2blSAdZatPEVkDxgB/PgaLOva
nypRSFRFMYwgFZ6hu4gt7iAacqw+hby7NZQ+KiM4e/k7aNdx9vqd5UFc1LEP13em
ddgP7XLFnarxPO2Te/2GyWM2WZgQg2neUfzYVlK3C6POP1dxRd77VpJrbZGWuitM
q0kKq3tJF+UNMM+dbFe00aM5wKNZDFj8K3EBriVrKwFNi5AmIf6H6mVQX3O90UaN
uA8gP9klEmQuofLzNFB+eFlVNrp0o47sFxQj4voxf+Mg7qLQjnypRWWEJzlPia21
IMMQJjuxMTeGxeR2Wjjdw/0i52UxehXaTFY8Acqv5iwiwtZHer9JBcmDpRqTr+68
M5OOuuMCfaZYhfK0zxGjoKuRmJbE+SAaMBXwc5zf+GSRU1BCCfy73Enz8wtFpkol
pyZSXOOiE2llk1vB635cItbXkTQ94G8p0rv2crCHbc3nNwW+V15wFZ/0nuhK34q7
mOkUOfMVlz7FJfTCFRodpxsaOZneAjJ0g5IZBtIJuNEgmP39qNEL1kPchwo6/XLt
z8IhFUHWaN43A7uRRD5zucrTvUKmUu2wUExg6JTcHzuelIpqmOni7iUSaYF7jGb3
70F3wZhMS4f5aD7PbAhZvNiU96PeOcTMY0Ngpv4bPskfbNAqBDH8cLH+697vEaxQ
UbaOovmLPvAU0eCJmIn8relXb+JdhvuydHKCNPuEks8tALfIofGedmkMO6nHlLS1
xPdKVdWpqfStAQRsOWA2ZUwG7z+gZnWoViyJbs+0KStX2kVvvBkqB82z4zjETV1P
O6Q/geAYQEA/j6fKFhzNApeJw8n2yG74NYAf/Zn6EDh810jdRf8xARc2ATjH+PYH
Fhft3bU1mvjxUo0azRqrxwnAv7cfe8I74D5R4N7rYodMUUq9qlLTQ9EBMYV0DECU
DZq9uRNse+QVhECRAQOV9AlDk2TGbxfA2iXfwsrJzjKEWfSl/9sloCxqraNOmfyw
grbha/ve7noZLLBV1y7q5pUuj58Zjk8cTo5J6C8WBsPsDZN0HJModWKt25XRM/dJ
+81kmuHXM/3rGsdpkXDu6UpWbOy80htQW7C3ypdRbq++YDJWE/qJbXa/D6Xyoc5m
UtkPi3VoDFVRN2LHhSxQMrkZ5OYRXU5CK33Fbgtd0lpIKdjA31HC4ehKOtLIH09N
SNAM+lYWJJXO8dnwAi8AkXU4p9EQmSrTqF0J/E3jW53abnpGO72pqqKpd9nMt4Iu
DGCnN9YwQNsx59x5ULNJITqXa4RhZhC9iONE9x+8u5iQreMHm/4MS3NQvpuAPvqJ
GBXwrGCFflI/KzJFlwA2eIZCNWDeMk9jnfiv4Qlts34e2pZ2pcEMMaClEp2mY3HH
/SMnQy4IeyJuSOkzPLMllWF5QAJLRLCEueV8ofSBzvFtCrM9Wv0D3+SliIKejoeb
8EeODC4SUe1bZN7BiRhBlndcI0cS3JUeI4vtAjIF0blmz4bxdpTnl/tZAW1DTx6A
zUNzKCbTWSGUE97Y9ptgZv5BpwWQVEJGDrd4vNcE2IoNRPaMzJJavG6mywcxLVf6
kIu5McQOl1D9mPRQ3x4usvC521clKfLpyzK20ah5mrk08mwClTqz90NIDBjThgrX
MkleqIxzgDxr0oAr/6D3+K/doAu0rxRl6q+JC4NG4u03+gooB/81sCJNmhJSUYis
FI+YHOEB0cDr28J5kF6dgrg4qbSqVICRYkkUerL27vOkosqv4nAFcCtIgNyhBjPR
Mb9vlG/gdY1EL/Ts/98LVEsMXiRKWAdLfSo/whmYaZoPxFxUwAJI072EAPPoxLoL
dcxZGMpyxvxbJ4Lb+nGemXcyN1HnIsdYWgHRdypcZez4M2KUiTihAswxNr5QJ6bC
BSZ49/VAJRYi6TZ30OIkAvBCLLauXWyFi3gqpVdnL7DVeQIpSXU+YkwzXn/O2Enq
Ag67LmHdO6adlQcy/EfRv/SFQl3Mi8JkjfQgKt1cwD0goPnBDuWJnzYXN23YEB+D
ij7i/qXQiJlQcxm9eEUCV+lAIBtIQ6Dhdinbm8inSmQ1p+tVGXFLGai/txvXz32B
if9JFsY1qUego3zgTSVNFRryFcH4vC5GKv1/SVKNXTQJ95u8szK5CV04ogIC5gKa
Ex8JjPho8EC0oBXtQ2p4syE6cXUkrasIAMhdtGYKE4ZRPzCyWUNXyxrsK1Xngx6B
ZdJeGd9Vb874FvJAch7HFlOBVkYvTvQPMfOTqCc/BLnOKRqFI8uxM9f8xM+g/gNX
Ymuiz4dcryde7fb/KotbpyNUTQWjUJVgIYdwgxMwp7Q+vaCBi7HsXfj7833FMCfJ
Sf3BJmA5uE+Jyh6z8LQkAFrF5r4xaT8ODpT39V/Q1QoWNOG4yzvT1HEzMdCvN7Ed
bqz12lh3wzGPN8IK47nahyljX7IaBrQB+SJjnpz/v5QwaYY32JFlPF3HI5OPdeCy
LjK0CCvhHSJ9yAoe5w1X+vraR6+tJ4DMk4wWONypZHbTsHX1S2ejxgXZBAK1aRLt
VgEW23WKP6PUKc5uwZR4E/ycAlJlrZ2mnqW+WNzPTab5U/1BN/sOvuC1XOfeKjjq
doJndNcbY5ImyMCaO3EpMUdWdcsiJIbUT6/UqQDw6l45Daz+X+neTpmLScvLhR6j
Ltihj1O0q3tWXYZp7Lk6Zc9vqQwgt5xVzpIp63X5Uuad4PaFWIYRe0ZTMwr6umn4
OBfIVx6p7rF44yZAQ2P7R49dibyFgfWf0LBcAswVxndzRRNtO36uariEt7Jmpo1D
G2aarPoNs9RQkdzPGI+NfXT1rF6iNL+McQeiGizPrBY+YrAKKJhfxu/8MeV3YKDl
N+e/RZ27RLu3/yu3+lItyuqGD0klyF5eGvftjOFQjHiP5LkHbVMdVACL73DaI7RO
Ws9jko/hQCV/vX/J8dOUPsx+fdnmgvckAOPo0Dfcsayynsn/giup3vwA2vwpUDQ5
4ASkSEsaQ27WfCwA7wyGfCou7uRTQ9Ky6TyZqtzFrFgtwt6kg+lRekowz5zo3c0d
AHGB3D+8881rpeeGg+W/S46I2tV63QRUQ0BDh6gmKke87ydiBD+Q8iNfne5R0f59
v5jicnzbNKxihiitNbRgsI2rOezI0xwoU5DpW2lQ+CjRJSbsI3O/SsgQTAOwr8gE
2IoIP02wWA+tQxqZA3XUyeJQhpv72CmWy5GvmyrpNM+YzzM2qdZouTXgjwgF2jC4
Yoz3+Fjpq3XrlNU6eizP5BTcxl1ARqb2BLuPuV+1ZniCV9pdHtMBkerhjJ2kXb8y
U1ZK8U+mEhrjB8Jo47ZyK5feJR5bv4aRBoqJ2A2Q/dNfcEYot/eLpeM8zjlBplKN
zvnlUWaspJ/vlZRnfgyvK9oDu+C1xczFF2InTseEv+PNcpMMXXxGVHoVjjfpayli
Hk7pKF2rVkaMqQTbOqPDr7+U3XVrTRf+MbjNxwhoNXYn0XTJ7dgib4a9L+evw0mf
iYR9bLXm4wscqL9GmOX9BecWJK+Pe5+w52KzSyDRyv4YGUyxosTf2cSDGrMoC6CI
JcIaRN6Guzv5CGmLwwP/O0CKaNHsS7hgPPA2p46bCql1/qPNl4BuLsrlNNwmqDH8
7SdRTDeQAnkST2xFU9EonjC1UO4ZXLmb8aAQR/xE7LX7V00dpamfaAuy3v5w6Zth
Oo8oYaOgXBs1Bdlcs2QPsBvN+J/lacdDU1NSv5n56xV8s2LMMo5Dhfye1OgFoslC
UGTQAAZrQhd08fEII8zBrtR7OQqsfy+4p/F+T9EwCsBugFCyNLHsFH3ZMJR+GQAz
Dqieb/gT/g0stcqpm0U3U0ZQXD9yCOA8DAxs2kolb8nKYenpVam9K82QjBgli5XI
kZFjlY1i380YgFu0yOyQ3+qYln2dHKNEgb8pWDPmwFE184lWlcRO8zZLeRyKjhLU
erZWiV0B0W++LT0Z986rrzP3tz0Pz3+zYKcPmv83bHi689vljuu5Ezw6ZwZTEMeP
X6cr+VzfGMq3DwXbhg+Ge89HdXJijfqfeDoajeUFaNlwnKzycECkMtGFjsXLsIc8
tNPCtl0EiTESnItccz12n/cIrC6K3G1tql7nmbYC14+TYGN25M+Y1o89hc0t5FlL
xG5AAdlAAmopp9EC8n56r0FTlzR4OteWVwlagDWfm5svUD//hlsrCo6Xn4EP7R5S
8q/bu0PEpA5l/tokxFKEBTHJLFzuoXWUncGXBe2u0GjJDIf8dUY9wH7cRiEc3VtD
gJBs+xksFrJKvd1tKih50Dbfgu8TnyLJJb5QTLUkkvPilQzliByVjUQkgfLUOnHc
lDNDnWAckRieD8HgFJVtaAWUWFPsA6OMWMry9On8snXpxMHeLtFdC+oaOjSlkSs6
x46qG/jauPmgGrorMJSprCKWorxKqlSeceJlx0kOi+APflNsFwfYvEaQao2K0/M6
43CXNsp7Jph9MpyvSTd2KNS0G4PKFtVGXswmo12GHM3hNaym98nHE1hQAVTwEKcP
ZsH8D2XIcDHwDEehY2qW55FX0AbZJHanCxb3AFpLZsHz7C2DxsqYl9qLq3jUTwwc
5l99bnZddiuA7NEQTAZ+3O6yvdh0O2sfJzBLqSzEeUNPO8xT50O2D7HmUgEL2cd/
ldKFozwyJIJpZtRvpKkS9+pi0na+gXepuyYrotleh5EP3Bzq7qyncMXpa8Py8rjD
U3bc6vqyAzdYuPjt834ecmNiZVeAFVGJfNPdPku1b04YOEKDooYPfm0rjYoNlvem
R15cFCf+Oo8YXToibpFAZY/GP21jG2/a16PcyAs0MKTR+YnLR3fUP4XaP47Zw8FC
hvIYJbzHQpRPF4917if7vkS7vjqU42SfD69Ko6HVbD+oeN/UiLXGRl7M1xnQZ37W
JeQqyxAoOVvH5c32SKu/CMwd+dGi2Al2tQ867R56PGVcjJsrGd+useuJAqnKEaGM
FG8320ZOEej3uI/Ie3FzX5dL7XK/zIA4Y96vGdiFTZTx1JdhfFTrcqKbXqO9REFL
xvBuYBnxXKKX76Ea6MabwtV5iFVlDSJ238xOSBg9XovfozGJOANZov6emMzKnZ/6
iQH36LGK6J1vKPof+z2557AyptyhyI2y8xZspK2bSX/wxmz6XRpv4mS7CBXH9w6y
BcUWZ/1Q/yGecoKrDNSkU0SDCfKS+QrP6TubrF/doR4Jodq9ChLMFJSWriz6psiT
ISeiOg+XvEU/mL1jUi4OBjJmBfIjFbmZ3DNeb4fnGvwPKk92flOTlHR4nBwm3jMy
WC2ha2lSc7UsRVdbqAfPUnbVpyyPy8IJ6OTIK+m42iXt6GZ5P9FlV7614bb9sABk
lsMsfMW9lLO6dFQfQJwz6+G8zIUSHIsKT0pnFuo9up/+FFlCZ5JavY8s+yI5qEDH
AtxIcJTq3Mjrp+uDvn8N7wBcbn4plvFiO1KW31uKo8LiqNJ+UFC6GopGhscJSanN
Y3NUE5VChgrG2SZE0NLXdrnZnwJodVKSH0G9aiuAoVIhqziuioynuHEO0lBVHa+K
wrRgqVcjdeTUHgtK9AjCnPiVpkjn3AOAKBDqFw5LuqcO2aLp40XomN8bL63UE4y1
KAcSCUmlm246sZ6iHBJZZy8eF5CtNJWCoNFEKP26fZExbbxGMBpstjQUyNlu5q2I
hb8p2UjFPYHyPS6+ov0kcee5V+BO2panAanT+Qg3rtZZubZ96tSFAk00rGhFv5Vh
PtsNUCNpuUm5qPVCCix9Nl0w4uC+DRnDQZSJCjf7bEFRquXwP/x+ulU/WdN5C0QW
mtd47fcCggIGk0CWveM3I01xmfcyqRlJGzI/dA+wkiYk1qonxNtwOjlUfzhUJ6nb
RztnLOmBK385RgbAOXhrtDtJ53qhoEuqXL/nqlkOcBuV4nQeV4V4akuhUL8EFhOR
ZJFywuLiBlqTdfAIQVBLfnRLNyhM5rs1kzJL5TfUED4X2DhDrCZoBRd3vlQy/sgU
QVeDOP2J2FlXXSZT8uHMUwjuEtTVaB95ovoAih+I4SFeYvn/pQmqL5hxHNvdV7ZG
jKoZd+pJX5Xtew9nXf31Bk17oDsN7L5ajPntQEmkp1JBz2xoQVYFr7yUmMu4bSG/
DKgoN9G5UGI1Jmzz1XrFdGV0g6JkBCvH5H7rltvfmf8UCd4W4/bwb01ruY3B7C6K
iTiol1Qt5Q376YEcEAiky31eW7178samSmi51egCPPuCAZ5oC6a+GgoXUAyY1nxw
rT6wH5VuAtSj7iySNhNGSqvY3oyFs42pIgMO8MU5uNZZ2zwvqlRrzA7m8UKJt0cE
kH4MZG9yono6OuMutkUteg2HQ9LHhyc6TPtK8pmJ6oN0WKWb8V11GVbCh20cXAhc
L3YCrBAh/GC9VXuXt8luiQyjsapEzfb0QBu00EcwyUE1OnsC92UDd7uBalu5qqh4
GRzkA27Jcqr1ZBMHSMWktkZLzMQoVnd6a4UwdiEjMdeKye+MFhG1uP0IqVAvhMao
wcnimDQ6Be3crjb4cgA5W4ubtS6n7+0Qk+J1NA043PDKcpUroMEht1hDmIAjSg9p
dfisgtygmPwTUiIRo59YEyKpofRJ0GogcvYYO9YbhPCUkYGOfZxPs+b2Lb6j4OJX
5hyi8JrjK2tbIt0uLy4Es8LbErEoEjl1tdewvfY3gofXtLqqqKIwApvs/6CsnM5Y
T3C/GW6N/4yefhSFpOHq4zucYFeiF29PkDDm8fj+MmX/2FeYFq8CUCaU8kMEIAHh
F9T80xNgWWZl+1dqcHAQIMwapIkl+pWQolcVUuIiab+Sl6JtqM1NO0/2B476axcj
xNvBxDPL6+x9iJrl+0MD6P3n1IBxxhoiGc2+1zwjsQUPws5Np5f8f2iCR1tgFXUA
eKERAtIBlAGDE6Rrg3MjFqAlewZy3f+xeKKr6MSb1TkaIVnZbiQI2KS7E0Vavfgo
mjnAd374muho/EDod0ddmhBfWl/Ia8IivUvafR//VSZyNZBz8LD6djNi58DL1Nez
1rC9vGhZhaCjva9S5gkJJAoQqNs0+Gxwtu8ECZbntcx3JrLl9ohTvSOoG7AVPtVl
fMn4wcIEGgjBfLz9KAv/k6JIYPmD/S4ls4TUqUpa00WbQ45TicnucRyHMkmH5Qaz
pdf2KLrL41jVCdSmwMtIibfj5z7HGQckShDpcsEfAR6fuwbO6vCecmDFHMoaUKWu
Km9d5xxC7RXLKixpCUyOxsuhYN5bUR75KX4VWsORwh5mczHOKvMa/hM4StsB0qz4
AF2CWysx3AjG3TFc7w/AVzCHtKsfyCuJRKUia8EeRDSmNQfCZOCJHsMMsX1I3xpj
GE6MHCqjvZDoJMH034j9GgV6eSQnPct3VJ3MVlJ+KR4ApMk3VMbCgRJ2x9LNPMaT
s5knQpmsuq3SpjRSO0wbwDjglou/TYxeBNcoUQ93oYw5PB4QoK726c3Umu+2R8O0
2bjRRYBpErN4TEO6CC+DHZ2imIPz0/4wfMgou8Y1Z/aW18S81FK7M2KDzcYhsyZK
ihweJ1c+mIxwj9LhJioE4cPgvErKynjs+lmr/an33x8zc88+12ehV13DKHGok+Wd
ydVDdtnw2IevXsgfleQgi8BLgDp78DSl1RBdJQUATRrnKQ9NOBo9CQXp6UZNT6aw
wpY+CMNzjE1LemIsDE7m7K/Ddwo2xgbosoi7KFt1S/8ERj+4kQPvzrpoIJ+VRK4D
acYk32COfi5xQIRs5jSpjWhjMZve6CiK4vRhV6IK8rTb8FZwyAPWc2RGrnipXOGq
r/dYfdzwCEV56+DGpWrRGDuniIP6S1DfLufXNjuqwixOHaUsTOUOFuNJS55LAYYR
Rr/cLuzYYngol3pFIQB5iR+m0Ow3SXMe2bi+VMt1kqbECSdd0jBIrk//UOnPtJL+
eaTmvNJiNCdbJK+Wt74w7YJaRSZRCJqxV46aKuKe6R/ME7B44SFGmGBumXhI4Vky
mKHBWgG3gP64/wc+eZi7IIxPEtWreUhUMQXqpZLrFre7elZWYpBiiF3sGzK0DTju
AinyhVMLynlcO3/D0fFaWKQE/EyaXZVUV0hy/a9UmD6a8u9rNcDa7WU3nLBnPGTP
JYIHvOaQHfYd1PICbdhLBBGHI6kdGhrwD6fx4J4/3EcOoyov9+W3BHErtTHZfHkt
AxF+cI3dvzM1lJJxrcqDPVJISpRsjAPhDqh6Bqe3UuBRkr8gJPaYwYjwUiFBhQcO
xLf8KhI3bW6+1SHLgUtkRiWFezYUe2zfKpANPFDQM1n6B529prS/uus0IS0FQyXB
YmaFulwkZWRPaujD8ci5aDe0A0dToU3Ka54o1wm+mhskOWMEZeGpIPsApahQmxUn
foA5gnnmyxy8gmJzpxwSxLhevSS6/WHXOnvMycAsMJYVWNIzKqcQhXCMe5isef6K
p6hK6WyrYqMduo/b3Uv8UQW389vC80fpTObDOhtCX76qcoB3oOd1vASxbtA4edJs
LonauvAX+BQSTEyo9wVYMq91cA7/XIkvQsFXmx4nPsarKz5FF4ek+I11EDoZkxUD
eE99JrkcW93F5AlRMznwi+URzGRmbuAVhDHrXdwRdCPwr7I9d0XgtCEG0ZTrvKKy
otsh+hSzb9tRWNx1fD8luuTAJ4ujj8JrLBjfzRToOLEbBRqEyNzvwPfKtADwq/7T
P4iSrW+28CaLRv5U3zkGWRM4UB//308X8XU1BjClQgiPTG+GGWU7ftTRVE4MaA64
LVzRSMiefziOG3R4a1c7ahSxl4eDnYo+59VjQ8TXmLCtqMBR2lvTuLbQRSjiW+VA
UlXdzBRkrYmcKCIF7Zyedi/ifSOpadOw7mWLLjQF2E4pXWpgQP4ajQn9Bj/g8/i1
Fb+1FxEo9brc/f9tTPve/QWiOpl4OntcRd8Fc80q/IVyZxhhmSpeJhy+TseQjKFU
oq59yDVPCcSQ6dWLr4YCzu2bgyO0FPJaFM8RBTobUe/l84hKOmp4zAuya1hqbkms
+GDhduIgEf0zNmPhK6SBiLuzr77FD0S6YcEGXodr4PRri6JyMb+rnphi8JIZIUSR
EK5VvdyiPQSjMTqD2amCzbeYXDhjXqF1g3Cel5+rY8Hz7HdZ5xKpvYfoP8InByEf
HNUVmFdav1YVC5KcDjMskbnX9vG0hzuSt3LsHHRpoH+AVHEaYWvfalQ/2F7bKqsE
utknJjC+0D0j77m92Bvxa75f1pHFpXAOt4n5esxlaq+bAAhRg1WweQ19W+7TvVdV
OMW1qRgxo9KGFE2X6vwBm8Tu3yvRJ2sSz5NhBQrK+jWobI71RYsDDESchvwfm7dX
TwbfgvfxNlyv8SlP8kih/W6t1/xlHv40ShAKo0gQn7BUyNEELwjRUp0/8Bt4gb6B
YF53eADOJ6D0+h1jrcf1o8zrXsAIycAzIz9TLxFyVaFuemY61zPHVZKx3tO40pzm
zrnq0kFLn1KvxyS1q9JMGJFNo8j773Ld5KBANz4P4nVbeKC7mxfmBoQM7zOnagRQ
4weYAVzTKyiy1wlHt08H7NXgOW8kJV9kr/OoIIHxWI5+vtfdi4Ei0eFBnbR23z/c
fVZ8S2lxh/U8S3eKQ3JARBl50PHc8Irt7avW8/6L5YcGNOUlipSjDS7W87scg2xR
sEbNXIapCAkne57nZ3uiCsBJpJLCSBIM3iP6fIEBKUy1rxNgLQoqjEzDhvKM0fx0
CgIuqJAYng/1fMhxTYN3C+GYygzq5wWIwbg/qBPWiHu863RCARkGiY3zP0dvSEDy
6af4OKX7XlOfPl1DUnvd74rR3ngWVyqQvWM8ONKR9EjpUpGQGW9SR1a4QKl1/h8+
EuLX4YtQCJgEmn0XizKd6DCsY966HrJ2D0qfYLXz6oU2fCf5iQ6HWCh/oeHEWy8B
PMdTXtId7FTastUhjvE02laww8Xauo+hhES3K1DTvG8w309xyz+k6RIJdUPSx8+n
pnJ4BqlkVg/gvztr+HqTBkacIzjAlmAasD+lAiHh1GH4yuK4CZxTB8qbMDHVk9WH
EgwRF+ZMnvOIbI0fNgAyjh1b0wGlsGgZrpakyN+NDbwfJIGB42oZSIsZpfvlN4+V
BL8z8XhGzTgoXF77Xkkki+onEkIXpyOhVXzO/IQggxFv0Y7FF1DeNBemjIqkws6s
P8r/rSSeOiDAHrJL/mIUdZ4Eo0JsGKO5pJKO6Up6HfoaZEBPBFKXeG4xq1gHGnOi
VirU3LyKo6EsL2FbEnPqMUEcBMCksuKnHNgw7r6NqDRFUx6PVJ9Ak0jctHNIYWpa
bx1/MdTKIuIkeerPB+MnD34bqllUVgtZZOJVkVk9ICuxVKqV8DnFMbCLmLoAUMTK
oUr3YWMGCwkNvVe69i/SiqweExU6VirytJ17Eqh7SyYkGqa9Pj/abnl6LYrfXcl2
Lfj+tDulB4CoX/Jc0Wb7kG2jn1Uf5JrqSozTz8q2lZiEzgiFgaaBE258GB0BsINZ
/+1Oig6LQIfCFw9b04KJfiSymKAcWfMYmJ5S44knWmTPu61vJ02HOtLoabny133o
0e6H2/KKTzlOxJvg6zRJbZYbB8hByHAO99mmq3cwoEEXnQXBw6DKsCgzisU+TMyF
pGhnz/ncPh+P5iTUcKQ32PxTCNdPuMKJo6yH/mh26rRMbit63YvLWdQvzWcuypC0
Uyg0Uhmp+FwyIae1wdAK+lOAi6rqPt1hDn3TsR/cPi5AIv19ssfvkVO1NsOnfOiP
2rYfmL7OqCTI5zDD5s+5QxVtZOQ3UZyUwet1/PGdnDLOrUmbNTuCAAg5gkUDQTU9
SN60ujCI5nCOVhyPoEBi0dw0Xgsi+6AGisCoateVMdo0Q7hnU6yuE7M/K+X1+V84
fVZYocsKziYH1yqG9mCRSN4O+RagCrheCE6v6JlTeBEITraZcgHIfbheyCtjkjGt
NXjpvTy4qG5q7kHLW3VKDZitKozA5KmPLbOlqpwiR5lhAU+KkX3n+JDnwwhDev7l
p2a4pMbOjSqYSz8GUKgOWMP4b/r8uD7dzCMgPlY7ruNUUoD2umMrWbqah8eBuxJp
1sKinyMwVo8jqRKrw6kb8O99l5B9sKAFMhE4PVUvQyWMpNcdG+WkzoTSZ4JRgfXT
woWYZP6niDg3envRo9mAn+KGBKuTf0mLMxqrXKo8nW8NFfw4mbDXes+i1S4/Zxkd
DGCvyROGKX9dUQU+WYm+YJba55MfCh50Uj3RAu6fOH75GPHM0ti0cy9HK1b64Ndn
hjiL2Fce7OigfRxI8nVJUTYPRAJhO9SQH5tFFR9HiH/RcSA/ip6K4HNt7U72k3ea
SAdIGCERciQD2F5hVcvw2s08YJG1XdpAs6Qp7o5EH+tbe9n9GiIhzD7T3h2ZZuKR
YMt+RYmkONBu8mzjd8SFDy5Y6UTn4usi4P+IoBlIaE24cjwc2RIahLUtxjogecHU
hpAcvBiCJis+AcIFVQ1+qUG2j9Dv//5WMXDFN/0EZMf84N5VN7LQLZGm60JDZ0+O
1zhaf3Tx0dbVgOHbMvv9KqK7R9cILK/8qQMRYvLoRNKbZt6502PD8rydzpZV2vOn
znfa74Wtbn2LdC20yzmmTKASrMXub/BtcbkS+dK35kXUehAr6hSdGiG6XVq5XCmr
axbI7M44/SLZOo0gYcmnn8qqeqU0iXcGhulOZ29XBCaExY/AIQwTPb0/uyMHZA0w
N6alCwikOSXNr//2gbpYVKiTAuScOqhf6IHjW2GkPViQG7oApd5+pCvq1sR0/VBJ
CXfXPhw75Yfsw+QUSyhi0nZDtjX4PjCrufwcMMZHqGx14tgH+lQuQDbFII8pmOK6
ZYPocBu/rvCppDbk4jGTVCChX4z8TVzr67oh+rMTKW59TAR22HLyF4lXmsINI5yV
D6Y5zRuwGYk9ly72pGsouadzUeFO/3yNd/Z9kTC1w44kqXfVPGk1zzzEMDsSwlaf
pCOGOtQptoA9NMMDgKL5UgBh4eAWG8wAD2GocgkXCvBvv0nCbOWYv5sEoe7pPFGy
LPzFDTKZryzf5nOnznLmOJOed4oHXa1CcJqp4UOKzbl0HApoAY4xBqiH2jceTTUO
zemOw2khokyVSL/BuNs8oOBuObTpdHvIFh24Hn8E7HhneHj9HZVlpVOFfTlBFRvT
sv4jwMyjrJCplSqsyWRYSG/lxO3RCSd5y+rsBmh/uOI603o2YzkJYNlVlFz8wCHk
Qqd2Zkm3R+BFHvHTFXXrP0xkRdZu0gGbbCRX3h2gxyvt700bWuLTsq7ZDGmyYzu2
049f24ft9nGbNLsCNnTtVzWaxmilJO+2+M/nyHnySYGY5u2FxCUKmq4LCSeTrptk
P42L/imCCyMpoUHfJFFxSmevraPqk3V3KbaDadsSuFBJoslTVmD4KJ++yXTFbAq0
XPLXMqfQiAoLDZ3ut9Rs2cD1XKDOZ5TOAOU66HafJL8QtsqBLye/5ooPDdgRNzw8
ucCH+5ul3M98NqaDHFWJhyk8rPP4fZaX1yyhRK5ZqmTJZKb8jy6aJULErE/cYFwt
fNCel0z+F7e98RkkpvCAgMZOlOUTR1Zz0FdyJ6lQb2PU7hk2WM3J7vU5P5uKmks2
SCmN18k3Av4mq0nifiB6SbckBC13Swz5cFGvKq/bl4/+0HtHNJlPrcbNTZwnBoJf
Gvz12vlXewGI42Wq25eQuXyzoWaOdSR+NfRSiJtLXPF4RXgwk2Hj6d5MsKFTccGk
41MpljfxwoU/w5P2w5kLtXT/r/0pQhVqmpylmTaZXQxAI/7rN2MiNjmTMInGzDdd
xE8O1XDbCGkVU5s+Q7du3LKbwFRWchoVIx9Q/mWN+aPg4oJyTkKtRTQBfxwbMd94
Nwn6UiXqk37cx89jMqwsib0MuVeLhdAeBXrhhFbzJvOqdj2ntKyXCI3LM0WpJ5ni
ADjv2NLtLsC65UVhvjc779Vv3wSUT7hvDlXb6htA9cll86E0SuTthis4W5WcPjLb
DjLL37SneRrVymXtMjZUuJ/AJdVFoQ6J7NiKjjgP+nerT7R7ngfT8G/5pt3NRvpu
8Zz/mGnZGjbyWn/JCjqYjLRbkhM/C1FK0+bau+yMowWsIjTcMBDuNk4iCs6wgNmW
CkT5k0BwA4HJF5Ghhm1aItmPCd1/xYMZRj8mXgQHdyCx9lgv55mC8jaDpW1jvrHw
m81ViSXLuBaheX8EjHn9UgqCms5uo4r24V+sE95/1M8JnkFVW3gEsCU49xeV+3Gf
SHdvrBtplDEBcpS8NnBWU9gEsnGVNr6kk6dw91j0s8x5X1h57u74TCpw61rjjTxO
1vtEuRKqfneF+j4jCjI3SRXQLABk98Qks5mvvbocqaYlin3+KseJ+FxA4wDbr0In
oqJraNjLqAWQRmBRZaRBBqy9SR5zlsTDMW5kKWzj7p3tomByp29ZWl+J22osTCeN
oXmhPCeweF01ah9UB7vqU9cEY+LBVXsFE9QcUcMwRmEHVAn7nrAwTqD/fX7m27W/
M4jspYTWVKTK6yautlGKKUFpjwm7+SaCnyDPVpCzRe5ivVDsIZnB4UOTHwuVYHu5
NHZrPF0TaDUpIFnOzTurctEpQdSAMTsM4fYYyUtK6BPtp+pKpknBtyCEVHrQ8IdI
AE1j9khpDGCn+xqyat7+/uQATrhD5KVxHhUls5x5CtzC9aZmTA3VZZxppoeRgd0K
sHrh/8L1HPj+bFQpRyrOkTih0LYsw1behto3ndj/jSua85x3iyM3VSko6kT4srAr
FJ0k/G3bvC6LQf/YDgxqQqTpVnsNn/ergogXkTiOj6YoX/1SUC8Ku8h9kkJrle5r
5wcBLO6J2HyioOT8XDJFrIP8Z79nLIwEKreArHaVg4d00DttBUDhJnGI4yF+jwMi
vleuGSaL5jrpSGQ1+eYmghvLvReoq/nXMOQdpwZaxwuHO+pUYbH38fMgYNOad9zF
aD5dhX0S3NNN/tESRGcj+kmfzMfWdPziosIivR/Csg/R/Km9xY4gzTF+cO6x7Bgn
wjST/EgghFrtV9/cnjAqrQ3YuB098V+zvI6Rl9k7aCQrSySxuwQ/4x+VQHI/LDqK
IJOmi4nlimuleJkoaZXcfFes4wUpIhdoVMW94G1caEOwEAq8q+gv1VLnPrGX7/wK
FAdwYfmH7qFBBmejrVRFqSGXc+0zS5DVdjoUMUCnWG4yitnHOIYZa2IkcGI5bJPB
PplcmHPonzxjtSteChBlUKwu8M5+jZMsRKnjnks8kvfUnybnul78g7Y69S9yEYZf
XHGaS/jnj8qP+TsytigGykIN8nl3nsMnwAPp/GpkDj3nM5PofxtRwnqMlzET+heW
tAEY3eBK8NzKDUrYX64jDrl1gWcy8/cQxWBYQwHtpE2+mpkWsD0Kx/kNKBBfx+Ci
9Xf+1q2XW06Y65oAITIuTla15/C9pt1m6TYdM7Tsa/jUg0+a5MPsIBa/m37SAwwy
jJ4ffbd3hV4U6cy8O3O4HF+2in34U2cHRZcvpKUquVXmZSLGum6+WfwXv57K1du+
i/irVBucPCmVAucGo5q0WiCpWWthtG76k4wQCSxXocIMAkmuuQ6N/g+PnD3gf+rW
20kWlqqISaqCjFNe6ObTXKx8Sm4EsyBa0lxAheTM1Das43RklCo4iCt74w9HTNX/
pBJARlnKbtTWR3eUnxi8+zfXPZhpjBfrJyX1gABS0p5MTG8DRC9Kt2f3zrgKDPvX
TprzieB8CLsfYvL9MQXDfsLIX5ojExEVedXbNhMOqHt3+h7qFmznq5ZUkVEYFJXv
i5MQlKP6iuiPTqrKS+Ipyjr+cpry13KUEBuuMJBwscbQOsI7+MSrcC6fZT0IzmKH
w9CHjI2gM+i/w6OuPIV3/t1/571ZKC9ObG4AMqQrHJdu6TwlbjOVyiFD2dsgqx7m
NUAGwO+k6QHJhIQWXZFhZY3zpUurVr146OspSn6ZEsADLXJqLJTjBzY4xJa8c0Re
wqkDkbvuowFW79CdknX0IitmCswjrtWDAhkZOhI78JEMz+g+e7s0PfIfJ89Ot1Je
F9Wo4/olE3thCWAIg+TnKCkXgjb8FBr/2QQfCjCVnzu+8muN4jBl+CZsw2hCJXeR
MiJWHz6/suEKcpDPpEe4/LKW+5yXaJUylfrS2h73n3wTSx8cCMuavjQEGUmfmoL5
Z0E2RCUOAppbuJc5K3iMQMODvpIeNUx5bHPIix/L+4RDmhyhOaS7KLo34Y6cJSC5
PNSdURTcGLcZEkfFS9kJEnoxx5+BVGsjWcLwqIwt2IkNggMIU++qOm7mxb/khHsu
2cqCY99+oe0t2AjiHLwphdf4ALvGgOa4khts6IquDDE+yASe7iB/I8rSxbX3mgtd
HDoANge1pWqo4PoIrOhWIfqH64+bi1z8Q2BJcQV0jrx3jkZLIXUQfdWxFymf71hU
m738fWWIaH2PzjsxB5ryuIH2q/lZagVcYGwdpkAsEb+HA+zj8VcMudyLWshg76lz
S/Cw3Ra6N9XGabHorF4rActIXI/rzSIbfbAGXrzBjz7CmhDABbr0PnVFYj0jsnoE
pULFdGy3WonFqteQSY2jPsYIeWibOl/ZJ3245sVPbxwEDsa0GBgyDYcnXh5Vx3In
Kz7JahUutJ9NHcCcrkAz6SWCUTZxIduHNut/VRWHXbz4zlJ1vmJ0D4Y3nLnIuCJW
QqLmb+4M9IAm4XEV6Q4xZuYzSD9MpKFjPJjxXFsbiaY8+0mznsqyW0CcmVMSrwtn
uQuekbIaW7QjHCsIVI0H3v1y/nRFDyHDP6p/RsOWWZYhoZ7dWn1hDuvLxkpqkOj9
KpPwaqH3sAvqMABugSIN74gvkFcVpH43kF3nx010jjuqbwcZu51a1GGkCwfrKoRy
uVGhhfotmBPABz7xaEjor9FGp1QVEgoTDE0ci1hEei8ZXTxyKF61MJtc8fneGvze
AqYeK2fiZAiBM7zVUMT4ZO5PTM5Z1c40BdO/A9eFwsnfTjx6aRiHZXiln44U+nwM
hi9J4gAX1r0qha533ZEnlsYPGbipk/8DTQIqEdakdzzM71LWoSCzJAxom7kQIvbG
o9Tus01iJY+saZGeLReX9y/PNb6zVeRETof9jf6I3A0IOhnTLoUjdwkmAV2BA9A8
WNy8UE8kanAyYxvv8ef+3Wfhq+GUST/yOgzyYocuxu14fVUfNw8x8phdeDSKBH/G
AoYl0qiSvbCvbyXlyfhW0VQN7CpKshIcyJqlA9Ky0K8OecUX5tBH3H8zvcxSnWuJ
BCLIIoGkVyDqLwgunW5KMZHvrc7/+3xwxuhx1EwpxpYe02xljozn3anRT0KefUi2
EZ9+q1apHg8mikpD7/1RozFeld9ZwLQG6b6t4a5VIJlQ8GtucrVpwbDHDQHKhpUu
lZPebmbHdOvDsiJZHG0zul1959KCoVXY2Kv/bz4aiKF+MVbjYG5w4190HsHBUN96
yrAAK/sRPyCLu9t8srsccnML4XS5Cn5cNbtKjcLlyU4ajGbDzSCXXni85cOddd2N
2y4hjyBG7EJ/kVypN8EQ0Qj6/qqQUKIt+Dxbp6NTXjIsjL5O3606k89SlHwfM47Y
MIoACShTc01V/q66vrueF72vJDsS7xNef7OMhRVZTOI/HzOgO6yXL8F+0GtY54hU
3WLolz9WWs9VbciLzIDOrm6q63nd390nO5NtNAYYaS93cyR0Md1kN3bDUGDYIz2/
7hyeEQFGA1E4CqMO94U8mNRjgvCPmQ4YwF7omcNL0XT3cBtSUPifECs0DsdE/zDJ
tbyImn3lmgnr4Mrq1e1MxQ0hMopIPlcjtOlPK7X7888QjvaG2zfJIsBX1OkC9Yd4
MGg7Xr6E8Cr4TP2gqdgV7JAoMxxOT85/c3kt6F0KhJ8eYe29dG8e19neodw4h4qR
tL058LQ81FVciNkfhYB4ER0K6RuxJMZkmzqYTwUibms0yXFGMBWcpvuwRwTIMD7r
g6TWFuxNQSY6ASuPppjGWn/gSUSxglE7mYtIAwKZRjaktroRl9JkslSJDM3jMxEx
O+0dpopVgRovEQv/UxT/Dx5AZiPgbW1Kcsh3+b/XCGhfPOLb8yOipxB98qvMo/Lg
mqSjwmo0AAD/zSWDHjX7XOIOVJivfWbaQieCw/hhDT2zedLbgARJuHeqahf1NhcX
bT9AXr95t2msfvxhSpq0s7sflmq2VWma2LBOrZrm/F+L9N8tzZJZKl+0wpGtxsgU
1SqEvXZWnjRE1SsIHs9nczQ2lxw6NfdifbwCh3obx6zzzVoiZ2X5/rqvAxsu6Wb3
1hgQ+vJcULrGUZJQMgqTEe6eoaZGkiyAn1RrumSXPOS12xOX6QID5r+SXsCN8i9p
83BttxCcRrdb1MlqiidHpm+WLCRcMSRt9Py+l/vYLpRBKQTJgLk8n33BU5Fpj2yM
LizyB9K9BnUcaQwAhHScHj4i7a0u/6ybIGPybDrWlmFE4d5uMsq8IOCN5PtYC7OM
ADvNaeTu6e36KUplZJjcpxfK9itRWZ/suoAx3ZqSbxwjaJVmFibY3ry7k/7zJTin
52Sg21Ry7HlbRb/mMFzX6/9WwfHlA43AluheU696e5ExEiEmU43pdiJN8w1vQWbl
5q1oEJz3oxvqRO1gvKJQgyQUMwmFOx4Cp7cI2CT6XD2xhaIvMcqhOnLuPCQ6I4DC
Ls2+FKn8W+oVo4r6SlLI4JNMGq6WnoiNU/9Y+dt654VUXburkWYBhwWI1KL2UyJG
giREn93T3AM4JAri2LyqgQMsIQrrvGvOpV4MN4x2ixhJxEjZCPHVmKrn/Zbbuk/9
zPZZtH5lgAfrk1ZF4eHHQA4YvxMaLXUCvvj/CQIjRtoviGU07nUJTTB4uedDZvU2
AlDju/isnNpl4HqXyHvsRXEBPJ732eukl/3Ht9JKPZmg1CGwgNWfSqrnvjq/x1rG
kfyk5huTbkqByxBkIj4UWWzUzrwngzGajHmg0RMnPtz2JMBb0kpA0PgoyYOIE1CO
/sfOMOZQzwfplqAcgfKMPZMVm40CGqhODZn0FJCzvHVxv8J1jvwDFDfDwZmeJK/D
73OHYLCVawoA1SXzYlQmIGCj3tawm15uIdubhpmlcfA+qjnEAsjW3f4/DmhViufa
U22fvtngciutF2l5Lnt2dzrFSqRcwFdUr7lcYjfnrfesb+n0WE2KMbyq46QV+qUU
UVCY/WTS8wPJABusQf15s38ZcTlZjLTzBEsR7Nb4D+sZOfYGVsaL4PrkiwoDrjDr
OQu09POvYUvpXVUDLg1Kk5vhNoqe4qMtWHo8FOtSE+4unHktSAXDVrQTIFXTKtst
kR+OI7gNwAomjd7IPbBocU1A0b4Li0delLc0dbd9S1zjBazSljM978Tx09kgXpJp
OpNxrHvuBiNm294nAISXfyM4uuPWo8Vtglshe3BCC0xWL6mS4w+1XhiRTvAq8VCb
h+A0yz7lpYmT/RUiyuOXHztL+DYjGGrEnXeryZPfzPQMIDlboUnKEJTtAdE/oh5C
PEP+yYGzTlErtnyO8SsQiK8ipuQddCIrASzh0yGNmH7CIfe1maMXGuiZioab39N0
dts+j2+PkdOqi3jMMLVzVKtsLG9+0TUFFF3UVYtdqfaBOlwNExb3WKPePFGyPnTT
gWMwBabbpD2mHp1kiZZfumpb9aZxdbkiDi7BAFOzZvW6qXD5cPubvFszt5HQCLU5
atJFMJEmIbV211EyJtjXl97lPrMNh4PoHTXlHcfOxw0xsC0f5qFWSVG62c5zsOMQ
RKxziRUJYKPM9LGIfW2V4gh2PkyJf2/V86UFs19a8PscF38tsbq6p3qNVmdcCHpz
mKMBGqACE5KhrPa3I1Ihs1XB72T4VKlw7OzfzHBo7YB3EykGVJd/oa4zYme+Xt6O
vs/0nZRdqaJ4kvXha+W04hr/J46vpPiuPMazolHHMdtbGyJD/Ozc3Sn5UKK139Rj
gGaVf0L1iitB/vf96EPEfSpVSRfymDfzDel/R2+jED7rzy3mBfHv/c/258FCY6+g
snfVehvTznZpDVRomSQR0hxarLhJpo/5IDmOjDFEpyhiol2l4hqT07vSbYJriX8H
k73hCAJVx8acTk81PBLs9V2HK3ZGJTMOvB/BduODUQ7Uz9R6W9dBvB7Hfc7mB/x9
Nik0GgHBlO8zcInMZYC3dwTVEcc5CtZFbUYtBwueeOGNMjg7/UtqRrOJ/wDZtfjA
ODaJz/pzq0cZpB4ISfd1nMRNDVwjDWfVO75tQTjQy+mIPMHjyl+VTcg7Cl9i9TB6
X9rOwj/OUIOlfTmMO2h6bDoMMz4u1zMdodT4tJryguq2fTkBa71Hc0RsLtve0V8w
lJ7VCw2Xc1Ti87fGSXWKbbvjwBSMtC1nFfrwp46PY76jxn+9ot8dcrq6nMAjjlqW
hH6bV6WgM+MCtFw7zou8Uunh7Dcpu+NBNpMQUYlfEXX6xTVOfS7hcApWdy9ODi+b
h0DGDv6AAFsKqRXOnByv56I3kg8Hu274v+7BPGdCF1yjTiQvuoqkHjr8GB2Sikqc
iRHAx2MPqPK1VfGDxSfPC9DSEz2i75HNRDn4pkqUVPi5vXR9OZwXaCGf3xjI2a5v
TjUje0qfLoYhexNp4Vj6Cwt2Eua2FY4ntYVwT203HNv7YOafNswXWHtW8FR2YuhI
UJ58vqtvcdYV33GXWmwV/KtoPbK4qFPZX+qeizz4FysFvt8ljwqKkXcRxN1T0HhS
xgu/mvB/wF/A93zj+ov1Zxo1m1u+ue9xghKGCkm4l3cNezci9cfV6j2CRWChiIxy
SdKdLrvGfLlNjSicw2/2aKn9DTfNfhg1XjuslfG8KOnglr6KMYVlU7NBsbvICHqh
Gkm3j6pLDHGAavLNLao/daOApw5oKeRn6X6p6If0vzdppAS3U7STq0x+GHNMyi70
q2CfwZNoPMN1jQYJzAwe2tjjr/6bVBxRIc1Rl2zM335OXLHg/Q2duL4LB9HCmLze
pZfgs653j+o1tfjQHe1Q25uuziqzr6WpgypjEoTTlwpRAG0+1drFaCYnxVST7Qqu
VDR8s8CJ0wg7cWLT88zD4NHrSqE+et2kuU54o6CUSIZslWq/AKQ0ZsLUmwNoKJ3n
GahsoAh9LmMATBw18f9HrLVT7T3prrnQASTg1cLuKVjOk/Ij5Yb3C8DSsLAgKo93
SF3t+R7o+dh7Sk0gzeOvZl38vI4uqhswnoDytw9SpWG3iZSeVdt1e2zujMnLVTQF
zrkXOnJHd6zHFUDaBkyKMDrBLgJyilN9sf/ur1fiZgXi46un1Im79lqGZvpoYfLb
PjJVqHv1Y9nzzbOoY1gfP6Ueib1KcldLuJOVyfDmNXZEJQrMFX3tQ0WAEu8E7lbw
nRCW048c9yLJ1Ro10EtgLziTtTO8sHTz5x/ZyvjJ3rxEM6OPK4mpGnx1Ldvc6SW2
gQboClCJOx0qjwBbUokGIntaHW1eC58j6gqMmmn2vO98UBp35mN7GfusZpElac6O
vxyLavrbCUOPLjE8CKusd/Llhy65kTCfmnP0bkE1Cqt/UlVfNYEBO6Olb5Fx8yYc
abvZuXUNTFiu5HaPLDuH5rUnBiZhPP7nXPhdCfuT2c9lzO/KAdJa8x0Zwylhz4Ji
899W5gkeEW4+zxXlDnsaXi1f4XomTwVkvXzlDvp5AfRqMhmlgfgaUBw8nkyml+iY
8G8rc3oWzt3Nj3EdaoOsvw+VoM0O+s9UvWj5mdvUo6H3t2vFZO2QNgl8+2xVzJDV
l4zvUHNEqdihhjZknW+xlYiSB872hZXWLBk0KM5Wuh/eHr6BEL9RTHB6FBtRl/oc
XZODE1Qtm+xpyJ0Q3RjcVG+hibNegr/YVqQdA7/gGAxrFJG+0JaOIqkoWflCVCKg
to0C1kIdXldXWqx0Zbf8hsuLw0sXCgCE6CO3K3B3nKU2o2yxEAky7j+mZcGe1Ggw
7BtGmt4S4+urrbBmOgWPNIoDwtsQKKlIVh+BCtnE3R5SSJILCdNDsdxatLkXxbzP
sbD3zwif9HXG+HMLPBqjLrKppiB7kWutQig1YAtR+rHh0xnsSJys8v2ra/9jTFuj
xeAWL2amNC9uJe8c13MSI5lz65EhYuLZ9GlunJhC9kNCv1uPOdIkCJuIQVyn8cpN
69s2nowQRwprXuSpqOYrnN5jA73Ak4XoNu4LOV4Q4bPx8+oCwNXCguXxmGncFDgg
Hk4Sc6v0zRraJ1m45KIynKKtdO5KKqjQdXEfl+/N+g+gshfSv3uxYiHYvkps7yPC
WSXGgENBWRzNv4w5qkt1lxrS4vcR6Zk0YEbojf5ykgX4UQDv2WZ0xabOhmfzRuIA
nwzngwM+a4P00WTipY71Q08nrw0Plv+ZvT7/SOBRkMlz/3fsAMf+pP4mXZ+vQ7Dh
cNgEpao3T00gJQUIk+5zUoCesSr80fZsa+PCS5ak5CIEqRadSbMmfewaCSJ5Eh2d
XYR31T40zgo1D58aQQPiGu4LrthdyoJllGepUtmjOIjaf3rCAwXFEm2RFFlQWYfe
fgAjbr0SFnfzgankMcT6QUW2p9Vc99DqwYmaB8y0LgTPFGn3HsJT3uEqffJqMvgR
5PlKAQvYrPdnDMMZfjKPyaS+8soND0JyDxaxTtNJfa4oElRdAAijVLe39eUaPqQb
ju2K8mzNqS8U1H2WVHnTOimFcq7RI2IYGwF3HwIuI5l6csodVt5MZPuB7uQY5So8
iSgN9aLkRNLYOuFLIVUZXpBuV5PWM4nP6dQrJa/3/18AV/nIzpAsIG78ggKaPmx0
LBcvVUTqoJDJbuOM/1jg+62WsW1MzBtYmAnk9/RYtL6ojhLAkohSNdAXGcRIeBX5
9pqUwKz8iL40dgMHEpOaarpYXUEEM9OZLKahhbFj51bOoubZpmrknZkA2w/Y1P+j
zFYo+KcxRD8SZ9jzzYernaJbV/IeZye3DE3Jlersk2/tOqRKebB9RuJBpqBLqdZJ
Q0dqyVJOqyFHgIDSphRNQ69XiHudPhuCfdJX56AgT235Ei9bEYtf9q8m/MJzOW/i
id23MfL7o0Toreh+U77tQ8S3awqxPtErYc8OsXRkEwGXgE8h0d7dYxqGw7RjWUiV
qws9TBRPiVoaXwCh/LTtDy6TRXSqp+hdq1vrBfXilIfKSbVk/d/3ctWMg/jvi6Fh
+6wJtccsavFwCc2n0UihqZT4Zs6KgI3BCqtN6ZLGWqbcPPOGYQw9gnyRlY/56Mrv
zXNlcTuX/nz2fZ/j/p/Ulom2va0Ea/rGnp9vvOzcSZns/z88FnmkhljNDRMbvMs/
HgP5MpjISLeIY0UFzn4dT8A6GeGLd4FRaCtwxRv2xkvd01WwybfFQlDb2ZYLnexF
B7PUCZDyUeAC+7P3WB1EJ2H+SlF858CFNfHsqJ+MBB3dwj1QWVcCCyZcuMuNzItL
6kmGHcHWrP8jUwT+8Zy6YypJy5pHMXerXylZ66Wj2sda0/bw2FI8jutuWt86oSIk
S0bRcA+z740UnWvvW4H1bwJ7DtXnFrQaJqmhfkWkw4ywYvpOv5XOJg5dMqMM7ZE+
afSXNVyVzXI7HeGcVZPtya5TUEijgX39gYPKwX3ORb8waOvzJD5D6r1DIOl5MUQQ
yHarDSUPCCpbEs9rXZwh0iMolupMykFcwUtR7bQhUqG2bBMQDqvATZ/3FQUhbs/U
PglELM2Cp/GXk1TldUvWgZTM2go9sWcJSQLklYwl3qsCYpDB5nyRlg/OiNkVHObx
+JEHwkVAMRTAZ7Cx/zO1p5Pf9rslmCSqG8x0hRFksb2YgjS2eRYw+FLGq6t5DFmh
eklEjCe2EJ2N/Tk7FoHjwbKN+aZ92KQbAVtb3OsY+aYHa5OKXqJBBuEPVL88wziy
x0MVaM+IDH0fYcMEBawif2jG5gKFMFXHDvcVvsSxtF3lTIHdbVsx6S9g2n9dA0I/
xuZTHlQ4LiPqIjKg7aB1FsrNGWCDiCuhjqWerfF2QVYY+GWfLUZLk7LxBSmVJ5qh
UXQ+k1Nq5WPwt+zknt5pR+9x4cpP+Nw72xkTZjUtoCng0p/T5m8IGedS8sDologo
iQ4yog0RtEA+Gv8CrCLmoUbDe3tlT5AfOBc0/oUNDNz7pGu4eyIOlHo+8tYYlgF1
uuQTfP0XPshcpTS25myzc0PmOygEwjlDKMizgaGWAH7ufOLoPZM2p7RyzDjlvzFq
79LAbVtKIh1o3cveeNq9lciLg1HT519itYs2uMnSAZRHoLUJUzwcr+zmmKYRbzzD
ppu56GaXuOtgIwZalVgQrv+jRKzXFoiCfZV6pRjsgLbP/hvYtz8rrJHm/AThmEss
9EfMr6VfL2YvtKLMLMyqOLuaMKwQcPwrd+71xVBqa+ZFVEtniK4Ev+kwOE2Ag/k6
G6EYfcHdKnYspohkyTRk2BX15irlvRQiOQIs1DBEvBbpmAOFgWXHKjXHyqmvBkzc
ArkZBugduV+RKvq30vgLKX0AmV7STc2+ZEF81WzlJRT3wrX5zOHBmHolHtu3bTBP
fRJrb8a7icneOtSGghbqfUXcovOVmnEti4BOUflTthhEyuo/MIIDy8vPDOkBDvuf
YUiLO3xuPWeLE3wp97gNQaSP5RGPaXHKtczUKN+jJpm/Eu9e+jnGhds6K/QKw2bx
E6PIsdGGlIVq9jXp/c6DAwTRoniZZ2/IN2+00Rj606+elDSTYyZPxNBpj/ZYayYx
zHdaqHGjF5Kg7YMtqD4OqVfQrwVfvIkCECuDjCnUMyeys99UnbRX22EcCzWwPE93
jTUyhFaQGBzp9vBkiVAGNzb3uBDuFLy/GStFVq68xe826JezGvg+TWfO+g35i3iN
XMCvy5givV7XKG/kQ7zCrDlD5TOg3rTVG5ct/sqeJZZzqOdwIVXl/xtJhXpf+2lc
bfzzPdM4zg6cTdyVnJ89A0CnL9uHQ62jd8nLwOBESzHIik/DRXixMMTZHhHvAUCd
QvCGlfBr3soCxcXWCW1BdvC2Bh5FhDxH4BhboGoOEHMtt67lB9zI0zBejJPDVJHK
dUC/pD9Paf5krj2aPTy7ic5sldGI8mrSehqUeoNTf6HEUKm1h8RvaWkD4WiBkau1
t7DTk5GQT54J48rVPf0fMYZQfJ389cpHWkpJm3PWsufGaAE8Fs4syS3ip0IN16NS
naEOyRshJf2CL+K4rZ8GtaubM7vwwZNiLC7Rd22EvislhbAd3N/umFI3RzKbbeSB
0uMMqqBv+apNp2Dk6+7DfK1U6ZWt+9Snr8JdDuyudsjsIwH7DHgUBIMwVpUgbQSs
TJzksOIh4WHZ0GmynJ5Zd8KU2FtLrhKIUpOXvtFWF2u0hTUJpJhC3J10F2qvrWGk
GJriD/z7EK8ijVpx57hmqqSXr1NR/EQjVxSv6X0XE5cqdyRRkw1G4CQ+1QZhmJHz
PjKoqkmevjYkNnQxRpXwKc25M1H53WClOYz1/2g2T1ngjMlCW4+mO8JnmZrH82tS
t1aYoVmKXA0Pm0UNhjarOXYMVr+q88A2MM6Cp4xWADHNsv+HrFmFDSVLhlt2v2Ih
7mnhwVYrt91hmeHzK8tYGQrwg3B2ptdI8J2J2007ZyeDEz7XM1YUAHrJw5YcfNMC
Lsx1qBvoRieA0rI44Gpk+Crnkn7OQ/943VvsvlvfrGqVQtA4KipeURscU164qFpU
1w6gGgp/F26rdJHpF3q3w5H+dlB59mMWNNhGt9CP0BPIT7hNU93uDe8r+BgnfLod
Pm9PYJqUHmvQXbqga2KR0jDeVgVev70Kz6vi7F+s1BTmvR4KpiahQ53wt7pjCcSO
9YKl+zqhcNTaKxNBSH/vrra6qHk57TgZw8I01GrfSe3tMtX7Eoh5b499hzT79FTD
FErmEWuecRblgFxJfEwV7A+f4NdHR3Ew6++tGfayTMbY/99qoQz8R1M120iCIiF2
dITxmHEDvKr+7jhviO1OYsEA8i+jrITygmFg+PUIq8Yeu0dxz28gueAXGuQ0jPiQ
FY1c9vqDCyhmegOSNLvIOE6d9YAFkxZA8qmVUoMPQGocyShqVz3jrM9RTgUvnAIm
fQz/YNP07X5zAo2tUix2GOXciUUGG+NYiIBeq7U7ju4bAPvKCoarUcfcLyXi+3BC
cf5i8p7WxelxDLeyfUaEzoluRr3sR88RyU6pbHcUgdyuhxKJZa1ZZ+6iabOWGK9G
U+zhdUUrOKuYpey+OcZTPsbcWaR5n4ZLCWSVDPW49YgjjDkuUcNpi3wqeoqWTFE5
dojWCA4oG8bgc5TQehwEMRu9oRq+u/5Ypzt7t0rg7Nayv4roxKhkOzEM7cBIwtMo
EDB+wUE+qkTpTtbELUTFGOtIIYkMZeSJ522SPA//VziXXjCqg5YqWdP45q/ssomQ
9p242qHpY7FjQA4/rwRMK0n5C5/za3nt6jbSBVqbhWEIsekzSRedzVMX3f45C+Zc
d4HIRUrxlMr9dwJ2d+XYCjeGvmDa/gtnRiyFbTJSvBH3UxOFVOteRRa3zwtmHboA
lxuEslA1K1NLyVzUCQCQCcqa1mzU5cGicUaa5AgO9cIsipoclp2UvgV+Kji7ddKn
DWbXdHF55hSZfEhsfiHCVt//gjKypTRWamgnxXCI/tlSGBC+E3iywiVP9NeLhGmJ
MhC2zTVcXJLx+E5o8HTb8zB/xxgYqhiSWxSgcmfZ/t4JEfE39vvV4D438Gp83BLn
vpPM17rjWuS7wcYcGg1DJ/SX2ZoJrrQvRqyZQorn71Z6qqyqitsXK1Odwjgp4gSD
e8McNSjuKqybLGTGx9sPeh3+9K8O8XCf1ztwVBfTpMavIlgjaZH2pfMyk2xitsGc
B2vNIcwF3eLDLzdNdoecrcRQMH40jkZYTEj7JnhzQUL3X3n1cdBJF2R/G/Jz0qmy
Qyw9BZVhCupPLsW2lcIhqfLm2Gs2flqXgMvd9TOaSul0osVA6ib7v+ATwxGaQr38
lWre0wHIkmdjZbgs8qN7tziyAjEwP6OdfMEJ2mnxKweQgtbGvUunc6zJgmnW5Wxe
Fy3wgFGKsQyBMiFgG8uA4zYpv7VaBkchiZlLR9FltxmwrW9iCBzQJwhEqnW3ImSp
B9BwsMsqtZsg4VMIFiqwHaMlmlUglPcttP795SxT9WRadvxi8leuZcG+YPl+nyhh
c4VJc9KtR8jJYHinEaTTGnfmrC0xTrKT47H4m875M16x8Es6/g8tGxdEqcYQaOhs
bJtdEejYFm/oZxzKX5zgKiX8Sl+DZ0AkKQl3xvVMlbas/JPScxwXl0YSUnFh5v5R
xMt4Zukd7L6Ky16uZpY9z7Rp4Mu73GU9qbcLAVdThj3IS9J1VowiPOfTHk09euTk
Ofm/lXfzuEcGzzuWx3HmuddEBuPnlwe03xbAPl+RFC+Licwd004AvBj8H4fVG0CT
WL2qjZps895eVnfPFVV+MxM2W5Pnfz1WePgxit2Vefv2xAd3Efv/0nsB1zhea7OC
E2o/EHMIlaKnPmUQSk60nwyw4WMUSozXTY8SEYnKoqmbptfQDuG1VRIwD3RkeXuD
j3OGztsLABjqP3xJw5V4nSs6PZF991uaZmhx0zoxw7ml0STx7mbmxO+grTwEwF0D
x9Yam447X8wFWEotT+8+tqYTdxWURqfZXb/GkqqCQUYkuzFQyl3jRLs37faiccUc
jbAE3ss+gs572kXij/ihypvVQanR0Cn8GpAEE1c419XA6+o6GKAjqbRyIKBZxGVI
iAweVjbIVLdazPpEZwOw+xfxk1/uoYi+SxEVwytr6pTgcdeKc5IFC7UQn+pk7jMm
sJEy0tD7Z5ehjIJiKSUtGuUgOPGmcoDFn7BBLJpwiuw9XeOvfxuEeUJP+EcbNW2I
xGueqIeaqPiF9Py8a6be0HNSKhK59IdKT9xESS1eG6optr3QP8yenzgdhOtwcAz6
INOxfcymuGxB9vdZf20ZdntLPwyQ2n8xkIV+r06YSZr/YS0or99gxUHy/F7i7gXR
RopurL7pMQmlocfkjY3MJ21EB5sk3qtIeE78RNJAmNhtKtNi1BrZwh6cbNScDV0p
LUC8hwkb0qmZX2L7C0/zYu1X9amPlL3kxlrmEIRpC4e6JKI+2EdtnjTJYIophf0W
yStZR2VKx1gWhl5jWaWOB2pSewHkhywYS+zIQR5t4AXsfvibX0esRWexYB5sqDI4
F3xGIB4PfZEBlq08z1E3GDBBiyTzdJsMptrxmSdN9nYkJ8DITRNDsOlRRsDOEpRr
do2z4MDoYjRKtpJzZ9lnNaOFB72N4sqyhwOS0vPPddCAfOYMd6zaiTDzr4AEDz/8
Dl3NYqKnlTAnAuJ3TeBiYbgH9cy56+Sbzqt+l3my6sj1vvx8t6uM+zKJB166m9t5
rmxrogJAvOop0Ermz+wuDtrx+Z4MhxjGkzAbUyzPuELjdeGuAa9zjW+Of8GRIHta
usjZqSUBq7jlsAoZBgK0BPx0rFgUhBIs5N4nvrtZaAWXtS1wT9SQL4GNWcSDFMAb
bs8b/pys/mijGydWQR7/d/9RF/HEb+GmShxe9cY+DyO2llTWg2fTF3VWs3EgP066
ovKqXTWKUEqGENV0A30eeQE6RrdQffJt7ZEEAzsx9kOf3LqTklrK6Gn+2tKfngua
q0GQvFarMYXpGw/Segigr7qbHXLnSPsyF3yGzMUHlWjEDlGEfDlHon3LvL+Ij4a4
LtZDDvGme5BJmNyNj6cTfYouAg7eI7qQEzYzeaMGF88mlhneoj8v0PdZlrEn4xBF
9HXfQSjPRc5qBNC+fQhU1LTo4+V6+MGXB1uta6YinGjRnocSK6qYG4RxPJ5pkGHP
O6TMz79jHfQQ/2908obfJeCts3xxTyzrXX1g68oyUiOlxe4ZDJaD7tzW5raqcXXp
QKvxLgsml1XgJ8I8Ftlqy5Tiin3imYGAiOSLB1U8WQlylFbDpBQBgFn9hp5crnDx
LsEhWvlnz+ZJU3jeRWc7ELBUj9EkalMiHcQ11HYnyEskledc4cP9ET2+XsowdRXU
MxNW1OBB3Jt2xDdLKpZqpRYYXeLBJvAU52vq0Gd93bgWN4nFQKxcRZo1nTrHPEDJ
CMZlYxzwiD0H/+7Vs3rO3yBMi8N1ctdMqvo/zsxzmJedoaMVO+GQjFnIRRJ0RO6N
oXyrI08a2ZBvmqIPuysEqcTWqei8Rbq+YY8/jNlMqQTrwpdZefHWZ/mlqWePr5E+
Ki4r8ApF4E9mIcP9jaS6W/4OtGGonXFFgUzv7Vomd94FTNeZHAQ0bQBXty2JR8hm
pjahaRFuThva1y67+s2edkoREs0tiYcsbDaC6AqtRu+XulvyHvv5iLI7XuR/tTwf
lTmi+E1hedJ7Fjt3htK2GWvqZS7C3Wd/DslPjT14g8B7D2odA7V1oYjWJYSR4+Q8
ykyAxiXBH9rHyVPkFs21IAM6Hzv1Ptbzi0rAAKOKrGrprM+zT6v+djYYeu0qRcSB
DWm5ayw70Hrw5yR6/rQluGFJZHVuqjZoO/q9h7+QKkjtcGx3SDdhX9K/R3TzJ7Ch
QDIKGt5n9OO5rqzZGdthGpwoLfbhQUx1az9l6aQG/DiJceuyURONXoNeiAQ4044E
DxllB5dz/BYnoxRs3/QrdT23VmQcSI2o4GUlgeHEU9CqC8vIrSQ91igeCebq4vI3
wPxHYDNXhWTSWUM6XZdfvjhR5NnLUOPjuxxyqBV0b152tCFpBO4zJiVoY01qJuiF
EjcikILf0avFtjmlRwqUURzijHjx+KBSEh5RAVkFAiiF6nKVFc8SUd5n/4UerqbO
pLW5uexWunVK7niZnpcURoPjMMSAcSStF6JIIqCSDmmI7EROIaee3I/VE+/d6aXx
aC4Qm64ym8V8E8JwRZoVKuAXMAMVwZnjsi/75BLvAAtoma3Ucj3XLVCTXnEYUvHM
pVN0+V2UmoBHEQOUkvA4AsO0kYIvQcaIooNYjqxjyKGg4da8QkgVc4BHVo53FGHZ
/c8ZxKOZ0DAYmc7VYwcspu/t/ymJF4X87FpvilK+i2uSHYWpkpI/fDMRey8Ml+zW
pqnvB3Db1IL7FNKeQr9oyv4pTE7QCCPXDRv6itHLS0wkngqktlj4x5Fv9p2mio1W
x7E83HQXENxol1ED6jVq+C+GcdMcEwIlGamccIdkLuagVoOAK6CeHwuBEiF1x486
s/jvgLb4g/OOK+629U+iP3Dkredvfl3wEL4g6TKYh5sxwBO8xI4KMkPoR+lPl++2
k61ceu3xHWp6AgqyHj1JYu4f5UmPDHkO74Y66PXQoy9/Rio9PZos98UljWkLajtp
urliB7ERE4guoM6ExGmXSCtwPXo8Mih0qApIRN3TfcHRVS8RnB4QPk2daf6DSKVQ
4GTyCTrsBjUdoyLSTHJIX2fuWR3KVEW/SxlijurclOCr0GM92Btjr2rnDmyW/a1j
kIpRbXPPL/uxPtLGlFjtkK+89gtYrVdKkTON2pcki133HM4K+y/Gybwxga0Cyvbh
q5T9zTzPETspxQu8nKdDpAajutoHOXCsBTNux3gO6yWQcUzuEmRfMjIpNKYJzXAK
N4uqwtaxzti1zLxFUKMNwP+ZVvZE0OzytpEdmHwLIR/kBSD+y3xiudcV3MBHWh9i
X+ARKdzenZXIQ3hYaF+lSK9N/Yab0Q4dZSj9MTG6IYgr58IacM7MW97NvMnqTSkS
vvLgVFtfeNOToo4RVeZabp/euv5ae6pgTqJpK2mYtgFGQaa+AeS5t3bujICuxbu6
k/yXsaG/J5F+K2ej3pWGQwhkfn8ZGqsxiiTMhN2T7yF3Vm1xJpXh+e7z+He2p5KO
rJSjuvSvIyCyM875DxqbT3N7/V8FIXC3DWTnbEDa9cBvDAfYadrVN1dT5iXFGaLM
wardd+j4ncINRyCoZY4VQwzYzk2OitlMTrFIDv/UX+v8oHAIi8+gcYd/jhiKcEUf
qGFVqdfZEyeKbpiBEG0FsXvlk0wRLRH0xLleJ0E3sADi+jzojJ0PoQlR0tK/OgAM
7BTTPriKxQsjUfgjhqEtL8ytkxJ2BvI6gWjojTGk8M136yMB92POSsrIsZACUEwW
uLFxortlGaOGIYS3JPe6z/tQHctgbK2FnMNUevxyEAWHtQ4ff6fRsWBc9+rKrIW/
9qIgDhNfMhyIPFy1bzxUbR8x2gMhxDmGw4IlTK5RO+aoT11/5s/XApmeWja3s9a8
wK5f0vF93ttZVtTjsHPFDYKQvv1VKopOXV0wJ5ghBDiz18F3nXz36LD7rYs9gxR1
e5ZlnhvYMyd9UVjzVBPrUhXmwx97W0mPZtyiikhAGlGchhrqGwxpq36JuCfYrs4A
zPv2pLzg+Rtyd0iqNAPqc7z/HwPPs8WSf3Zxxj+AZZObr7PxM7ydDgrLuzXm94M8
23cNO6FWxzt9S4ih013cOkZW1LAXldbLCORtusqyWQYzeWfpIFbiAFZQUDm0X3Fh
PNxuJjFo+RfkD9EyyiP3+ccVsHlw9gcNpBQJQXnDB8d3FbEoTNNXhOf7ui5Tn5XI
h5Z3h7CtsZfEoIyjwvs8vmuQ5JleqZTPYTCDDqYYIyU8oSeR34BsQ798pH4J+VMW
JC3i1sVIlWJ8xe0vqYtUZlpsF4HY8dmsUyD95AV4pVcFZy+q4iHgPEp+CgWFECuj
H28WHm+I2dNicuXfdZw1hk511kBAoM4bFcH58wX6PEU6h5uzw+41zyliu3HKC25T
zeUlIXZQ3IQNcctQ3NFZUyZQLN+NF9We7E15FeRGmQH5i4RHSvX4xvXZe4GQ8fFl
utnMQjLibciOkvs0qhIKzXW1qzN05YyaYwBbFqZKE3aKTUU8m+6MhX8NjNacj+zf
idH4q6mxud10+agcs1ibDrnAi2ldB0i5PO+EkXdQQHhv3YjJqQKKXk3AB09k0nUP
vptT6r03tgYvdiS5ooUNRYQCq8/QjWSGRDCV1qvdv+S7xmz7iuSUp36Ap2eIYVo1
mPoO+xwV3OLdk4/RZJBYqRY3XFwJ4P7T+qbcwHzimBw+ayC8EWJypwcReYJq/yUD
2/D8NY+gM6x2YtZb8pPRzY+5uVGrgGPkFXQik+TVY9Sbl4AuTUcOz16zBBaAlGSu
7U3Wn5Vp5W94jbTpsyE84uyqLyRa2C/lOgTR+3Za80L0iJr9yDqdW+dsPiA1+B1/
dkDdTpDEvMrr8zLI/sBmoCleAnIpCE40klykCBMQZDPIbmx6z9gFJN+6DFCyXlqb
chuFJpyYrFkTVG8gjmC8PEAxauz3TGj2kH1yikSW7nmwsGjPU8dJIaYw64+1QmOC
tXk2oin6wBzb7k6XfT94zvdiwsrfCo82JULFocdT/a5I3eFkdEURjnsJo1H5qWiA
gyfgTuT4ZnSAPwAsf5m0y0nF7NP1PBAX/V5xxVllo58QCsMTQ1JqGefupCsR0frC
U1a+Vf+dVkzHm+KTtRBIHBNF2Qu5Z8hPlLIDfbCwk1eGRjZVz93Ox/fZhQoHBNxu
PCm9dptOq+MtFHsLU9meQHNy43M4wmN6FGF1No1V8Uf4QwXZFBdX4pclJUikwlFa
GpAxKDLw35g1Jh4W2Mx4c6KGq9gEVJOl5AUBQS6p0DeMLz+hYJn4qSUfaxZtdJpP
Kp74Eb3k+NkQ844dMh4ayP7vitd/mPLrokyKECRy+H4uXUNivg3Jgoj0aONrrTnm
en0/l8Ot0lTNUqcQ1rOYYMHiGJjX0HFWptmcJlvA2W4N4/Ny61rVam+JiyS4Blk6
8RohzFPBcPYs1yMP9ULYTOpCWzTR33YvRA0+0d9A0PCbkCxiIWQJdAX8h6b30zkY
cTIC4muhCTViT9KEFwqAcothMdQhaiH17scRMhrUNL2b8qqlQH4ZEFhjzaF7XIJQ
YufXnEoaJadUaEMZKSSE8pB0QVOY1fKST/oCkwGoPXOF6r2dx/qQWQYuAr4O8VPt
5QJOulZZqKf3j/tWFM3A5PPV5PlbFzmESGwGBC1eQRnWNTwwdYnWhkrvextNe9Hh
DZrwe7Wk1nbqz37ZQ2hFgxMAaDTiYLdfRPrWhw9BLUXmSjAfuCW+HJM2cOudbO2T
b6BCLYrzfw0Iwn6w5MxS3RfGP1RH68ExUXKCX1HTCO+qPh61k57rm9A5TSVjM5t9
2lAmNjRaoXjMQH7B1aYI2OQkON7oCOZ6DZXYxLFF/qGwymKCaIa9CAUQDZuQ3/Bn
NO+ehFt4y82kuryjY/c0soyiUxkOiMINWqHkcWrkbwBdGVsY04G0LaRap44VRq8I
4HT2MHybyMY0jAChaAhW4YDMF+Lb3hP+nM4gwZBrmlc9+Gb5ypevRddG3V3MUBuK
iIWWjZ6yWJYRHSXBDshFdK2PJ65jIEDpy8BQIYgTLawEm3SYWruF34CHktojKMgh
RCp0N+J2GeNP8m3v0YGLKWGjWgzN4YN+3YAv0E+ITfRhO+esYMYEAVEiBgwxKT0U
Hnng7ViEYV0WnI0FI1q7APpLirqEBVWZTVZpYi+Te/5vY/U+JV3od5+zBIdnIJz3
GmZfdM30963Ls8/FGsUkB1TWO3cOrE3kd05ReVFSzfQvhj1fUJq49ipdw+Gbrhew
aRq47mZc5knwrT2jD3U0hHl8U86LscoaZHrL9sA7K2nVirzcY0jDZ+c6lYUvXGIj
AgWN9P3+Rwis2WmhbzVFLN8fzG/l9Ebs76+pTdy4mS0+4BWJhRtA7cC0xY5qZw8/
ocMWffPm0bUKLLGGt7P+zOuDgm5ZL6AlWOXrzLhTCW2lEOM/O7xPT0QcJCbl014d
6uHP4WdOsJSyUGzdlzugsMBQcBbebkENVL25Gj/ovNQZVxAmw0vB7P2Ac4P1UnsL
+sGL1lXlFnV4e4qGyNZqDtgB+15OVuZRgVwT1wT+u3/ikdqdv48xRlIEpkmWC3zd
z7j5OTcPE7Nbe9Webo58EE7Mu/QwgptdL0N/FvlGx6G3jSeVh+Cl59r5BhaUp8jt
FqFrlPMgCD4PxpYj/T+bbgJNHUFX5X35uRdoc6M1mbTUS/mBhgIsMoXQTnUs4aDO
SyqUt1iVi3GtHNsgcEXjFJ4Lb30ex57G+LF5JQwod3rlhcJk5j45dihLwiYgqCyc
7BQYOuKLB/hBY4/ifAw+oQLBxQ0PkjaxE56b3ZK7U6Vb0hcG6I1wvGkKaBcrOT3Q
Dp2AOuUV52MiMoPqxDuAB0WQQ+w6tzNXaUePG1yh5+OEIljegMSu0hHimFuABCGp
U3JyBjeubJBzJAvcMDH6eZFWxSJhFmPhWtCpNM7tycU5qic8yzplucKrV6S9cHLF
edXF4Ji+ZYjwLEAMMXD/GiGmqXnb+gRJIBhaVLRNov2KSu5Lq9Yy/+S7eVvY7JFZ
65g9Ja/7TRivn6L6wUUS1rojjo1TnkQGkOkFHPmDz9tNWXyi8dKT4fPP6g9V5Yul
Hba3oEDEHsRaKPi0E9BAkd7xA5wxLcVzSfX5GF0rqeCSNMeK5dVh73ZjLzTlFnEx
A/X/K8/lt1gl8grUZUSdBMP7MVNH9xN1o4ZQzjNsMOiyK+d3LaphdFE9jgLcEP7j
kER++3LCic28ck8mcB+2a91R3zKkdPYVdhzkvmlTjXT52w05HVcgzhLk3GrIAOeo
gv5kfmPjexzFiSQajA7CGa9/OwShf1r0wH4rSykKFZVp6AAXCdDsUG2OCDi5Yy39
FwHPYeRdx5+Y0238E97qTgfi1MkjQHeWmrkG9anBNPBfsqK7WB8pToBG+s6I8bV+
uebbu2GXEhdYjcR5+NQ+NBTsVn6wDd0XaJo4pcV66mQTy5vs6oG+cttA62eKsMZe
wYimixAkps3meJDG/ovnT9oYC3TDeHL8nqWKjYurm6nptGZnYuXrPYZmYQBkwJRw
TXU3diPX78TACfRiluBNslNll9sAA946qCnonTHp4Xy5c2zPDcZDFLdAP8hQsXUF
OLDXF4GmZctWYceheurxutruDY0oLtt8grqoOQIfp0zoSdAxhMhiNs0bWysL2c6b
vgXTWoxGzbyEeMPU9UclC2x7F8oHPI+mED0fWhUQMz7p8sYFM8iTVpbQxmUXroPa
Iay5WDClZetB1fC5Vr+wfm1xtDPRux+uYQApCRfrNyqJhESCIGF5mS2GTVMLlTqs
hFwZDl3NlvViPdN0NXNk/icxI4Y3kfjOREzRNmZnC5tUvG3lKgpK2SCCsqGwXBzq
gzzyxfDAWrvHV6S5YU5Pz1Z5HbLjeuq+16DaH366/bWWW4DA6L2dsBMDuamdkuhF
YDiawbkWv3XAbSLh6YWxudOWidFf3QwskuBNeVAZdT1Xno7fhnzKpaNcxznFFZwb
Uexe0bxXjRMhBSjBuhHhRVvxIenqfTPi7rkTQOw42VVaZ7omkVHkz+ES5fo1KfVW
+wI/Nb6RR5hQ13OIjcZXVu8xcr9QIuHNf7nLD7EEwGgig7kTX+J2MTZJiQhNiRyE
OZPC5KBJVgAG7SMONucEMfsHrTPkWxQ0yAw6Fg90FzRK/wNO12PphuLWJmCP+SSY
dYwH2nSHeaCsRdLq14nP70lLofK7bNedZ9YNF08b5YC+bXEb4WzLyViqCSqFur05
iZvMbOZIWumlrMfhjBXUr63OA10svi75sjU06b2DE7KLwVkZJIyICONDzmyi7Oyu
PPY6CNKh4zZoI1f3Va3spvC9LAB4BAanZsY6/HtRFqhzTUWhnkQxkd/n/EKzwoBz
qycRcSniaQpU9oADgrksVzeYaiOu5MSkZfgcouH0guS6BkFNuFR99y5/Lrnx1i0C
MyPRFdjj9J6lFAgA4E3bKrdI450jCe2akK7E8K6z/tLmOujPKy8oB4L2zdMloCYX
IdpzCcdIEZ+6z6dZ3W9RbwgUyhkjCz5T0UpojSwdlgtKZq6hJICpmyp8q4Aa1sIA
M1y4eTP+jj7tBkoekHhAK8SyZ+effbymeMrxTIdtGqNhGsO/E4ZR2qCcmbcI8m5Z
CKYVNva81so2+9y6Uy+/QZGpMtU+M1pwg7McQLEbrKiQVPzSzy8yZrf25grC5BqP
jyLfO1fixprEIdRdswZjgeDwjNtBoNmzIIx3eNNTYKQgv0q5HdWUHqmInb2pucRh
+4AQJmPEQbH5YTKAGdRlSsgRMtAhRengMuBWkT81bYsaW+DRyNZjOyUm1QsIqN2d
vSo95v+KwH7HroPRpfUWf5xuWZ+ulFN9jGFRvsiJCz1LgUI2yU+/jJKcUcMcLKKS
jPgKjsJzf4MsPS9Jm7zXp69909IGcbaunlhdR5vqOQMAOnyJ26LKhbUKurObWaaj
1eWHP8cdMjvZ5lllUwZB8MEZZhXGGSuETytI/iWrQ81neSdP89Ao0iVDHHJK1QUs
FBSX9UkrPcw1vbp87N9X2RjnIJV2aNIg9ZhYRmYlPzLr5oB8kaCB/ea2EzQQ0nyy
UkeqhTQtFz2l4T88DTzXZfH+ITnOE9sSKDn9ZihtdjVEcxIjby86z6u2/2fOXUum
03V7K9MhAvi/7/XHkvozfVwztsvJxqO3c4GbEdRiPsrvqAUXMTw3+fORPh0XsP8u
3ybylnrolyi7grI5BWj/ZyijBj2e9fuZilUHnAWVOvFuI8w3bseXX74ICtbGj8bq
g0hfjqhfcBkqAF+NM1qWoMdkHZkz8wOY+RdFgq1pVYA4lQvlYZttB3PJ6QJq+TQO
XCq9rT4mJm7f+SysuvMLfXU70vxbUaZyxJ/YbgzpeSh0GlkNNIZCg4luJ9vUL5jz
3u0EAZbecsIBNMQe9bKGsExyoXzai/R1tL4CWrh6PXvQlNkDdc3CY4nF/YQspxj7
QYmQPoeuj5vw7sofBl/GOTfYZKpZb0qCCMUX17xScwTX43PT614DyC/BVTOd3Lte
HQ7CngHaCYW+SdSJtOOxTNDmtndBTLa1G9THY4VdeAs18e7zJec3YZ9uo2JKb6iL
ofTLh/V+sHCLNgyE9GVHai5bIHCh6w9HfIzRvdRV4AUP5HEwCTl2uGw3I+9X8aar
oHJZDNQzc8sFP43GUqZHEQShi2z5phtmGIQ6ufLnxa2+b/2beswZPVqUZp45Vprf
eR4ccYuMZkgnhwMKbBt/635XZQlfQ6l2u27sgRmyW6uUx6qVF3cR17H/a/j10PV4
1Pz2HMY5vBCWcDz17gBPsrnwlpvZZmF2B4/KtqFv7RTvs3SEFPi6yIGTejneDZKn
o1rsahq1qlmglUMCZ4y0fuf5P7xKjYqNJ8W9g4MKPrsQiRrYIq3nh9oEk51V6Urp
YmUn4FFtoQaPMiymEUTyNgG6KguEZ+LhKjbmXCHZvCmJJilBG8IUgpREWA5rN5K7
ndYFp0EpoU0RU8OgGC+uVHsXySfVyK+SZmQZJRcymOwpm3vWaq2cbQmvsqvaYc/d
a7aw8/B7JFUy5Ru6nu9t939Ny8Llr7HeFyjokoDWCYm1F1Z3VK2s8Eg/xaXrr/Sj
zDoZeukBhyb9lRDcFUHqQLMYD2PoKiYzAunva1C420/TMB6ktBnHxpo6BPQi2G4r
2velyPxiaR4e9oToTD4K4JtS0D2huOqpakjAU01CiaajnCnGmqlFwtjg2dlIp2ws
/GtzSN6h8KhWvajPigDvGVA36bMT6Rm9Fs58zmLGUgO13DgHd9Bjd1mLcCy3tv1g
hob2vosCO3wAIXBkpC7lHL1LrfXdMGziGtFEq8i+1oF+PIuVOyEXwc2Q6wlxSZ8u
0B34edYx4Tkb7ASY4V33VuiA6uSwo5zv4vEGdySWOa7RoCrQ3ADxcB7nYvwAiYeR
+myxskEhzT/6xgD1X2VSPlqp050MhqlKG8qtiQwVnoFPHXYL5bEdWzm5NlQ0PCSz
Wha2BShO9nsXy7Aey3yDVctb+jgGn+/lOeVP1qFVootsVTFVP9qtj6s12ycnyF+z
y/fecdhBS9DUCjHG7zLu8PCLHHyMXdnXc9tsnbkASjcr0KBx01q3uFac7S1s6afR
aKJjJHxqN+/UgxujvkRa1jnktTefMNUglJTFHn7EbtcR5k6K+2W+idFqFJflizaJ
lUzCsPJJQmhUxzyCJabn14EODZ5KwFHSJBV9ZfxoHWDxVt9BYjeKIfC0fw2+gKpv
EUraIlJRD+yfvKnVeeTIySFA3HSDv4Gl7+8TU8GANy+u2JZjldnphxKeL1Gkyaxc
/ArP/U1iCdcwicBL7BiHP6KoXaaSwyIhYTWVRms6d7wBdfHCUgzKVDkaV5VTwOPv
/b+iOj9kMFefs//ftP76vRtaaortGyzBiOdncQh8GqxX5LNv4FoICqc/DNBuVo8Q
+zZ+g6qZnku9GGnx27JtR2tBYvdXh+9PK+8JJHtimY+cvtbJBiJDsrx9oTyscXaC
iorpf0zPuWFgnKm1bspsjgW2fBVdMDOZgo9wTR7vcI25wTac7n9vEOjVcjzoiX3q
JhRoWDa+tjOjh/df1cZQ9OyPdQnY5HyWEJjUn4NJ7ReHmVSzyOXtr88JQMQQ8KkS
BqxienpCs8xmRc6qPQMOa0IpSjTXwOGdLzg0P459vbTks0s0Hnyg/8twvkDC1qej
5VNb/xq5FkScp0WmL4viPMXJEzeJN5dAw5sOq3gx3QdEoBJ5vSk7UxFKQDbMY2c6
aHqlHbHz1ehBfC7p6bB0uK5ogKyhfE0pMAN/EbV2of3krq4D8Vzt5bQzNznLm/j7
vEQrxhTVD4/Pcj97R6GJ7eOheIdyGc2EI9obIB5aSIi5Gnpqa7HLqst0d4J3/Hcx
QgQ2FmnVz2o0X6SoACc8ImI2JC3IgjTWUF8WhC7vtDYyKmkrdsHxN2lE3g7uH4zS
miPthPWJT0MTprcdnYn+B4Hb0e3QNcrFYXoJBhvArf8Y49oXCICf2UQJCp7MDAJN
N0nrkOmu66sOQFAbwa24fus61Y/WhZsGgNV/7Ew6Bd7REfzWDbxQTYsvzf8ffrRi
qa+xp3MtkOtCrJa9Pgrp1fVt7owIdh8od54VFmyVrMc9YJHS3zdWeq8IEDdLFbT9
rV9gT2twPB5YrbNwsUqQ+nihj2ZmXYl8QP3kS7Anc2J/4j53Vyvob4cZNHegZ86k
iXM4E+vWFhO14UIrvIOKgHrdM7FGfAt8c9+f6O+l/0UNVvHZykcZU4e8wnna0SSN
W5+zeXCa3pJmeCKvbOHtI/oiXFvoeaxtBFAhEG3a9H6qHF6kXtDfXfTOy+pw+Emq
QZcQ52bm8vldSE2D5rxl5ctl1Q+Y9wEl5DkcO4gLtlT1f+LCE4HuHjArMPXYh9Se
ZkSxWgzE7OYXGmPk8TXawFLtP4XAn5AkO+NXADLXtymSxX7Y4r9dm+k9hdU2iMUG
jlcdsZeewYP50/e2gmLkiz4bzMHjJHCilKq2UQ+Txtdi0zPje3SxUU2Eij8CLRno
4scOmHS/I9hx1hwzkdhFlbRsMk6deP59QD/JqsP2ovdBEEnioFMj0oc/6iFohu98
Mo+yafVDGtt7gjaTjgpYAv/+hVi3+kXBgJMnlKf8P6+cyI7eDUhiQ2RCeDsu3Ufm
Qmey2zdUWq8RSM5ElI8iHn7NvSRMn+zoyzqrf8bunB5EO75TNeOb4zpxxRZXhRIZ
Z97H2okHe9yK24TMpvJkYblYQYqv7PT0R7in6jskBlC0f9PqREVgUeIiyNsEJtif
DBW/jDisxSYCWtOU4eNL+C8Qm33i7DhwI40Lkid/ZDue25RLWz1PNJliRGTdtgVw
3KyuXM9mXh9a9faF78+9gA7AxN3ZhFfEHdCXzAVcOxRLcKhJTjw5cBlQ/aU9kuvu
LnlDw7bjoPffSqcEls32G5Y2+7fzRi/KbRzmWNmahSaP5klSTGk96ss4ij7coxQR
pILgkFPCW6i6Kar4KzhZlP7STPz02ltTV/1PicsKZnYzxbD8LUI508yDn7e28N8f
MXnM++2vTHtc0BhkOMz2P8pO6FEdm5ewx84qg/5KKJGd/DeCUnkTDYOl+jdIJ3NC
Q2D6e/n+u73BC7LUmTzA1ReM5JCFsXdd3pBGZqbrKExgcS502zPvd96oVPKtdnFc
OMNQkNR9RwUrnzr3ueyU22J8wlPq1wqw+5FtPh48Oz7lwS2dSe1FpNqiICoBCz4X
MhPZdD4aQ27HJGLWiq1A+ybLTn0kqPu4CDA6DGtMQEAMohfpOk2R9BQ2Ir9KQBtJ
oiWFgPtIqaWphTRENVTHMv8aKvIQn+E1x49D88IayGVss8Z7xsswQMMxX5eYB2c4
AAqBUbPowzDHaDGXG5rqgFGmXmb03+fLbyySf1vxI50Xhw3qg9g1SghJUFtviHZP
NXLpzku2OY/1cOrXoezBpLVFGQTGy8n2QEQznGrdrtORLrWmtrDng6ikaiBDV/vN
m81mcO6+BN6FaD3FEEkZUSq1ES1FmYLG+b2QD+/3qqSzffbbZX5+M6+tfOkSUhWt
ZripprXiyrA6HI3bzSR6Db3b6wMk7/A+9XHCj7HjY73PbBfMf3OOHFgOSTffy4ZY
g+sgln0lEWxDttFk6GRFsbX1y+0fkUjM65mPYptA2j41njOTVowOEKxiOFNo4/Xn
KxJViylGLFVjgU/E/MloO3ON3IPf9X/784P8kDyX0uzALTPDad0MomEQrlDNE6P+
BXDvDHxmJexvKKTklCoYsUun5+9ISJhd8IFJZpqpVTmDJWBIfNlB9knBAZ69kg6v
GDjnSYBl5EQK39LtbGvAXuf5XmgnwCLIxOZIzm0kHRIFdnvm3kNK6sEvfJSsvYxR
QRb105j1hpkBGS24i5czUfzh6t+tdkt8ri7v/8ZrMoDnvtfz6t8W+PpdcZu4B7zh
fUbj3OFRgI0u3kQCohyuFSZaOroecOcWDjy1rmmkXAMDIezSU8t/dETYphEJKf/C
UkbDM/1vnhUMxxGDJPXA+xz68jqYtv/fzFZrAJfpfE9R1cUfgohclL2WXpM1W54X
uTA4asEceFag2iDZkTiOKdexrz0s12xut4IpkKQPOjextm1qwZEwP3ffgBpdzFPV
tIHeQVzRoCnaEmhb9V2zgWNDHWfHsGSldDcGICJHJb5KL7GjA2HXUIxjdPJhHRWO
JcNbKCX2Yi/FT6Qqt3dY8T+tsdJ9zZ1ZL0Fe3oh5EqXM64SnNps7mpvgAv8vZStZ
c5Xh6AEkyuSiTN04kvRvyEUpZ0Yg0Mo2+Mgdb6FYV8bof1ZUvRKmVV4WBRXNd13u
cdVIYiqXRnEsn0nU+aCul0Vb5vqrWvXkJSgl99SelwIdLSHQ/GsmQyfRVEBdgucn
BWzFr4c5RjG1xrqUzbb2au4dQS9LZAXSGsKRk/XAx+fZakTk2EmMxvCVz1F81tJm
0RLAQJFk3BSr7Kba5WB9U6goGmifF9UFOBijV89LFtbp+l3WyiqEb2MLKVsWmZON
bcg9S5/FNsHoPxS/GP4znL0IMchrk5v5DrHKismQYmzNI1dx5hOyc0jgjEGzCK4W
iDrGzrrlskJeuvWSQcYH5BF+Sckha4kAQX+Zm96p3opgnHB05suPvnQuYtJYaEKt
5S3U164AdFY88aK2c3mgeHAih8Q9+o0Ekmiwhdd3kdC9RiwqDhX0fFOuxI4D8av8
Hs7RIwOqeCNNWyV6wQ4pkYp+AiZsub2v1F1jzrMpAEIlQ9E/etPda9oImnrRPyxl
QbN1IrKOQ0UWApXY8jwAZUqFd87oWCfEou5E13N5YVmFt5H2JLhvVvYT7bhpHIiZ
Wle+0J20zsJxvShoBEuQJ0f2fdylWflhMyFRBYoP0ROKP0sjeBGVL4WsAG/9rWL5
/GszNtnpPEJKiENwBCOx9d77hKsBUOS3lgom5JzQrzBmxGPCutHHe9AbxY3TBLOl
duXbJN1si17hLBMXx0lz9nJT77jJyMqZYwOpPUK0mspoRm8TAmTGZHCEH/zpQSvd
KeoxeGANrVIpGidzLR8Ut8keJ1jEhqjsXns5mXYaZFPkiWWYqLotEicQscCKM94Q
72DebXED5AH4wp5TxzlGZx0kX5mpyTiIPf0J2lH75yJXftd/os/VKG5LImMHw7KQ
xZmTlfTMgh87zPF5HvvXDFA+t91reAq7ClAQXR/U3FS9kKWWM/fFijvbZilKSZ93
HePR16oPE2rs8utQSb3Q9ZdFla1XHrqBbtZiBqm/e0ZQm0Xb5iUuyXwU1pMJrMOb
/+LfesptySnw9uo6vGF54bqxf372r6AhCmH4otYCuc7BB7Z8U5649m7ZnHCCltZs
KS2YJTfleyZuJqkYrDdfSU7rKNwXcaWYhH8FOlEhjgCWGPja78MT8WQzPy9x+wfB
KGEMUsCgJv1w+rV34TsfAslvQzyMMx10fFGLVaLfBnaW3jpbWiZUD3yLPvK8AyMK
L1xWEbVIlYucq5EDfPujskQibnuNMjqPCcoxX2b/3zV3EmwtrGz0YKGbeQPQ16Xe
+RDBl1Wzv4N4JOMtmr6Hcd/Cc8VpXa9PD6CAzFg3Q0e3gkge8riV1pXkEvqX7VyJ
GjGn0GLSao8dynBDn1pk+8dMwYk3sbzknBsNYddhiXnW/4d0znOzvy+Yc0cndSBT
14d6T6HYA3wNQhnFNhT1at48cDzath336Jm4o/tIr/vnpw5YGDvTqEtZ8yGBZeCD
+jpps2nlYuuGnQqmgZBCrLx/6bjV8zVHl4ixUUilW6IFF4rcE2+VNCL+zEl5wQ9s
nraFrnQJrbgmt/D34oubMdd9k/oZSNtdeW0THoVdcN+kJjKIW7AbPyJZZXLyA3Bt
Ur9OSZiP2NfDU+8w3/KIWJV223q/sZSM353+mT9ciOkTkOwpfmW6V+gt4H5LXSu9
n64aKinFEvBfRq8DvFDAZxMyzbAK9hGdiPfso74PDGv5vE3VVeEwuEvh4vL/i1Bh
MLgyMsvMkawLHWkOxaoGPpQaKvB4n9F9CkHll6NwhuvVYwqvlqSzJFPPVv5oLYJk
3G5xiDpeWRzoU8/IR+4/buKROQwHtQBcuzfj04UH3EUhpgJDxxjrHhHXhA5O6VSS
O+kcsbnVsjg2TtGD8jBqPYjHrvMn9BDMbawOHVaeWJFV94WDqc90ZpWZ+qcjkWaK
02zjJE9tlUquiSZN6dr+iIulrvNKwpUoTQ9I0Y+F4qj2i68q9eHGoTf36rZYUGoa
PoIfKvvtakCnlu92dGB83SlcMQO0bBoC3Zng2xoezIrKBOcJ4QamwRwcPIsEqA+O
vXRZk+PSJaoj1/XCw1YEo07qUEh8WbhBNwoZnigi1oHFQGiS6VqSs87eXBCfryt7
KyE/NUtA4NYek/jE8WVKaNS6PTgxJm9+Tf3vTU4BxSj2cHBcDb7U8PezEqJqWsRW
+DdgExuh1jmHPb41tjUZko6BjP5sj0OdB8744DRWQaM8EZ5g90TeSGjyY3jF6uPy
ZgywR98ADuXWXBfdBDb0O8+mOpLpVnYhdh104KPiuLNQwj5/iJk67CNFRH4EUc65
UkSNyRzbKXqmQHJU275VEHSV7BXI+T9Uq9n32qV5ZQoowLMXwqPcMgBnVknXQT8/
QsJ1mjcpcs0b1ELC+kx6uSvC5ZpNVyhIFfJD6WrRx29x1B4t1tMXkrQqazCgFmw6
Sz0TBGUCpyHm55SJHcHEXT6s0UN5g5fq0HQqQJUX2ysXnNHXA5kw0zGtrN4RixqH
bBOBCXtMYdBNv/WYjW1yW2+Y8krfNDSUxyrQfOqZO6K4N461iFxnp16fCN64NhB8
lVUK/Yzq4B6QDOnbmvjzIxswrdvztt5+sc/U/U175q0yPW0SF8uX5ZJ7+IdyvgCx
gu1Cew99Nf3oEVP/VSg8ICNf9VFi0lqeT6+4582u1weRHSV8jIyNTE6wuHMxLZzU
Nupm6fV03XtXD3m/oDI7jYWxKafqFpcnN+31E/eCELmehhDbpeOxXM5KD9zLq865
R1in8ImULCTkMnliUjypMoXbuPhPa89bWUIpxTGxV3OC4cwOm6jF+7awPhSgdjrx
bdICYbvC0D7+DlSIDLZlcHLy+2klrM8a7k9wKsFKH3sEV+3xCIO/nfLjqcYu+yDu
PsN4JpNcY7koRvhN2B96eEIZALbgCD1AB83upAYecm4YUuMF4t4aMqWXECsdzYJq
MqeZ5oV9F6lwDg3tRfxrQoZMPJUsSPCqulqN0nkPx/NLjzCk3VGMhS5ClfSUGejV
TR2atFPuAdiZ2rupexEpoj+K5A++hCGBqyavDoVlvANlHi62w3HOCulBXuzX5Nq5
BmVaaD/EY+FMUf7LXbW+R16xu8wAocFvyLEb9WtAwbQsZ9gNlqajZoOZjhBFxMUT
HRrDI8UC0HyNzAVbtnCRm+Yau6fXqzuDWCNpN2pjPuUqI4LRvlp9KP9W7S5QOrBm
SEn426whNNsX0XSf8ZaiYdnQkkLI0nchSOScq+ARXynHuNilJU+RlrGCPTf9v+yp
BpQUXCcRDL62Z7jW4RukGZXnfAFY9W2j2GYL9l41GXVXb2xi/MGhrIPlFVftzqgv
J00ecbflBghLZkFQDb+Mvt3yL1c4fkUPHWY/mTR3Wwv1mn2TUbEfQ5eys7YRYZV8
92kluXzU+7rwBVkhkmDrIN5gG6WZR4/hhbIml3i1rJC1Igc4mBD0ZCQ0NMcNpDg3
jGM0qs7SRt7xmeIsy9ibKBFc0YuNRR4NJYgbVlaQ4lAVokDnMChIaueuQA1tR0DG
zRTZ4vXb/27sbL37ewX1yPD34e8yEh7ZORb2Eqs1/xrf32zQmwrBpkilCC4SmM2l
jQ9LrdP18JSr5QpoqHZNSkwFterKuIpc77iIzWsZI7Kj0zGxRji1sEhucDrCO5An
bGsgqIfOBMjK6PKLKKoqp21kikRGSju1N5uYbvhRjevNH9yzJGmAY9Jvy1P/vCjt
qwMbLQr1/QjUhLKIuCV4K5/kCPrVJZlB2bPgNU5TmrQI4tnsvF+U/aBrChbOpuEr
cHSxWuTFY6b/8YEEHPaz/d5iyzX/l7tcVcR2ltJKREBdD28GovUOpOjLev0pu7hK
tFY48leUS4NTA7Q1IFzMrmCkQUFiVlHEUY8Me37halK+n2yS/5QUJg13D33Xk6bp
HssAlZ0tn3GdOeb8Vs7LB1uLL7gi4hoyCTyrPdI0HQmZdq1Zn/neTxjAAnVv6BEs
0L1VKFueGgY8KCkeEJiGp64L8faovMZwnvS4Sq2CfBSJoGn2+g62mTyBq+K2o1dI
QakkxyETDT5xmbTd8SwqCM9x3S6cRpOcIuN6WMZXsuVE7M1eA/BxNjsiO6ZFYOzU
1Lp+H7C85XeEK2iClmWz7LWJUwHpnrot6FIbfe7QX8q8u24ZOe4jUWjekKmrywqu
CyICxLmB1wlFvRXL+b88FlCQJm/l6vVUhDAxuF216fzv3BS5M/MX5w2paBkxKumH
QZy3IvKOsy1W1bb88IPmAK6iRJlkHmVU4A3M4yqjcHkIjWl4X5Aryf41V/p62muv
Y+mu9rvyvzQYOT2lqSKVKCKQwbY0pTvtZuio5wyLRkcrbb606czwTDg+QoG9N/WO
lR8B27WqPEWtPn9+y5xXQTugsYrZOJiauWF4v0vveEJ7KTCu815log7kLhAUL25L
Bvuxkmj+ohnsywEvEIZKVj6E56ZbWLjVWaEpQU5tXLtoE6I4SDEvloqrmjYbhQE3
gats3ZDoG5l0ubrAevlaHK470whOiwMCBh7MAOsIUziMnP9Pk+HOqp+74PO1xSy7
rEpFv4DP/fl5wANhfXQ8FLCAcV/4i0GapU5NIVhgEDcZU8dDQ+5PyWD+V3T3/wqO
jEZMagBnDYWSNqe0yMKuMTKoV359hZxeRKDc6CTLT19BkIWVQsge+T99cwR+wV6j
OHZxm5dVqnTYxJpR6arhK4DOCPyu+0kS4DmkAl6VK/3sqt5BhjOTqml+v17o2Ba/
Cz+tjbXYXfOHbfUTgYen0QGTgQGQrvUhCg1tw6z2UgHL18FXqlP/KH+MvmXweRPT
mH9hX1uGjasRdqS/k+eJflDFYXUq3hN4ZrGagy58XNqxqFbC6g0VpbhbUlLaeE2e
2VKqF2iVmETMpkOaM7LsfzfB2bF5fycxA4l0BnWE0ughh9MzxoO8K9EmS5kbHgC1
1QsyLmDoz+Uv7u9d1hz6yXHlHIP4ffqUfkESbH3CmyMxc6UWumlX78BueiYgX5nJ
DtsNGjh49wwruiLI2+0qICsKcGiIMY1GKv+vb6A2tPOiEwLfrlWHeg/MAHPiIr21
8xZbq6cDvWYvSnDqJB5Lk2GnxKQMGGEaw2hDfK32Hg0zc1AQk2Gjm5PoXCZCPp/o
fm9/KICbkX7rNHpTcsdbJSyYbq/524gsTgntw8otxx6wxnQQl/h380yMelyxYPkp
dV4+k5m7PXrOFndCfukfDrkKOmOCHO7Y1oQbbMa0K+yHx63l9PIJCWQG4s1VpSJO
yMeC7TkHDGQ2pUvBw9l2izgipvDfeANARZNjU7uwEfVI9iOTrYddaWgkliqPlpIp
NFf3Os8Lm793Qe6ZuPJz5k2IzJ9QDfGgTBuK+KXQhTOZipVBxc3ZenxEJVSOwxKj
jTNSJTK8W5Zo/VzqnW+jEEabIdBpPurSHR3wQg27gYmI6o8CrSusmzcKeOaB7JWU
e4tXXclzlQyhDhAEk8GCUZGKvoWbY35cPU+8tBzDv7h00ByVDJGyUEa5Q0jVux3n
l5KF5uLzfNWgY1pQ9xO1UVnvUqAsqrGc385wqldI0o9btpj7X3QyR+JcbzBQC/5M
5wIH5q4wZVMxERxxK4tNDOwCk5vHGn9NwH4LS8wfg5SnyaKXQ6TGH4zgGX/1hZSI
ccwplBv0bkjMpVViBz2cAqZI6KhPSjypKWiO72TETCk9eQQ8wHwPJIrRzXKshisx
IL2PypoD7h7SFlZugAzryAomlPoSbQpQupEfDgJ1T4m1YEXTpAyRXlYjolXlXYW9
WN4il+XKk0UwSgOZZhfNrMjstjSrQEP/GgGauYYk3Jd7+WP7BB3whgYGKUQOLIJZ
7ZBPdH2/ENEslAx+XE31kysy8UNd+FkgB3AuGo1KWn5QJSskUz5jupwu5//Sqzi4
ra5ODE8OrV3aPC69hoPEAzc/J32iqbotXjzqFeqhmaXv41TvYzrXicdmBC5HvIj/
tXK0dIzGHd2g6ITEm/bl5kQqOFCvR139tpJjLiEhYYz4MN+yLjBPbxn437wcgsNP
zXzqy27b1qyoq90lAhbKnSLrNZvLlLvfIkDqz82/stCpTb4ZUKqpywEl8KZSOzCa
SEFsxdYZs6mO8l4EygoalS8CjL626tkLBx5SXkngmZ6H2FdKbJODZx4yfRSmLt0r
wW+91yd1osc+kSYgxeFLbefaPhDAY1KyB0j/WcGjnMkApWv3mjXbpQ2M4ncG82+K
ONG2Boil6JtWXOh3oKSrObErBAJOYf+uYmgkj9UAfFs1pKUlpoLUGz0ddPTEgKTx
qgYTsbdXAXC0WdmWflzD3PUrTZhTfkAHKs/zZQTSviHo2VANb6W2Ddl8tl+uECM2
gb/H2UT+oI/ZjABcxFGmULtGQB8z76flkO+LbcvZwEzD9bFU1jJgY85XbD3BuqfH
SdzhnMoylo0UKHLCCFZUpkGTUwSBvisjFs0dJCi73Zkn3ZFYEn7/E//xJvixYNoV
fxJWoTq92neMJjIAx66JIzfVUXZ3cxocmrAYts1UHienJmDvHr1aRoFvLIY0Fzzj
jQkEqowEX1oGXGzD4qjbLbbawVtG9bEtHm+GXw8bBc58dUw08Pl4SsI5KxQEf2T4
iJ5OFGsmVTt9KXpRjMdKIGXMZtjYQLnKHs04MOhzNou9JJipAloI34wa5lnOIkyf
f+6J9Ie6sbvtyYgBy1RbA3M2sFtwyajd7czFF/O+ZHlTj4PzzpFaKu+rWwKmDHXj
KLzE+gLkyAe2j+I09wS7rbgV+QK7f0pc1i426lBG3vbbxJBdPUc6NgVx4aJKbYVn
VyTHGgEFK0oY6U7qtRhZFGmQ7hhjVfgOJas8l6N28uHzpWnQSQYrFypSMYyOcaah
u4ozM8k15TVdMbIMpnYErojRwdhhAeBNVIolkEwvQ01yYIVecS41pXDs8Q4+RlR1
V8n8meQHesGxcYUav8Btl2MVgv86Vgz5ypFx5jpxydevMWejiTuOKgPnZkA8Ghnf
dhaZt/9KvEJJOZpBpg/5uLt8JwmfedisTMxs1dOKxpa9LMnhi3HZhOzzE0RhhA44
GQkjE7ef37Nn147R38QsbojZ7AVhCSHbXhkGTszRk2GR+4A+3JQbMkbV+uG3atAQ
nmHo7U1TNTJ+1x4GeFUaHWCvhNVfJ2ypvEvlfdoNA2RgGOsLexF1KoOR6O4OJn0Z
n88NVKIYHD1pP5ja2eP2okM5RBQnsN6mVLKoA8WwSo9OyH0/WkY/jJcMh0cqUvAf
FTX6GmwtftOj8nV8P4u1RzGO9pjDHNpun3rY/Sj1cPqXZjlhV7NX6g3Q9cE5eixz
wIb2O/+0EvQoflTLCmvKglzu5D1frIEue0oiiatOzgy24Rf5xcfOXtfGxkOK0ByT
CgyXMza5p5NPW3IJCDhbs2o7t8OsD5QeUcOvkR353WgdEKrjMnWe02T49TCyPiVB
9eXghY6+TEyAYmQfb0G9t49zgnfwqQ7NUsYcBThf2WRzez6FiSqup11Krg/PiknS
xghInzQYH2YATIGWMmUZBi73tegcCu3munzlnyuQUE+ooCKq+OoXWPD678RATl68
jJDGUMRSiPLVO0e+tGrHUhBqWR8vxZB/N1JrxsvXn44Qy81ErWBF0aK5mU7xYjtn
j0Pi4URKTYyOwot8TW2v+exWLZ/Vbmy/lPfz34GRpPJkjGnmgPo9Su/xkU0PhXi4
5pEXVELeRiOWDrhVwpUC1+9fcbobwYni3AQh+9wVr+VjOAeEqq70iq0DUAWgOK9q
pS/fibWbDIfKTFwG7mG01qUvNpoCdHA3TBb0nohPAOSSDoGs9F6zJRZWOxw4c6sS
TWxwRfL3io3nHYBDTEMEXgKOGTRrGa5HfPWKT7xZkU9jVM2FYoFmOC2PykNdYcnp
XS3DypqM2/rT//obCpOEniTUJR7xPE/SqB2MNk8AAmEH0+G+9BhSRg4NLcLuyFaf
D7KjDxdVdA1hjSez7fq6JlYGlAmZqdAQh2DG1wBFyPp6ktKCCd5d00r4qvXT8nFs
2FI3kqBVmgKbelgBUc8Gwstt++SKPMXq+0YVSAME0Zp3rWctlBknnKuBY59Akmuu
q1u9oerYrrbvek/5jVG2FfKTRPaQcRVx8UGbtmFxCbaXGrdJY/X4JAgv9kvXDv1b
VN1EkanOJCovM/H3vLACdEVG3xXCFwKr1OnaDg82cDub/b/WI8r9/TLpRomcqGiN
gpTFtARkldbDjabvAZJ3RrP5pQqsn47dhd70XqypCNl8jJQBSjdTRRmlWGVPIYYO
QkrvYhfu8sn+o2oyK7xPk5XM4XRaCBmRr6Sxx/aR1aEmTwCNsQM8pguH/YNmqi2m
yvAsg3ucAP7ba3ewhBUT/8KOMek1d3VBOV91L+6fUJL4ag8N5/hdWnnrLcubbtcS
he7XpIzyQH3OgjXNpsdqv+j4i2YoYYWFBcFaPSeQysaB5aPPu0L/F9hivvPQYx1l
7cZOZAf6IvfWA2oUDDMUpDPrVz1NOalfwFWI0Gx3FesmNBv7wYOKl+PpWppIlO12
MhIGI1IiBC/7prlPlFoMurq4vaAZC778Vjba0yuV8fGLUQ+hYOBKzycKFr9JOHYK
vFSh5xEFM2UsqGrYbYsU3tmDZYd/RLUFoK2HPQ+OQIUTWDk99fNgllYA0Mtl4A0O
mc8MCgu54pVc3wVV26/whG4GwIh/YVW0DPd4fdHEGbVUV1L5oKkLRJz5Jpti5Vzd
aKXnIz3YRL5VCDsiAgcpA1InH01XzNFz7CsQqx+ltV4JMb0FlWIKZDnlf0irY+Ju
NNIjkQKpBdHx+4ZN1qmbmIQLs56VHiVKW93tz+N0Cz1vGFcoiFCYxGfB5N/MkgHO
r5GvcHy2MDplmO2SGVQqRVTaqf95vDEsnzA14pMVtgOdpBBu1d1CN159h7Lvw1na
3b8L4V6GtX/pua55gf9wz1OyACgob1CrixeAynklSbJFS9jsmzCraFSXYfYu50St
AIMUpET0WExA1uLB9i+iPQNXlNCdG5UmWCoLzKaBDchC+BSpnhqpdTx162mAI8uh
jYLapeKkRGoJZDeYUX3bDclpLV8SlGW9mfbb2lV+mDANO5A2HiLYYQoJ1q+Pi6Ni
wfdPwcpKXy6g5ZdmKhAFHWm3HavU8j917AH/ZRsnqDjwMyGTD1CLuJx5nMRGc+1F
55sRTxl06Y4Um2YgsDH5JgFXD8Y05PeNhxbn/9J39Ht6BAqTIFJHyC1qY+Bnx9AL
D96yV+hrFS/Aj/I3BjHhMZMWDr43wURIJIWqfH3QfKxMTqo1SnmW8Dcbl11zBDA4
/f2jXG0yp+Th1nP6EiOWz5fv+VnNLLTZe5fwg+N9QCHnVEn+Gr9UUnA59P0mymsa
KYCctCx6p4NIyHrdNM5oMXcE/r1M3vms9H+GYxf9ueeUB+Kx4x4NRrSith+Iy9wQ
3seHVDmVT2v6rEFLQuZJao61WR/Tqga2Lh8b0ezv0YfDU0VvRPFf7z5zNb+uoFGh
93LA1TAeULHz9W+Bc0LW4Z7haaHbFD0zVwYY8CKVEbi2CK4v1BFhJTRwANVdfk8t
62EFpnpLPVajig8kQsicPkJmpFLK9fhaisZC+ZLddaoSPFAHJIG7B0b/iTdQoYUj
8cZM9zToOk/0Be6ycTRPFY6y8U9lIV4kAXD3OhMCqFMsgJrkFxIVltjYRbT9T3TB
jMNaAk2Rz9lVqP7/QS2MlH/3Vrg1jFYGfOo9RBVozXWfeGYarKL8QVqpsobt/wwB
2z+WOU29qxfXPiw3+AaUCdxMJrg08WM/fSTddvPK+QH1iVaAX3tkCCPdMsMmK/Gc
3CEjh6JxZqrUfgfgxSrir8aeC6X0lY4wGuwAG4z9kSJ/FpChFmVRbaWCoSIyBVBe
uV1BCKR167YPnxo9KBWbDb4XTS13qhzq4bHD5rVCvcl6sDc3vTg02RQ3p1k9wJCt
mWYZi9y+cgPWKjg43z9A5qu3YFa5EPHZQvT2t4eyFrI3248W/Qi+48NMX4WS67Lf
Q4eKN/BGK3xKNeh88FhigOlFXXmGC9DTdM3z3fAIxPRPEO3X6BwOXBrxDPKo23If
Llua4+fRDzggV+MjqS6OFSj4eF1c1TB6r6ks/ZiVH4MkmpwLlZR6lAf9qmopz24I
HIEHnSXLxZsHCI1dHK/vO+MJWYwioyN736QoizAenyu1KNjUDl7szJDtbfyKC2yZ
NLQS11WNJzEGFNn//VcZmV3XX/n+adqLlQgAl2mvxQY14peGBVCLuk+Q48KT95jo
ixPoUNz8KGzCnGt3sFc7bvkh/HU/pDoQXtrTjB9xi6VNhbHXLifCaEGShTUwX+Sk
xkNkK98U/FwWzuCa1f5YpMWeQudrAVzwV1lmP7AdqTUR20rghk48V5Pv/nDvHabs
9l0ipCwiehl35FdLiQcJ9xEKu4zvMGqXWXXKPkINShS2P8wo1PFEKxEoIi2yRGCm
su/mnqh7iPJRW0YBVdezJdVuVglC560EUqRIBWQMSkK1/MGxgaacKak7QNLvug+j
RKxWj2wLcKP+SUdFgd+Iluq6wSw90tatfjY0mA6olBiMg5AJ4MloC9ft+P1TIbbg
miJuXCmyGpGp9VWBnDIut2d2ZQI9KHNWIaKRh17mi9oIem5GoAqcpse8K11p2m/l
ruCv1vy/3ifQn8f4pld4AnIRBJDGkYcxtEWLley0VDxvgFKHq7DePR4dtpJFoSyv
nJLu+TfAl1RuIS/gjoDhU8SwhXao9/apD97bbpkoh+FAgGaWFBIEeX9U6ivwBh/v
uqHbEFUbijxkGhxhleczgW1j5za1VOVVJ9oFirnZ2gRtOBW99SMOjMeQRe54FYVw
e5VZqoxd3e6EWpTtuPU83ShpHnKpoLtr07/qaGe43z1Xje84CuBbxfsWHG0HxmkO
DHZW3hWJJ/mW+jt1LrYmKEC4wtpXy2Fo/cruMu7qZmi4RLU7XBUmf+XnfFVxfs1E
1rbjIgUAnqyLISEc+RJGBRCQeTaPwCQPNzdQfJgVi3CXDHSmYnW91eQTCFF7sqeY
zA9Wo289S1EpnazXvNi2b8YpgaJpfdbIX5cB1IkKxE+Temnn+7G8yt0Sz0/yzIP7
VKmCEJYDsm+1GFCrA2zRWAbD7cZVlGhNb10UTq62pU29Tuw2/q0+HdDN8tuhpEVW
jIWZgMbXBCwlQg28QaLEOpDIm6JsT0Z0oLtGWAyVX4Hj81rc+/JPnZMXNTQ/rahM
/U+KeJAVzefgUSsskciWk5encEl5QYp03znZkW44a5AGsQB+77TNOjrPcdtq8aPO
RlVmZzOngQ5wApLZ3a/HH2ThimGDC7Jq6pbH8twgokFuCU9Ue0bbJrHBW2QeFOaK
Oa1Jz9V3JFqBQIEPMSv/Y9B6/GQEZnME5GbnUvQBzsUzX2ulPIGM2Gby7vGd2bz4
Vp830+ildAoJM6G1U1rx/Q1WK4iHoTM8F9yrtP5WyYklezEOMmMoKzh+ig+DXzS2
k0XHXcoLobM8tvj24FTgCqZmWhV79X+u8k3sPWyiKN6iS3wENPIOLBaazfW7MLsd
en4dMGCStTgkq/CaWzXUBEduen4iZ6tMdNXAiKfqq/SROWoMH+ezNzNOZQvcNNl5
BPYG+3XN3r5Fg37wriNuNvFhpAg4Cg0VXl1/n6hwN0BCNhMiBmPrqPTaJ1ZM8na0
kIJBmkMeRT5led8lI/fgedIiwpI+05Mxv+sR1kjlVh8F94DncaPOU3q2YnelNag9
z5ye2lGLrmBgdI6SmZDNi91bZo74xPFxwQETYymbDRhgPqPnY/4y4UjaX+Uz/Eg/
u/vKiR1Xt2kLycJZdtuWQTlj46ypozF0i0bL9gmwKw/iEbyAcia55/l/pam3Agw2
amCmAOra/jViYeBr8ElhlX91rDiU2FTkjee2oSZYnj7+JsNxMEWj556GUp9PtfNC
GM7y7yxsNxY7AN1umrsna81UNIrEe5F/5LgELKu5jhm5ag3nCfh+JGZM/b2niN2V
k2p240rbeS4fH6Rm34+3ExMYuVmN1EV8roWMBblspqgo0qUBtoASX2KLQ7Q8taPL
blmK2w97ZECSmxaRQjW4tItxiaophbpEqzJcmZ1dnLZXghX+7GleNMQaxA/YB3m5
/4zuMT+ntr38TpCzleRLPjqYyNQJIQXYP2uBy7BkD/uF83mxYgunZX4jyfeSC+Fa
VUv+rA9O3uR+OesRWE16VrZ3+dVZUDqIPoVcUByz+FVktnoGQemqhi47ex+LUbHr
ISVj22s2FO4ANU49pLwMfRUUA4HIbypvHxFnFSboNUvNrKGe1nwecQByQRYH6GJ4
//t6U4QGAIzjo2KT+FCfSs9W910k8U4M+J6g3d2w1ig0d/xAVOMqq6Jmx+tOkjW8
BujHVKUA2KEjLnPyfcLg8DTzHfZC0iLSYq3PNixGtlZVyyHERaRNW/K/cQkPvoiG
auZ7ufZR4l8cb9ZMDqG4l4I/bkZx/JbIpt0CYjp+LE54nu732N3uNyEwv8WO9B6o
pUq2IVqy+jAYtHesLYht9LBapI8dEpALTb2osvsi7TJmKAlmsuGOFSJXdRS/MiEc
mVp5g1JxiV82eD+tbokDB73NxInukNYefphv7WiOksGGDmXn04MVJfqLeOantNgB
XxnD1dEYyWvoCT+DwkA3r+I/Eg8Wx5i/njNAFScl/v0R9KeINevW7Q3FfGFwbw3z
y7RPqUYIIREMjcf8VjxEMnTMUTTFWXHPJRevPNFTW0oSC3tT0mnkoxpikA2uFxbR
aKODj/POOlq2aYhQW5PYrRrexy+uCeNzkNsW2voGmHFhqhRbnmoMxFgvxfvyU4t9
pQqv2gXxUCG25YO1jfFMUU4PHHUJrR31rWzWGbA9oJFGitqRQrbUxytvZ9sU0JRB
nFBR2s9CPWKj27ONFa9/lwbZKVXr4dAtkt99oGxhZ5mJbI7whvDl5bNs5XYxJncQ
knyUfH+iO5y/37saDhP9JlxzazUH2KzfMaajlZTu9S5VgCXeEVlFKUNFLCn1j3Jp
vMb+/dkcPRqLjz7bM7t4DGfM1Bo1bc0pDwv7vRIth4IoL4a/j1QdyX/CtE4J99Le
t36qYGXyMureOajzxcqgRA7bA+6R2RzEhiL3YPPAZvxiJV0X7+P6SzYrLlTKdc14
WbMuS1d1q72qz4fouExMeUkxgaTGT000AbXRTjzfwyA5rGmr/M3VvUYyGqojLqQs
r8OkDUNEcVBU1KP6d1N4Au+RNRViiupQ2kY/05kUz5jRPs9h1lyH5qikxjlwS0mw
tpIiAiaroMPySyt72Uo5AngH0CEHLrWNdo8oiLEeNrYn3tTxYgzg1sWWO7/y1WK/
LQmddZ31WOolWJ/ZAK09XmhiQ8i/RgtUjtcRPfN7X+F04DPDhi8tPKTYJFmoZ2TF
jOM2sfJuw1WQNQKdx0vDDcCYCrJIJUjBKrmxfr48Rx/1hRU4z7KZg9gMEZASi1pS
k7RK1ZFRdXcyl6K+9NsGYeyZ7uD9EovsOIH0P40ONQRWnCjUQ1oPQABVKiFHM0ha
4bblBl3v5f9pF0c429Dl9VLcgVfWZT7g/cr3fKZbn3VxxLcK09oeXoMjUiJ3Ff3m
C9sVACtRxFs+QQ/PRuF4WQQQ29wUQbfvnFpz7x/UOOj1Uh6fbgjlVMmBGxq63NAV
20bbHJscYkJVoS+6bgYmRtByGho//iyUzbMn8yQ0KuG8CvSNBN1awm8+IX546nZy
6BWnDrrTHLmlyx3YxElAEOlT/1raxP5W3X7WSWT9owuhS4LM6CEbhWwqwmJKvzTM
9BghPFBDlpnXaXaMZCGJqe2B78TQ3M0JrC4NdnaokB5KMPtaBx/+xuWcYWgC43ra
ehAxVSb8f5Zv34/pR71XZq+CbMpQ3u6VhxJhHwAQRf6tOE2NoU6nDInmuXhQvXvs
j6nv+4Dm69ffucF9VzygJPPUS55Lyn/aqtu3M2duXctx4WZ7pBkjCIatYt3fkpsA
Y/ve0dobcswL3XLU//Is/4M37iuM1Jma+zmhQ8Fvr86al4XY+KG/CMJCOgrlBuaJ
RNgL1n+BfsbIpV0hICH2j/CL0yCUZ8ZdPG1oCVXuoQeUUV/NHLIMDToHGjv5bCHi
QpVXx3yQGzdobiCjXaL6eygPKFmiPsV5bo1eviX1zT5NJFEERg9Op+Y8PBmRgnBA
IBtsnehtMze6qjjOnSlb84xqVPS3J/G+d4RTbCqmf4IZ4XwfWJK9JzztkTtVvp7N
Lv6zfETzTyckbmlqNeDWCJ/JVJlUJcMTY5Ojxae+g3Q7xbTbgCBft8Wu4zPxlC5n
HwfGkhHPQlOonNIyyCUEvR8cQ4vAYvA78KiaJj/t0OIkXdhp2H+Laz7S78wN3SMo
bK5G9ZA8QY347A8hAI0a8JfrlX9WE1UqE5KAz1JXa1oQFu6Ei/DQYXL9UAGBzCcm
PBfh/3gJKZqVzWWRIEfMbEzaOH4/fkv9ZhQmRRuD5Z/fO7AB9t0Ckb2M5NqUk7dr
oBV+KZdT7VJWcnqesLdiicPNk0AdnFz8PVre9gfG7g4iraEJ03y4zCUiWpuTczQo
xbVBAieRRlDki0VxiZ8pP/ugIiQIrkY5uOH8HSvgQNcQ2P1Py1GTElxs1OHicHFd
yPqDvLEyWLZ0l7j4KK3yR8S3e41k17rlX92lrHH4mQVzNIkXjGMQ5hHHc6W3B3GZ
vT0yXqJk0sM8i+YFHL2a8dPkqPHAOzIioRUJW1YJW21N9ePudfLTB8FK/2iO1y0R
t28M9ylaWrHj5ZqiUJapcIRQ8ROPmUkYmRomvf9Y/mxGco7qGThTGTzVUGdowsQV
bhAeTaO/EkbAxXezQE7g4CMMXRgfSi9ponrcv7pSyuTCdU1MfDQybT48yRqP12s/
qGQw4+PtK/ymQTXc86iYwygbfffKMi+lmAPbhC+s6xz2GSFodRx403HcITtdJja7
erEEyV7E2XkwOD7B149iaiQfHoOrtUW0gDjs0p40BlJoZEEGrHB+2+tF6REYgfZ4
73Qmi/9j41+XjDzLMRvOoTV31ZnGys1NBfta78vsjrGH6oKXIh69IzbXv+R4GiwW
IY9/JtSxQdA+8FgYK9oiCw0bgTCVFvMl7364y8IHuxn0RtQakanVIXsyeYaEhyEb
A6KJqP2ihUKi27Hrpf24JUkushvLpILk0lMtXahJpcxIt06myalj/bffnd24Ffws
CzIqC7akphQA0zrK98q9jbYMo2m3uQ1EaN+3Qsa0Q8USqpeawKSwC7wCt4BdVYnn
boon1iwTb6ES47ge+RaaCFzltrFb2H4NS3/Q5bu0l6BtwBgvdXTmTISSrN6JRpjJ
QL7pavzuTvWyXtKyKAd7NK+TjMFqKD9CZTSP2VjfvpKQn8WlFDdIW6iV8ndnHaWp
vjA9XTiUM3cEKhM/PyLwk+Tlbl7k6+j6pH37iZQr1z+/NgiFH4a5s9F+lemPJIGm
Btff41LwRbDaVymoiAVE2qejUqTk491lphmBTKMU5iJ0d9bnaaOP50ASScWRq7He
dwyx9SYwqXBcNHHQpqF2yLBemRgTvRuk6bibpaE3QpcIRMlJ04gNLE4CJntzuhid
Xh1h+7/oZGB/RdrBXTwKWwRfGkzfdgptrQRrtd4yEN6UMoGFDUwCFVZRWJw+BJl0
Hf2phsSwhzoWNjREK3UfUpYVgeGamCP0sFk+QiAXUmqEggMbC/h1hlf+74t2no5R
pQeORwALojef949S92Rr/DsxCwurcg0ZGDOrS01rljgObmfLSeUtqxAZoyyYbwV8
IV72dQPOPDuRifBotOoA/GhQJJtuxZNSqNoLDCS/shy0+h0SFzl4tSB/dYzxHEbr
HNZHcLln/1Fuqdl0w5YGa3NadcLCwRb46Log/OJ/6rI8dDN/xU8tGs1aWZAzvc6t
oqan5LtmzVHd3eHy743U8a46Ba1nI3i88YKUTtaPDZsknP9psWomp7c0Q/kOaMch
FPPHj5gZ8DIkBmoJtHtPZy6ii+Yrudb7p5FKPLSX3t5SiJHhWX8n6X9Fbst9ti8V
UwLpagL6b4+9votYH9CYemPD+q4ZfX1DNaZqKQ90+GyMypGOUL6aSfAmsTA1bHVY
PU3mLrsiC0b24X1dcsk1XmjgoJjQHbXuH32aPSYNHQi20Mc7UOiIRiyMak40OvLx
pA5e6EmOso/V19T2Ne9rgVIcKVIa65naK1FDhRTY7TQiLBocUmxqk4GFFxjWIQTr
D6csbJyiUWjXA8IwMUsD7WwJTJHRt1xSkpMNBDKrphEtx0jjU3xBTt/4pI/tWQfc
92YE7Db/Yv5k6PohetNI93ro9i6UCYTYOz3alEo/LgfYbyNTH95Aq3dVNUYeK/Ae
PY8PdVqfWA5h5e47A7xzoWITpUUVsuRvWU+LilZQ9jIN+Cipy+R0hWj3vAQZfQH8
yVqnoEKk0ud+ZtPLQ4OGxZb/rCuxATFUWcMkr4/FUl9BWZnGKpKcCPJzuaxEAdD9
xUyi3eADJl5/eRS2DP9u4Rbego8KK4Ru3PGHyH864X9PfXeCvJpk/kpqaxD050wo
i3/9fpgizYGWnAXNDgXgWeOPCFrnWOX0mJdV6OkIv/SzjRZ1FmCX4kky6+cm0wjq
A7cIxyUKyyNW7mJPoTNv9eaM2WIfkMqHrPLE28+SAUuk/bVP0RJqmmbS2uDD/3fi
Ft9yhViBZtZGNuO44FbDcUvGFAoZ/I5FGopWtkB0x2/0tg1Jm5faR0jV5+/aOylx
RZPBKTNuizmBNYx5JYit7Eq8mXRzll+6Duls7QF8hUdfm+xR17aOm1J+P6v2USlQ
kcUfglpHIMWi9o46Vu26mVPEz1Wq422ywCKJS4lSupfZw/Byp1ro0X96ADUlATxv
6nACzBnIH7i6EyWWS/rGypf8ghKsZuEwnswGeAPe5iVOn+b7QSIQbFhr7YbRVZKE
SInAp6U59R2vhrJ9L85Xv7i5HE9m77nTgKg/GZLCJmQsCZSMc9hP6faib1/GWVDr
06l9gutLD97W4YKpmaTvaijhReDqRmI5kl643YHrm0XHnYJ1kJwdBgp7llLg08In
WeTT/yAD0I3/SHp71V2H279DFTJvEB2UNivJauXmYQ5FOz5HLLGW+OzrN4hSbCiV
yNI6UUgp7QGI+951naykX9RjMyN3eanyi8HfgmTyo2qKyq0uWUcxg7pMapbEAG0S
cldhFLRIckeejTRWzYpksH2/3pAprVvnJcoGGfVmDHBhq2+qcVOophQpA8AITDH2
kW8DMoAIPgX1RLr+b2ROszk9Eth+XSqCAEjl9PQHcIYwo8HSTlntv1RHq20BAfUg
QF+UjzToy+lYqySAsr0UpIN3Usb2ojPC6U/yMQBIRo8NEygoLPOnvY0kZsq5Q/7z
YQcNSWBPk2hhqwhvPLsuSMUPo9OWlyVWsn/X4l6dl6b8hVa74yyOO65/OI3UUVu8
f94LWionpuB8LQ+jfrCxh6Ve4SJjWbUg97uhffLEHEzLP24ihv6BJPCRuX9HZrTU
Gexjp45FPWRh1v8WaZjBBMOkVgA9K2I6JrOn8frnkN6oCPw9NBgRxPg+o6A2dIsS
ToAzwT9YuuiBzUw8+zoOWQr7NEpWZ3YoCbI80g9oF3BMgEOzqUwgysA5lcn7ZAFN
hk6Zk9Pd1zJMwpGgP4Lo8ylrY45M/rmMgnl7a3PWHTylXFKrbQccSLK6CSUIeJ65
kgOcRzT8Qpd505vO8MDF1U1bg6o+MRxmePhNLEpYVqXXaeCXMnVk5KMfm7Escyb3
bnTTtVkqdjdXKSey2euvNDwAU9bk5vPP7B/brqj72CWc5Ya4a3HBIXpdguDJeX9S
kd8Wpz1QCD6iNz1Kc5c6VorxKDWVZww2UZ+9YmNdoc+VUHZuGDtODxc3N4KHrJ8u
cevdNi2DkD9aeIJNCkzXAiy72psT6EMpMzikBoo1imKgxKHLMg1EBVemr28XfNMz
g9C0A6Hl8B1X95WuMMwa8tzPi1KQFTgmhajIFmyPVUVe5DsdSZPSmuFHvWeXRPy1
0HFsu01FyyOKikrXcjSPfGKdfwqTMJ/GuE/OC6NFP6wxeCu0GMhpgwIGVsv3tthy
Qg9f1nzCmYk8FaTOOzZsBwcJVrEaZPYFEPlcjuGQcGaW093Scxy2sgTAqeYbMTjQ
nOrawmFZM0ZJ0Yq3S4y3eKTyQaX0HIem3wNyF0IY9fRoWJuaM6bYPqHIJa6GOl5V
ijdIQrBd5pCVyG4soHBUIkugNoqaa/5hzUxvCyxr16hPlUhVk8ldRTzha0K//MYr
dzC9zuH+cSBEH80Q23aVMe+yy6atZd7fuhnnHx2+Q98yQtVX/HzvdR5SYHNxFzCw
I5izyT6KhkDd+RN7qC5L5GZq7+w9Y0rm6ei91xNVuPXu2inMuq3W8fpUJuRwmxSS
JzcDgODpeoJK/r+Q6TnoIXVdgmFPIWx5rKeX4SxompBH+Eq5xER0wMGPpbHdF+lW
raEkAra8PJsNeXlsIp0PIej4wHmrtsVwKliSCyb7DifRCbwFawrGd2rZMql5ip/v
VeWVFiluHN1/ptPa23R0BRddcyTo109OhJdxadnKhBeTQtB70joLSnt8W0qVO3H7
Sc1S9V7wl2Fv1pVT/vCEJhHpS0CG0rlS7SzMCYstylyv4oJe3kEEINKxTdRTZJB5
Dbzbdk5OhDVkoGDO7aRa9hjiRD8uUpW9Lk0rhMfuCRowuKFfQDNE4CvFgzKEAWIS
UE46JGCfYgTPalxDHLi+HXnNwIb/J2vhyW35J6z1x/OnZakpYg0JqptPD7AzlVl9
qfRsZNPmbvmcCjizECs1bnvcHQC+iFpTUDCVEvttnvsBjjf7DUyXWG53jAFB+DjY
9NiQepH4tlB2/lHItOXMpCJP2dSpaWNtszOJFW5bzSGrSrjdNLqlS28oo+iNK0sQ
wCrLjS6moHtMU98bjqPp56eeVWMwHljZYljCW+JG61F+0KvV91ArFIMNSAc0UvMb
jbDF0VRkEv2vhovhrVWyuLU81SBQF+O6hjSWFdxMzHZ1HEDY2rWD5gaCMFHFBwcW
OKFdk7vU0bHK9DGjlrFnHqcI9hOMy8pjaxBHW/Pw9sIosgwOyUYyrf4HC1bSGA3n
JnEpc0foo1KnREwsjREf9r1hFfQDRDLx4cn6/UxPuZnXzFacgWF7emLNtbw4sCrf
V/kFeoSdAyBg+6gM9HZQFOw6+xRvE2XT7Qq39dlKA1cCY2UADV8LyP0zfPTg1Gq+
UtnBmjtpN+5a1cF0Ya8x55EmttTGdzOD/2sQbbtp55T4Ht7t4Qe6dr9GOGWnP67c
JGZs3yq+nuEM0AqMVMK7CPl1MO4m6vUKwbvARI7zlb6Rh6Okp1pDXnE4+rFKCqdN
gDYRUFvEb7gw9GXfn2aguO7foPSJ5HvkODWGhwAVBly5TztFTFIUeHYht2nvPs26
Uh0krLiGwVYZ8Xx/S1GoLhQXc9eXFN72Kt3zbWgYYjwLhiLLshx4hJQ4HNbqaJX4
a0emIM9umYwXek/R10O9G09RMIq+LW7s/T41/Kqav2spheSFD1Cs2qlTAI5mSMQJ
7PdPuWVUx9AuQhEJPJV8/rGL3IEv2fI1JkKwQ5OpMZIqlXx/rBgglJFD9oB4lCjF
3b1JhsOmYGe3//qmzcCJ+v4uBDNWKO45acqVIIoyb9W8luGRXZgJY6+HPGPKeJQy
TwbPSxoPbHg3pDO4AopjO4givXwch5Q1j6N/TWt2vaWxhyDeBkUJ50aTOD62bZoE
jR32pFAQSXDlwSOKustxnL4yq8Wh444qg+3Hbw7gp2+Mb4UgNiTI6EWcqFTAyZsQ
g3vgRlpmlLj8mMmwNt9uaN185hix6ydgO52ASMCibcB4b1Mi/sgwrKkiRSVQLRDq
hqG7PspVGiRccVWazMU0KBaXQCHpBAFAjy8pc2NlT1M1ptZTaUWR7I2BcXCJ+lV3
vBrImvPZwTUNbQh8l8a9nfq3HkjFQsXmTi1XqUkumV1cnKycbCV5ndonv8U8ZU6W
GKXchxk126tbdM7dNWsRJMHnqmwSk+Zt6+V3CUdDEfOav1WejGD3SD0pcrBRqUqz
Hgk/7/rIA7Sa63L/qg1o3QKOIeiIbtZZRnM8z4rWeLV2SNTh7tGS2qsLD6lkeRea
t0VMRiZr4T2MuWfGN2US4QhgNN8xk9wOCMI/enxoX4GnJxd3EBzWYmm1kbJp+VSx
Ti5SMrH7QlK66U0FwhhU7HKHR0EVlRyooCxO+cjz8VKzh5P30VG8CqM96VuHqqQr
DXvrHDSRjw7rbNjR4dbDw1JhYoMJ6CwfMAc2XDCeRo5kyPHD0DtAtHbo/eeVWJOV
ckTKrEQXaFeDhGoF3Yq4kznqyt+QBeJHzZF4hscTbDSmdQsSmOamewl0wt6a/VLh
dl03eqmJdHqRPq8Oq1SzE1LsdBYm5nZyUaeYh9g/JVJUKT6IXQ5T8maxb6LcEPDz
RqBOdWVln2VU8F/Jja60HOVNDxWdUSA4txoOSAomCm9eHfxFds3z3+t3iTqoH2tR
JKkHNfABtBbDhpoOswbqZ6hs81KLG8xRNKNoytDMeHvEmXv07Lw9xJ0C8ve2d6YU
WvAMubOs6cAFK0AvqQA5ACofABbdPIHb2fZdnmLw6M9xiBxZebXNZREGf6Ktb3vj
qd4febBLldPjDfEo2A/CS5IXhzweumxzZLWMh//8WfffnTO5CHseJq7AradAcOum
7nZAv1jNzw4aI64VcFWtU1J4ruk9+hePG2EKxuv93Dp4a5rFfEWo2fA44HamR36+
M9ya+wVjQEO+6k1Y4J63uXAIWA+OTi7ZtajFkzdWi15Oj3A8l8HBbk57Vfq012oj
7ZfgylGL+0Z1HdXifUfDgwbHwmfUnJWdJ/RFyUrIEnf5DsK3OlJgxnfM2b5I4QJr
1gxXxB7ytlLi9yNsm2zxBhPflk+Nst7GIu//HpmEpjpFbxMx9dk8ebBOPqJxpCfK
uCzZrt+k1LK2Vm2TXFoL6jMp94uduxlAC46nEHpqely2vsfdB7c7KyM03/gCT+I/
Ej0DiugW5NfUlEqFOzKt10VS9dNs+HfHfRx69t32Qbj7dCirThrGawWGAnimsWFy
ve1TgRVBVcOL+Q+onomOv4t+Ms5DBPxy8uqZtDApJz4teverFjGkhjP6C2sG4fSv
wR0e6UwX7ABGJcNWt+DtMbSXYlRHoXi8LOrf8TsbBXWdR8tPsH9MUieFp+dSQPa6
X2O3AHFI6RC4pktr0gLosJwWQ8OqDexGzf27JvrcZhvg4FZKBB21lWSDubO00pBU
iTbBelG3OxkW9HOMglUEsU6D2hnRC5LfIp1459qT1swpd/eMURGQgH3FAu/yeE/m
uGy/S0Djl8GyMnVKhIM2VuvpQPsrehwny1UHHchMZ4fw2j38eZRp8b+LNMNDWUmL
75TDVLOoC0jpf0pqFu1chpSZkT2JqmCKI7+WTYBbcjJ/NQDTf3QhnUCa3Gzzi4ha
JI4VSCjfYGnB9us7Yi3uzD6x4XBAVsPoFOahZAmIDuqS/UKuY9JdN8b8DTFEQt/O
+zUrFO35mie/TSGcCGQqgVDNmzTBceKmCNhrQfhVj04rkMcReuW5a8tZSddRu3PC
OBKc/PzLjycBBNscqO+x10aRtGuhR+nmmtNZO65S0Ms+1hgLrJSaLKuxRt4IGZn2
IP/4vbeZGtWNqoEbph2qYqocqe1m/VyAk9sA34wosDwJOm71+IPwtJxZPAzB+4Aw
ZZzYjPccvGO2+dVEMa3Qr8cE3k/TBidELEVb8U+2H4RSRQd08S7VPi6SJqoPaE+8
3cydrwg76mYsZo6WX5Sl1D9wT9UPj0T6oB8qJCW3VEhNyUlSD0R1Ug8nFFOoXnai
rFuYjm/v141tKMF8t3Ua+N9YsaHj7HE70S71os1RQbyEtXkNbWoJGJL7tFfQ34+j
mvyH+tDPo8dIWp+Z5Jq1JYKO7wRNkqJilCFH/xGHZrnnlJk1HVumem0YRqVxG3NF
ja+N0mPYq4GZJdLu4FPc89zCLiqwsGmGzaLdbZ/XUePjoU4xX8+gE+ev66pxM6uv
OPKQDXDcWGARACQvEi8/ppsWmtEgJXkD0xsNyeLZEZjquOjDiLPp6KYhH12zEtPD
RObpIWXMizFWfmmjks753K30MizE1ZNfDUoRH8dtu2Gdv/4iUQL0goj/jWqqmMlQ
jOOuoFHjFdE5hIfCUGIO/mq6p4SctQOzCGyFsbchicvYJVUlJF12vpo/4RPVwezy
9Z7zRAZ4EEiI4xOt+Lqb02gR/3MVnJlfWQyB85529s33XjwugQxfykDtqE9/ruOf
K4C9H0qSOnav1iFoVrltO5VKRbqWgc3mCjkb1o+scm8vzmFWskuziHQH2adIUzc9
ANSqBAK/Hsi7vh0aaJ6CyjqA+dWwCy/hMXf/bi6a0gpcnlzM7zJuqass3JeiOWje
UVfuFipibYbLOPBw1ooSHzQulGK79OZE3h7DBSbLlHLsl6lkSwq/aSWCu8f9ChPB
Izebr19KxYeyY8LaikNHdpqkyg5Zq2P8DpQs40WnY0eU5LGTK4Lw6BgdKOjSPx0N
qxcJGbvyJTNPNmo2njKcJGj1z6cqMUPzI6wnSpCoqNRMiy/W5pJIkaY5xPupAfeO
vAxFQ50Y9p7c38Vve4q5ILL9NEX+rFZb+xbUpVnsszckrICbAOw6tF2TJRoPwqY0
6pT0gnRoGwNhsZXEq7QhXhLl4KX+FErroddzqMymuGlTaydcygj5dEUW0rOjvTZ9
TJSaf3aaMayz/5bB93tNWPROsl58YcScX5TzknGQlDplzjjq8kJ/VLIz13NdggJW
Ku7grf1xeV3+DZUdT8SWXv1zBWTHp0jpRs0bVKtkly9sQa05GHuIxoDIa4gzZQ3r
rOo0vyM+/Bz6vMO9AD20tT4kP2l9RJ6qVnXEC2pNq7oIydmOobGZ6T8FV86sAm3v
UybfeuSGjd4UpKX2eHCdvyT156+8bayo3jVttbP8+0p1hZWNEPHveLY3PhTdeo3r
YAZJU7IF4XDZiPThsaJd5FBxKBY7YK9OjX2nMg+yY7KYP62jeMmadSaipmGe/4ej
5Tzfb5EhacYRmNkXg2vsuk/ZOCzcW+Ld4hDC0+hncn/d+txSXU5PJ7DkW3zKEnEO
izbpO17/0mo04iZ6GyE2v7o/93+V//yBUJSY6p2S3pyVkS4/XOY92o+KfUdC6PqN
r/ixbUjsnlK+LcJrAw//R3iiZvH3l5MrZjIMF1Df5dOWhnoznQ/pn4Rfl+GRV+SP
f3k+AbLEfPkzEFkuKr4Iu6WkgUr3Nw0x0Tvf4/8kuOmqIgpeZk7oTzigxnt9AlX4
qBUW/1pLTRAZ1/BGwR7H8cu1ly4Efb6JeA2QRRKVmgU8xvbBcupWxYW8UrIxB92P
wxdLbxfnnfEqMW7Lp7uOFuRBQwb5xylgbyE3kZInqoT+rR1WcvXt6c1pz4g0P+ei
ovroX/BBNBRvOxW/MCEJAIT/vw0QndPSBa71ua04/RNnKAhrcukKib1s2uX1oTQ2
pUW/rGYGeYOv92mEKOMQrLHkgMk3epma0U5YkreaazSyvcZAp0HPE1WL5txIBtvq
UZ3M+Hfkdo1tNdIjJc9L83oSNH/RQhwPrcYyOf9WNVfTtLeIsJfWwwGL/ah4TdHi
1xNQXMPPK4LTD1CC/4zxEFzPtQ5m0cUaxjaCY9LR1YY39HCCytuqIoqpoGvaN4sr
KgOWRfUe2wJ+RcLwahumaDGlA0Iv4mJoK65pD6SpHH/7GAcWoMapV1Q5yCaoRyG/
12Oc8DlkFNakj5BWpjI6DIoDrQZrmKHUou+AG7G2YzKxJGp7WodixLhmw386kcki
Ou0FMizcp4E6LdsWP4ZUJpeQuMSFw4HMxaI1kE+VOrTCzRGPlXq/IIWMnf7V79x7
5ulVYoJ1ScXNhgQN3F4YOT8iAoQPkUBM0JsStex/dhU8225Y2dqZ1WWuqyAlHm4u
dK0lOY+1Z0U99nadmSJAguhHpbCHMZJ5fGd0u2HKzpQpfasCCpf6CHR2Foez4uID
S0Th+x7MgmPmRtv2uH5PxjOz3aII1w6bSOyq894MdOlLIjkulnbHq7rvq1cNcqNy
z9byJIpRnQNQERI+Cc45na4GUGyuJKNqJ3hzW0r0McxdGNnVXuTdQRYTR1My6e5V
nUjWVDnQ6zPls5YlNqIh2frxLHS3NPk7GU2f1y6YH8t0fHQVxxgFN0QK/oCDmLLL
8+kxaio7EzjdWz4cdIwCb31GVlL7cSe1fydyNA133uZiyBUclcg/sU3p1FaeO60a
QdPhVyw/jX/PtLmkG2E94r4ISEV4WmL/Tcja66Y1cCaDtp8iJj84PJGO8i85wW5V
7khA3ln3QCKhLonmm38l86i+qhaPXK5LnMtsITqZf1Ua32iPol8UyzMqlxIjt0QF
JBpIyeG182O8cz3niLl1gMWNZxueEiAHu4j8EsCJcZPRa4Q2uiic4TyjUDO3wxPQ
oNlGvP+pcvzYl4jVniVfQvviMV67d3AmI3eQXmm7zJpjeMEdj1ytBgiqsDfqnsum
niDEJFzbgQYfCDLAmKz5XJlHjyceidCo4MW1RFWCYBoL/sU3NTTB+Yh4SRQ4IArn
lma19HfY6TCO34EHjBVPpPiVziVzJDZLwa6h/+e8X5KXGDU/Vx89/Yk+5GBW71RQ
mEnXqUhCit0rlGCSGk06XatrEXLEoEGbt5nYqbsTxWLpvcvs5qQW+vFY6kXe3LPp
BD3McbqZ9yA9+lTNGubOxaGBN2LMRXEn/Xn86RB8lMar40g/zyPCMnxGbPzfUmW3
S/Jl4LTCIhYFRvFWFbpdVtmDoDQfze5JMOOMZ+PNe4OZkNM+ua1EqW1g0Z78ESXY
YKQ90aJV6j5/peBBcETWA8TANxAgH4fmNtPv7hKhy0GVYG1AIcz/R83aKQbe6uH4
XskhigtpvBGqejSe28r0Ju0tDMiPf8uCHXSkEkwoFsA0nzDOHoWhotoYlIr9mfad
eEjuI46sPrG5jr5lpWBBnjkdB06D6HIpgvW32locrSnSJ9lqwpaysyvZCl9ER78E
+qJqATOw6RdcXji8zzwPqt3OMppYuo38tDKQpjUdCOB7JlMA9hwUvdMMv5rQU5RQ
91CkX+Z79F323k+8L+qXZsVO2bHqAXlWTJA8Wz8a6WKMVP8Hi+rTqGfLTLrVmimV
4aqW1SBkOVMoz3/7jB0Da3hT7WrFC+qGi2V9ybw5AaUiQi97U+a7QIz+SAvfK7sI
PFNKbWimm7ZPt/NrAthkyMKm9fAIGr0SHqahj9BQMyAtI6v7NwTl12i3xp69Zb1U
rTMrxGBN7zzmN+Xb780N29X+Kz7MTqX0uXny9kF81BPVOwAME6/NAOemPOtbEFix
6hvXHDuUMt7RVjvvxPp8tz2cvXB73rK5Z6F49tmmrjuzYYJkytkb4HRU0m6fUznO
MGSiFf8ypt0djj+Aq/ayPogO/lSV4FQ17NOUTITOzt2aVx9+BJbmQzMXr5zsAp1E
83R0fPTAD3L/5MEMx5kHYVoCkCZh0buLlaXaWq/H1G1o7hTwlVTYJzTP3ODRagwT
gH4+Qi3FwYLQjpQydGozCsAfG8NPlcu8ppcDe5hliG/4TE6J7roc2R7GDVNisUNi
EKPQmsR/Vk7N45cojHx9HIx4G2u6+wZcHNRvXm8XhQsVkJYxnEIeHvK27Bb8yNYA
Tt7P1kh59SAwYC3Bg9YZD5Vwcp29OklRDGSKO4baSWJwGy0B+HydnkdHk0DbxaoD
+jUrUf2qqYH7uaVeYORodhZGFx4nVIkrTzFs3PmfN8pVeAg9/p8Mv/gjG/2svo+w
VeQh4QGBHcjV13EObeJDvfkTiYLuAE5zeykvkKkH+D7fHC3JCSpar+R/AysSFbMA
f0YfUzfc/wGrLMcEmz+Eerg4sm2n6/qAQ+L/eXm6M0chS+viAW2VwEkDe4A98Yll
9VX7nlIyV9HORbenrnUWC5wuMB9HWumRK7q8QLmmpEQICWcFIykFOvhs8x9feGEp
RngE0GjeY4T6v4ypIryJIRX0xd0F3Kj7STefn90ZMi5XPE7KaeDVW3zRQR7nSeNE
sU+ULtFVIKvG9S24kk1gJi/Fe1TEA4Tzwx70ADMBIQuysE8o76ikX1eVxehF6EQU
oYoXc98xDjMBJ0up21k2UQDrTp6wl7I+bnArZXU1fHJm6/Shc6WmnCeUvdwmj1In
4XVmzIcT+4bx4fkdq+HGvUkUG/x8WJfWuRi4e9nulWjjgewJDaOEvhtb5ovtK1MP
0NY9NZOiULoQwMpy6SjcNVTr5PpTnuMN2RYJjZczJOVpyogdMvelmxrWD+FY7V+U
nyagHR4lqWhHCjdE1Ab+b5kD5h3a+FMtw3Wi9KTVafULXbsDWPmjOpjqXGcnGpYd
LsffZXc2vrCNCa4bbz+yse2yNf2FT6GE/Zi3/HB7+AQvka61BTYxwayam4NoVVwa
qPx6kILIWuC43Oeug3YBjwPqRa0KaAvs8efOXxWIyE6LcM5TEX0dhd0xJVDhBxFS
vyXCcRSKvg2v+oJ/l8un1nHYNxb3QoHEWswnBA86inkMVJPgxm+mLzle/bdJ7Y6q
QbqyNM5u+/0raDLAu56xJ/OoUR3nUFSISxSgbjqbCci+nfHio/z2HabY/nFFG39H
auWMbi1FCs9+AOQJC6SXi4WcyobpwHEp+VrNhDYjirddIH31jeY3P6hZsPbksloV
KNr1W43ZzXyl9AYdA2UNO+DsWMRgHbzvy0ZzLIPp5UCFKOBb7HWHlfDaEPK2pxQO
Xvv83c7TCHlxOOxxrqIURqEP7efhZrJ7rj/IIIjpB/M8WMGun77BDFjx9txj2Cjm
W1HjqHn/zIgSN4rMKLDf3lzWT5dpoULqZ7RtjTflWzrz2x7HenFsppzVaoVn6KNm
ky0zj4bP6Eyg4oALds/qF8XKiGhs8xhAzo6tjU0op2rCu2AE0n2VS5AP732YRdvE
QMq8GVb2WrqCMetP7/28aavDQGISDpweepdnP/qz6mBAYmOG1oMOXrIJkdEdTjei
WnaAY8cMVjr4cN067rjkXNB2wVL/yohG7V5pe6jkV7qbyBxSwRtsKkrGGIbBk+0E
x+zDZrg+UzrP4jpXtTXcE5nz+0SFk2zRYM/wiyAkiELegSq9LJBqjhiAQBCJpdOu
jzTqXDm/evvMsY6UD8fmnHNu8I/wAKQqSv1J6KJ1QPJ3Bd94Dl08jqU9lVbF4z/u
/N+dqTc7b19Zr+R/mSwmCo4ih1Ec6Y2Em2LTHYa/Aawn1eSvryc9Jn2BBqnXwrqN
H95q0BKsznHcFNybnUbIhecIcq7Wu93wAyom99xvAIHjPbQUt0yf+Hx8gRap13my
q2pDN5klyWXOeBCpbXlBu5TzWoIqTHpMtg6aaa83H5iliuvNZnJlG3PiIIjEukvy
8vumiAd9YB6GfTjhVP4KSW0T5oGWTjDSxCuJNbWFrjWXS0Vz+YRUOuOAv36AY2ff
dBq3Fj42DEhU2mg4H0SortztWBFGaRO5MX0TQucfNS+7zOX4MbXSp/N6kdlpuL7B
ExNIv9gZlTXdACX7nPpx4xyQON1eVrYp/BoPbloVAqohkxE3dDLpfC1lXPTh+flf
gFxP6LZ4Xt1IE3y3ugCjriBWFJTRgyAyomFnrOZXctNeIlY3PYtYuu6SkCzl9kSM
wG6EUiNL1yygYiGthEeoMRE/lvSd4kkKp31bC56WsR6MaykXlhrk/harhTiwTl90
IUiNpxhtUrC5Y7o/E/V2oncjEF5C/pgs0CUP4aNHYXpni8zqlIWZE7yvzRuYMSqv
kQcJ3eRm/267+gh0Xhe7ABL0LbHQ31Rge7xDCGM71zyqB5IOgHtRkxVNxGgkcAhp
sDG8bfkMb+J6TUcvCYbhiZFYXu3Vj9g/205ODt3T6xK/b/ZvaPtGqvIxNWadL/2i
W8agJapdKTYPS1D3Hq/WJCYMsp4oBYWz8CjoVcEa4Sercf1B/JhXX3tjCPHq8P2i
Q/2vp+U7/xSIoDzIWx1lKhsrqE4d0mJbb68+BC7FFsrbiHB+tmmi30LAz80urrXh
k4d1VJeEFpfhYmHjURQHTFDNS1PA1Gp/HBiWsuc49a9VezYRTJd7W9a4qquaDzUL
6twKOob5/GGG9gF/HykhIK/h+u//DnvQYUXqghD0KzYPmGp8xBNQV6Ebp6SiQGMq
EacALBVeQXsiG41bsYjcARlR91gMqs1a5HPE47IMNM+Km0ON5itETfrmDxXZ15Lf
+IUFiYI2EWMhXvkhnw/fAk3pdZz8OkCKytyKRdAW+wBtuVIrgVfWlnXKJtMZOBYn
U/IoT1uus4w7fNxTv3ViFMvxF8G4McPEJEdK6CyPQnlpAn8l4U63mrmnPG/QCaAA
Qn+PJXJ8IkAhvn/ijcHWQ0TLko1cCgD/IWBVr+XLVvMsgB+J1AcsiMzev/eGag7Q
ybuGsoS0Hzt4NHTXXDjQdyztVW1PJ5vwyDwpgZbzcRx8CHgJ5pDWhtqh9IuRZEAu
F+MTUvu70ObaektulQfP6gI+dZSjnDQP7I4G78/XHBzbLE/97Ozzzg603+o1vUTd
s+4gb70EpRVBXrp+MfhjCUiDbKi6zAgyVBIvctcIw6CpA2/Q3tUu5YxfEtCS5qtv
SLuG/rVfy0nJ6fuqiXcXu6EVqq94nkqC7ZXr4LTWQZgTcNHFBzzAsJ+Chfj2VG6o
pYOQCMJxdgPbfz4anwN9dO8x/rSD1ENxspLCAUApxr7IOIjTVaxZg5be7wt3mWcD
3yHLdeLbH54kGBSt3le7V06xNR7+3bAOTBMyhlC4dRqmBH+pj6EhYGy4TyVzNbrV
s2AbVqxb6Du8X0Hy3bwhu+pnyuSN75hKuDgXC5uDJv6O/qG/nx5DdvxQkyuGaB45
Ui00k96FMBApK4P95gn9bAb+L6OSgLpvsJfPvhtv6ot58xGukoHgvcC/fI6wu7oa
5TKnRuNlGMy5Vgju/QwIVhcVUapi760K0YDfLIlhnXK8dOmTGIR7RbOOqZnFI4id
fpMDXiBed0IPY0cFHs5oA+ylniqiy8zpHF1cydvnjpF2vei8wX8VMLJaExg6GANW
vJtG5yAiTrWTU586fgh3Qmk+XPOLdsHy1hojMi74a8wJtXlWi+kc8vj4kKgWYFh6
uLzzG/GbXy1w9lSAbQwxuffQpQgFZk6kcDMd1epGCnaZvzlyxb1b0w9rHg1mfvru
wVThx8kfnxhnVdVhrn9jPN4tVDk4rcenDoALDr1Puzc2hj3OW98apjeVBpMtaFqU
aN/ZTdLcBvQfnyBm3MaUs8If47R2xBPM8ZP7dU0HsgIx7dl9L5pGFs0Ji18LODfA
/bryuORSP/g/LS1/F2e9Kwvzz//UKdAEY7jEheRcm5NNQyaXJpWaG2im1sYKowML
y9/QSqTfsmldAv3P0Ax/njRgQQPwyiHZw5n5TdHZWNbsUUiWvwYaIoCjmXn5IfeB
2ffp6BVdEu7xkI4JopSOOju4Jz+kTrsJCmOtOLL4oyaEJX9TMZ6KmFiH7RoR3txO
gwDB2Z0kM04U+BXOm9hPtwJAeLPqU6fiM9V+k0jPtxG0XCHa0lmP8kZXkaIQJ6rb
WwpTIV0hhUVzuIlxY5wweyWeLe/mJWL+ehqU/qhb4XSrPPt9gSHu7ebC7FEpgigW
6iRKgkKjvg2CGpMCIn7XGbjRBSf55weZuxIZE3apStXAhQJzdItPtd89XnvTmedz
4wx+9R0auTVGLv+YPRr+tPS5dJe+udnwFKwXcMMkukFswuf6r/kPNP/B0Ed5lr3c
nlEF86dr75y45ZhCw3OOgGsDtvtnrZXkKOdpseQPq7HWl3c2XO23J9uBIVEO5dAS
wgvtjjmwkBio0Fwq/1ZZ4loOnBIBh57c5OHrZxnDCDz22TTa5cS1X6NYaupn2nRR
KStPA/ACP3X1QgfYlmVjMKX0dy8ci9vqEhI3Fn4EMwcwsPXi2z9M7xd7CiDr2t4W
cpN6DVJxpXZYc3Xp+kAsIXRt4qVjrfwD/mDL1Mi9DyE5SbFVImq4JIEv7EnYEwsO
d7pLvrxSwxgGxSDMtLuYltcMy5CuzEGzrty1hGk+FvWoc2ty9NCC6FVvI3jfvcOU
KLIlEIs6EUQS7Yj+vYYsxwb6/lENxZBpBOtBGy4zR5YV+EPGrzM0V6uT43LYPnxD
hHi7AuFUOw9MXaTLMRrkNkZgKVUIqt+wDH++u6TLOMgPgnYgGXDHTjQI2EBzIcLN
j/wY4LclYEPRb9CO7JuvGAEOT1SGTPwaFHFKAZ/av1UDQe7/5H8inqBDqQw6rp/Q
6/ysuyT3Q5id5SsdtHdhFcpgyk79vGA2WmzViJSroD1TmORWNjeu9NWExtaiF0au
vHZT8TOyIYLJnXtZ+bwBBNrmudJ3+KbEEeSjVsyyCbbVmDomWHWl3GD+Z8hlTV7w
2p+NBDov7sip+go0M92ClB/xNDmijsgKqI4sj3eNdNKxye1aa8EYmFF/bx0iag9l
yVpqARgEgpXwlTY4wCzR4k1wkfWNW150vfLaoQDcpvnTeDuxbsmPpLojQFQErOjJ
D5COX4eu66AyWVQrBcmfS5XigFtWMeZlVzwip37oMFQ7Xb2ufA/67FNVhMDlGdso
XI9vVFsFHlB9ndbvmWthA9f9RU87S8kMLymAKPUfKal2C7W/uPq7EI6E7m/gra9O
hGPCl1XB6wUG/NUbOFvWhibBF20ZLHO0aS+jJKbAlfRvCrXKYASZk3kK+p/yLpDr
sI30jTcZ6wV/6yytEXyU67Th2hzShdgODRRLkdSX/AwasD5mM11VX9004SxuQyi9
pGt0nYsdWZeG5zJToCMfGAPlX1IhZfFnPzMqD6xgMCNd2iHSLDLM+1djgnykMq2T
vOCi+yfTt5bI3Cu4po2ZP6PDWDRg/64nsTmWmswgmmOiWAb+fu0XRbDyamRp43u+
QShAsYRm5mU7jvA5BXUCTYAlBxgGUCatHtXY6S9+cgbPewhM14kXJmxOd8bntm9i
gRqo9VKUS1RKKLaY6MyNdu1fOwdx/CCQXQJsK08gy0YMhhfWZ9nAUq8ovX6v2H9x
zldxaGb64AJPQEuybtH9ww8xWg8wA82DIHEA/rv2HD6po/XQxlp+2FeahirY/JKI
qcbijm4Hh8g3NH4HmLD2sQa7QlntZ2J7gGIIfLZjMngwpPiDxLPx5yzKhBS6hiaG
O+5BWQ7yOptiiTnUzheAbSmNMjO0T745WqVFnxhNz81rnbf0oXZ6jMkMIfDrGTiK
sepan2BrVpCqogBUNTRYR2qwevT89CxdevYcgZrmFcuZMsWAq6365I3uNBHQG9nz
5GTtEGEHLbcHIZTFxCcKmfyggyANEPz8w//9X4a1cCs/ts2mAKX1puHtzLlCOAMM
Uu1OVosKkV+wESoI68bqw2746MYz3vRK5bDJy72bd/5OrKveYnm4zo9Bck0+KF0r
I2Z+Dn8iUwT87oMFCCOOZw0NhNCpkSj4jjN7FUtXPuR+T2h4XwIJvFsnZuhq02H6
vN+QyIVB/EncmUwczDip1T7Tu1iptXFr1Aew5i0u6Dzs0BbFSOaFbZeCAiIld3My
FLGSvO9gzY8VvSkDXxi9Uah4jatI1Gn30TS1sacJ/Q02dA5eWJE1nImjmESqxUAz
/RTLq9bEUHyZZeYoSwH1D/vS0z4n5CAmQwFCFL1Jy3G6rAtooM4UOBhY3qikoNl9
teuvzrGO+0YxDJXYd/iJwWiJXsNOPE7W/tqxtiQ/57zTGR9JnlFWYpdZMC4Q0koK
OrFbROEYoi3w8vN0w0+6EhXgCAXyrGxgVO3IklvCEBrYBUR0VrgITvlJfwmXeagM
vQvSpgUs0L8Vr6lAuyYRdqeyKpE7SxQAGRU/G2nYAevO9nM4qNMd8vGdUt6gOnb5
ex9eeBSEUdllhdBk+Um8YdLVfv06zEyLHVaJKS4xz6fsKLJ9O5XIq3n5siTZZvCW
GwogxIAAEfblmkUjqBvjTcT3eebbqyERDA+H7tO09L2GcNHQPw/su5+h7PIXf2L+
gYIGCzNn9xZmvcyyWn0sHvweAk0N4jy5YUwSa+of/npVNcbM0/DnP3t7ahkyXrvj
ZmfiyHWa3+dKO/amop6LkMGXaLQYpzSst1inEBWeFFLRa084yDiXSDkiqyzN5Rnf
dd2B9Ve4HyBuVTkAZ/I0qp6RT8B4btzFtrqR7gIyceN/m/+y6OUCBGg/aOxxSIGY
HUx2ABpQqhQ8QOvQwSJw2YDPP9oLj9AxiM9kL0LjqMdyVj3+Q74ke5RnmtXe+kkA
LuKL51BNBuIMow86gbULtlWO/P34ProyuH5fpPCp4gpc33XDlqXzkmBljKHNs2zD
A4lV9CvGjogO0NO2NduHiHgeDKfcZ5JKfTEZPsBrizz82BKwtx0VYzC+0KYHj7D7
hWaLEAQ3Q806o+jSuXSZXzlhAfiT0FFUNBJbeXIMNMaAa+A0qy2hEukCfUM3jJy4
xKUeP+Kuq3A3/ydYjnb3Ws0IIbwDGy7iiHIIDJsLp92DvT0M10nWLT1UiS7ALdsK
dwW5xc6elUFJQRFekzzej6II0Ohyw5EGus+eZGEaaVTpuI3deiBZn+gpkSt7CASD
XrNkbZYgL1KV4CIZ2v7lX3hAKnGHjIlv9Xvpsr/VVe+w+lUJKLwPwOg5I5Cv592h
6fgPtZd2/OOBEUiC1mp85+bfdI74Wq/YowmtzYn4iIp8DlVMno16LMq/49W4E5iA
xc9aqR/cJzvFipKw0CArDk4cXEnQsokFBDa1z2PhfDka+valdBs6kNKuAV4R5ACH
1RHD/O8H+QMmNtT+t7i/3ze04yQqD1/IPkNXOvz4AuiZJu6AyD9BCUEJVuWjRk4m
UbeGoOaprNuawkLxDY2fz1Jh6dZvn8MALOUMwDoaVTMW0lJQQipAX+cdU4tht4hZ
N/GXXAhX/o43YB6UIbcuAdO/tjPWeO/QIZRyRvjv93j0wqvcqOi5JdZqFddn/jgw
GOWAVmmbH8ZIAjxu9l611zgtm6pgSelCqUhrhMY/QOa8BsflGQ49hUwRflQG2PKC
s94ATKIOh4VJc8k7C/FHoUGMXoQ+0jwLN3Xh9lfR+62wF1M4YwJvF0Fv8eu+KDjY
p9ZX4ChfhkgqnZNGgDBGZ6VOZ6LsfFKbLI94Gn8BhrLcPS9e+ANiNvd91Nnaevm9
FzMOiPYkSc7xnyTeODtqIZZzXb9wYyj6HX+UGOo5KXZ14x93fOVuGiOY4aDWRM4X
iDBf0o6jGdFht6jMaYG2tYR2zvAqPQwEG9W8nWMpTMeIRpB8QiLWJkdWm5E2FfP4
6m1IxtrMYVm5T6tRUGYw269NampR1uhwHFsbtiggOnohGhWF9WfzCrRPvIXNiYSi
ax72LRYKYs+stWScEAO0YXLXXAyrvj0YFlwu5LF5m+OA9wV9X/vi0RLVxDGacT2Z
0O32Hib9KdNQOfiHsz3UozVUn6sWHnyX63G/8IjQIaIkh4bG5hMBd/4IRokLDRaM
3V7r/pmWFXGULH8v762YX4eBwlTgGpla0OuOpMhj/H4NNsyWkIil8ZQMhjv447ab
bTu/Pdp3QUURrNlzSR/Fut937QMIlJ2VsSgUWXiRu2ipdsc0IeEr9vCsuu+uSFiI
UBPi6TO0FY88UgMczBtXfB+6GLYzRDfsz9WkajfSmTqb/Gw48NBOKCmTeAmG2mvV
rjIBIibQJLfWrBAl48uV99/oSpf67OkXrU40aKDQQkRxhnfFLLHcbxysuztMpqR5
eEwyu7+OOTw+IyLj0guC4KAknESsey6EP5gzYnIEmVjlWRSsaDJXDRoZ7ieXPFJh
sDLEHa3Tu+jYK/D3BJbsiEYDRfxTJcQjikWY6ST+8B9mJzQTfpcmjrTcB6D4n5/f
HyDH5MKrTveFxk9TmqZmKWfLZns2HyKIwBJYiT96KYOlI29T4oX86d61T+v+aMNl
vF1CPpA6z6SjBvQPZ3oCmAczDlI8fOlst5DoTI7yW0J4VSYzwREF6Ga5BoZyB/oV
qx8alqHdYbqJpoekoeVbowgbRN6qA4uPdwrMygESTgpFMb9Zl+AVrSOv9ZnbhUzE
jVaUgSWYEoOSKP3VYl8fcerx11YYjrOiBLR9TYWo9wxEiKh1lu6pvWvw/fCdqRXh
8VNpoKAZCuSSAK3iRnWrblzfbuEx2p+IvPMMm/QzroiDhYGheXJlOM0jBPML/MPy
2DxFTML6C3hpNpS6kjkbdkkD2tRpaVHSpGkaSitmXAhk3zWY483C0GlzItZbsUQ6
4gvR04BrLImfqZK9WUf2XEmYxk4XDeehqCaZ9Pt15OdFv0BcTQRRSycByleCyWWw
g41j85tdU2FrGPbgssfboYGXvbMCecrQdE3gWqpzPDcd32NHsQcYwK0IejWNtaxL
B4cG156wwYMLzipJ3ct80z/axqoia04o5d6pssfL+euy+jBIZ0hjKqw8SS7+eGh8
nNJgvOp4ewYvQy2CIGqfV6OYr3X94Iyz7iXvT30/gbnajBGiB9ytq4yqa0RwBJ/4
UkU1wcILNUgzuaP4Zx81Ka/vOk0FOuQbov1pVgXiIui0eprKUJQH+GMnGD+Tjs/w
WzgnybQZoo9dq6IoHS3SAnsNGX/olwMxMADBx1opTdyUTFg0970MOOVALoB4vujZ
UBWXvTobjdcttaBu8rpMmbYAorVXAjzZ2HgQf8fHrf4pM1+s3e1zvtHMAHrjAUqD
/xqfByIpQHkXz6jujmM+EOhFgvyjnMmCgXipey72QdODsKdB+eBMMmN/mAIejERo
bd/3dylz8xgGi34hhVNSZlLusg+5I998vMXIH8ODRNzMrQgMcm0g2QpInii+zOTM
NAxxWlQgy5Q5+3+o+42fwsocMeB2DnE035MenoHIOiFONUIYmdzP2CxTEPokpBiJ
IGVjfJaQfkfm3CIQcp+MVjW+AncDywt/vYttaJbyta6sBP9M2n/geW0sojKvHena
/VvDyIOs+mrlWZ0yx/1ji3+xRmYL8KaH2O+x5Iw92NODG55nHheJKiUjtyg6RgXB
ec/VmrpqEJ6dXFvIo+IwN77mYm0Q7Z738DUw+mMP0YA+DmGy0idi0NDlHEES6TFz
YYDAKb3gbaF4026XIAhyKCMEFigxgKQ5Jw6cgJh8bj+5B4s7x8Si1Y6sisuD8rD6
dKhraKXGWOjnA/ZzD4miidzioBczGg7jomTyIAAqo5XLZrwOg2qPlf6NVnEXkCw9
S+oi4fLT/coRJzq5taUloQAACNHCmeyxKxwa0Aku/JlbrP1WtD26TzSiCY0/Keb5
6AR//BYI3M3T0T3Ngat3Nyctws/hHczjhuVp/+JQHg7hbT8M1wXt4THB20bLHkkx
WmW8M2I1zQ3U3HvDnD9mFC5yr+W6Ntp925/mETWXnx7ceptAL+zmgJt3Lh7P3ccT
mZw/75RP/cR1pOGQseWgbEF21kqEi4YRZPMTjLFwZuiyDSyqeRb73BZ3fwxCK9Ij
oPW9R2tOKfA+7p/2H5Hb4xPWu5EkpMMZ8oNlBYyLEHdhs96AG9up1bqp9GYghwew
01FCjFFpUr75wSF/phxOY+p3A9X73NVlCx15xaAhKVmt10SB4TnFbz4a6RTr652W
jmRnG9Vo13IZb2inlemmo1/i+Rlay8RMuXLd6qPMWcQ4MyXmjgts0fJ6g4DRT56a
LWDaTxZi6+1GpQrj/Fdes99LAm1tYUeDJ1rRGuFohVT3h6liA91JcUWnhkl7Vy8g
RCev09GukRKFKnQhkeBb0X7qloFiQwDF7qiS7TBtRla9a0QqWg1o2oiiDwt1ECc1
c2mJWGZZGWg/SvW5OAxKpn83sF4ks5ADTtyCsmpNalBaxzxBoKl/czDYjHFz2wth
8fM49QfD/N9wHjFuEA638yRs/h2dqssnA/wnp+Yz1kdtb8IA+GJkUweYziFI876g
qU0NOFQMt0EyciquuBeeBjlCEWs4dRZBwkfGQz8A8AI89m9GW8iSpnvMwOAVVg6P
hnwgMWa6jmley3wvpDTKvJQ3KOKga5YUFumS5FR6DY+OsJfdMquohZ6cjmbo6oe/
UsLrSgTn36vy5mWxlHVi3xdQIIEBzRO8sP2EgOF8rFlgwTS0sK2jb/OpBrn4a0Mr
0V+e000PUiKGHy4lbaS7cXsickkcZ9fNE+ik4my/iG5pju4vtoGcmCyKubOWzV0p
Y18OdK6yCRy21d8cDQvPnL0iBs1xgQYsUUopzhcWC5mUffCRUTE0do9Q6itV2lkj
Uf+M3tPzCuYu1jHXTBgr99+RDA14QC3fBlvUK8T6iPqerMagKjHsOVLcdM/spzdp
a7g5oVTZgi/5dPFyxYUWsIFL9c27Ewc4D+ahYmCVFKle1w0x7fGTINbFTThw/t9m
v1H+qY1RIXTAT/Am4Z+YmZ7o5GQ5BNPjGaeDaV+cqyf43MRtz8rpIlyIUSkGqQur
5QQnjWof15OG5+J3y/ZldkYIQORfIJEtfmA0VLlb+jun+aEyDb6RWXtodylIzYVy
/xlx6lG6TVRA0CaeGQDsimQsMIwHSBf3Poi2J5Ujgw4AnqXWWTLlsg77xYy5eXil
f6WXGftm7TYQeWlozpI85nF4/xTgIt2+QRD75GMOd7Ljfa+fk8cQr0N7K1Jxz2P7
FEhZEwOt5anKnYAOe4TT751woSs2yamDUBCTcJ9KSt3NZfLa7FrrJNZuk0lHanoh
iPpBI/TF0Zmc3QiHBGxwDZ597sTEZYAxlPZzaaNhM18ZdvZPKlTX+38BxfElw9oO
cV8uZFTgQ7bH8B+laXS0ltyEGL8wERpdXzLd8jt/BpXWEY6rntBDrN5kTQRTID9t
2UY9DXp5SD5mWJU+487hGjE/bEYM2oOQgj1R9Toa0u564njCE2XiynL5KXnlYjku
NAw+4AZZg1LDAGuEdTxd9/NM5Mae6/PGSHgO/mXDCO/kYinzfKJiwy6RIyJn7v3o
uWhxDSgXaudBSX0Unons0tVR95UZ4N1IpLWxafkyEJJEcZJNswrxEyPRGmY9vvuJ
1ap/bZUNgb/ZlML8VRJUliFVGeOHSTbJQX2+JQbuVgRDZbDAJAMHCnRFKW2WOQoS
/qiKzXs4FFCFlOqArk4q9OSisvP1mLRtTJGZchhMPUGi/tHoQxrA/6zw+mxMkT3j
zMS2LWQNDvSvMweSZLYHUfyLM+XJwLWznTN77jeC2HTsrfmma3GQqtcSM831rUZs
cknqkIp7iLJmecaVQqOu9F/NujWPW4MmxlQ9pWZjTKDeZ3b2T0e8qjIoYIvVapxT
7FeJJbkXn5ByAHNVn6ldp/7JNZ4NzPgbNp2n2ENImoFBOAILs40axT4nk4hor5K5
nyNnCT6Ee/bYUfLn6PBgX39WRL5VRslqMJ1X4Htt3myE0QTtlab91jhajPcDIUb7
tFg9QiLK5LtmkdlFtcNE2f/dpfP+Od2TAm11p9LkyR5LSaJMgIZIfuxgnDNq6A9y
0G7m/YTq5yfLcSZ3y+JDrQCKbiSx7F73JIrGVZh3fCA/Y1/+AfbaKqjKKlWwK3Sb
rXbEM/UC9iyP+3zEM9IVSRnf+ppFYDfJzCWwHGjgyogORJ/fibrTkek+dSaRS1Ej
wy491bvWGcs8n/sJRY4HiqDSOwfglZUcP+aUYyFR9QKQrhQiVBGsW4uaHcbnFruj
6kwfdhfFU/R89bTgic0oYDIlEAF3KkAlKjxU+ETdgJZc3LGYvGAAwiodcczJxA0T
q/OQppOCfpfBr3fV9YeqjDnTjXtSQn6y0aIf07gvYWJVdef6BXJLwq74OOlItwyZ
OLzh9rSoaeWazeKS5Svk7MJaY8uMgNhp0BlHt/kD30WPeR1ViF+oV5+hmr96jARn
3oB7N0MGcXZ18tk/5qI6Qms2hFsCL2xjjtNoJA2clfeVcjJZQSTnZm3gO3ihfAkd
t058C+fu9j8IN1aUlocI1mqWBdItqgW2yUrmxmlNKgPW0jczhy3N5RGnzuO9KYRT
o886pOsXW1e1mZNzSu945jE/5DNVa7ALS2ARRHAL6tPGcTMCbhlpRjv8nG7up8rn
9jtzx0d7bjqzKJno0eJFKp2YLDPUSbAwyoxPPJWaNDpjfCmK2kS4DsTkU+CRE6On
c8QWVUntB/kQY5Ohpf/qSlBmh2E/UNnpbw4rli2c9eBC9jfM5OZgM1a9MtWWhmyH
3xTFOG0kar/DhnPK92HRRk2RtrfvsFltmf2XfQsxH8+Tz05ysF9rKz3Gm8eKzF/5
l8o000ptgaEVV9deFa63d3Dmh3Hgw/IpzpcgjItp29eq0F6lU3R+9g8WOKpV9NTd
Er5fYdazDGBNCc0ndBEDNXFFy+i9i9yEaEMTOhVhksReh5nwXz1gw4gLfj/qbzlv
49LBKeAFoAM0uIrtkTq3yqah4dlktbB/dER1RIHpQnf9Ari8fGrkD3YorPZgPVn0
WYZxByokXRh2n8LlE8A5xCz8W4022pCEaoVeZsE3+Ma88bCZQzEghKWiqJNVV9yA
IzzcI4vNiPtuVdeQoKEvkfYquubm0JT2gUonHEX7U2t2xKXZbC7z4/inSbHu0vMC
NytKwBNEGbg39idtts5ff2I3AXQ7IjzxlPHzI7r87DAEMWyVVaTs4EtLoio4SXos
3yHENTrMuFdxOlR/8aEaB2eblddtgKRJlxHv6lg8XhV1GSqh0Cy592Jy1eGAJuxo
g/NQuhec+KocLQ1Mtuevk54qH7bU+xVvF7159PkGgjfQH87/UZblsB1huBk/xx7K
AGcXrEoN32efxsN8bBB+U6Z10lG/NplfToedG9r2Vi7dwkRyKM8fhmYkKhYx5mAt
HuhzfAJ0F7bwoN+CcRXIrtjc9oePtaWXKcEwyln8cqBQchz1CicOQtkJE8AWFQMQ
jQMMF+Dl4PPCCp5ij4aTtZMgL7yOdKTGTtNNDAUwf4VxCU40YXprNX4i3vkmisQa
UiTqa7/bHlyQhYViW/idcWdD2JtUTY+qq6H9Z0/sEfdvpIGuwQX0Hc+Q+slbts9u
MDvMOXkFnXPFp/QZwgua207q2W/Vu6suRpEYSZ2KAABI1AiUmYwSTz650BxEfEkY
3qCSOJF20o4xR/vwGTNZweG/hK7xC9qcKkce3VbZ2WlgT2NPAFMBEWw0Es/drFAH
ivIYxfjmZUKvR7XjDHF+y4c+1G05JrLog1Q8CXktKEhdeKpNjwL6r3E0YFOR9Hvd
AkGWplbjpq7Z/1hLziAD4upsaJh5vRVV3e3AYf8zOyKCwjqE8QQ6qi/VPWATwGEz
O+xHRmej0ckkrphD7qxgc0mu+dpWlfgsUI3TEPCS85txChD5E+ubQv9itbupNM/f
9h56v/qCm+QjO/mloTtn/12CPW2QSv/bywjKikFFBedhkZDgme5TSSRFqvDJIAo3
oO4zF+xjh29AWwpVZ1qF6FyTG3mk+yuzAwQnH/bwSMIZeybCgM+NgfFxymlDIJ+6
JpTvAM+JdzIyaRJdm48ng/MeTsARlrJBSEqIDbEtgxLFXLp2AAcOizpWaVE9rJPz
OUNo9LsMftHtE1TzhO2fa5xhhSHnkIFOkB+s9JckfBT16eP5tSD0cRQcmc6UqoYm
YBMxq9idHEMvVLr5hX7hmAg8XC2nNx3Gk1AM6ZkY/ll0K3Y1SJuDkkkca+wq90cu
sjhwpk5vX9OZywaGET1IhXCwic+EhAo+J6DxCDnOzPgUecuEsfqGSH7pnVjkh92N
ASPk+zN/4xFIJu1A0lwta/+KVBZxgDb1THl9Yfk5EhL+GOS1JvhhtE5fMOTOaXWD
jfozvoJYHVB4QtOKnV8siG4V+8XMWbhflFt5kIpULRVj5Gbu6tx1c6ew5BbhV1O8
ZSA3sHCBOVk4L2mhQL+SPhp02IfPYtx1772zRTfROfDikENDh4gTV3njPFh5qDLp
jTorhlw32HdzLI1YaTQvyo4TVkZCHAYK4ysqqbNPm1FXvOjUF3sReAYQnsCQn0Wj
+pHe4tZnIeDaOHyDSFRg3KmPKzW/xn1P1lYNFRm3iOGnDxqP+DQFrZeiN/xVFehF
rumEFh69a90uIvsgEQ/69dbp1YYghRF0wuXwWshwsh1qevux3Hd2ZgfXSAcZwwL1
8HlIVXQE5HQoZt53mvyXSujQjQGCLqNKkciJs2Gsr/ay1lSozr44vlqsGE4QgcqW
MeFZ1xGQlAFOs7U+VQaHoaeRbYsY871/HpU4hSSghzmLYj7E3XMkXu5nSDDE4qvT
9ljpkkaxngSJZRch9dd2yObBleuUudJ9Sg/5WTHHkID9hqvU1CNi3uUTJi8oH53M
rsunjg8Z434e6VYZMTFw9XN/7znrm2gE8LLBPG1JCE7vaLWXfSHqQsjDWIlwgc/x
mWrLkWwiNEnZH/g/d44MqPB08suAsJlLzz9AqasQj689kmZZuXHnoUVmRjoQOYZK
9RkuN5XC9uB6MbLxKXQVgW3hufhrv52l1cVJdZWDXkoB9XRHGKcYhR6GYAIXmK2R
ytwatZxbqdTY907e2FXQYPAjqPG5kEcw8CWz00DCYozOpi3KFjrbHv7BmKHeBM4W
ovDBzH0zcUZz9DjgoD4+dwpJiI3YPp4EVP0T0bwBRfhTBwrI9oPma1ZUFTrigXFM
5gQB0fXTmGkAwXpuUC85sFR9WpGzyMUI/+uCQGzBXL72W/q3BcIM6BhtgzUQ4aS5
tjpvcyzMlt12JO2JKoQoBDcoGYNvp5+69VCFfS5P6SqEcEM3VysN1JeqPF77DOXp
Tt7GGT8sj4tFruvlDN44wVe5oCET5NTHYMN+NoGWGXymD3kW0kt6U3+eghZxRnq1
U5/+ci9N3PujXeqlswTrKFtsLVoTSK/SvFNHN9QFyDIh22cKBofS3F2w0taOZtWV
/s64Gb8gYwicslQSZD4o+uvDn2dSX+XQ4tLd0rpVsrOCaNvKHgdSTNtX6/QjUtyj
kxNl1BUxHDX5wx0cTufmi08ZOE/4ZwA3A6lXwdVfBuuBSUjCn/LGDjVV0DmnPIaK
zRlSiT24ZqE0KZ2rRxMa6bPsE+nO6bAUgHN5iCTjAmaRbB+3wb2RUywiavf966Zm
Ug1eqPvk50Qbn/MfQxs2DB/WykOPYcFpLF0ZRIb/xGpkEwGkmIEIuAMBVs1oTKcE
dKk07JP4J1W3A+hC6LyVFoFYeoqRL90Ne9Y2Ez8LVxwh6DSVcSbQ/y5eBXuk1mdd
6WOlXy2tDInmblJrzIQgr9dHaMD4vEKrzZBMhCJZ3reYlZP0CF30eVJzG3vkubug
Wq7Gy65lYIBH9Vnf+N9O8F7/g5U4OwrNN6FOcN55bXnfkBkit0QnkfmIYX4L7W7B
jbwrExqVRokWq8MYh5zNgzLYlwCQXDV2VlfYOUNLyBQKMdov0eBaRoL2MlxTkSpQ
TyytCvddcIvg7aKCb2UhecL5N+RHhsmKgI+JOFMFb0AM3M6op1EQQ3R276ogtZwr
ZuufqJ79OnhlnHzvQRjZx8gLb+QRriMhy91WBmp0HNt2yb8/obJrXOGMUOx4HtuK
nctc99hchXSH5f9KXK74vwL6Z3J283+gJFVJxLnyv22Bmob9X0ohONHZXAQNHtMp
Pt20RriAwVu9d1YnNXs8TpPsnR4txxuKS0iSj7M4qYVQiWlOTFLSP3AnmithdyGQ
zu1TN4ZoYqIBaM03K3d1YuyBPN3D/xsUP+wk9qIC7WnbsukUc3mBhKCf7KtDyzdf
B7q2Q64DiFYA2W7AjAMhAcLaUlRPa1PsOI7wWqkEJli/LBnUdyAq9PMOvICzLkqH
Cv4qzKXvaXNTbPK2v1m5Fi4L1qcoA/u4b0d6juE5O+pGuW/WHoGsmf7MM+vFpsmn
1rcxNujPoEj+Sl5OH0tPWX0Si0O394JN4Y5yGn7J86WCszhDR68P2nF6Aldksvqy
9t+32ANje/xH22J12ZMH96iLO9Q5dUCh1rioqc1lAaq19gDrEZ3l8TS2VQtUD6OZ
CZzctq9GPB+GICDKidXpLrQ7y8WxfT+t5fDI0C/HFBr6mklXA5nmJysMer06Qao/
D+KsPV1TrQKTClbJn7rdvibF13GyhILs/iC10zwve04rvvi1cyLc4G7OAvHMNbvT
uBvXAIxeVaBjr4fyVLDy8DSWlizdexcVZ3v7sseSdSBbD0cKDTjckZNwbjnESTTA
EsGkYrAY0dA/YCwGc53s1LemQtR2oKnmrQHkpEY8LaB/RIeDsBHlsWDPPexUq2KG
msO6jgU+ckwRyv+Qk1pChU1IUB0hPath26BrSu/QMqdJ3/nH272IG+5Lu/nwLVx/
ymtiHYYAlmqvuUsXvPek8bhsXa1OcTjVKGY9SCF8Phg/nCBAlkzNUAek9EnXX7XR
0ERqV1ltJgn+K+II90hlmBxb+8xiuvtLsHLHu8dnzIBXW049eQgYTRJRI0/irz/g
eVuqSsIlGqitSN47rbe8eFKInjhKFuar4pZ4bvOWzzcD6D/tt3dDhOMPDjsLSVI2
0yAZ8h7ZW0U7b2RTMeJpYvqYDwKuNDLYp8dEusApyz0MBZa92+vZfulO12yrs/k8
Bltlw5pdxIEhzDmjTCzaNOW77r3SjLW9HY+FAaPbbfC9zC819mSrwBBTeL/mCcb3
3clRPKDRa+ooZXwz+QK4yB3rewnqSPl/LN0kjGTSli6Y0FTMvXAaP6EuqwwrB6C7
iSAalnq56o7vt55EW8M62C/dYFuimrRjtN8diljJNWuIPTDw2gD7RDITg7gxJa5E
rWU3uBo6IVjAhiXtPBwZ3vr5RWn6tE+pzeZrsUG32R2d5BBb4/XH/b8nzI9Jqu3Q
ZyglhEcid0q6vC12OBwFRKxKvqk0Z6UPckUcZVdKVOj7fuAkYGhQIAHuFGc5MTBp
HaGsD1rkR3ZkIP4/zG7ocb1wLIfzC+Hn4ogbSxdbXG3skSR1tOBUiqhG5icHUDN6
AEW3IgY3VfmYaAEGdBcNKhhSu3nT5wQAYNzAIfDwCl0P0QcnlCKv8utI9/OpIMJ3
sF3p/NAT831FGFEf8c8Uyb8rYeeeILtY8wITJOVp/qRubIwEvsQjjOAE2rNL9aDw
YySeDvMb3YNitfTODMB59YNgXfokDVVick8fy6TN0cc4xnDWvN5znFXOj5in+czT
P2kKkLtVV4vGo5Mf9wWLGvRibAKO+9PCXvihWgpWvBh172DLZGSkR9Vm4qF5Ocq9
fQzn26RS+pE9H+83GllSyXjk6vC82p1C5izx/KWLK0dM34tniNcbKPIfZILk+Uz/
Z+hEtU0sm9MxoYAT4m77p6Bj9BSxn8n/w7UQimGrBRoag3lmZI2NLKzbe1HfWnh2
VXy2iRAddZuG0q7jw77uf+P5WqxvaZqnP7N2hAPJJgUrAeZHxMOsa2gpY3fXsSRP
AtONbvvNSkiHw9snHUO8yDpsD509Vnb51PT2PTV0pFl2q9dgPSjL7umyAJHZ6Gy/
9OrW49ucs8LNskS52L+i4peJUHVDbSqLYHcfMR8RiGXNHsYiYatnJY7nj1Qj8pLZ
PNqMHfNtA7dfKrY3BJ0VdG3G9gLzDz1YSK76M8pyYqR6/BRG+ETHtAoVPvNVDVHm
+Bt9MreMgZ/41b9kD96k5zGLbl1S1ACHz08E3B+2jEoX3vWHrKNBATORVhS2wW2p
Wf6eayZFssYYEFs/Epoxybp98QdKA01Zq3vq3lQWslMBLnYv6qyqxu1trTIcmKOU
MueX33byfrF72i2jd/UYyG5REFUSgshvH2fi2iwtvZb2P7E4o+EI3J5ZDVdssj7b
zpA8m9oRiFM9HrETbR9mAL0buuhddzs6TGdBj4m31YwNhHufh0qyfv2/h7YHsKQH
EqJTOvOtX4HYwm2qQ0EUjPSQGvhkMRCkxqjIhpT0uoZWrQkFaw3+4G41EstTc32E
67/4heDV8cOqPejv9H+uXAHP/ghTDe+tePpgGc1CWk6cD/nt7KEDoQCEermWNMUr
/VXvfbJnR2GIhWGTUnQLoK8mF639P6DeXG4Oa+2D8u9Lvw9qgGsz1cHHcQvkRsn+
0BHsB+xoZ368hAzd0FKHpEyeOhdkIJzw3CrD59ZWqo9Fm/f+Bgc+FezumEkGVFjy
4H0qb3rmodIL8hR59PwD6aYit14n+03yy1l6UjRJelTvLpTPNKgAURSEthL3Kix0
exRAy0T7s6OzK9CUrEstJ0BqG+LS+yJ92rIYs+4xXMLgSRr9xyAhZzWZBkKzKCP5
bQS9tEXA4FYrmCq7g6hiECqzvOo75hNRUkfI9m14JxrUed7Gl/C0aT/s9Dt9sd7n
4hf/7E97AkW1sQ1vAZLsHg8wF2S+OOhA7Zmx0YqcfqdxkhxowKBARJU4oY/pHz3Q
l+t0oo6ABDIvS+XuyXME++rbcwc8SOZOO07UnHC8xzzNF7D8AblH7qjKmZvBbZWu
3T/Ct7akyQSfCSUipKOGSy2mEAGWw+Osa/d4cmXt7HNfYZgXCq37CK2JPwvX4J31
6quDiohQ0isUTiwndzpWUNTnvdc83OzGHQ4MsydH3zeRgoKdlYLzXXPESfS70uHX
Z2M55AdQ+tOMBHTso2C7TWTUGUsqfRT9fi/emHNwEOZmXJN11b4aVZowRJO9CeYj
2xZ2AWLZPzm/9Ty5gMVEg9xOT3pJzP4YMcjWtIzS7C9aS0OujQ4hDqojWACFrU/c
HoVTnnxhGdy0rHhcSvrUqogArcDLtYyuVlniGhz1CndzJlNrwigtRCZ4mEi9p2Dz
hZYSiGffMWaYEjTWTC2USnlJWyfDDKsH0nyEUpBwdcAZ8gS6W4KTuZqv65sm6lJ2
o1/2Lk34DnfADq2BTS8H9Wka0cLmrTkawn5v3uzA/IrEIOhDQ0uWpc8POm5RFm5z
jZIVImLLG+dpdKh90i09dcgGyt0IIPwwEn+k40eUW3+u987P6hGIDOpX6mRf7T48
U3pOJ2P72ptDiHNpDtZHJqSlS0MBoLllTVTqkKBMVSK6/f9ItjOOCcGMO5WsdRs6
8VquiT6vG4z9/KxaafwZKjBkvRcSz1i4uwznFHdNlzXGVhy0SnJlRQKy9dSvcPtc
lmOdALyTBeCMxlrwJiH4PfKotLY+5Z8mdyRegxIy000F09Uu5dkt7VZolzLU9AN1
et6esRd1Df4SgsxbkQgUKDV6GxxuO7v7GW4MKbOk/VdkoFmHed5iWa7SFM3sgMVq
BIO3Cpv0b/y5Pa2UFp7Y//a1ADj/HGKUuib+6+/E4KqtnbVsJN6FXaxVq7NCxh2G
lcuVV+I1E6YRxAqA6Uis9OKR1lFumjJvAsyrZ0Zl/I+MRPOUlik7ugaDth07XPBp
ktmGnW4ElhtPMBzXe220PADCXnAK69vjUOQfmqAdzKyILSOEJvyFYtcWtqbumbTo
NnNeu0Xl2G4wcqjhENkeXUsmXlMCz61eRpamrcmTWIk7mvocO3sKzsP2jGTo09ii
108vdH7S4o6j2x3Vfw/lrpr315N0XuOWmkE5jwshERSGEKy0R+LVIsOn1zrpQAaj
8zqboma7FBSGcZHmOdsUkfM44BHsNFNOAzdidm8N3rFQoTXrcuXnIOjH+QsZKtuq
nt6g+OYjvRx92QBcq/9aIbez7gPztzK1/27KcHy26C91K70b82hB1T2kqwIuJiUy
ZydFXSqM3AJXhdo5CS+c0AU8snMlaxdY/C7LkkHuwVmQ2jMPFSaGb5zDNkSoIYat
fAolvvkT8sDaK06/MY+Ylrkj12X5B+HzU+5niO4rpUd/ytuXp1zfLBvD9tj6SGux
hxRu6mg0OyW7WCWyIPljKwuaOWJsG2UVufBmT7tDw8E/nIlmcRTwzolKQ4UbMBtM
sO++3ZHZYEY2w1aMJxgHN8VoixtSRmofbR7oc38kh7HS+9xM6UnOAHK3WyVfhWCD
84MSV+Acia6+Ql3eW3hUNw16c6Ye6PcU7c63Yj1KcGQ1Dv57Y8lkijo+au1sXup/
KTb1Xbrg0i+6d9kVWtB6uKmH2wb8jGF7mK+SDKqo2xnqueExNC/pRlemgF8yYI29
7uuWjQ1sESJhTz745+bmbpRh9KBdXhLs/Vv1Qol0Gw8X7L3zKzk6KrQ6Prq1cLBX
6AA46bI3RuSs7JUaJgAvmqRUBDxu3VUk0rfFg5YU1WRkkxqnuGQlAMX0vNg2Zlrb
DiBFpmVo+8NZQY9p4JgJhl+Nuai1BIlJfk68Dwnk17LEEeqhLtoWI6GNldifM0mJ
BOfnePu5bc/6VR8N2Vvgj3M/8kUgsFnHc1prUlRYkcbZzoi11/CRZ/wYlZTgKp83
UO2FNuWqQZFrv4vQlTjlLlzyfzsUGTA7UOipQJZC1PSZdJHyEN/1ozx0Ancjb95I
hjGmUjNJybwApF8lM+bm98PWZgNUspVXJqInfjqHVHdXI/aDNbFssyn2ar5ZPO0H
mmUWHVfBqBW5TNtjPdhCGusfnsOaySJL2AVrSvyngVtW0yYVGBebZ7zB/nauxfqi
7KETLtykwb+nyKwXUfhxh23Vr8bIcM9BSnjxqwlYYwPjWhouKURYkfdStVrjrx9T
U2qsgg4lbBa1/YJP7UUNjRqwsuxHrBr5y85HXW73h/GnvbJVxPDUjUEuWlWbXpOn
18DUmV3APIe0BePqoGD92y3eOHTuA/fJULEFsW2WhKwS0YB+pM5aNZVae04mAaEr
8t7DiE+co9OhnDyswOqMcmUGX+RZSrf/sjUi/BHxnMs6noOLHHO37sueyrl3Te9z
400E3YME6eoVYThBVTe76dZn3BhVySwRmLE43ndf+VPIXpcqCIIvf3zxSqwMsupo
GdtcgMh4XqpkRO8o00nccli+196jbut10BXuuMWfHdChG0zzJVVqmJPhod3wvkpJ
X8P55z6ABErXEapTyJyfexpfLL3kaMDluYRakMerpWNz12Ni5G9ALC+kb5TJVLf3
zXokmMLtISmBxAXUYzDjZ3iTwgOsD64+HUMmnkedAO+nDX8XdysF7Plk/RF+U62c
aRAt8FG/3yE0Pr9smKduF+M3yXJ0kzxo8UETB3tg5llPlVWXIqP7y8xcaROJJBzE
T8V2geW46T8UMtH3BVT9mOpyOk/HzJVY9lPrW3trtEdiPGHi1y71xN0QhOwSifvX
PBfM1dWujVALZzxUaoaLAsr5xTJrv2Srga3Sbt7bOpHNzdVO1eittmEB+J1bFnPH
X6Dtbn4HWousBuI4N4Yoj271Dzf6WtCVHUbeo4sjh4K0ZPyEOUyaZdj0s0Vw/Q15
z2Fma5O8LiWQKcF8Wo7rw5qnkFXHw18PZ1o5e5NOF7rd0ZX3Pto5OZTfiZiu29+f
EQIY7wmIvC5dOYMAix5gJjCJa5MthYeU4EzhfGamwt5szEN4WEEJeiW/JbmT3M8J
5hsMhviNb+KDLdkbiMlzxbsM5pRT11PP4qVUBd8F73j/fZgZoYWZYFAgijApmewp
pkTjoPClhueZg+Ioxe8V3mMEccS1rzXpcqVw5ET++wRqF2jDaIeogsBgvS3urw4l
qcGyIDqXdhrnwWSAb+ZRFml9qwm9222F3rjhM6Y5gD3OYkRFEZ/ZZMS7H5nUGxJV
oFy/is98Rc36G02F8tAL1LObUbEy/9DwCde2O5SBYWz5kIS1AunLrvsAEfJpwhXU
9nV96qDeD5oa5xkX0rsGZ6sQSmtzMunMFGfBzJDRlVOM4e5qp+nG/xoVfrDDk3e0
F4CexY1LP05XAVGuK49r2rdgdJKc8j9w8q0/vg4kI+DZROi0DnhN2Qm0+y1mmDwo
3zDuzGI/j3B8/LdTDtt6Hsup/WLFlxsmvhrEDNaalhIf3DoFRsCtCrzRJ8ZQlubY
VyefXYrQ/vG+g95kM/uBmkhT5qfLfaTwiwQjvMFjHJ9k/sIwOz5rL7maY1Eaf+7P
KNH0LhHlkdzTqC/b803hLbKKIPvfQqEOnaPZfkUUP5LdE6WYoqPT54haYtJKaVv6
WYCc6jtV2AtknpgHdmBxUGaTGhewv+Voiz2pgeRAb1TdF31nU3w9dvgKd+OwOgjw
JOkefhmYsttSbkb9SANX5NmZsIDiBkZOn3xmKAT0TlvkAfzdw6BYnxv6BeiOs/Wo
A+cO9mNlnxxXvkmkIoQM9e5Dne58ygtQy5hYaBCvrppjuLo6p6FevmvJrbcSc/SX
9Bh5eeGpG3B1KPLSXiddlvUEPrVRndrgZ0n33s6eDUvkS2vg1424r+jsCcgQDsZD
foR8x4R7PO9EwNxu78AzYVu2S4KaG23qi+opo7i3Oovl+i4a/lkPGCb0bZG+FyVA
EEjrtwiZN7uoN5u+A0vlFhXUZG2gvr+XYrZw1LEij6wuq3W0FnMQY+satgfK573n
eC4MvZLkVViaxxmA5VfmtCdpRjF7L7m2mlt87IzQgvWjFGpOHvlH1hU8I/fDfBIF
hWy1ydgytQN2EuzaWkFYOEpI+boJGgmTPD4EN+J7205PUl99BydSCTdeTwzHZPAp
CsBpcBJnh1tmPIbU3VG+MMtsO2qnJ0jIvzZH3SJtcyxyZHnIdIVGVsMfwpzYitfu
9muLdhUECvy+bdGC7iJDBheZYpzAUTS3ZLA8ZtpRzLF+JtcM2qZlW8zoTfmpF0PP
fwYfzqD3AswImtbj2CdPCeGncJTJYPIKSSVs6400pe/QRblzzIkO0Hsc5vTRjfuP
wvZFeQBiUxg4xz6KJZXdzMYMr2gZJCMzIKt2Xhq9HGZoMzya0CjA7EaXR4msMxst
umM3VbwYctaEilz7dHVdNiWPVUhECJ2FVhpHMmPoM+6lvVlHCCfTEPWJSD/niwCx
kN5iLo2+NhyepRw26Yi/PcelxPovGLXzf4NQ2ZDLHVQ5K6Jw2ndHA+bOc8zDstMh
mM0ccCjtSF7uoFEHnd+cdjkQHAvNXMY0N1bvD8XqSaK21OdxL3HMgRZWipQtjCTf
ew2wYJrk6xuyJhpMllmc8xAZ0HcEXVhxOkExRofOXQryOVaE9/pP58wrRo5XaVPl
2vSbII8KrAvq08vLE77PxKCBXyuYh5kYx2qhC8b5BWNbDiOPuPCm+HNIKpyvXNz3
KdElt/6ZIwJO4yTXsQYp1uHwTlvRLy8FKTFBuSOuhQHTpecVvQRiw1RmohnGlifN
JQ1RRqa95uv83NR8HxLYCHHs2wHTsbcHIOVsqS4yfveleHCC0IISBma3UCQDReo1
wuZ1uhLgCy1JHF5E5ijumQWI20IeKbcdlBZIEcwVWMebLObJIW+clTjwREZUiJgY
ks8FNl4r/RkBZSdwxjSVqy5b7wXfMGAcM+evLsK9bVp1lqaclG5TaZVAo9OwUJwC
bWHv7mdY3suMUwdbVn6KXKoR490dKIAeQIJ1cOaVFdpqxGII67yl5ooV+oCRU68S
iiUJC0Yt6mN+bTqVoA+pfG53yKF/c438w3RAZTzDlwIwSRQLIpnKonbULkVQMTq6
89RAPfHebMVrSmgqnsfymGelwbUk9kskiJh1FwkIWYa8we7bcCC5hPEAZMnOISKk
NPvYZ4cQ1lDcCCkkRrHUsyvUkpEGEbhI1ggeU6k+xr/pTAOwU5SxqnVHdPg2VaIu
gGn9AuXViNar+NX2LNSSR287mWZseRviPDoW41TWgLRdti5Agkvpxn/QDChsixEg
O8Bmc0eekM/EyC9/Nh9nq1hHq8M6LI0hAFcPjL/PKb08exgJkzL0uHH5ra5mIMnK
yzbFfdAxl9OcnCoqm9/6ZD3F/aK2xP03lmp8anMq4Z0MvCJ8vzn+ROaVLvKNfMDV
b4OrupMIq3HVtzAaGIPSJEa1ZmxCD1mYrvBxMZvK5sADQBjEiwWylJ2sjDIprpqD
vWLd6jDnPdfyuyfnh69qVfQGcBRndKvzlTtS1zz2QNeLElWM0QB0vZWSWV0V7Sig
+DPiTVvzmZx6P5R97VF+UeIep+X2EGMiKi5iGOH4UWtjKoVvXgtU/5dcZRrkiC4o
e1sPNTgOFiGMKO+oHRt77EhEjwa8KJFe/ynA8lYntUjeHQ4ZUy5MCuD5HngiKarp
WasSmvttgaOTRgF+3ACzgu+i3reSXSelvSAzUp/KS/D1HzSWq5HcqTl3sTVYYOFU
lCu9/wXQfrZRz2rS756BSsfYjp4psPM7oxNmSji0kPCKAweXEfcBbbON/6nA2TrE
GUK8WoM9JKdzJRNI5FhpHilimq/K6cOZUFu3B7crPvnKffL5YhSec3sYv148ilt8
gm6FMVWyoAoPqJqLPzzpsqaSwapjjllzubUv/q6XqG+dUyVinQW3x13prf9+WtaZ
AkgtXOdBVc1Gal+hvSHxNYHBe+e4RhNFVLASVxf2XAC+NsXELb7MB3c0st6VAsCK
gUBQAs5j19aUNMfTWKrIxNSbVv29rfz/TtTUEpqDpmfizAsyrLmUsGD3utJKo6aR
mGQrM7AC2glnXbOkLp6YhhKrfATU60URjX/BEAkDoIRXG/3Uggdu6j6ofTU/9qn5
gjUPO8R70hPNam0A20H4jE4SH07sheku3UtC0iZOFC49Ian2wpcYEnXQ/DhxnK8M
oIw/1EluaZ9bpXEKC/YYzQG6yRfIeqNaImbqEXDYsXCi0NvLFj3B9gV1wg2tltwZ
l7RQPWROsdGMJETWBpH+s8NYQB61aJNKnxJSVMsQBUK02W6HRXBUr+R6rJZK78Jc
peDFYJgEQkqUSQzaFt/LqFspI97fQxIP02BuqU/rT/2RaBk7sTwqsR8IaNbzN02O
dXaqE9JjxoMAP/B2CtP3Ukd1BNmTrtisireuGvF+03RUkbYM9AySWEp/wcvvNTZZ
s9Rjy+MLgOO+i4HvS6B/aC7Zs9zki1b4gAsjZ2coUTHgooOU2AWE3469/FmOpIJ0
e1Im+DYDtkNBAloetq9c7RAlJc/tdV2E5D5MmafpAtNNd8XkId2sx+uc/pQOHWzf
YlL8gkH+ri284BvPeHNUxcSmbDkiVcjwYw0bxCHjpkNc8Zhu1Mq0befmEyeaXa1y
opunG06bIpXKuZjdWwjG1kYZUVekUr6Za2mY1aSK0pDrnJPEnqsa63GwXFb+X3Uk
rdNdVom/SpXgJpqNWxX4LF2EwvF5eEB2TTGR0EWKjNmc+cxFYGx4rLuWxWoI8qjU
Wp/6dTZQtCjLikexCLixWngPvcPMCYgVFyERKGTdeJYLX5VUE23u5O37evAWqzD+
HPQfq1t/IyqXqeNw3/tAefZS9s93F11cVvtYl29KCegeiCQZh4fV21tbXVTnYTji
xxDD/X0L45QX4utFmfu58VDUAvsfjOeDRk5Ln36jMLbIZ+/j17CL3beM+F4vyjbg
LWAgQDdEZo5t9W3wKhGDrCkRNLD6UvNZfkDP7AmeM6LRdXbjtp6mNjGNVSEXkfr9
nuFmTaLvfbZsL5EhQFLU8t9/psjxWMiOhrxGrXEB3sM933CmvKX4CguPllkvbVbI
vma5azjhyHXTc/iUvDWmriYZE0XV5FEjRljqR57Tm3E/Ng5DsXifWkN1msf7vFeJ
iayqkcbKD1Uvq05cpBfe7w8Mj1n8SC7nq6bE44DWcOs5VAE7Qyrxz4fcw1dqVbFY
4DFhCONOm+9H/ktNIm76U7vc9PuOEeMI/cKl1sn0vYLIwgxAXmTCnuBvRaO+39dD
V+29uALaM70u0StwhQYa1x5t28I5Q3bwjgHAdlDGMW0+E5SOEIs3NgblLwXrTv34
b7/M30vgL81Swak/Ux9Gk7a7NjEorwcs14TuUP2mBVB+GvDkOSl7z6OO1nvbEcwW
XNfrWSSJpSk/kmZ7iBBw3imSCFKC8xzp9ZpMMJ+MViyjB6pu6KMPkpOsrfOxmXD7
FtQDuVmXXZeMCVI9mRLpPXWphAzcqt1f4LYqaouzhbEXPSxCBBscvjE8gbJ/5wpO
Jk0LejIWpXljcJC5voBX+wg+wQ9jGGWHbsTWNn+V7212aPhzCAIeYk2yZjeiooy6
QJ5vBcLQMg2rw3pchqBLz8IIcZW9yDMIMtMm6zYsBXcNZ7qVczB2TCGIU6AYsFSn
7gckfm2A9+67GsqZNTlCxXb196Gq0U/uLpLD3h67cJOfCnKUy6TS+yNGqEIeudX9
x1HRUSZ6Il3bOYeGUs/nJhU7nu6EhK8sjftKDdspkHaHCl8C4gCfuQ6N5kvT1oZb
0I/Ew0R76t/Hk0jcUH0Xbm8AFQY72TKDtxT54OoRhvMwdBsTm9p4UrbYYKsOjC+e
03JApy4Xzn6Qnko3RaDgKE8ip4R5E9qOhScPHbmDqswMEPA5yi2Z2px3Ufi2z5o1
wOxzUUkqSUtBrLw65GT98fdFnWWtl1tUzfg7GlWM2mltTZRbIfFVWVixW2zyJ2Kj
+obaJ8keDMQhw8B4fJqJfgqLFxVxs2GnErI+qMrforRerr4oagd12imXs+2kK1dy
uDzudKGN1yULpMjAd/rNWt8uarMuaLSuys0zG/A5cEtj+NM3rZEyyGSsYxSAS5HR
WniAM1vdKpgqdAC0KVjFikqa/6WNHexvIQWnRDe6g69W8wR2Yj4PjMKAVuJAVr/a
9HECGBhLrZhnclqVIX/uwwlGvhqkcw8tzFzIaVB06jZHiBY5g0TGhjKneGPLAXt3
1DmUavrwjrcuvN6uwaxzp+1sStAX+sNlBlf38+hAocZJ3X13lSfFC95YbekeLdPW
qghLU+b6MDyaa2NJ/b5qIHrjGGfO6R3XFcWXbycM5v1H2I6TrFvoWJ3ZmDY7A17c
RbFC5wT2yBgg+XPriZRItyulqMOJB4gh8yKQhgd5eANCbj8l1qPJePZNtl8ferRX
01n0S4SMk8TOmlOvwBBwm1LlX8np0330U6alRwdQgYOlZWZ7haBsB8UocmKPYT3s
BfVHcLjsaTD7hmcAD4Pd5BRDnf2iAhxZronJOEq9N6RVIr9PFHKlWLPIi1Ge25RP
e10HtxoTj+1HZbbofUDXFyrECgv8g87TjHm28qWqHO6kcsVQEzWRCDQhOZ/yQ1oU
Tkdx/hXjx0cOipl5RKqwzBThBqQzTU7uU6V9Tag7X9LApQ6pezjGwerei6YIw3vm
+UvwR6meKmmnSAo/gv+z/Uy3ZBH3RnwzdRy1EEXXDnYo8ffWy8qM+K8ApwUi2M9s
sr+k7nTWchiR2HmWuP8zUrrXe//gG2vIPCkqtc8qYzeizgz56Lnqa9J6V+3h1DLn
hjyiM6+HsbNifmzkY0qwC7BohC0vwXmIjpcUr+zqk07HUihEkaoKsj3+3rabkOxs
RRmY45PN1SJp+S/MHY+xH83BppT/y+bmjC5Rn/pu3jiDbv/qGLeVO5M5OtXFDtLZ
0PJLUbkoNhzLrOXqNju64AGQsUmfzsg+gs/4DzqgDFxAY/ZBofsQq5YxpR4BC9rt
ANEeW4el5GLOzcXyk4gxyKfE8wB/vLhnzN4/TtnGaho2L0qH9d6YNOt7tO/y33Da
YjZtWZo2ZoMj/gAZSvxipqZI9ODux7fnwF15hl3UXR7GHtrdBn5z7VYwcZMi2VN1
2m2OCm2ZxNUax00rNTZ48jqfFSjGuuA9feG4NawOr0M4gObQ8OY1pIwOyU/gg+/j
+J2Mt5ik+K8MW7Fxl97foQbXjIluUd/r0g/Stsbj6ghO4OK3FAOf1k+CY6V+htQ/
ny9dGNGdNat51eZ3K5kIMABDwI5A2e0M7bx+uyt90fvJeQvpiZfOoq/odh7hVWq3
EtFAO6SQqXCGPqrxVkaNFGnm+Lj2bc6a5qzLZcv+Oqp2NBDMRedGpdGoh05u2STx
Kpb3pR4OjEsK4uHPkYva4ivddv+0Ug9vEVbWcVEk4i5Sl8DR6MbR69dxlBEdx06R
g1FJkgyqqaODE5RHb5Zo/o+zdtjEBcNOTzH3+2D7xM4PSALmISVq1nkrOSJwmv6p
Vvn7H2+hZtgNBUQuPnJC7/bQ6/NCWi+xn47WZiwTMpvt6EwqhTu4u21o2nYzPSlw
euZJJmE1r3X7MS2GA6g90JSl3jqLk7164VlTRM7zMQIHiL/yNfjA7tnW6gpDv/kI
FhqiBPMEfdX4RTjytLcZmiIv9GzkcKa72PG18Iqv7p+BlOIFdtp3K++Gm/91qYiF
0Re/CvhRWj0MptIrmAykL/pP8dmV3XAcYoEj/D1NXEnDoy1WkeRBer0ub/QS5FnV
Y6K0S2Vu8LH8cZxzW4fOmVd8dbOf1mwb9OH571m7GsEPoNyEcVTm1KQrf6tKZ1Qc
ukEv1e2O7961rPCZrTzgXEEoO71qve8W3lhBRqDPzMRLkq1v7SxhzShQq4gScZYa
iaGumRgcTPitzSgGwup9LzbJds87YnLOiQxoTdK+vRPbVqEk99hWbIW83hZMVMFO
l1doTi3yLW65oclRJjt0P/M9lPa0UJWsiHkCeiaKy9xGX50X782Waml+cvv489OM
AFf98E+fzgZBvhOdO2bBgvE/HNzGPOaOB9bgtMruhw66JWLLP408/Le4/Q0dbr4+
ZxDW78TqqTbMgYYCgBPmxgPpZ0Wl4Tga5h+/8onhpn/c8uR1jtJi3uok6dwgeiYS
E9X+zy0OV1xtrmKH2Pw9gVIboVn5gsqzPbyC719PlMdeTsHR/iG5Ag0t8J6AFEZj
Xubgdf5H0cFWy2Az22xKpY7CqYHgoC+hCDMsbsPu7uG7YzeCfGBfPcRVi1SBjlgL
f1B2FcT8E8Zuc6aK7dfIVe3PCzljWROEy21H5YPG8NRcvqWJjntww2sawB6DV3Uq
vuyt3G7EUBik7vlNnE3FRffNnwoDU+32ZheHzB2sIWGXp/ZGqeL6VhhMk25mMLF6
u46hugQaDD/bw/WuMn4X9nYAdrHXBjoqevhsYksG+vQ/5Vj5MgzcHfw8gdmDeWPx
qalnlU6bGu4rpMfYXDhtrG8pO7DL9w4NzSJ5JLMDURNyQZ8jHHhLgEf9KqnirVok
6bsag6J8gle0pHS5p3U4ZxlzRiaJjXorlBsFU4bkp825eELosFv5E58DwIz95ke9
9FPGIBXddCwt1u4BGxdNu18rcCJWT4hDLlBxjZxhIAWggISt/E2qf0RK6fSNIf7P
nLExq+GT7iqfZWgQJo9CsKRATZy3GlSe0egxs+B1NhV3XrFaunyWy7mDBGXZ3r3M
nELhULH/XPpjvzuSmXwzBezZCFWeTU+WO4SSb2HtsuTO73aGk/1VunpWiMwGGKyC
Ek0JBpOXpOppST5Uefp5IbSsMO/St70keGB2ZXAwngjX9GN36o8KKr0JrjVIDlmH
FKpyAxt3EN4A5cyJafsgpSJsUhYErzRi+qUrw6MsISHCFfFp0kD1rCn0rLN/xTbJ
T9efMIPLdzol4YE7OZbXYkZZfZt2ECRcgOKJYKchr7by+QinUFxNBCWgKy8PenEI
KFqXIInO4dmB2qVteCL/6z9QDyND38EnW90eLkrjxE+dkMXyYxe9c0Z5OzFnX86n
eA8aCTisetUAvRpI8pKZQy6u/ms8/SWo0zb6mm0mdVTM8O3P/wnd6k9N7HTApHZC
//tKVLdhraO3AfnvLUcai2WQpjZRCIt12qCdF8Y4uQluS4MHEVRkFqR6ACAebcym
eDKOUYICl7Czw/oe3hCDGz+lSobY7pfBDjIMXFTfeSnVQ0PVq3ZLacXdKLuGKbw7
+11azx78CtzU9O/m7WWzs9iMIzupej9JoDYrkHqEtjM0SiTUmCeya6jw0cOZmBo7
1V4AKbvr1jGIHVkguC9IEUSpasfIObfBAf4WQS7ijpJPWQkMEtmPUCLVM9Yqc0Bj
tcv4xrojbo0VMWPU2rEMiBRBqVU+4k3NhhiXSM1s1qH5wrO8eu6LBC6K16xVdFlx
O6Bw8p6i7UCJm5W78t5mJ50ZqaRlHSceZvXA06WioYRmwjW+ZFf5gNuitjpj+2Yn
zfVznlgiricVcG1ecmL145Jx3mp5GKR2o21wWEKc52pEforg1JkgTPckDAzd/LcP
ZzoMdRxiW+KyyHr7dk3831NVBwZO4Jw0y8v/esRyx1NlFlxe073kiNxktm7FPTKH
IhqdyOEvivctZHuJimw6ClrGlcMcQS1z1QoOsFgRjbzsizN3SD8CylP++KTAcY46
QZUYbuqeuunnRVHvdbsJ5N9iZ5htLTOBCWYh18B6A2Zv5f63aDVm4fAUejPXMPEp
Iin0bm/XhBgCdeSPIIREaOmkn9ZPsNmo4H02FDheeNpyWdqslcKLqTrN6gPsUzkE
tt70U0kHp2WEuB95eRA9RA6sVvJaOXhdOdCmb4tHa78VoYvNZ7vRWkJxW99KAIMT
WBAqVyn4Tv8MFwiKCgpe1MHNd/DPAXAtTvNdhQtBUveJyEhNKUNnHSL4UWAI/SEW
6cHnLGmcEsygxFwy1LBTWDQTT2HZSChmsJNrIaB+Lfyc4lMnmO0t3r5rdJx5WcDQ
524Y+y7uMfuse6b3KwjIuLEgNeK+e/yd50s1asU16L71k4JnqqP1Ri7QL7n3GVR4
HcvERVW0Tu3lnAQHPlZteSYFZ8cfBW+Um/WTPb3a0rtAKwRlLTJBIG0tb4TH54Aj
+M9CLF9LQh/+ID+rLV2ls6nMr0uy9xhHM7vgaaTnqA6sP8kfY7lIHZKSym5emCWg
I8JILiZtMmKRcDCtEpMqIoNQEgZrhqbP8h1+uJ5Sha8kbk81f0PFB6S3GBA20kOd
JV0SwhNa81TgU6mp3hmmRmuk5PXU4o+1IZq3SAPCr9+Zz5PsAtkOn0KD5RiTDpe7
Wzqn8U96XYXkuk3wUMkTq0Y/FZ3DWx+dyfa905CXzezpNCAgTuqIZNjJ+KZrkPbN
pZGLR2mY5Jayiet14Kba4c+akPJdpBwYruzBg/DQWInoNYRILenqI8hFtWttcWsx
QFe3bkFZOK7UszYOTJaSwWwG0NGfRfJzOpxWeiWbsMDR9aHqlRtSE8H8uhDuwGew
J6+025Z/G2uplV/OEmpAmo003qx1/AH5f0wj+4/piUgsF9sHqMVeu8+6LPkqLYaX
8k5fuOQSSCEhorSCJilWrmJZeZ88AtuyGK2zH7u/PHNc+X7CxBuhKUSjrcsFWzFC
YoiH1UD4newqlOoZsMiKUgBPv05DJ//Dp+P3kiHmmpHrdTpj2JV+oNM7JGDFZbaQ
6Y5Yqf5ycFyVsEFAX9xjWRIH+I7fbJg/BPyNhXdNBBRTKMAOGBvq1r+m9lzpitZx
7YVKGUM3U7OQITlVwlXRlLGlqlhsq0JJtbSjiJG5IuvjKaqEcg3DTjrFI4u0VTO7
YpvBDSkq1Z3X6wQR0NBN+udmc3p47ohUrI1HlRrNL4e0E6+5LCEAihQNVar9cogK
6yminRZazA3zwmgCECC4TaRW1xL15Viax/T/7ALY7dCZ9fAIcBQWXTWb7tTRRqF9
PquR1xAtFtqF4X47MFUTV+GHcIDJ/sa9/v2AMivxjMsDi++1x/P736VJ449NsJkO
00VM2oXX11ANLQS3cUkiEx5LwE3Zqw/tcfZIc9OD8whxjndx6x/pLl5acGx5i7cV
frf9jfEkgXRI6HzN3h6602qX8Kx5KrI3OTeRhRlovYdr9dZJWz1GuxxrJcAo20XJ
mmtcIFHlDE8DyzTJFMuwbPVEw+wCs8iTgb5kymBx12/x6kWtgZbU3mX2ptp6Lojf
pq8IwdsGSiK37yv5QotNZaEbL+aX0qorY+i8z0DfIydzd3p8i27fXLXS69dQhflF
SEBKswFLQS6H0NAauQ/zwJg5NHijDhLzuqlrIXEb+19Qi9yir/J3S6F0wOUnpfxw
h0AnlMcee9fxARbC9hADMhZ1o8gCVIvnkaeRGCNdswH8lprgPjcBUASuRbJYka3u
jx8mjq87ZBI7MrCput03nkg6PYqo67KoGiN24OB1i9u4W9kj2R3AXD8XOfcwWPzi
Fpib+gLq4o0qM3XaC5UYuZNztWDKv6AtGWVDZ6jRDbvjh8OW/RFd1VYbdlUDkSfi
RoFmaF8bvigSwAPblujvraBUQDIBw/SoWpuksqH4zEX6Sj4uW9XBhiGVgWYKn8jn
J/hIUAEw48AlQojdV+r+Vo/+K4oWZzxaFjXMvvgNbVsGUQwcZu7j/DBiW6If9MuT
39ICBm0t1hhBVzbq7spN4OfQce6X+v2FVvoTNe6LGvipqeQU+P3tLA5Rz4RSWluI
l7KMPQ7XOQFYEtRusfOV+0mYTkPE88Cii4kWqFDGn40WvQAqF73fdc6jh9tbyE/Z
C9HGwNEZ3pDmk+eAYAr/Fb2/fOjVXJDclcmrmDxBiyqz+KdTpeo/0aCif1eBwBXx
+UIDf1fKpHVdtvDKYQ9CMP7gx49kCB7JoNy/4kvkcQSxl8FidHskh86ub5yhK2Zv
bWD7m3ZWQmImGCuXYtJ8lcZc6HQLAQChNIlgpckNeu1PXD2jLejpIrNTGcrqKBgd
kNPXGOz2K/xnxdcMQtxfo9IOS3QHbwy/LdTx02OgnhJ0JPi/3bYOGRkeZdVyLIdO
bpBYzUhypO/A9aWxARzhTLHxIlbBk7zuLEoMoU0tMl6xP2THh2q/iHa/gwMv5KCK
lAAfzdxA4y9VH/SLeKaS5JJFCPiorQFrrWqfklrNL5khUomdBl/uadk/M6zMGQWD
yKWhtaHCI7HVVpHuId5rLJpd8tpTQsqz8h2h1Wlm2x2XiqL7hpYFLGKLojSxOrRM
lIhT9QyXDlO8uyDQhB6rB9A3UqIjjTzrV3w+R8sSIGeTwcdKax4Htjc9HQFijEKu
Sw+BE4VxkkUvCJ8QiBMbOgw6RY/RJAcNnwomuZTEz2NZDr6A4XEwrC4fJSOiGmkQ
DvI/8RP+haci4wpYc/KHRAoZT4iKnLLOiWCk+QdGCmvFcF+V3oGqMwpDyfIMQUoo
zd3pcEz6/ssIWY7Elv7qAiG5tRXtmPG3QEnkQ6E7hE2VBQe1P2zVVmiKMKTo42dq
DhZnsrU6jT4/xZoJnUiuVtaiPKr09b+XswMG3JeR9Gh/Ey8PgCgBS5NHKfljpnzH
lYh0top27PaWFcQDkYsRYKWrSlKRIHUcKcTIhhXzbcTUCFZDQXuOK7QN5H4Di16+
1mjUGYKlhOvf4a4BK8VNAp0f+bKAdHfXV8PEft5bmZeA49weuXKFgJ5x8NdRcGzC
WGN5Kub0RAE0eNod5GmMyD35iBbOtqagHlklKYvQHuf0lDpmYt8XvGVJuhmTd7Fi
Z/5Ou+XBdBF0C90ihxWofWJBUj1IoVX3tlKuK37YfQgPvXAhrc7iklM1FqAeQeTX
fqAVQqJY1BYhZq8/yMgpQjNX5Hme9yqVHTmk5xGXAe54ElTJB6KgRrdOZCL+MYa/
iNIQsZKXKzz8KAvqNla9LotJUfsKhmqeGV0ZgGDAFoWMCkGJqZxP5kJBDph741zQ
Cv67lYko+AF0wHYiNHE1MMAjs+DbhbXNTaXXTJ9POvH3T+J0X4mkgGe8g2pCvRp1
uNc8IsW0kJ4sK0p6YdQf9rbMMa5SJU3u8m+yuMYN3rzAUkX2JGsBbvrZmFdK/WzK
6X4lhDfFo1JjIjfhxvPdUmQupqsyuf8RRJ8xYgrGXCCEGhi98ShJTU7ZIU/1fR3H
LmXMVEWWfWlQvfqU1tI76yj7qPKg/Vxj8s9Rw4Jmb9hRVLSlTtgNkh8LB277EsT6
2RARft6vB9heSucyhC7WZ0Vw3+hET1o4TgtlNCrB/g9K+bTKoi/g7qSvEKoA6J62
8MJBtNqG5IgYR9EcvPk/rDqkPfQmnVsSzgHQa/UXcuuKCEIBTFVyxlrD1NUGngme
jdThnMOo7BCVu6XRbcJbOLse7/dSBoK95VsAzGjy895frNW37hak64EgnHS4NL3l
NkmJeMc6/PSOpf+F/YRxXVCzW89yNxxa8oZ+dDLxFHSi4RL8KeNdfPv86nLfjRER
VIuY0VC7GFrCzue5sfaNBakz81o4YvVvmxJgLma5/fZV5AgfAg3hi23zBRts17ph
5O0X6QggXxa9CFGirMOW5w5nsu/hi6x1ELpRCnfGnum+vMN6gR/Z63qA9Q7RTMjB
CJOc6J0ILKPjOyAZzrYHNeQOK39lpxeWcPoteLn7n5Yx+0dT36HOKtVvLHhLu74Q
PO7WKpYefLsvwdDHkknfThqilw9zBWNS1Dnk3VUoxijn5sXrT1dLARCOAaRACDu6
FSZEbLdx9OxshOBh3VRFxElci/iOyjn4w+OoVbV0peZ4xXtAR6fEucDFMbn3zhhy
gFauzo8VosWuA33I/nEUgTjtBhyKc0o0KGQwyrWo5VJ36vrratRJ/WyqmGKhDSro
Zzz7cldKUczzeJ5CPdbtGCLp8UfkeiXwMa6cQZSF8twLkE1mCSgHL3ECzGL7f5tQ
Df6JIK2eCGPrBNvd4tZgYqbRuigg4j/CdVDzJ8ebkQCPQJGZOwccvRgccqygr3Z+
+T/f5jsKQMAZSur1CFS8f7ciiEP8c5iVGJ8FpSqUpq2D9p2HEZ6BiCKRrytDzCL4
gPjR67bVFdmssdaIrPDEijmludroofnEWM/tpklNCpElk2X/3hyZnNnTQBPrlqQM
1yLZ3v6m909nQJ0jxaPJWGRgqDZwXZuSmurKYgVcDyLVUL32ByUSGfpCWKOdWf4U
dnG2X0O/2ZjTqtAvm0WojCXEvxUMcI2cG9aAMYJpoiCWK3aWnGJj1+KEO5sgbK/h
YjIUHq6hGZ1jswTNq12YuNqkpLeZ/ej05gs4vf4GytVvp/XJJj2WyJ3f53QuaWcs
gdB9kuVFMcni+PKiZ6yUTFYlV0TG+WKb22Ef6Pc3PaEHei+sQ4cMvaji7eoZ5myu
wfu31dkrrnWJ1Miyaxo4BFdlvlbW2Igk7b8gke6tgPtP55XgB64V8KvFHvEkPQMA
fBhEIDposTL/05ebJZhAJ5u4c+mgx5h4XGB0ocXUh8WHp1uPSenetJ5r4JIUm4Qt
nR2gmBIHPLsc6UOHxVKrhxwx0NEcR1Wm2hbjLbiJGPmE/mVvGUrlRxxEDCqgWOL7
WpsxwI1WVSLYgph6dFvkxiohK/fzLC8m7v3vockRtJDq6zlXlUFCnM/DWUgjOss6
Xbtrj5RdecL8z8IY9WavlQagpTsv6Djt40F64AtpHtjU2HdiHWvLQBI9Fz2tJtvv
iRD6fy5im07nJeFoqNqzDsD8vBDh8jAVZGpFesSqwaDkfciFWNDbEAtqbDQWwyUr
qUoPyp3+EU9FZ4HMEW4NLu6xO/HmQ2mGqxRiJ1ecucluW9YSuxPiVbvDOyMFFq1A
uFvmFaUCbmILVLHIhoCnQMwDlVRS4nnIGUucgU4zZJZ7rvEJPdBgFkXq1U7AIxvE
ku1fpofhZ4aVfQR0W0P+/hDYJyzV9hyZ4cG5CY2uzMKsTJ3qn7JaiXKulHYKk0ki
bIpg6NFgkfs61UH1BgAN+t8jQVaylGFOsdtseoKh0xiY2xXIyuRywVBaq8Ei/TRu
G1F9dLC4xkBAptrH9V+VujZDA637pIuWx5i9FwtSy7Y/SVELoEIeFJyNyy1YHAaB
UFfV4AVCt8oGD5xRsWICipjOhMsfXp4XjlwIaNZLKibqAQsibcBwiUxtoklXSp6w
x1MHrmqIY1Kv18GuFRvcszTRWuPDewkrPVYVlGwnLLTNRrM1Ga9yz/DT+bRkm30h
/cj2BpYA2e3zaPjAcNYGX9u8JEhTLBUMNcz/48F4G9Yrgoi/Ns4cJltaME1dqUyW
+Gu9fFoug9qJzYPe4QIrE68N52q4PUBxTsN/+uUH72kLgbYp8brrrJbVoVdKr0m9
ELyT4Al1iTpl/RsqOvxDBJa1ylnPjUQYxP238YCiPHtuQIInUSSALSVCALkaRbXR
tnH2qa+83Z412VzbuY2jc6yO282utwdyDVjQOoiUUYxd/UTktMzL6geBTGqJHZXX
FieRel1bCYZZ42F/4bcqPrlQo4QSEH9Dzltu1QYhGfbwbwL0OGtYjI/k2utnrcLF
TJXccOjwWjxKZz0TLBhfipvQOqUL7U0AWAL2jNXTnNMt/i4Tu4O/0NqgaYNolG+z
bZtO9bSfqiTTPDP2jP0zVgdvaR3KKoGytxwJeHVYDP6tV5s/SdPDGfRSFQgfuw3q
lG/KmdsAx0So96cZFHeUNk1ObpfzTdN1LLPGOMo26VtqpIB8jqva9OBk7kNTr2lv
ALr9v5ZOgBBX1CfmtFh3h9NyeY46TVcJ4ZyLEJH4Q86LZOJ2PWxOS9umyYpRN4RK
bbrJFu0dt28b99l6MCZd/jRJCg7OPIxqbJl80SWt5IEK2Sn4WLB8QJKWLHjbsCWs
AMrBNyRfFPcy6RaI8hCPCOj/VkuFuAgX4eI0pQxxYI6ef0rq39DO0hqw+8FWac4I
WkIspGII5mqQEdP0U946tWh55/Pv2HjgP+jN7tolaZMiita4GJnwYHpZ29qW83+g
FRhLAa8wWhM9nmjIUVoB8DhNd3ms7OW5nUbNO8pzXqmmSbMH21fDAz3zjyge446W
YRHZqiI4EIUkw4F9Pq/dS9lvKWwsdlfuilMXCzOT13WpldpbP0Ef3PM3lpyqvlbC
VcOJPJ0/kS+q9BXyCCs7dAr0aoAkutH02SnUhPN4pGhQMV4XVJZlJCT/dJkFCNfm
D2kZAu9ZS4yCQwBLLA2HHxZhDq7hztPOnqf+jzk4tqDYLgcl2ceioozgDPuhoKVS
wmrLts5RFmQPGJMQXPjZnCdFoLXKM4Lt1u22/hd1c/5Wg++Mur8ltPNVlVJhqtT2
K9hzeDCV0tXmXXjWMT3TccWhsSx/SEUE801Gr3FiZU2CBxWsvweO8xQ33ldSErDO
4WqobNJp3kCBU5FGppHPhlR6IFI3l6ZOfnn7L6EPv4qnIMBnL4MbHN6I2IJ4s7oJ
EsY+WYDt/Dmr7FP5tBE1st50ZNR25sm37uoMO55PTgIhSZ6JUZVbMB1UYNEddTe0
pNk94BdEd5g1fO0QGVNBtGoh0mOcNMx3I75iOp2dx9jQeS10jyYg9yZc/Nwq6dOQ
Dyysn9ceixSzhub24Q9RYAmLEuN9/Stm5uI8KtnH6LL6AKMNIQoKNPOIrD39ZafY
eCovoNMJaCC7jOTmlgGVBq4GZO7c99GzacknsDTEGJaHflJpKJFGGEV6jJ1bxr5R
tUkpg8bbStFRtWeAjgfSxffABNXVPQp/YgvlFLcd/wxEABSrW7THObZuBI+/2yLq
xm2zNaEhDF6aZgAhuvBivxZqE5SIWb6DtprppWLPa6eb4e5XSR6Zyte9E7ux2jks
8Fm3OLFT/tw22Sk2/7fa673DMNcxe7bXUuX0ZUQTYEICxA7SiHrfdiii39Yuggt4
lAsO3By77n7AbaIA58wDwk/qUjjz9Pzj/jmsvm13gazgnL7PM+hy6dYnQf/iEPE6
cyiScywrS6PxohZoq+uMFN7Fxb1EclwwuLxgAjnAOubCGz6GElRSTMH43RF0Fbwe
FSERH0Jyq0ZmPfO2UqlSmDweY33Wua81NpGexltP4OgZPilYu8LLWzDggRregjNH
dRCdu079RJbhWZoC1sCJIcT8BbY4UhA8sn/mVoRfC6onO6DHQfdwhFp8EjKhy//e
v/QQScos5JAWL+TKDhI9y8mnlmJPbJ8azBoJ7XJD/KiUmQMaKJcD4zmoEeVLFgMy
/IKkI2Hzy1xYaAKHpnFWkFwYnb5W2kRZxLoFHMxkfoK81/TzTUDQzx4bxdEmTdrN
R00SThYj4xdZau7ni7Rlni9o+wJLqoDLmBqY2FGWY5/Z+Pwg4iYmhwX9LB81Jzim
qaEiYZeInmqPQB4EV7wHDwTqOJKzD1c/MMYNAswE5ov6OA5vZm6zsF6bq1H2ZlN5
GP9lsdgHhJpZO4pv8ONh5IHYvOjNZZ+/ym4MbSZv27NMq4eKVdGO2L+gTveLk5+1
4wsOVi6PTx6SudzaFucjN3rL5O+dQConv3s4aOyr6r8LWHqvtH2dZ4LwmUsjIE/U
a769H161P7u/6FPC/5IuR8nGqsuxEYttXHnF2WIEpCF+VIFFSyE3UFvjaffwe1oh
MYkgAyy0V5lgcPHzyEBPAwxhQx14yEsOZ+BxHEK66nFC0S8E87Z7BKHosiGLMje1
Pmjt0zhn/HIjLBp9/8G8JVH7WWvow9C5jpI+npcC6T+++Eo+8rLDdNnL9pxkzG2J
1OwsPCTpt0wK05lBTlwFpYulofXiR68ZOFY2F5CQvwZJuHYTBillTTSqH/I6VmqK
3rRDnH52kAfV+Mg3mZZYQqG93gIKdlZYUCEg+BfHRcDcKhy8q70SK3aiGf+6orHb
Qmtmc2Wm9o2tBSS0m9Hw21gw/lJGIIo+Qb9iZjvl7sjae3nXGLt+368X4LjZs04Z
5axpzRmy0K+33hRTJD7tWmlC1cKibkhg4KOK568k0LBmwsnBqQ5XMAkY7hTTqtuy
7C83vhBxQlr0Yhrvi1hR4+cE7NchTah4ncWv488TBjRdR1YJap4KwO1YDWlwSv6K
R8FLKxiYoazqr4B39Xa2MVItDQFk4azMC7IuV8rLwNa88/np+jiQtYNFB5ccWv8i
nHs3jmyAKMTYmVA0sI6DE5M5Qqkf5OBf1p2aOROtw5hqzUBPzAe2gf8QziRkHqc7
quaaExxj75AZxuRlHkKbUforzD+pvqXrv8Ti3RfSnfKD3KHqy1VpE5NCjcKaui8D
7qXZhlMZTToolMcAepylka6WEOUfHC6d/ZmUdOyKTBPTz3QUjLBxK7dvKJ1djJRK
tVHocb8ubWIX3F1bX1raba7iaOaFfEPxH+ANaYPqwA5eVGlGHih9ZwtpexuvRicx
Cgpa2FltWFdTJljFM3JnYHtn+XJV+o/soynUf40m4no/h1J2ieihJnJRSc6V3MFV
VILc9QRSxs9LJZFP+CrAvVSv0/TinQdF0kjGbkXlNIfJvD22e2/jFn1QdKMHnpkk
OW7Rz1SaZibkGt2q1GYkcwV+GRRwSSNvJ2E9JGUKnp1T/DV2kZW0nbMsFUaEhKXx
xGLaQQE2CzTV9akqD+r25hay+xvYF3YpkTTNihVbLl40IVHbSBsyF4rci5Ap0ib6
WxQRJ/WrlJXTdqsXqZrZcvNVcNUC/5PobP2lKBOj6fZhBeZFpNL1K7kjBI+LPy+F
QmvXesMmQckIQdoEiKVWhd6ZmVWLc67TEWdlogBi7y8+rAc4ZPrxOEdMdXxkv181
V9S2K0UyiFRMGMAUFrqszOsUNR38UbX0ar9nqU/sblwL2bHdmCvSNSsQt/fsI+Aj
I4bkdziQ8fttrVflwsYsSm0zUdwv9JA2VdVoAKqyIfFn4rRsMGVoKbIeIW5+uEgF
A+wOXtE0AfCOMSrjKR0wYIBS56tJSZQnu/jNjdr/AExaTk/bvdmkZro8KCDyc0Ow
S5NuP1B6jV56mylnAaAKoswHvmJI+Ia/La9W6dOpb/2jrUau4aOQAjDLrmgSxeUb
pgC8Z5iJigYLoaQBYIZXIjSb5oEF7TsUIL7QG3acLwv9vCgfZ7nlMkkFQEuhF8a4
xwIL0F5WdWTH9WTRTaCetK92kTd5tgXQU5uoTR0GCx/qt/9WxvagSiAZB/OnD08t
29oNGJkWRKjKqiDCSDJL1/jSodOLpkdPSbzQD8acIkgMcPzgeegs4UFY7laZiKXQ
twkrCEuTLRjJgEl+IZcWnPD6jqNSrnvSqMslD6/alwXMnOi9j+EF5k75wbZ/clAg
cYbWyzoBB3BJAH0vfrCnPt7MTB9dpWvOuSZFZib4vK11POFtjeUhN5irRG6J8z4Y
U5lvDsOSAOkMjMCPZSjbbfaFbeFDY3uOC0eVqHfcnbN7Eyy1FOsAZYWgKCS3VXt0
AyGrchhDlxAyk6komVXFhuic4PgjIu/c5P3aJxYDYsZ5GYCGqOssuwpo3+kvC6YB
cLJfJ+Nz0BrmKsLxST45W9Mf+OQXJacR4mbM7He03XpP8ivcWY7B7zvDRkRWD3TF
0L/9hgy8hfrCuEAtJc6e28R815N8lrZfecbBs7VKjyRJaz95ugUMNsB23GPvJ2fF
o+CbXLoV/kGt6+42MB7NRAalEMuGAPNgUOfLlCqqMFRbk3fTnKPqzi2npZqGNXh7
nLEefrJW6JPHb0V10wd+JzoMHslge61Dk9uZPS0awHmwHVckvI/Q/51Ni+/q+ApG
76AZcOy1WjEdmh9yA7lnarHIgqzqX6XVYvjQ0QC76lvuotoa8EPIhp0EZnm+K1Mj
/Xlrsex2PXeAqnj4blHKlOSDui2xpz1BATkLzWBtdRaTDYjLM5Dfmuvqo6ROWRtP
uLX6bljcffQyqJwuqauG13SqXZOU2sknxOmshGdHwE3W+0hQrZrvipJJnTRDYRuc
q7wbh/mtdMDcZUFraCS+FgKbtmmlWpL5xQ3yWKQ80BG/dTcyur+XfPfDIeN7evUZ
Sg8FzwL9e/kxnj0pbysaEFEoRyzBa4CcqIEF/t+W9Asp3lJje2mA4HdjxYy3lCFP
rupGrMRhT1EvdfTUjsDSTax/m6VJ9Zko6cgpU8hirhycqsEFyNVIXwQY6A3BLDl2
zOUDgB7HI+oXDbK/Rcwfor8rUbQ52b88vVWm9DDFyCj/nvy0VmfEeEbDHE6N1Ioy
VNjbDvLjI2m5fZtJWPpBwxPRiWH+a/6+NyoPLcJFytdDTQY1EPCSAt79U03QIgQu
vDIkrRi/6VjINJ+ralO8fS9T2XS6BwVvSgXzWttYVDY9P3FnykiXzLT9uJQXxUBe
GHgcun0UkrznK4iXJJt/GTS5wqW2+oC0VAQ8ZfldP6+Hd/AC3ttt0W8HosDnM32x
TgXLhvriVPih4UCL1bJDnPv34AnipKabJ1m8XzXUZPof8U/XWct5N85qJZGDm/YW
3Y0p0pYW1RlqTnsP0nAi+IAOJVkI28ojIHFEcoMuphsqliLqzT0Icr8GsVjSbwdW
u8/FBBcH+GBwlq+thf5zy3osuZXfIDWH2d5sS/AJu9vLY3KyKs75oyrtnsmZarxv
TLznWZHgvi0SvKqYVbI871B2A6jg56RDOnbizFK9oieWyxeBsIswC2Lj0r5mzPT5
DIWuYmTtxsoOVy9lJBFEjnGnBdDASXd4awnCTjEbZXl7+WXWst6Je2xnWEDXcmTZ
185hXkY4HlRoTt2nUnr4RRkK7jyxjWqZT9hFO8pSk3RwP80jKQ0EouOkfS7Q256S
W7i5IhxNEogmPXyPKO/zUPWTBizZxSTqAB1zxY2aqBdwbz1q0cUlglMh3MS0K2k4
mVFVKWaKxSqJMsqJbQ/G8+IFoyi5BCt1kSDBvo0uVEiQCSbF12HyeS1ltpaPjZPE
ED1KkbaKs7vMhaee9RmALDmjUtjT3Xo9DVdD9ZPRotm9cIpAM365na/HmmWNPvvl
JK4KaeRA02wH2BLdiyT3NH/TVKHNkpngaOVNr1S63F/2FjfMXWJyckx8J2LF2trC
lCYrLE1CqLBvxuxOs/tbWWsGIfeEBk4qqXxu4CfC2Nx6zILrsCk2eMjhL8pcrFmt
8wTMxPID5836Dz7H/mAaANv0qVCewsa97uGgEN58u6hJ10fZ7knqQvj61RbE5zXX
r4I511pX+yTOxMXSJmBl62D7PAmRcfrR9puG70Lle0PCUzWvCXQVQ8BrVkeE6FBZ
oZ8+bi81Ruwg6jjAc6j2xdVKP9qoc6M7ZcZUyJAhGgURpG1MZZgvjIn2DUFfS4wG
crJ0K4jGUahRc91JHm+PeRDJ9sAAKK5dcCisJgYAPqMneaiBSahuAvEKMYofTU9X
7+IomNV1Rs6nUBi1KCI5hdC5FNuYbM6n9SAr+G8MT4wVFdQ8RxwtkHxb3j7Gr/VN
G4vHAQwn8qgDWmfqq5QgYatFPbiOrfbxATQ/6XTfrLppoar6HvqYvaQmS/caDc2T
RMF1g++dTSXSGcpTqhq9qqIBlQkk7FJLSnaJzqp1JS4CxYwmfvxmfSX40uompY/m
n9D3t6+OlPLnOo9RwFi/tOObc4mXnioJ3Tr3+ZaS9bAHHLPDmocO8XYVTstGvUmg
Sq/jxOzXsdlxuEx87jDoHF2yh6zz/hJ8lO81OnQnSykPyNwsegd8tSt1JtK6X5y+
tUYkQbIf67kqIGnXLkJb4tjNZ+fewsZPf6N7JLHn6cAzAZ6RVQPN5QrY10RGw6I8
/4Oc0Q5RoWO1kYaUov36NM40jXkCPsvIW23oEbrAhdOFgIkd4FBsysWUBAElD8Zd
yBQ9dT13lxSQcwj5SyhO5vTna8LbHs4F1fi6kC7f1kf3i3G5AUnOIgNb8ylqRNbR
B9I6onSJ0PToqsROA2QRRrTSt2S82rkqJf2716eSPYbCPAV2t84VA50xt3z0tFUQ
YIQyEHCgOIocygC0IeIzTg2QJyRCx41S2U7Ng6ftFrt/PWhLRFvrhzbygDLm8MQN
nB6EejNm5v/LiFLvyPgtWJSxtU7K68IJiFMcs2s50/vv7Nn2zcqGb/C037IixmfK
T6OFN3AfP8/lVlSxdFfkN30NbvTSH1ts4alZ5VbnXNkmnxFxJY8Josryqd06uW7b
ihPScqwnUwUa40PhTEDG7Qi+iVe95zB/u8+b/UWT8FWkVgEXXLinON8rNOrGH/fT
JZh0SCbuWfCABuYxdCBDRfJX5Ixu1x2epU8y9TLCPCXTH5P1APapSQwiPiN6gyg0
x8NGJC0QAl1f09Ne+ltUWJdQ529bIARq1PGiTvtk8YgwwL2hQSTaMrxnFMpJgYOx
UMhiDjK2cZpLbz5+XOw3qzB8SChpE352LkeG+WLOnOOVUZPq7LzmFuMJnGY0nXqU
rqeyN1cEk7Zr44P9LEG4iEGr9rmCjaLt85uLwgJwiOCTZyMVAFoaZv7zfQ3berO7
LOYprYZ6z0N1ETcDObr+Rl/QCZv49S350LSMogmOkcQQmNgjRBzIRX5biVagyLjc
SIFwJTqXEBJsSZPrDT3V1B1fKkPBYphNypzXx/yR2hpZ8+sAuO2iBFjPzrbO9+4Y
dk1COOJsFc+0gGKr7rY6k/h566sJVeYONlt80+D4eqeLcggBCfJlxBtmaCDietUd
GGcb27VQtMT0D+Vb/a/S6ftbXpkpSWHkVzPhqWkPurCtM2hkCnCqCvEtd1ECvxXc
fGdQ3TyAJ8hYJ5G+3TtdTknq6/Shn8blkGz8K2wGyIuThlvCatQUs9rWEidZI2PL
jo1R1zPHIhA3t3HyYAoiOiOsIPRzUtMqjkPeLt2neOKWZ0WFt6Yt4NpMuakokydq
rw4YbxyZe3PlO1SjWapIw9bdl7+N8oNTy6A1zk40w+zn7t8VCaD5aUoL0YhAYFgw
qQLIoTsu8PaNgqhQAADIDpFyZlM4RAxNAjSB156teV/121FmmMxd4nldJ879It4S
lur7X6HuDDZL2r6E7afcvuNQ34O4aBEfV6Ojf+gLuLLQQCfWAntKLV2wN0apt/9P
FgHzQ2LU3m7WO8NexbhNaIqx2fxt0YzoEKCeVJRnhFIGmDgmzPAdWykbBBe5vnKf
waGmU6AF1kUvXqB7ezGVxV2qugGIBaZwb/RJPZWMNOTk/LtCW+IZxoreCMCGgun2
UxDiKNPkPm/6vNj+fnZNn5i8YlFY3Q+6nXUwSXofpiKCSNncaxW28S95ZtDUzcNj
LQsw/zsJgjwRfdCxbiF00m5DR1OG13JDNXtwNtvn5PCctQCbRUFyY+wcGcUUSaU0
QoGccN3SW59sncIMv1RI/pxhkln3ZtK4AJRupq05OyJjuTnIVini3JD29GhH5k7n
xdQMq7pzZa0jd9nTuOmKKQGwc0qF23E0f6ITijREyFm68RxRPomFqJFJdUlt5R1k
CzraC92UvL2wGnjWu5Si1zjWY/1ZfAx3v2XHADz1SJx40n7Oob91wSGXHQUZIGUq
4RLbrfaNMKrDPOGpyINji3K+U/rPzGBkPCldurpWi6kqxffYMXrVLu3oSRm4Rlex
kN9kywqnsupWCUL4qD1y3ANN+tzdnjig5Q7H3990TMxjEqsCdwD6LMeo1e1Ve1Kn
3U4VvZJwNlEVz5GKwr5zofWUpJntPvsNhVvqq3xi77XOwUPCB7xAGuY5GbPmSDaA
hxZ9rmFjJPqjUIsQ8M84SzI1whmFSOSXVYtdfLXtpA/GXZ19xCaAMh2XVLMTJi0O
Kfu7O4z/VRWPLn6D/ZyTfrQ56PRusAnc6dpeSFDpJ7V/XS5f7k0v9MMdrmgzx5k0
fteVf1kSD4ZVMgWiMcOuKIPyxIEZU/1NmBMqOvfP04wT62AF6OK49iccH/jawx6F
RsxlJS08u+ZjPZl4G99tLA+77BIrp7aJTZlM3nB1t5WiHOUoPM5ecQ7FHZHMm9Wa
Fglsg7fZG2SSlWDS3OGgMo/1hAKDrSnz00PRf+3tyNmYMdpfi+F5HfD/Nbse+796
e1yemA6y60MPuodltIGqLSym6eEUrHBTS+IhFvSIk7vzpQucgGHOiA1pvPzfGYNI
G3uRUvQk0+KvnA7RugahnY5cQ3BxqPFkv09U5mERyvgA1Dmv6d+UxiWfTA4exIpL
6wMlhdZyGfCi4BSs4cC6Qk6ZqSbUBtkboTbcdRShKX4fXVrc+CGdBocVG/l4EOiY
ASfx4HSh+u9eenBCnN+gtVQiEv+Ihr1aVhNAEJtn39M9t25QacLmjDQLYpATYVcU
XKAnkjtKAwtDEqcr6ZRBueJadsMb2bgbOOYvM3QuWUZNIsUxWhNVjq8A2+Lq/rC0
3gpK3uTK8RtJN+DFFq+yNWmeLnymUZmJsHiFmO9UnAENAeZpyUjrmUZsFC0NOE9a
gqNVNTH4VdrDBc6Q8B4zMdOE8MMw94j6IsAWsge2Vr9JQK/ec6oVp4VI2mb2g2We
lzEZz4c3VCtpKxO7KBrTkJzaNHAG6XokVKZYzlllHBeaQOwDeo5mr/+MONQhkLlc
zGoIvxMFekVtWWvC/VOKeIInN9dI3Ll/ze/eoO7UMgoTZeBJBJ04BPlrf4wPg3Ky
T4HvzavauERuINkBjHxpK0dsRPW+52ZIkTMibyZSOh5SXGxSYG5FFx4XXgSC31xM
gTqr+XBhC3c93I4vvjqTv9hUmFRiK53xEIyC11sDiOtKLBHgaklAygxjm6qdzCAL
yRl9Xvh2+PNnjj8vj9+ObFJvD1sT9lN5zptHfTBMqINcoYmfRm8OuksXw2GDUSoP
F6Np4w1B2e8rKJSrtYzDSOgSDdbIVkg6+D6x8ou+VSIoT6YxF9Wzod4PKRbmLAGR
r+nnDwJYDTul6uVYXSa52WqLUjwXrTMR7ZmIzQ/7hZPoC1B2Q+YF/nLoDOOL8eMj
mDCurWP14kSeZIZpKrmgIj69TFdG9GzFrV3Ff2QJNgTRJxdoO88J18ajw2Gtk2mj
NenNOR5xH5i5tgyr0JLCSnoKNHCor5POPj8Jo6U+LeEMWxYQMPsnHPrPDHv6ju+n
LKF3tLcxUk4v+qX5CqLMhxVr8o5UCs/HreAU+YTWEx74B2ABa/xZQg7aJFE4Wm6v
rVa8R9g8RfKRhLeY00Nx4DHGaHhn5hlDbFFQeooPta7zoqx6afJtdTNJeFCxm15c
zjl2ljZaClI+X86KCu8cr5pGQd8J5V1CIHsTZW97j7zS2SBBDQTcCw/qucjSqIS0
VdYH93x0W6QtgZJ0vpuj1EFR99NpX1spipfs2gmB1WjeiPipFCEu2Wi8vCYG6lS+
CamFWRqReBntSniMkBNgGQFy4mkF4VBGy61GalDtZrpIyu1CakgNFdx84qo44m3D
GrkDNaGxJOHO4YheDv87I+cXsUN7gyyWzDJ4qN26lsRof5NzOvFH5w8S5xIsAi48
IIhxrmewTCvF8886VChzuk0UNvXcwhzESiAXni3p8Pmq+d4wQiXacvwVziMGeYwu
nP8xka4m6ClHHsOlcxCKDnLnpjqNXMzbMeCEs5a5pOUQb3OvS1Di70JCgq7veLfg
EOdqNmPe4eddHRGyLvze/nYo9zXWXJtqvFvW40df8LygmRfmijwhA47ReTStXZMz
R4g+/KpzuN5AIQH7DNOsNmsp9UY/wJIpxhwlObGGM1kuPABfmXv0pj/Q6gnJIS4F
b0rWY7HE9mPBJ/Nhe+tTmI4M4qizxvDb+T6LIu3k/EsQGSsCWJBXskpb2YHbKCcc
X2X48Rhm72TNCr4Smg9QONlTj9Aj30b6XfgUjMZhFgX9skSTeNPx9adFULtlAa+3
N8EoQc5yQ60pTlUNcSHn3ocmZ7eiE95ALWfPRf7jO64rVtCNbAEsD21YpU0M7E5o
nJ+L6Pv6GTS2kRb69xH2yU/hpuWlk0cs/ZQsuXE8XE4h7sVec+GVSRgP8NITugWS
0zQe0kGFerHLKLuXySG7lEVgOe7F4Az/5MUFAllmNx8bBY7nuF0pDBCmq4ZTPEor
MYON7Aw7ovSTIL21tA7UaWOLNMugpbQ8jAIWeta9ZPrbTaWWwDxg7bxakdYH9BBH
Q54JpbbrtlE+eznpH1xtWx8oa66SocDgo++0idzHzSAAVtiHOZBZPRktq0eDayz3
gQYWH7IKUanKCFczMVCwWb9EAvgmUZsOru9ZcysqvQmxs+1YRkLHW5as0l2vwVym
dONT7Zp4dbHHxqztF1mW8Bq/mehT4IltUVwor0w7ZM/3BFy5vnDNYYQ24NdlFcrI
bnPI+rYKlSjSMJzdcR/hxKVG+xbK0qX2vTyQxznzcIoxdRjQs6YWpaA6cdacwI3A
KZxoiQ/m86kkdtoS6DlXNQHZctueJNbEsxs3co3vMMBR1noGUPoGBi4J+S4PEpdX
+nHeAXALEPXKMs2JeENTTK5e2YcDvOSV/ISzLSssnRSQEzf4MMV5ssIICxXvpT9s
ZA7Lx1m4Q4CWMUZl/VYvywomF3iTX7NmspeaBlKDfwvndjWgzkhn5JtA2ADTaj+v
40ZQmXuzPQiG+pUpDBJnTL9It3LkOKzVfGsSCMD1nV95xY6zfRb0RHHqX+/mDUZo
yvWqVXwRo/tlQ/sNAcS27h1nXXUWV8qfqF7tJ81bO2tOf28CCD89MZGI0zByQuv5
fWqThmwCbf8dNk698g1IlebDCilQ/OPu5ggWehLhxcrqvn4MqjCAQpIjEWH1kIeQ
EysMHChkouxtX0b5KYraCcfnhw5B6x4yQihrs4mvieEpKsAMZDrqXxvoOdm1kxNS
Uo0mEJuzbKdEsWnU5KvKUFQtZKZTRLvPbG5j7w2u/cN8YfMalMZNcUdkBRo7tcRe
iUGYvRpmVVsyQNlXGhjLJUlMQfJIAJw8wTmmC4Ln3948cigeRLTpw7i2Q8hVG98S
iRr+G+74gByxVu5u/6VFODKpe0/paEyemM4ILAnMIVjty+GBtUQ/sgZDZf1btP2a
iAPErouMm71L8zZDpyQwD4/Tss4d6/5FThNUrGZzsp5mMzzmdTQGDE+0OuF1/5IB
0I5CIKA54v+7/SOPctwMwl9OYtJEikfj7Pg1X49irpGYEZ7zXGh1QrdF09LoqSEo
9MMiy/gksNCosWZzU1ZAnOYWKBliJR/LsH4Fo/zlaKOuAo6x1aX+enX3M6/qSWua
Y6nxIrMpJ64RMEpKBr17fgO+dmiJfTkd27Cn/M52hEVoiiBEJjQBv20DeoQgv8DD
5iFnOG9mlHAKaBbtJiSctdtF3gi+ozxEiMAvKQ1skPmLD4M1C+tK6V5Km2lCDCf9
/jJGAuY6pZSHvR8/Pe3ZBnPk6VanSLILSngefxi4sc2Z9AzWZlwnRI6w/e4ovbB+
K6Lg9g/j8kE/TYDwhtIbpxhIykxCSbMVN28vEbYm0IEUxXaC/cRwUNtj3y4KXeb1
jChAo5DHcmTdMjJaQYwblMfnh7FqAiuoDhxjuZbkPLj3J9Q4S/1tJAKUpNR2dan5
a/pq6clSsIFHDW4ZgMZQez1vvZ/wGOJ14Y1tIrC1DRzvDrVu6SvshCNchNHTDjK5
Rg+1Zw020HDMoiJSUYwxILDz6H3J5PwbB79SRrYcOvA0C5cM8I41k6fsvlmfuINC
XkfPYvrgaq+MsuLyead1MzGBnQLBwDqf6vw2FpdbC/020yJAG+5AzBVHQsx5bsx8
4HQh9dCX2oETtLdIQC9hTmjVbWzhK2SjfgY6a6e//xw8uUvsH5JBHdj7T6kQpntI
IjTrDLbkCEy8kf9Z1d9kLVSdCWrtgNHgnbzn1SKpYyHHXAYpEUq8PFyq0+/+2xZB
kE9VsN4bLRQZNK9Jo5zuIjsice+aLFQpxBFYurov/QtYcQh5l4fD8cLKMJWAkhiw
1EAXnn7SRZUqSg/FwoL+UJUmmKtSRdK+uU96RDZ9xLEa1haXexNJrWhSVY+B4iEu
sH/687Az97sgiphe2BxkRUR1b/smhmIE8RpnUsMrHJdfShl3oiD0jZxXT7gPYiQ2
VHh5h89aumnfO2a9ARdYdzjWojfj5sjQJ70mTheY55w+BDnjMe37XJea96fSXVMz
ewMTKFmuZY5XPTYwIIx/u0QLpg0qnqeLaOBjSi6OOGpPOGDTmxrXXMvE77CcaW9M
5ZLoOfHb9xHA2gATtc+S+01xsUNAbyfsXtKeLxQlXp87pF4U9QiVOj1DltupET4d
clVwy0BND/OA3Nq6Wi5UIOpgaLp16FdOSb4/MBkmzE9t+/V2Jtoq41KMhvsQNWv3
7A4U1MqVBShL3F1j8odgkQwERtxyp/9LdFWhuQ5VDV5bAU2/CQuNDGzJL9yPhAJn
5H979r3kXJC8AlCEHKUC1gpujfxwEnuClf6wMFpsOgCdxpyA5Dv9u6DFIjJd3BnQ
OTgDBjSc3oFFfD66vHCPwoi+Ly+nE5PW/91Mz6LDqT1Ebn2YUv4IATbqt1myHgdf
Xu79mcLzdgakfpuHhp1nS9LXsM2H0VvmK6acwNU0/IiD4HnjVW99N1tPDVp0I9+c
kbWMwCwZHSj5bIOuRP3R6+HJF29EM+sfnhVnosPiN2XsPOM1gmERSGnXlJj1rfpS
YV2PD7VsYEz5yM4iBGn126GNPPDk0Ck3deraR3ah9zOdtOE/BRAEgjMlCaEdRCg8
xUhVAHxonSWbdcU89gmxgfOFmKxb70djT5PiFTX3lyHf99orjq7NTNGTqcgZyAmZ
5DAKhOTXRd82YayJTEQJ7/szxdl7bWBbfVfga0ifW166NDPxhCNoUib4F6Gw7IOr
WNNFjLwBxtcSdgMiOi7imPIEsqmEJPvCR3Vv+Y4s7jYTSgCqiRiUmVgdcF0RCA8d
l0/w6PZQEGcqYHkcwMPhvLRy0Up+0d3zUWkQet1qMGObQTzo8x9MaW+K+T0r1Q3E
4HXn5ASe5H2OP5xDoeewhLR3L2rplmne5v1v3o/caWtmjLFrHUfZ2hhyj+VWbt1i
dFjbsF//XuyHFJN530FTUJ2AK00U0Uvfwuw3Tpswxs60IWEd5kBmSubYFgNEXvuC
7MLC6L5ONkf9fjNW6Bkombm7q1qPJmO7w06psjVc7UTQS2TSiG3GgHbQlZgRdwRJ
dilo+USuZe4twUqUFprj3hgt1+GPCej67lCqnMhJOfZ3BxJ1b6hejxyg2o3og6Ei
daS1XzbAL4GLkuWvbkGRpVEVaM9PsbMhqQyUUHyMBGD0miXQZbvzuC+axzqaPmaq
ykp8purBdSu0EEe83io5WwSPuDkgZ4MrS9he5RZAOKKBvPXh+I9D014oSF8x+KE6
QZp7MPxLAIZHNp55OukndTE9Fn7IKCfZH9xtL/rCtY+PHmHOGnOK+DMfEymyyAOI
giXc3pfj+CbaxKFvgMZTOtm4agdU7a4qn2DyP+GRuR6AHCwbxr+84hDrlz0CDmHm
XvgYwNXSIQt3+8GmM8OlxJd09f0/+vwUfS05npeziR+o6dvvECkDMsgcMMkd9Y5G
04NkMVWdkF1nj4rUzg7sa1nuHyvOv3TMbP3ixv+oo/Eb0ADQ6ruHKnLi4n/erzQg
TyGhNdh0U6nP7KLpR8xZiADlQ1POapuWgEUmQefhCMc5xsizFQbUbtjEM3WL35dk
i/w08peTNNGrTS1sIvZ0AIoAt+it76Cid2hOAIavKNmOwwHf5L8h7nJHm3x6zP0w
7HZWZ5qALXukEOSRDJKqmAfTzR3liEN8tRfrTjKkLzlDB3H6ONXKE3KkBx0pMz4g
lk5okmfYAMyl4yXMENXDUD66DZRQ1dq/2ouXA5VvyQrzBKrPhSmc1dpqIQF4SN9X
8ymwAm/mcEJ153VdCm4v5eWJ4lA587jr6itC1d6MbFZwmAaPJlKjGFEMEmmIon0q
fc5cMJaONnLGx1LF15JMJ01BcwwoL5mAtcG/tDxY79+FSSoXSUyMQlaUEHTxg145
e94jhbAqztDh632zPnVACwJXK80BBWGqAeGZbJmoLrQQIvFkjVtt9TDhEtEBEOZ6
FZhFY6ptrvcz9AksahFJzvsENecOJLDUK8Won345I1yv3Xa04NnFmTSU+dvph0CL
mZAjQrl9iMtlfsxVkUXEf+ncHN1UH4PoxvDhPPoMFObdD3wrwixuC0HZ5XB0PxSl
Bu3SIxoFoObmDfdjsU5DF5iUH8K4Kn/IKfGle3Ef8uzOISukLWacdQBhtjwvU/vp
CwFVBQWp7JvbtO8tdRgZ7zEwHFQT7REQVEYxQvGafvhES5Oa+ZSby9qh5mFjzUjR
X8I7L4GGYVGqDtzywKAIxAopMgcdG1SYHOBefNrzcZkGSwja1fgeS3FuglQw9zrL
Er2BsRTD7VMcaf3I4tDNRzmFDttEO0BqBfKV+f/9WLE3/G7SmeCGEkBgb+KVAGPa
Tz7t0NqfhhRNMIwShgmJCxDxV0GAgRXBJTkVJOEpPW8X/HADkP1XX+JXBbJ4YiWu
95zRnBD5m2KuXHDU1OUj7wST6pbmsASLf/NFi8FFus50Q9gmEFWHW2PLZHba+2jd
Ql/vP0XvMe2+bPJqv2tlTJoy45LXg9pMA93bcCvH9LUVvSQNWpCM7ie94DEApU2i
p5HPwPeFjSQnxQzl0AZdxvQiH5K/lw1uJNPMyQtfifaWV6QKZQvRr6+IejXxDwBt
gD8Rj3UkYa9hHdUxeeT63d7cF8TmFVD4SOAhr/yPcfkRSaJePE9guNRVEW1kQATN
3A8Iv9gwBYE2XWOhTDkoOel4jzMUdvbVAVSEnFLj1hA39PwaKq/WGKBVF63enAUG
uRAT/a7vDva1Mjd8HI5P4ZBvvKroclNqz3RgNPUIE0G9+U0j5XvOlXLfSAWtIxtc
fdpTI7LHiUOHdYW7ECx6Qy0iiYJtRSx+rcjCmRku/9NFx+SoeVRCpbb+lOfBYTW/
kuqZ9UUf8vFIuDiTUgaKZUe2y0D1fhc0G5kwB+RqtOd40mk6/Qa7ymJj55CQs6ak
5DXscHB8XwapwY7wWthrfaqom7biFa24BfkI1VUTLGwNE+9DDfilbi+nA2zYE9aB
bUPTpTuXdVKDbdSZ9XLLPOAg8OVVugLd3/XP+OTFAwmPrr4/moxhRS1ITYi/F3tS
JDccTW98GaumgXZGsHj5uJMkxmIFjxoYu7XsiEERZpwZ674iOKg32TixFeuWt9Ru
/nS0NPbbHZrPJGCJfooPw+lFXS6+nbNV75lKE2cW9JvN4ZkR5X5n1f9kos+20Pv0
cBhyRyKHkjuhwcSyiQF4ok09c4QBLP3NWzomu3su5/bo3jm2QosP+ndRyDclnfW2
vw8n8nVjqtPmBpnDdyeRmRKrQWNsh7nm8Xy39H3ysOZSAlQT7tPfR/E7c1mmEcTw
nkwROsIKHMDHt0eD0bnj7y363eRGTOjuoj7FQr+QuW3TSt6h441zGGDAjai+yga1
FhcXSjFTzkl1SS6gkSZ6RO+t5MMHn4qvn0QhuwHpiYPXDkZJqxz9JGeAi1ClnGWv
Fxaa2bMoXYNYwvnAOXAxsiAW304VF5E/X0C6+ktN/dDFLNYQsQTncWEjHqZEBGoe
aXPQfh3Aj8+CRX0tdseirWI0z1Ulq943o+4DBA/Xm72hP8Hx0b6wDadRVLVh7MCN
hddCrh/055YDbN3jV6g0LPTIjs1Ef8kXAxdrpwQfj1rAetLLuE5TaSK38wHtPQ4L
15m3bF7C7Gs00Nf7sxp/vThwMfQqJ7ZqbnJj2jHY7NSgCFI3X/yUvEB0usjY5Dm9
RVSq5QnSImCtWM8G+FA2wkRA+YTTS14DMzMC6v7lUVuw/8KcBHXoJXmZqtzD+HiH
1G34mgblxA/SHIvMw3wSZRWbeF1d390B8qFU7upqNJkF6yfz1N184l4EqAmu/0t5
CE+CdmRQgxbrrVneRxwtTiCEfjHstk8R7tPKy9H43bS3L6qzy9twAF3iCsd5tmWS
gfSiX16qoirdw7OxG6q3XZvIyqvAYwtVuuZ22vLOqbY31LX6L3n/bOXJWK5QcEAK
4AaV6NQVEZB25SM957SwOm7UYs2duUe/1FPzb/xHGRR2fY+h1x3NO6MuHKc3c7U0
K4VckMsqKXtnnq9wE0VytCMyMotwQnlSDhnfhDEQ21QeE/jOLhYhcB4mRsmOd5to
cInvcjzHAV5hNJx56EqJqxvWiOGfZC+Mpq4DkjbvH8Oa55Oj1ndAijHG7ibRYJhC
+uP/cHdtl+Ad/If4rnZm6L2sNQF0HChkhenTI7xBi13bKC5veLS6CRnZwDu9dF3B
OniJEw96A4D/e12XjDsM2FQqQZB9sGtU92pKagoFSzwkkSq0/nmYeg9JAbC5ZT+f
Hznis/l2gaNMD/02lUKscCiMN7/13MegDijtBFeI7a86ofjbp17q48DS456yLAub
jxtRVMwo/6twy6Qd9Q9yKBPlrU1LUvqg4lBPdylSc0sWV1Z4QjpkkRV4hPmeM6PS
I069IzAaZSl8b+jHEphv6GZTh2kuuu5agyNJSoBuwuHRXIYByvSh5SEmOoUm31Um
9X6q6KFKWOFT/PmQ8vVcJ869LLcAI8m3qFaeQYqaJqhjgQcwLgyyHnHMuzzoARIB
w9hO4AdUYShRKSTo/stE11It2p9NUTy8rShkzvQ3S4G7QcdCPg6UP8XUnOAiZImQ
tvRsIzkrOEGm7j0tQdXgz/3MYcbeF57MW2ZNlblC23xK+FIdVROghhHH3QQva3kN
wl4xQRkX4NmJLSqpj6f4WCWrCRO1gtN3PV1ZtzaYGYoaFgGiwyp2mytPw3Kh6Nnp
XEr2IRU8LP0nLysQnzCiicdlS/7LacoSTdzplG0xgIVG7pNSeOBLFpCzar4MdYa2
lLa09dHm05y8h7gxwYzDNaKX8mPZlErg8h7QptwDGk/12ACl5avutIB4mpZgbEiL
5V6cmI5dpPwIDrBplU3qcarQ6RdHzJ//K3o6G23pXB6ymohdJ7oa7IXZGRVPJNve
VNtgCsIuWPjUF7CKF2aoceh31X39+IRK5dOiUWm/NwHSbsH4OoRFfBy865loeRPv
10C9yDx7cQ4TwC7W1kCAthrvUGlIRJezZBCoER9bdQNdy+X8VfeY+MP5S55nZNSI
1W0q3eDZ/caoOI2IceWOExlRapZ5kDzcmYhAmb4zB5RhtinP1qlpRHn+PyOAdcsa
GuZ9zcYVCPyg9NxJbQMRovRJW7jpd5alGXGwXkehnVBNYZiiSaQoOzLXGD5lIg4m
pmgQdxhtf+r1ywNTz8TKhQ9h7maxc45xaHApDocMqVDT/HDFSrlvsXyCz9dAPcfl
O6avLtK35AZwYah0Y/kVBmynjnzu28dyUH439CyJf1iEIN2iDWzFadO+dkA0H9TU
siNlcJoAArjN5v+DjMwIBEX24ig3fQKZdmJOVotvDZimBlYyJtLXKfVs6fbtuWWB
sLfW1I5nfMwE0NxoL/QNtyNBk2RfqAACnGWAmONPmCAd2GX191BHTbykPVlf9aJo
jeT9xX4FDDZWu2o3Y44Ol6j91VETU30FY1p5gW/b5DlMDZpJY+/RGjDW0Euw3GPN
OweYk7KmlPPBnGLH9RHDs/jm5GmiK+73lPhKcTU7cptTQ14VmmRKvwbMiPhqZt/A
ftqgO40S41g/pieS2cAOe6nM3WevE6zocjAYxymr6GP4UEYjG+AaYyoKHbwR6/dM
kjeAKxBrx47knyCac52Q/y8AoIink2ufNsxtJHhfW8+7bqld3R8gcQuYotGWo1Ja
IzM2sNMygQ59aJs4nxKqMzOWTqiOZ+MmZQ3vM33ULoOLzGZZbiJn0MFWwdYoza1b
yCkcVaH9+wMkxi7Q1A07C/TGORJ31h7mvVemKjOSBqe+DM0BhanvBGJVNnw4JLWL
Ex2Hgah1cgScfgu3IUnsjR1wG6lOHajDs9i5MZ/nPGkOBHp3ueUhIaq3FUFsJk+t
+yInVIFWgmgD4meX1MuyEKaKH4zBfHOrH/aIPTvumvGlrvn6ZU6aijmShuDMhMbo
pDmV6U0kbZ8Oz6Xf7lNusnnZAK3tgoLUMiBuHOa3vvgbYRknzXOM8wgOiaR16MqE
8Ifpi4Kur7FhpzQrnYmKdmnVT9VaF/iSgqRvWI3r3iegOIFDg+ON9Qvebq7jRvx6
gB9csPHZUywUKPuH56LssW7Lxi0nFPCdRQAaTOEAP8RJlPCWM8dV5C5mBlrKQMj4
UAoM9QnZjIsDuWjnQizkrFvixb5pSoOw8D8HOnSRa8Fbp39tqZprykiCPOmU4Mle
L3ElRPFCgCT05debIM6rS8ICZeEkPbOuoKfwFfxJa2nPhdYRyZttRjJNaq1IIPzj
iS+qqA2jUsDlmU+pV99yF2dSl9FSWexX5lbMPvADf7TRyZTR35Vo6XDFFjVQ+fc0
8Y0q3UU1EDn/ilcV1Ksi06fwgHqbSL9VDLxBLRkhzLTbbcCFM4cP3evQjtDj6zrv
vEoQD64MB353PnVOUz/+Qwd84dFJDAbLTh6eX5MBs/xv6/TCqv8KKMQjEeqz3SMb
ptgVzgDjLz1R4jb5Z9Q+i75jdjHOVHHL2dO50XiRdraYxT7GUt/4HD9a8PzdwHVr
cK2rVI2uhwxzDEZaSaZI5gVjWEpEOSvMYuI3OKdyTwc4PKKMt0z461i21QabV0bb
RqeXEcgGKSvrAgFtQxufTD4lKZ26ltkToUaOwXnbekif5D3CWSwKlnmcBjCXGTwV
6YI50JlL5LNy5wRn2pKJ7dOjqFiQGi2j2EkmMebO0wvcYmQrVirPLjPg9UX2oDgA
qrfFWzioLrD1qw90KtY/3k0WBHH9n9BEB5Ti/0pLAdOmHi+m1frK2khpjk4DW0G/
f0+bl45pBibs61e94ovMwZXLkRkgqKXjm7bG2waIesucujJm+aIP/JD/Tnt9wSTd
OY7pLIbM5P8OXv/dm/wXvCWcAa8GFrGFg2U19nIVsr9uTxIoymJ3W6jCnHCFoX+f
3a+iL2LUc/IjdaR/+QRsfM3R/ynmSU3E56YcwkaCoy1mxIOb7ZwadoIsypUV3KKb
nmZjqOtxOfQrR901p/IMruVU/1BdHY4kwoEB1L5Pp6CeXA1j136Blqz4QWNDD1Wm
cQqTSC9/UT+k4xUb11Q+Ck4IpbadsMUesvRgsSZ6W+j8gb9E5uILi21hlJA3l8Lq
fbGTfQ0M9/nuw677f4+gsrIFSscaPJwCVRGMKkUBzVtIqK2g/QVTRfRyAmkbh7lX
1V2bOWofrkcBzojf6ag4mhjKJDcMmBuumEIIOTdvbnn2bzig/0sqope32ZnAbxQC
pygAuuAp5bxZssUetPphNQDLNOZl56E+BObSH7BRG/7szmwQ1Y0JeTDlHKQ1expv
ZJUxoii6ser2tw8lyUF7nhgvwedlnQ3sSCnnEwyUxRJmPlIr2it0jcbib4rAZzZM
b9tY+TkShgB0Fm7z2SjE/qrFDzZcTCF4PRtvDTjL0/i22wuwJvEaSkGI6N6ILt/K
a6FyduLlKnizVsc6X+F0kJjk2rq86Mq79aK9fPTPhh4Eas36AjVUnrr/5xyFN99n
hMIiEAjOtfyv5yR1Xsnqf0DMSO4rnVo3iN0EMWJC2GbxDFbVymLstlVIHAe2Uvqh
X4GkYYXeF/ugqcMHmMnaXSE5dnPsb7HNOnGLWuye/wlaXSAr7njh8IEb6+47e9NT
5tEbe8ljorePsytyDICWSBY/YRg1p2NBATaxPZOITzjR9/6ORT3Qb0iwmJ+YDb5v
P+eWSf4BZsjRfNAwDcULjB6DuSl7B885oiT3DeQg6nxOo8RkwIn7ybDQeOMH+gEQ
NfdB8T5/Y+zOGqlhpdO+zGMJnee3W2gGy7scog8m3x44Leer7C+WfTsJJLArlpmJ
IwWnp8pPoIs++ZwAL5IWO+t7lwvWB6txDfBvxsz0OszI7NePsdsG6c/TvmQhJyEP
lZdGgAXAEo75JodbmIbapyUiV2D4Z8qD9qMaMocGjV+oSd/qNZFLklkRvEMck0HH
QAWHaFo9PAtJFHny5c5BA4OMwdiMl6+74R9p1RM+Hr738VVcrDOY43jUowNI499Z
accZlp2e2hc2SIUM/DQmGj8tFn8R0hhDH5ij3cTX2bKB4izVU/v3Jll+BQT8VwPI
dhh0WAVcZEe7T6+eRZUNHmjgskRpbH4oEnmoYfPne9wvgabqOccaQS/x4xWAo2r1
pT5OAsgt39CBPJGIVgzQsZMv8EY0aPlwsyOy/82mitCtmrglTtiFjMoGuIg+XNM9
q63lbGnIPWW6+ULrolqDrFMfWvzYuSTdX5PJYNtdV93wnew2nUf4MuVf8Hd5cuRK
/3jxaOOS3nAIk3aE47cbrMqJpjR+XuoAD9qC8r1qGXh3bgRQH2hfxNncdAfFjITH
45gkrdn+UXArV+maWCUBogXvj0Uq3/OSIEPIOE+MriGVinipMJFkPP/U9dltVQH6
8JM+bePlW+ZUXw624XB1O8901An5MkqQqsRw9v2OPuXOvsmr7/4cg1KCqp4moOXi
hgC3iSv8x5Mn1S9Quo9qaDmQJrR78zs80epinhB1uR7OgTJE/Yduj9/l2Txoy85z
iO7G3rRO7leoM9pgqNibnibe14GUPORDJDZoL49D2uvNZcCfkZvSoUXHfu4Epjsn
XeU+dzpn5/rL8KybKMLTnBfg/cQu2Yg0Bk30xj6zIJsLS3mVpJSXGEwe+jCYYtGv
S7zHSCqlaVdIUtzcngg3cPDA/GTDkOPSltvqM5ZVhjxPFg0AhMNQCEGIcy3oJ5Vq
AkiK1L8eM42EmYWRf+wGH1QgEuZ6lNUwWrscMYL8J+Ub+TVcKAEisSVUy7m0eJCQ
OWiotGjwJfMGz/1hUHE4WuXbwR7Tcb3w/kKH3mIZ/1dr3lPMLOwtQudYQYiZ917K
uOG6c43ySS/x7W/OHdW9UxQ5Gr8jCUhCwlrIm2AtOqHid1YP8NJQwOrZHYFzn/hy
BzjoCT0GtFN4k0eTgGn6cSIoevtS/RMrCE+/pPs8dDM4FUJh3acP1YOSENm1JYns
WtFFhE14PQWQLIm6K++O3YkNS1ivHVukS/1cIMVRgMloyD7jnG9hbOwvzuIxRA81
Ly3TkavL8Dvp/q6MmfsxfOWDgT+rNbiqRf1nhV9lCEWlpi9BJcdqWRg81GC/hR/4
bxctbv7sddafJH+/4MJkBbHvPgYGdY8R8wb2eNILH4utU08I35Bg6d4DzWkHYAfU
RZP/tAzPvzRd/Ou3JggDasusY4g88rpddPNN31n7zy4QFNh8Cs60pNqJxin7mf/q
wnl5TuTrhf/w4Qd4ao8QbgOxN9T74/KLt+8TRVP+s4v+FnV0AEtGUQBR1j411UKp
B4NnL03uGK0Qvk1yH7xT2dELfbZBKO2DedjKD58PKzlJT0cC5vgFCX5pt2gCvbIY
Ebf+hDGSKWZUXlRH4Kn/1OKGAQZuGDHgT3oBKxGhRpHYhL//HUlTdx+dTdtvCgAQ
q4yjPftFrCq96+iQP4Z+iTbL3RZQjPdPCvFxKXKka1zQfoz7ieZo6J7bWojR2FNp
qHLlBbakRzRFumX3BjOCguEUgwAVcZoblSgLRyXa26X9UshQcd6qASFBkcrYARP/
L/O27QHwxsuoN52zrUqayY1N9kq8blz0KbLnBLqoH1MzTvWMID08aV7kwqUURq4r
iaT4GTR2SLRhEH8BKjsskoRKxpRL1i8ZnkZkJHVTpFKvKDsmaZld/2V5IHjwFtlz
ALVO4hCfWo7N/eZgJZy0aR745jUawWh2h4Tzu8JziyHKfPKdyHXPnTVzkMKiLEQx
S+CAgs7lvJ6Y485iIHrViMyC4cZi3YsY22bdKX78l2ZSO585xmo4ouomu/Onl4Vn
4/+6EwN95XiKXVfEcdbFlYL83iKkyXn6WxrpfaFL/SK2VsqAYRAkQSG2PPBLPxVn
bC1gS6bnANeuL3ES1qrOlpjI3GOSLOj+SSD2xBBDmsyVgWwTLqXQLIkX9WRfSOGz
MjfKe88ORMV0f98GMqBJ7l7tYW5V2I8wVu02PMmAK/TYP7Ms7y9QjDn+lvPe2Woq
xnU5+eLVpXuK7zQ0iDMW5376J9cpF71HdVp9/UAsjzy4b92R9M5o4LlI9+jRilAB
0JRSED3uFKiLaqvBpVVYCx0DdNo3rK5A0su4wn8/IYOY1BKf8oXyryaogJvzFt8O
sTVA/DeKcAuaZJbn8K4eoJ1B3Mpk5Jrxpf04iyItAohg4XTxei2MP/8n9iwshiG/
oxFd5jrdB2/JkvL13O26vpsWvcs7rtL41n1IKWAAZmnzxczkDchjqESAeoyghRJt
BqyUNPKxFHNYU9ah32Yo/YQ6AtsM22P7LdKV9nXXVLzEG3baUvSW/Iw5qCIyQmgO
3SrAOSax+a9YqTwXJRxesV+OfDWYXBftMQIxKAKH2DIu2F936ok6jRlUMrkKIMQA
1/xQCwSym5wVRiPpSiOx8Ncl2bsAchVOYgA6MB26DzVs4/8o7ScMh4S0Mrl2icvW
7mxTWq6gAB/vIHqkhEaDNUGgLXs2nLpXHwMT9PjQf+vdOaPCRyYmkof33V/nZgiK
D3ZGm6WZajQebNh6gzu5+Oy+3NxalPorarHeTOIj7mtSswrBgdYMMgnWDl9iXVpu
Rq8umMhvnA/JDSqid1ypVcEWVlqZM+MYtaFj/NcD687fw3+3ZKjqf7tpTtKqwzBu
0mIDZYo+RDxPIcjrQaWDRY1njkGXNDE4q6SlJiagQCb6+UtL9G4m5+QUdsIK6OFs
0FXd+MmK609tLmSZVqoZw6l723DJ47jOOv9WBFLGPAKdZBHbuezo2xNLMH8Gy6xE
3Gnh0XwgXMWfvd88dtZRjMs/amtFj5ScgZgKq2P4fZcdYs0LEqh8E2c3YYgwjwJ0
PJhC7AH9zDtw1qbnsKzjbEiU5qmkhOl3L9w+i0/slUPpNBu1ixsMau42NpdVJNmn
iDY9MmxNPHSISTC7qxXQI+LOslJhGTK+NQUMXDu0K9nI+JlIu0aq0r7ZOj409nKc
iGmogUr9/JPcJeQDqbVrjVQSuCVu+CO01DPpXWvin2kmPT3viIwkkhXFPdQQK3sr
R7LbvvZEmi5ChPHsrAoQ0k1zKvixF5jAJktYoKq7aqvsvy6xg8XblMvPmbFPfCmK
kgCE+nUZIUcVHvKH3Q7wY7boF14lqVEJBzWxk8T3W6TtT+/INsPtJT7cEkzyQuTj
RfoeHEcCr3Ps5nJULJKs72LdsIMwzcE3FLQCNfo8k8Um8Qv0B6MKbu9Orr5s4179
VKHYXzOHdszmr4WPeCwfgC66o2SPtBHg3gBofQbXtEnP2KWFy8PB0G6DVB6aruPC
BTz4Zc25j52V9BuDdGnoJejUBj26Q45mQoeuP298nFUjDMMrHa4Gojw3sLfXHCjk
Pc06rOEjYfAVFzaR4Coln4No5WzzzsYgcZo7+o6JiFJzMVioPFqaj7Sxfloa4wl4
XF7ZF2wLYN05QTw6Ml23ktvK8d8VafyUXNeBr0e87FoRMIr8PoUAlxfzwBRyIfzY
0nHolXGocGeU9XIy1p87D5VFLEJ/WPDtW5772wuVpfWv/i4eaZAK0ORBCB6y6INm
cAoFOW73lE+oAg/be4BOkYqZnl0JkXZGAetzxm0edwwmUogC4T7TM6W8KRtf7aSK
+a9UcPWe1X1/WskFV9NBMNffleXcjmjuR3tHFny5G8oCRoScS9IexQgTieDWDqxX
9iCDhR6PhVE+qcg7ECU9qi/EDzBKmRZeNf9WvzgI5zmvpGs4ts6pZKiL0CVaBwcR
FcMNfCnFXuuOaxurdaO4/NclL06MA2qrWc9hTso/8v8Sv29nebQ7KKfbbZ65/HPn
xFThlEvszBTQIP4SQk4gYvp0bvqk1Kg+G/6NbncR/H6BgM6J06YaGEejr+klvufn
B77DBm6789Q06KDYVDhfjBFlXPEfLWjfL9XNSEDe46hasAgPL3b+A83IuYqBKj2k
d0jQL9vKrZw5nnLNMbd6fII2JQTN6gUoG6wWq1ibEV8F29Jx59LUvgmgvPpZ/Smc
Id9huxElObeBeHlxE39t58ZzdmKrVze5wSOVtxGbAUifiqpwBx5Eqyv65mQEmY0h
NG+wYAwqqlxDBeE45sR6liFiBB6Wk6dldQ6uojm+YhPzBK3SvBpeJWOyjGv26pnS
pNCp7MXopF6sYx/CeKcK67GegWCzxrvX3p6T782bMeqO0xODgVto6WEhMmu622O8
MeU1EnBzOrXf2QOOQLIlsOlZf4CXlmk4gn600nyaAHe8jD619Vg0Zf9RIshKFJRd
b4OZaCICnTbmZNpbhjTkgXpk+90VcGSIrsIuwhl8Vaq4XcZPlr5TQjOS3FPCRC02
HERRMjPEtJvu42IwnaHjdxkGFIxLbUJEfB43dNLtunRFQlk6WW557fsH899GW0FH
9X3aWaRHpM0F/EMnK5Hz0dRudnhf8dVBYeSFY16YtxlitlbCPdlN6qQhs71Nay0e
hpFmmQ+LfPBApHFTqIt1pOR9hbggCo6GRocSPrymm4BTNhqW63lBm/lzkiBDDvXG
fEeHISu96FlD+D67F5f8gajXUF4hmdzMJct2nbvvWsQ6hP7UDTsd3PhyH6A+yI7U
7hcijtuda2e5KEucWnV4Qj9lSDQ3bk9OEPd6QA8DgfwK1+SlIeTDCx89ss7kiouZ
TYZHhVwldzVZbXOQz9u3noltPI3l4I6HSo0q5I0cHNacPHa297LB4CgXxHnQ8J00
AQqFBM51xvYi2P56F44m3d5j9JyAvoLPsB2+8yWqnHJ1Bt/Rrm3UdPNPWJkZXefq
LP7a9fd+IAPGSZcKt9CAXtyGnRYZ1K75gPC7W/aBm8EVG4UnB1yteReOXt5v1ldW
PP+pLKK4xllc8tsFdr+rSvX1EN3d5mpv/Kth9pw/LcDrU6aBj2esul/WKIli2tm/
F3fbpmijbqQYos9n8yBCJn15onGYKL1ArIdt4MZEC5eWte14TZPw7hnSfKHwElOR
7K1YHRK0MK+xt+5CA5fcdaEShxuguk8rB6I07K0GGgOUO6UgehfLx6slzFhaUh4K
sYIUW/n4RATsjvZQfZa1v+FF9mlwngw+QRbBflSVsvSBhUyR+P5hLMUgprHpNsr7
lkpZWVke13GZ/QQBgDJTEJvpasOOjoGuNPxBSGl6At0ddQCpQRAOyJaYqLmqF0E9
9K3U3Co/kpfyK8HbR2LHuXkb7rmD22hZ/NYgAAyakIYcLOmo8QyEYYokq499/O1F
+Jjen77nP6IsjPLJ17/j5uMx5GyayhmWMheyFaEnSFzDx/n+rZVPZK2ZP1YT9a9i
OKqlz4I9OzzC4RxoQ39mLXJrkoN3uFKGfKL/9ZO+145OpHdQ/wVg9aR0U95gZEwi
49BChyrOHXf244oI9badHCii4IJki95wcu7scd46b2kf6zt4RRRTuLTds7r4lrIE
3Xg/9nf5TI8l6ap4wRbK5xo6YlrGNaqLQlcptY+AFCedlKGtHFI7X/xGxY60gPbz
fLWrXyl4U30u3gcYYMD2vxMw8g5uj0CYR997dPBN/aLkp5txvDUh1/O4SItQubsC
KxMAkC3wNMUhpDLTVca1nBVS95TgEVdfLCIhECCtXERVXEyLNJDM3jbQAUhPpsrf
MgVaZGI1m+DuW0yWmTdCvQhP/vf//uVaEG+kzoOVIppZuP2fDUDoEq4L/KwkYPGg
ZEEDWdEQjkTEhSoAhBoL78ciw2NkKH/QfxUMoGlgKFrkqKS3BBHXMp+uE3qP7U60
xdBqdYFqcXkckMksebyM6PwBjKE8ibIWrh+zKNMhFappKSL8Yh7fFosLREE8ibMW
02JwXwYRMF9SDkEJp4uXRsfXyEz5VGek4KuaDomUvRp8MfECdTtnXYbevWpgrYWK
KHyTYg3hMtnpGYxhweLDO8NNulLyNH/3Yg5QTm8XhLFm9fzA3f2gkwE3SZe3iR4F
O7xOTn7TTb3FJqtBtMnK7RiiZUGuik4ANQiIcB9fdl4wsaKuQ3jUpPvok1fBu2aO
Euda/JPnW9sBXh77ztShGp7h6TybVk6qwiVrwYjwDOSyjawkYYQ3D/+8Q7+/SPB6
s82KkS2+JWAv34YDf1lAnIvFB/oJ7HQopnyyE/7qudeOj9heQhp6lbI9TFzU6nuB
rMdRjXENDyP5DjpOz1cSq0oKKBzFnkpDQTGXUnXIVWb6fAqx/y17HwftgZOxbzYY
mT0eOfv6AP9PwDfDKHSJZsD+bzlkSrh1J5YuJ6d4bZhAL0j1k4V/UP3TganLbtjK
ErdvCUrKLovxYWfRBYhE8cB0T3aOuv3ZdRCwjIN79AnxKhh2BShoCwf7FIYZ+AUB
8YTlEH+TMws0viOTAe03EduSOJaX7my+YiQjRgCS35s/kYGGxQ1WWZYFLngE2xMp
TcVprOv2fKwO1rTgNceCCTcGbYCjZoqRZWeIg37S4Cs75M/o17poICweIha7+u30
IoBr6Pb2Hx3VAqXvZB2pXlKgseQ5ZAZQZhulbeGqFmZj+1vYO/ERkiGUswU2QzS5
ln63zAk/5GalmUTCTylant2etwAHKYNpEOzz7vvIj5bu3AoIBr3+YLMylDG7sz87
MdTHbH6oXrkcylFbaGbS2jKfHzW4BYZrJIsHX7Rj9grH+OMnbjme5d2RRQkkqEt7
7kSTXB5VDi2zoysJvwXa8NOsMU5i3mPNthxse3t5SGWi9LT1jn4ChWo0fvRHAEg3
ELYfnnoLj9dQjua9Tni/WsvED4MTURyHfvJrL3WALlphsbHjSzQWOxqX6P1lLpaU
trHRyYnPn+Vhq5OqmtFyAVXbadMCJkPGtxRwO0SX5yH5A/FY4kGV+s45YAcjsxsM
fWlok8P2U5vtzNxzEPE+7xKJ8LbNTBDr+ZVh+McTtQ9n25+FSVoVVZrUvXulE3JL
S3FrN+QpLt7DLDdazINAixSFD0AvnV1Wi7leaDwA5Kyon20/v4+8yEaQx+AVQrWJ
s8r8VIgnkt7lP9dqWEZ6FYIBKO5KOjCc00g0u4jZu/BWBsxhqg8jmiIaqNjLG6kM
WgZ6iEdjEiqEOGgf0UTOtWcvOS8Nick56ibZ4BBdWoE2l1JS3NVVeucLj23p30Z0
8Jy4RkrOg5AyV2q+Q8gqslcUuYF7Z8KlSOfGr6o6kxHJJGwVoYharYx700eR3urx
JfFKoKo5vtke5WR84QRtwejrK1iAM7Pz07hsee//e3SEUHEu5KmDcnHVy5+avvEL
+OJtjI6u8V53uiZafkTVhgJMU46M7cI3eBJi9dsHxCksSb/g8GVD7XlE5b8Vi+hh
r7op7itDaSG2kTfVnQKFRcIaqHEYmEtmmY0Lu/ToBFyn+DHP3fG3vLtI7y3yGWuM
NRS6D6Pqa1tDg5LLO+jXf8/509z4VYh8gjRJ50hT1ChzlKCcHiyo8+Wx2j15QV/M
K3LcgMKLFOZL/AncjoW4Ot8wwOtsjYgIuqYRGRNB8cpeqQTe4ofyHYsGQ26XN8YV
tePeet04K8I5Kt4NHOwuiGbLLXcwFgA/jETcpAr5RMgAIIKOQI3CT04oFr+Q+qOn
wRG8oxY1DdgSIDmwh+xdA7VzUVfTn1Bs10woiKeHJBaJGp4V7UOwIuy7QYcFka85
yYvAELcXFj/K0lM5vBjlYiyiK0yU6OMVUgVjKnY1x8GoBZVlbrVHCMaUbIBTsleO
iKDLhyPgzXT2NmXcQ77ukMNzk3zbvyHK2D7Gfgob8IuEySyZEUSBZPkcHXJZTeuL
4O/4/RMRnqbW2ec3KhkC/kkUaeOrQGOp90x+CGN6LsGkKcWbNGVAAVeW+QdzjNpg
Pn7WPaYxPf/vg2PzHGel7CIjsIt2UIJvmAjIwgV9Sw97YbSCg3PDtMPjfSbqSWbX
mpouFAHhfXXXSZcpK6aZDFBR3rp00nYAY1zDAP8PTKwzG8+x1AMTuvMqYsvjVf+b
zevgKhmovLrTRqSML4UABOHm98rPGX+cXEcXDqKjvvEbQN8zNYp3Du4vdDw/R4mo
Kfz078iPLeOh5cC8B6v/wUZYWG0FNrOmrMKYAQYMMFTdIbqOELFRjsgBOgwElUY0
2XF2PaveIx4a3cjXUCb30F+bbUg478BAR9oU/KFhRc8hi7WsWNQnjCyLNahd+ZUW
AFDLiWAasgKTXrdP/AsqtJzLj+RL1NYZrqLw0Dhs9iISe67xA3FZOz5ZJx2aFGy8
ulq8p8NgXMTq59wGxOf/pd//AjXbAxcuYYA6p948RY/dBsGBA4a92jkT1sjfeTjO
KIEpUIe5ZIHoNHLhGWXMwX1Xabvdtf0yykiiFsyC0n9KVKqGkEnEi8hEhvKZ+Rh3
xpfrW/WG9Lpw+POeRfzHhK9rGa/EDQqLt8sMY+0BPuwr/LI5ZgW+tbZpyBDpByGK
eFGM4Qh+ANZWmwSlK4vif5cw4dm43Us3M8+TUWYPZdnYp0kvfKu8yCwg719+Xg81
063xGAIQqlGVP3bo7pJfoUv+QCRGRERhknN7sGqbeiv63XoTSflKKdbAeZgjrmkU
M3x2i/N8P6K8EBQReaB+t7eb3I2IZwOPD2z0/5VVYzap1jGKKxpn/40cV1Qcq8Ct
n5yjbJ7LAebZvBsv9lpXnwe0q6XKM67EvCp+YgL7NgjyYxxiWTtkaA7eJIdXkxy5
5uUSJkwT13jItk28rOYOfmjcgvZTbq2HPxmPcDQ+fAciiVcJicKsuJ4mfiXut6xh
iSuhtzfwEId/mI72yUy3C4PNSoRqpqAYUtMcyLsMT7e5qxbnk1FIpr3dS+XyRhKB
JyeOOgT9jPLaw7npkZfNz44NJ2gbpQ3gja5sFfpPyy3DFoNGVGpPzIfTY32MifZs
GJz4HqhwRpluNpupm5UQt7M4WheN46vBibeAtxrn8NPG5A3BplN60CqTGlkRkCof
6RitcwUBFfBCDoGNSRIHtplrsEhY6K7LGvIDTcI41TTwp4+7UqH2fl8ILxPxboOl
Q/NjZdyEBmkf+yBud7gzcWpi9n8Ha91ezpx9LKRruCSi3JV75+73p8gKejcXC/Ei
X9H/SBsmrB/HgW3GObUpe2RWc+QtENfAvqt0csZ22EOGXHjPaTdbEqF6KiTRUT3l
bmZ4TTvq0z6FOFSRXe2kmpgS9rVG5G8y/aMdCJUTvH0/zEf9hdKe+dP2yUCMqADx
pUxzZQm/UzhqVXEgHnIk3CZ8ODHE+6plSsaJV+0TpxSLDPdhP8XOP2m4BQNedIpC
oIENh0joalolrx2/OapRWKGXAOAnncaFciwqVNnYyHh0Q+uc1P7cemVaPgYHrl4q
rfhvwhnwJmJL+PrEijBGD20sTMhrjZ5kiqVq2iT+eM8a6QUuxpT8SAP8XcYsU/Sj
5c5FfHCG3hY38+xxuy0EG38AIFu8SH3tABaijNBHn/SlJJ7x/vPlMN8wHU5u9kJC
MWQ9qvHwWBP9eCJdR9NmWz+qQ4urfpgfWC9/WlsC/QYl7D77jVqnFAlCmTF53lJN
hqxPYKY2xyS7ChtZHNA+qt3NkWp2s7BBhjX4IojrRW9sdZhETe4GSgflWMCvDPqh
zibLP8BR7eeMPRLpPGioIad3WEaftgWcEhVC6kETEmoNYVCL0D6WT5M2JmyJkq0K
d754A8dmQV9IHOIJp8tzAmJilSHzekxqykmcIzywGYPpF1VuVnevuipm485Fg9Ho
Soa2gSD7aTyXBa49hhXC01DGxiC9AXSoX+ldluvlduQpreY3rFMdzZbdhJKuENHJ
l9HR+JPan2wTD5xPN+Gf5Y+HU/p8owPmj78V6wQwNO/PM/6WlYcX5knOv/gblsZS
VcJYTHG4DIzuuHV9rFJNd7onexyumpGLt21et7w37sF3Oe9VQUgmN3ZXPIaeY7Kj
4gqgs1/5rveBq8esUT1oqRa4/gGp44Hz0IRs1vogJOD0uc24QR1P6wF/vZNTBiMM
IxeKPECD8VO4qCgJ5xw2eRtPmpM9cns8OYFDplaZhKyUAL902L/y+k8HbQKo1rh4
+DJrrjJ7jciTItU78mlzvl0xu2KBWGaHioesyubUnP+F7IZ4mrPOJGrI0fyYPqAg
qC/ZGurTSOhMqNXfJQ6rurMps5mk7wn2c0WQd0O02NhmqCY1SXWo96S3k2CfChw0
U1dtwIOSEMHGqjk7XYrRRTWDyse/vtvAZt5Kvloosb2rS9mhwYQVCQH3UvqEy9Yo
dgCMr4zU3+qhdE0fW+Q8PfqB6+w8WjXJh4jCt20VlKgpYHAyG83ADOPk6Uz52VaU
pdN8cRqRbQjXAJx9y7IY2K+DWvM4PILj6jfJnVg8dcHRyuay476TRHSMKopRAHqq
XwPcsrMi279xPWAoHbtbtA1nQJoiuO4It4Rhk18JMsRDE/+EZ2TGhItStjYLpHbB
xKXEawb9K9ITQM1xNI431lcTaUdV+5hJMOdVhSCNydqVGW8ZAJYx9osZ+VvO9rdh
e0P7u2InBDt7Xs8nKKXCVW2YdoEoVIKYDjLmLIk5UtE5F1vokjmSo59FZySf9Ze0
3WeHgyyqPNxoewdNscS2Garn2GMsNaKplilAX+7kgkINP3O+o4nWuMBE99q+BImY
iYhZxVH+WwsTmYnHR/WXyP+6dsQ/qojntPZ+hj3CPMsj25AwlMxEZ1OktYPFQ+uY
4yb6Jc28swixj9Q7CkqgopULQZC/2dMCuE5TtGTAJrGHW7bHgDyDdg8W9Lmsb1xp
+3sGGipl2OcY+W5Lj4TMYBxd693rwPQK3R0FdekBdhdCM3yrZ9eItuRtVZW61ubW
GNRfn8hlLpAg/9w/VQCnS6koUROYOVoFpWAzORyLkHwCG0U1MX/+xQhhJBE3GOy3
LLt1Md+HEignNM060K19eZQ8Le/ypy7MKNrIUMH/TC7LpQNXWMqit5rFdqtoSq6s
2/Cp0hy/HExQbFkYNH+SF4b13Qgswa7SlwHAYPDLmyiBuD790e2JOTEV9XFNpAH/
E20LDschICViB6eZJRxljd6Deoh6VH06P6k4OzLucbmqIPUdnU24tR+WavCbDNO5
FGqgB46V5wgwNygoKZfuvG6a0LKVskP/O+2dtK4boGruz8ULhXRHdTlZIcdYSSux
t+R8QXKfIk9yep0xZrNjPiRHsMVriAD16fxlvlLWCXho/NnUwhesfLD/e1ub4Qvv
TColfV6W7Mn6xiw9lyxq08PgA7/qH1VjY2Q0FJG2LmZXrltvs/Q/43cDKZ9XMCeG
fj2S4HRc5tX1zVcpca2Oxzh3Vbt65kSy7HQpHyWFNDAloUSyDYlBr1aN8VpkgliT
1Dm2CVSQGsWdEIkYd7QVQf07wgfFV42wqZXSLG7EVZczy25Gu/D8IIQ4JH8f2jsX
vJpgztbvwzqutmPK8S8HyefcO9FaD8xIYZB8OKOOfm1EcGKBb3ZrWKzqu/4J3u/H
0zdsN7ky43lf/RkR1w6j/WxkdlxJv8Am6gxjIhkToQ3EHdD3H2cbMxpoCAyLZLdK
/aXYJa1jwqUNXVYKb++8WvDzECFhughLVvj9LeDTMS+xSv+LN5KXtK9ejkVXvY79
h2Z67XEowG7WbCye84kb/U8XITcY2QYQTcJ+ZUqE7DuVKoH4H7kN5GHSG2trjpkR
HYg5qlwXhRvchVmzAgyh1CVfQBavyF+A6/7cML3M4jaQNcVeF0w5rFkXEjFWkXpN
Rt1iFwvtBdOXYsto6njsrF6OFyxqt7e3b+E0pq9caw83vZBfhjagSdT9124TqXCU
jN8nqsUrn/rFzEWdryPVknXP0O1nay0ynZHQpJ4ZBbqy7RsE9XIEhPwVkQJkab9a
+Qi+J+pQPL5lc0JlGDQAriFD9I06Sw3Yy+KkaFdkq9D31JnSEEOIBBfKrz0buj3z
Ku7QiSbuIE27MaKe8f6/M4HteTHqJCvdnb+KAFFZBBwawgOnlN5m2unDQx7HNrbD
ctcJ9hObxvpsWtbfM6/HJT7JOFACOIXftA8uUMO+Q5BHqpxWQZgG12J8090ymdqz
foBYlPN1VZmJOOZOv3U0qiiDZAsEEe2c80dhm05UHReClkouDv016uApBztlQ9aE
tFozPxjXICZpgfkxfeI+3tftuMug4YQLInQP7j1reGLIx20J2WbiRlpJewcgvPsv
a+beWDSWD3H589L8yfnE7r9rO9C4HGfQKNPUhHpVaNiTqQ6Wo/99LfKCNbK57aAV
NeHldhgZZ8/DYyCZXyXS9WuTYQl0upzkRKIQOZEjY5JPEqB2YkWMewAwVVJHJOWE
az5fg1EYBO3npbNe23Z/rsqol7gqFOprqf33449QjbkHZinTWrPCSM4h6ixHaNgo
bQVYmABb5goHn01JUpnMPswmBwBTKZAiurlkfFncF8nPCTsHldcdXDnajyQx3yt9
R9ty2BKFSQWBqOJiYTOkNYHpRtCuWDBBv95KxqRcT0s0w1lyXKLW1k6ztZHudCgV
gtNOT0pPNPdvCzaPhgf2Y5FWoCgZXM/w36hxJcIXUcznErEc0C7WlQoRaFmCFiUj
Uf/bkE643moHbUqOhw6QgkFLYc1Gi3VWe6OpZieCvNaysefynSddUkXdLunJkDt4
7vaCjT5j9DdbZYId8NFg/vZrUT+cU7JR9tfET9VXhLqzn5tTpfo331QCDo7fvQQQ
oIQglzR2AaK+eQCg+1k1Y3olu1Cd8TbhxTLljbAC+6X9yjm0+CoIvYb0m7zxdeHN
nTR7CKNmm+/LqChUs90u/iT63o3JsMnO5jqQBd19Qims9zAToLB7KyFvAa7WxQ33
/6mCjlqom5pWZnk936PvRlbTxOvPwGzspH6kKJKZwZ0pEVEgoHrXFC4rH6BHUc1q
SceUN57ebbno2uBUDC/ib2rfrPmwGzgZbYZwSenSBdu4DF56FGARQ9nXsVLQSCTe
OF6qqHbJ0cs0HZrGxhXAvRwQO69y52XOF80UzIFcU0fxMEA0EB7muCTke2WDhvmY
bTyppi7cYES9egotnuDBo797jVZw9KKoVtJit/MgL1e8OOvP3lE/4BAsd/yEklBg
4Xd17CTOUkC5qY+a/3V6e7QBzmIOXSCvP1zstmMcysfvQvE4jeN+g+3lauIkpuW1
EoxqYRXCuKgSaVjOAlONPc/2I4xI2qRJNHmo76WSFrtE9kOZUJrDaF+R3zr7mSyZ
xX4+0+ynZf4474GvQqMJ4b/ecWcK+1gLs9jIvE5kCgppHkyBOBf+V3bfBngPj0f5
ZBBP58zTCfupflRT1qZt5bcJEIO68rvujZd0dJosgoiAd9iVRBCYgfS1G31ChBo3
7VfLLH17zV4D/DTOcwcita8goIy3smXMLnDL9B4lWHyO0DQJjAjn+g/M3ZAcoWZ0
mo44TjvJCjnr6mdIhfJPjOS07iRKbZsPinDqM/5B94c5GfIct3bwcpvhQqPaKdmC
VRaATwnCVfkz7T+obhZh+Hnl+LioBAJUx0GqxJ4EILtmOXp7l4TjhTEjCpL9mS7l
M7OD0+oDd/zw5lxMXvGRgJYVSy9FGmdtFN5krm5QLjn/M+LEbplJWLvnX1wbjdw3
WDifqjr2kXYXINbwfCezN6TnoSbP7ugMwMUUybvcDUDxgb78fTLraB8EoeQWyuxv
BaecLrSUEMRFYiNxqkwsCRyV3tocHYYqaNdwwFwsD3rh6p3An9KW9SSnP274QuoN
7FN3wj7GAkh3reVDfwbgsuJ2tfZ4Yr7OQ/hkH0EsBTue9SZeTOf6hSr3ON4emqmu
Tupuhq7j6dbod3WuVxFrdbm/abaY+rowoB1tBao5FID/hpSQxw9MsVcOq6l4zIAc
7t5e/yRApOlChwxeoQ4C/FglWrV2YywgtJa9xbjTb9WtfcyFm4IX/hjMSzJNbV0J
WSa9bkDWQHtVotxbC6FHJv8N5o+R/krDSdcu3q9hROqQ8TPH3qkB8RKzWKCKzNkh
joRRXnr93OIy/3kCeAz+k8pPhKBMNA563Ha/QnBPu9rWHYs3TxjPvxqiUeUduPdU
y42S9AQhIrNL0mHbTRnEQ0z4iLNAN39HRb/e8yDdpzUn1ZifU4ox72E6qoNtecB4
KISZDUwW2k1OkSYpSnoNtBM5bUNZZsH6wcx22T5+/8rR+PQ0Mq96UnNoUqpOVpsi
aiOqHeAGe2o3UUoF1ub4/L2SF0LRE25O+Y3W0gwI05ZF531zkhtd3Fg/L8hloqQd
bAZMISut3JI1LHhuRBfesvn03+EBv6FuHSoVhyoPuxPPS7/+qzCh9nxwuS1KTQL+
89mVr9ZG7M6+W5ox9yYpPYc3DF0hgm/acMs2ziEPQUa+k4z588HDLQPCktqlC0vg
VLAL8REqUKYindUy8rC2sLauRImcIHlSU9VsCEpjviQb1SywWBHQV2F/PHMpiUGS
pHdNmcBnZE8SFH+sfn7p2SJssHHBgjeoZVeVAi3FD2ZowyL2uPvaqqqC2tOuL9SD
96Tqls97z24Eh+gNZGygFST6pi3GsKV5+BXaEZoq859YNoZlOGqpIjlWqqTJcOoQ
m4nRnQl39MYfJJDKPHbDZ9IzE3OykpH8UmErRmE6SC2hgO5i0zq6a33+qmYygXql
wYV0EbIBm9eki927Srt3nhtJE9lYM/KZyST6R6OiwROGmApbL6f1WCVbI16tPMUf
NywWgjTjp2cHVEuB2g1ttDlpRaUkVVn4dfMLzxMhSSNzJuooyf91zhaVm4pJgxaM
uM/DRhXsqDLKACO+FulrHYeq4dnJ/ZJp9Oo3toXILqrNcf4uHUJMpgdemr2RRdJX
moU3I3V0w/s77CSyeXstdv6MBoDrIUoeNePrkUZSoj1Swvt0o1Y3P5UjXjxPyHUk
p2FrFLUVMYSQIgKwFGAIrbNAiTKRevc+R/WTsx1dh+S1XDw3dsleVHJr8gk0v81c
Sy2lQV6hvxuy4UKO0do3u+/Eub3ruNml4pyVOsbzraeUqunuYmug3sxQTXgFiDms
JCD6q37qhEV2ovT/W157noL8Nqxd/tQkA+KkxgwJTPHokU1LrC8KgLvpX0slxFeF
7woso9RnBGQUSObyGkvVVEL4nlefW9deahrd7nzmcX7idSTu+z9m5jpBzEjNl8hF
SUB0JDmPMo6sgi6nGAULdL2p6w5f7LLZLltYscxiabXR9CVBeO6UCer/6jc+AG3V
Dc54rw/wiryFYWE3ijM870Zv9q0peXCS84C4fWbbiq5DoV2u5J6S+EvBvh6pzECT
Zq9niGT5rAzZ4CbtL8FGsRuPGbRzaGx0EPtHSzAkm2ePl+dTWKppJ9e8JK3KNdCA
y23IMVkFnFmqSgU53k+jSK+Y/f9GQCpRwDcVdgDvLpobekB7Psl3uxLfu8b8pAOK
Vqz5ZO7oRbD4KEiq7As9olEQdpYTh2CN0CY10wEqEUCLlzJJnIUeS403acH/7gk+
1iaROktYsOsifkkiOhdAAdyP6foQtw24OHs29WgtrN2qeeGifFzuebqe2eVHlDVD
7e1hzRioY5k25sRMMJ0VNkAZSvTvonSJOcCM4axNi/8YIGxGklAVbzpHgiUFgEss
+skF8FYVmJf6nqPaBDJyNBLKFIn9wD8JjdYtm7SJ3QMOpGIRX8GLgHnEftfe7vJt
dmwxq1EeouRVL+mH95A3LyeROJFKIPDNqKuF3ideEMSspghSq7ym7MZhBETaALPn
rcsi6SXPU4zc7RuW0AvADjU9Ccy2VIH3ZU1BcrJ/lJzybkLOWmW4WjZzI8RppAZ1
iOh0Dqv7P0H+in5ziN3QXpXPOd0I8Iuq2P0nHzhGxdMDPfTnNXEO579kOevQbKfN
y+igCOF+/84fzj++A+vRb+Nc42NXysCKKT6Pshyv0GngR4EOLnQ70ZEQIQmz3icR
P0Z3rU9QHk0VhIEaIyROc9nCfsGULXpcafwm8HBhUkoFUMmqaFB8vUnhFbrG4tdR
DdrwHw05Y0XxV3QOMJjnjT7RA0mJooorsxr4bp56Pwk2tSXAkEYQV3MbfQv0BnuP
Z1GVLLiKebg30RpAX6uZD76zFerO7RuuYaFIkSIYnTRHvvwCq/8HzEyiEaDzRdyU
qhCgQg7Hl5Aezwr36HjU1ly+djwkIsWjcCMy0x16JWJOs4bWvfeBl14ps7P25BRQ
BW2vVczoo3POKtWV7jHCcMlmOAztkLrnGaiGopYaE/EI0uoC7iVq1WlvZBgaDEKr
cXpmd6unkDOCZR/lWaJS2lnQhrXgOwir/htOoKgaxv1K8PtopoYvg7CJmZuyYG+X
qbAQ81FHO9tNXXlqRZuUbiQXY6YJQLcPx7HftxcKGwXQYVgl/SuSNC4ejDaHkFAl
Wd5ecG9w+4ijFW55Os8Mrb9b5jc9BQYMZA5JIqyqXlCiT8K38296gTmQ2YB19jhl
2OkzZ6Xilx+I39qH2WQUd2T3QbyjLmt4+jw5gFNN1fgTkTTvyxjShzuGNEJDIXyS
ikk84pEvsdnFfHj4HWnCZOxLkms/AMG//+bvmlmjWkRN/kxfoJxsfgb3Urd2+0FV
MByX2XTRsu3khzcsKUK2NAQor1dS7asCiXHI8F46bpo5aR7oBZ3H8/tTZbal29/I
t6vXH9dBZ4aj0f/xeUI65fxbWji23wV+m7FZ0iJZNcN3rqam52QFd6jUqziueFb8
X9GKh0IS3/qECyVINVYoHsScH/PYvHRNFZkdmCA9EoVNHimOiGjpNbIyUJwedYLC
PXS2ByYKVlUiqkPSgmQMVd89QPegiWBJVDMn2uth3Pr/a+q9Je1Er/ghT+bUeGNu
4+uP1PFd4/QVawDdbGLYpPQlVsNv0OqGXW9cTyM7jhVnerNRIcY2Y6fxgW2EGn0p
88BZR4TCQVplMWU1HQlANdWCKsIrt/o/Z9c7TztoCzkVw3B7gVzsDweIXdN9UT5/
qbkc35J13nuJK9IMhpGWNb3WyWtvna5uPxSWe0bytp9NGlXxNDQS3vYaPAtCQYLo
L0NLQd07ZxokoDGuYWNYvPGYpVWwI4MDqAKZi3VyETbuVRXOcpaOxN3ZTOL2EFPw
qTfi5bxADWt0yqRPPzWHUpbW2mT67jSfcv22x4EM0hRkBE2XrK2c722HesJXu9n+
cYN98YtoZsL5jVZzNlmFrp8XhcxWNeN6SDyCcXOmWC+UwxllPmosVJWev03HbN0Q
lFxYtPxDB70A4mFFF5sad0Y6K73y+Za+ZmJyDcvRdj45Q7yni6BLYpwWRIvSMSsR
jRTEfbQwPlgeshPYPWD7GSML34hi1wApqvT6qiavgWm3m+Kpy6HOtF3zp1qKGOev
ZoP4Ycbti0HE1GxKOzEzKMf5t4AiHrXmp/6o9dVC7WctaOqa+xdQGKnk4s6+PPrV
Qbtc9MQohXuISLswAjif95HkJ3Hnxezv6ibtlLlt4pXs7Hix6nobWeSGT4+8AYMe
h/bMKl5lETGu4EHjm8T4lAxqrDW4w3jI9hAwqVqJs5RPOE1AtQdKPldATkpOFRc1
cKiqmCkvNQheh9OztAnugS+wKD4KF06U9pR+XYIEtcdA6yhoS93JiL+eCrX3Yibk
vSFaClc919DZ93wWETBidbdvZCQWEDv8FO4o2MqpHVA7HpdmVCwOHPOnpSjhwJf7
tVAATUAd7YxYPwcPNzoqIlSU76USpEhwES7Npt+73FQqbdBr8gy1RExMGxxEPcER
UnnV6DnWLr19xu96og7rCBH91cRW+LDbfdPWKhzyPtEuKyyAie8B6eGm42eVp/dw
wAQImYtoS0xuozmF5DNqTBWJobvd9VPReWR+LD0I7iQXdeCLWFP61scvxcZjfGL8
llUdrGjIVRo3aThRy5Q9Dsmw7joDln7JVs6BtiFx9LignlyF1tR5EbkDHmWKVQ0G
R6fayV0K7XjBfHValWV38VEtwGJBAyghV9SkriTNbxFXJWwxmwoF1hrm+ErkYnWp
v6dGfCCU/UIg15TfUn+hBAPO/CHd862rV0j0ke7wmIs6XfUInrAmkSCE514cbcsf
9rmL6ZL6jjrdVAQxnem5qQQy7U55Sw/icvcX4lZ1A6wSWiW16Gbi6qRtTfu6v5pA
eODciaZXzduHxZ4by9nXkAVsfLGp3txEyJmAjNV/oeJ6ME+gwJ7xyDpRFxUz6/eU
JtSVbscr0YgdFqMJiimJpuvZv2IpkBDBMI1Rjj/AczJtrnjvYA+w9ajnDrzWYXF8
NvPI+pi/n1kWoh5Z1sqfcCfIMNfS7QJXrdR5PpHJMbD/kX+I5sZUnIGe9IHdlKrj
tOXsTv2f2OP+8z+WyOlhMy5Zcw8ohqfmPJzILT8hMhVVWYk9ADbvNMu7JpIpIBrn
UsqBWeXY0eHT2jDNAvhLQhv9TWfzMqT3Ea34RWLBDj4Ti/kO8jgv1D2/8lFqmoR1
wRcaO0WeI3R4MAjzKdVu42BwbVe64g6rKIiX4f48n6TJgeN+wafx9I4msXSYN35a
q9Z+UdFEjJIC3K5eYmCOhjH64OHZgxa6QJtv8aBYPHbHMoP3Hfy/+pA/i5/akZBF
avGVfx+wJdMaH6semkZMd2yQqYoZqNWSlgk9d9jH/NWwnj/1Zv/j//iq79ZI4N41
Nxp8nPH3rGg0d4j9E8MMfRGjpTH+Kb8WcTA3sReYRg/6z9RH96P0gtBj/Y68zOyE
++kwEcOvyykTi0r+l3Ri7I8DaYXctijRkjDHLM8wnQdI7dAaxFfyD93UMuucEm0Z
D5IMhKgTJGGPoRL7zeAV5W5VFQm+g8gOtXUMwTFEkPnkaZCTxxPDSCW5vZwEsWFq
2/HmpJ8Z00/LNY1axvIADhq2AP8A9OI+kLWgtGkPnRRJyq0v/29l5TBITrAaJ4fb
79m/WYylrxm0fcFsQ6XMwt8gIx5vohZbFOsMNXGunM1mXOluHsIVZhsNH5oOY/+z
XTEJbr7+IUD15Og4q1TLEbU+5l3Fj1aK1UP3Jd+eLvAhPXLRsujMbcUwBbgV2pit
TqR8KRrtF3K3a84sZ+gO1Lr/WyvUCRxQIV+/najUcM0N9SKb1nEEmUdCqf1QFgwr
VK9C3zh+UjRXLOP+B+X8cUp1imipux0g2PVeTl0ckA6W+rFIyuUbeIKKV5MYCZJR
fGq4dedjpGNnXVsGZKwU0zlDgdqSru8GMg7np64DgqD4Ox7S7jaLADvUrUYUAuaw
nfr+RE3U6Lj7zyJarjVraKcNez54ZxO2A9n5IIDvKMEwu25spsX9BYDqwwfBcfp/
ag1CKriPW1ju4aYP6cs173acSKyML2m7sBws+iuOal3I3Bchk2cqIq5L/YaCxbq3
LwHSnq9dyhGRdnt9uwI+WclIMA/rps1Z2VX/Xmbt0402itau/p8m401MZZDuYXvV
BafI4QeylTWCIaZHZUJGA12rGydOMiFYhBTsqvSA3/g46mGvI0+E+CR0mHhlAExy
FCOVqTRcMS9WheHwEQi6Bm1wmur61uEXlAs+3CWX4N/JdYbNBxHx9eFg2bTKAwac
xwkm2zL476unL1uUM08iXwFXDymPUVMnYQpwB1gy7X7P84i09XpU7MJUJRvl3/c6
ORv0FLvgGDkzZye0wdyEXkLpzwj4Efli1NphmEfrcDZVbwcrx3s5ES7f6845+4wo
b5+1RcCLIp5jKoqiHM+BH/a91ZIb9lQoOPIr2IVRFTy1F81AIhDRoEeobmKtbMpB
7MkXptTk/fEpl3EIMbJVwToI6VSUGf2JFwLTl2zdIG1nODwx9Oou01qdR4vvuOPt
HgGsIr9lmgLBKtRAy9JZdJHI8N2mMm6N4YWCWNTNN3GjBWbCKHaKI1FCicKlKfnU
SxsEa+Cy0sLQYGWHQ9sNaZcCGKcNpjEyrsMCePh/3AYJhgdwxBl37iyKcV8DH+WG
MGw1Rvt02ahHj+ZQD3hZANeUIcIgTGO5K2QercgqtjGSUivQZuxfn9JKp0T2vgiZ
300fgAu0ptee6xBFZEAZiz8Sh9iBTL+jI8pp0liSHGfa19cAeGLdi0EL8CEmdCZe
nNsCjyx6y1f2OFuU8Hf81u0/hsXmo/RobHy3VTYozjLnxh4l9MwFYQuGSjkFDxKZ
3rAiTxxlm/04rPfR+PoBJ4+bOWAdAMlgeq4M/taNYGJwFuH+byJdaW2jKXC7/02b
i20jKfVlS9bWFiGHAgAo82gftPZ9SXTGxIHNtHq/Qky05BPK4jrGT9uzMRDBNBGN
8yTkqdA/x/XkYJjXuLAY10i+o8akQ/y7jKIvPRCuFG2kgi206067qX5lScDUbpFt
iGfDzLo+JLvqmgGtaWPxzms04p6Q70L76LRWcW43BdgiGdv+Okgxe6MXvaNb/Tq8
3pMLG5sE3GHEUapoCpCXjFz9ED1RPEXof5deeHJCSwnvzZUA3PUhNZG5nPHfV8xH
cnOgYjBd7tMWNulZTrBYKpZZJ5BDi1+KlQjZ4IK2QpRIXk7enB3prVJfcj3f7Phq
k2fR47Uen45DboRsSudF1+6mldcnFP6yvVONziseQuskBKbyIxR/8AVklFtPmcB2
L8Botj3Y9ZSB0K36Yh6ss1s8N/MY3yiBagTYnhEiwTbURgGSmXeBsSWhNH9pEXZ/
U7LFCmKUdWD7cg5nFtejFFFbLfoZ/SLhxbsh4FtF1xUmEPSC09F2plalrv9GKM2S
32MHpj9bevcxK1tXCUUq+Zc8BFJn9E+iJtRdWTiVd8iXX2A3rwsNC5U2OoaYku1r
dAhwvpHYF2v1oxqUVGXl2sW8lBPM8KYKS0zLXoUAqlI/gU6XjF9WSckWC/Qi9Aw5
u46BdXANDfg9uxrRCZ1XGvufnGmhOibfNwJqc/frU94Hv2klNBvIOc/bErJnFd7D
x9q1wyBbe1io73tmIlCV9nZry6jXR8waN+Jsy9dFc9mIl9LoVOyHgesZvs3frHhg
yjDsQlfydXfTQhvdTo9FsSCbkuphcfKA0vyF5A4qNoEnZxYoU5peZn3GeuOECdGI
AcgY/iGWn7aJibXSgldf4VFmLmw3cErwJfDME0a9gY9swQ48oEgUjPZIRSclnRbZ
UyQh3VaFIo7PT7fbOGHQ3YBGCfQSIhYpC3xCELX8sl8SmNhme4VmG7DvfdCZr7nw
RMQbeQRf29Z1QGVwau93Xo8wUWKJRfV4XA9WYjTFf/fb8k1pYvAd1c0kWfqbTsYz
gHb9zvK0Cjo1nZEo7EpC9mB43C/6XNxmrWSDKBIAfeEbRAtXDm/POhBU4qlg/FtM
gLdc9j4WYpGN/zg6Vnhe+0vx0qOFIxJyv17unzZURNZRScw3B+D8ijhMO0WyGhlN
BRvMkpuUnIjGzVH7+hDQWuVNTaoFq/m88a43VVPMMkThg5svPRLRVIg5hRIGhMQ+
0EgM7kYNsPnrCdJRTK+8yFWdiwsnMJgQjBIsxmdr1g6QPSiipcOgHlM9GyqDuhb/
11Lp9eW2VXzK1pwkGlXKml5qceF36jjOEKV7ItbacAI5CW3Jmj/9Y7RAfrD3iKI5
yzOqWsVtckgNFi3MUzNaGVbKU7Hn80Gnxf7CUtoOCATFjYV20wnqiD0m+Fb2GvRu
1aTmgGS5cMdo3ws2A6RdKF3bycTiX5hIL2PcegpngYuwpYLnFxe27HvlAYLzsjBP
PXvMhKWyZ9Nfo/543yRSiP//kg2G5TsCmDtSfaZ/wCDNJRscWGI7dzcDrx+ty1Tn
KIaC3W4DaFv35NVUOXRiJi82P6lfYH4y9QSn2d2hPtb/qBwFIgt5Ic5gNfDAP0TW
skwy04+HHjTYIWpk1rOD8RCB9kbRDjJK9Gglj8sDSsGC0KZiEPVKVe62/6QUnece
3585IyfDtE6BDXdZKU5F397XaiBuigs5AhHydc8GIFBLbO7RvlJyPcVD63zZAwMR
vVbtuEJmr8GFnt3DZe+CTk6lKdqqHe2lEaUdadZROzluPE502fHoQSezoiBmFVys
CumF2StSCD1O6fj7dhoYLjSSJXq4X1Wy+KqHr5aHVkAnoWoJdl1w223cXBQhUZpJ
tbooBwO/WZWR1fbbbBqX9ocgnuxcoBM+0rzVoFMigFvgsm95xUFs3fqEkArW2dxN
R+eqllXNIINVMZQfdXzzy9vVa+SqAPGz0Gm48/HzgtI3JHG1mKFrKPtakEggh9NW
97q4GycDQtkT0ySLtOTLYTasN16PHIYewCAq2lQ+3uDCnoYdMicmiSAYuJWD+gQ4
+YuafDbcC753Qml4FHUcY8QFFjig8zZNpZjRDPbJqoCaDPLEADkOsexjopXCfmdC
UbWdKGy3HYBpMiRknnn2G8eXQ9ycKATG5fBnukrqUrt2cUfG6J+F+Wi1qr8Uk+G6
h17UFjOHUX73KCaimzbdqLpjJmRSFUBuFxOHUs02dS9GosQQoXKVoTczbcMtO1fN
ieSaYVh3BbiED/t0jOh7JD9Hzteu4O4fIeKXwsRBH6X7Cd0mg7dgoRxo+3mfug5A
ekGo47MoRSKMJRUwcpuG1zzb+NmQx/pvkhVL+ZZUYZr3xlEPc+EQHfquso25klt6
IiPMBsvM4JihAOnKMykoZ6IEwTMru2HyW8mqiC2Tmte6k1r2pb26AXAPlqsFrTKp
hAp5QPqMC5UGLFaf9z6AF82Q7loTSofOTh7tT0a4cqXl7XITMv2biUSWx/4OMWwq
0t2fzOVQdjob6Rd7INycXJI97e6viWGJxpdyNKdcZDR/HfOHAQvuWfmyDqQpw9GK
OslWsKFVj3nq+euO9BJ1FeCVyFQPiKvqt+l2bk/17DhY14LR/3Kgp19UtO5+kWZ1
DBa0H2Q1V4oDgr+wScdZSKswdPaUprLfPxse+cxrRKPgZHUxEmZDuujFanBNI00b
SZMfP5TjoUxHoIV+YDPYx0yE5w8P79jwxnBm9c+5TD6anYDUfkK/hYUfGXpuzI/0
AwzK2SRnbN/GV1c9PLycjUr5FA3EVQK0gRR0PLjl0RlfLzd1vI6TFOefE4JXYwXX
M3ZJU/8NCtuQqd1R3V92Q57hjizS2cIrH5y8M05C/4VvkOwvunfqYjzS7gIXYEqY
ruLSak496sr/uQ3YfvybQKxLUxMzSGwqlOZte+dP7pIUxCrEuKeFTHsnP83DYaLa
g/tpctHFSgmTIQ4+OqmNBvmkHkLI1T62KReEoBPAKNH6ffRs4P9QV/tW6fslWeZU
zug7bseqdPzdTwCa5/oIuYAw2VXz2aMAOR+z8VzUKtI3YyIQmEh9LXruFn31JoXt
GMunZj/LtSZMtixR77KHEaTMFX+FofgJUjkOua+WmHhvKGVEZXKZKVSW1DhH7UwZ
KTE8tM7Vwha11NTPwGxrWxvN8YKe7YJs2JytiMrZ5P38Vi6cC1qFncv5NPLO8bVJ
qqAaTceESqqFKPS3V+ldNYwVDkAdF/Fhg85SWyk/XBfq0M9g99Ppv9bnLzK6lIj6
h479XaO6l79iTCnAv1flwF7BNnS/HkuUKvjdH/OKnvr85nzoDjSNUZQnUoj+rCeO
HJEV+JdakINdYgpEJF2kmsBOzFVQN/TZ+H+Qrh9jGkHiaXbWSj3z9FK/XtCAZrSR
/9QYyMGNKRIwzb4nctRRX2pwxKEZxPmtJobvdOM7fa+SObdW6shgJXEg5nhdybvT
N1mP/L7WJnbx+gHfuKKGvdBiMDr041j1CPme0lP0a3/eZyBuwjtyqe+5MACuZef7
g+nQAvNbUinGlwlnjheZs1zs8a/DefwffBZ5mRtW8ccD1LA+YUJCHCHLUFptMFUA
OjW0UvoIEwovEEfjm5FnRCFBxcQvLXJ0R2M5wqdfudKO4AUM0DfoF/FG+qaWljAR
V/DLZBVErF71R3/dPMKVWpxpikNWWmo7igipWsDYM5+FSI6SupYNVflPEYpEbn9G
68ZOd/ROOLSIBMly1/TpZC7F9zoHdF8w1eOid8jT0arWB76rWdhhJTJKjRbEkiBf
Ra8YTPlDaj1cMlAsIRS6gjkB1j+DtwcaPMbZgF0jFjfJhOPJRyHsioHRtxrnpQOD
tGMaqgrPDw7NspcKEXvonfiM+1utZ4j4kuylrqPxWazshdXARrJb6z93N1Koh1tt
Ep1S+6SM54Eh3Os59u0tu3QziQe//KuF1VLRu34YaNxiicS8BqtQQVN/FUko7Fsx
0vktGnot3ji7TjrgfrowPTAwgAaBhx/iCn3Am1hqnCppiE43ERMFU17tDLd2da1g
XHN5mFDpKeWUlRma20TPB3IbymDgWY/pCk3RoWUdR8gzlmCudyxAE41N9a+q3MNp
JgsM1ls0eYjBhm7A4n0rj5fHXxHvd+Wbb9Za07qxexZW7UZpz5fpyVHMSHB8vNMV
N4f01gwrUUmHnWifO+VyD3XUiQAY7Js3t4hFuObsb7ETTgp1FXQbsb//r7GfEEmt
4d2IQT1R5zI1PIu/lmBLhzIaoxfFMTcHwUl86es5y94UyDTNKEu3owcrEQ68YRFW
iYOgikKf8YHRDXSbl+6Q9AIU7VOs/s1dKRnq+ioXhp9u+AjGwIwYrRXQ/0IlzTpl
06A7FRRkY7RX2uk21BKgdW1oVWIwHi5wNLnaDAXYqKlmDs366PF1c3dfmgGq9z98
e6B5fxhWvap4N40+yytMvUV2SigDlfZf3KpAvTsBx6eGUV4TXCrXHGs+MNVLWnNN
f7nDRjamoFG6LuBuwkHUQU2eqB+gL5idrNS7M9noNCOHclifR/X1AMBCI0cq4Tn5
Rcyi9nyCXWyIEwGd2iQsO+Wx7a6PR8CLpm4oW3C3kpaG0qr5fgdnzu24bWB6M9vg
XAilRWsHBPcdiVIP1AZ1og3JgVqujBfM8BfyK16kNJN4Dj2jIkylg7km7nqzO/gF
p0hrA5pL6+qZmG+pmxasLfzf5CSS3ae4cz2AUYxhmFc2xFgeq/XvtkUSKTg+Nomr
lp5iwuIot8vc1h6yDhlZFMo6yxRbfRaTbMVpGvI6a0uhHrgKyfZj7AOFvqjyCqks
jt7FScofJTvk0k3oNPr2XuILgTlLz/3EkHbGB2vevmlnu+0/b4/y9Xda1tyhghCM
To9mS4xnKksrrSWErzSSVT92eUtIlUxqhGjcpB97kRGm17dCI0g7GunODOOSSJqh
UoxbC3YNDMBuFS7qgGN1RocIkVmoLRE3wlRjYCd3zRj6n+YzFYSzzQox81/UkELs
/aZJ2he6b9JDnUkYAGTgzOMCNrpFsPvl+L53/WS+MxnOw5lSpiwUPQFQPknLLlqU
2R0Xc/HfPXgyNoTYxVqvoITrri4V9IojL2HpHh+fAAc6N7aOjOivSz8ZlffGWNta
kO3W/YrqJGH5NrVgcKPK2/q5pmO+vG0dwB6Nx8uuMcJOSIXqx2xNJi3+aC/TuNN5
iiS8xvU4k9LIwoN9oH1V8CZmkKzj1R6RvEjhO6De9VkitPmcr4tiOyLutVJQxzI4
HuUgUPdWNXPc7TQHHkgtzver5GmqD54z2QvCykHMcTIHY2uo+zD0QD36R9GmTl9G
Zo66WBkIuqkYO7xAFFK2IxHrAvvmrRRoYuk6uwI0uF00vnVJQwP3OrVsRQqENiJu
UkQLQwNhFhaObP0JvrwwZBd8j/u3AD2s4urbkAR9bWJoHgRKN+u/uzZua3Wc2Bc7
0YM3Apfwfj1cJ6qLV/d6ThGjAijaKmoqhCU8VcYV+WTDtpwF0H/Qb8MMPL0qFAOD
9CkkHnzcHdoyyaz4AISAZITSdxny2XLGpDPBBDztK3anEkFt16XPTxzeNJzqkE6s
QRo2HOt8lskcJf5P9i8Z7v7vJo4yLNK4AQCB+i9TEfHWN0n7uqjDmyqXFXNPltAl
lgbkeve/4f9sNYjKc7FFq9zFu9JDrdy+rYu8CD5vzVvqY5lb9e/ypT/rLnt8JLi6
i/Fs8Gziq4xF/jtAAfNcjAN46KaFxXxbIL9c9PNnHEWkL7y9CBZxZ1m+7U4XP00X
Jp9HVeKxZ7E/75AGpEF8UGcT+YTmiYPqja4HrfmRrH3G2CMB0sig++ObOHjKLahy
YuK+TKqCH4hmebBNooup2jTLo0HPK6f9Db9EVg4cwzm9C/UHE1BqBOj22IpX59rl
tasX1uMLmpvhdp920sNSWUu1II0B1biJpq41TP3Z9ItRVmxvY/QwMc/Hr9xuLCuq
0i8j1WNZNqlfni3Q2OvepOlF45NXs+l4hYOpRuA0cjlUwPDc0sELJc23u9XJKVxL
mGxSsK3HFpZvM7NdrEBoovtNPR6+khPv//U5pXt8y5fuUMfhEz0EVDsPvU+CfpAu
Ovo2bdul91Ui422uBJmZ9veUfOtjJMPJGwlkZXnCyPC7BDu8Kay4qfsQ+olVTG3B
kwipim2XDgXGHowz8ortmCbz7EuAmPHl1uBBzljwnkpQLMRg/aqkN0yS0gmV30WD
ZHg0hOF3uGeU4dSZFARqct4qoSMQ/4Kdg3VjbkcSt1hJHxFGS7nouIC/9NbO6qvv
OHqWZj2BjrLNVyBE6cCQuglgkB6Hd2WL2af2srsw8gvNdrk5iNlF3YvZ2VP7RcPk
nsiICoD0zqKQpwy9vRTUP6GOrMlvNjfKt5Kz3B1rYtga3/Xviic6VEWThWEuxSBA
YRNP3saD5QRwjBaD1dtrIJ/ZnXYiz/tNRPe9HZNvjT0NNGDOPUf6fOivuGho1V56
rJovE0NXmTDZrRla2vZZR3d43rwpoX143/CneHQgp79vuE4if9qXlD7HC2uFii1a
ZVD5K6XY/kBSCwFcMvNSFoQggsScThadertjONhiYyxtBia7beXGlyw5Trlg0ggD
LRWUPR0h3jyPoHKVVVsH5Fg0XCSZ3OjU98hwi3ptHP9M78q9GyDJ3c+awxlYOdqm
m4f7bQU3ZeCmj/eMVMlwRjVwXxetlyNJvhU/LyAmLDCZTP/cOAsE2yjyG4JY0dBU
Qo/F90smbhm175i555LjUx9VYmCM3uCWmUa6i1L7nA0fsrrq6WxCrDy5jns9R4Tm
JO+O2Q5uaJ+JRAMEcbCZ2Bf16iudqJ6J9I0ycarD3gbCcX+PUOOU06O2SMynxYN7
vQgnh5ZhW2SypU1FVLViNtmgtdgtzVwlAZnoy42Os+or7p/C129ITnPg+MzxUbJ8
cGrxIvt4evgoN7+VBzwG0KKwSOKZgnzjM1NPql2g4dS+IM/9TYkrH7Vt/VtU9lCx
l/uTySp/t/QotPLGZaCuVPoaD55v0b34/75ykB24zBLbB4Cp4vul3h6HUgSnpKxq
19i7M5L6I2i8z8F4dCp7aJKNMN0cbEcDdWcPBn2BfCMfTnbEvom1hh9psk6CGVFL
ACgWmXDN7D043lgpIcP3siGXUN523RctCl0dEIfsVm5DJ6iK6A6ecmDSou2xEkJ6
SCdG2tRdjfQXVOT7uAupJ1ea2GGeNegpNVnYxryKL8VDQRRnTJx7txsyE2AD7S/f
1B3xcbr9VuulmUrrLpzu86yAUUIE0G21YHJJRY6EoNQIaYLxzNaOI20/uggPWHID
28rZKvYs6IzixhGF5OVENNveZO9OnY2zY6Paw+SVmxSpgQTVeLdMhEcJ5vJXAGIt
bHSKhSLBJSFTrQHGrWlf9gASzKtuDlj7/hPi0MaWFVcpYT+qMQ5BIlrWLTvS94SV
QCDNePiZ5+bPYvNPWG9vDZZu/o1gMkMJeLnXqW9Lw6Ff3lFLuzoLTO7QYcrAZViF
JJwuN5Bzlc/SbRU58FCRDoMbGMM4VlXveid9PfQ16Rrw8Jbsh3WCnAqV9yqSB/EG
P9yUBkj83XTd+Y012TBn5Okzh37UcWW/mWarWGTTZHSuoyFnDnIWkV3v9y8Z1H7J
ptFAtlzRYGwVp1C4L24al+5uapYl9HVNlwRmH0XTUBHBUCdkne1QrQZX5Q7nQ8Or
qgXll8p2b5K6uSKD2Nb1fTKZc/DRXhmw5lctOYDKULH7ksPSoxnq1h+g3E+7JW+F
/nGiSjVVoK+VE5YS48InJ7yTQka8LGQuVnY+EDaxVA4tBQ+JgkV+ueAvlxfvWYiU
8fod0vH23cjbEhkWth2enTY8RDtMXhHGiDbdI5ruZf7kG2RMwEBy3aVcrN+ejXme
zvh6rIFgC0hDsr7p6NDq8lJX6PYlH/5ffW73Hf/npg9TbvYbyqhawCyXK99Uo5oX
2HgLivySXf6jYIdaeoekDwvtTKtDpzincnVuJ88qmqCVG7L3S2iVPV7Ojsp99o2D
gFXhX1ZocXtN6Uke/o4AyIlmTfTGRdOmqrG3BCBFfMqQw1xKkBHx3xP+lM8uYDmS
MrEk2kjVYlGpt4QusR1oMArg4tMMOqAh3ACPvJBM6Ylgd2uJyrF2magPBmDEoAGJ
+sPeQPJ4D9v5bWKcwoympNcS0JkR76CkdqATcqcyTpdjdb15d/62CnhXMugkYxwq
0vB1zshM8E9IcqXpXRsTs8fG2dLUynjmdlLS/Xh1XTVmLbUJi3dpx4LO528Zw15I
qF7FdKPBwOXXT16n8hwShIQn7qLK+3zpr+365q5kBy8UBYhVATq5h/5Cbb7m7DCk
i/lzezluzLPMUD64aeFMTAx4TcFFtnAlu6Ee6IAGmTbPldnhYU+JBkYmS1qDIliK
uDyFvFNy1IwdwjVqVEEYiqwMDdVWYbEcU20z2wvnco076x1uoUPPkvuEX2OnihKS
iDvO5GUyeYXysD00EBS21P+IWkOfT42lafFyhSkSXAvAJs6XWVGuH2EkGB7CApo0
8/qo4RFnO+fdBFhOp4Ee99jI0/BayDnFZL1yQ/pMwhSJMOA//0LaoMLs7eNVMro9
nsS4pLNsJ3vjU59qGCzUChPAK/7VPobVdze9XtlV7qRZtzGViTmd7RNthPIfLGum
D7HEMBhWIidc5d9RwkrIaD2hBs375jYD5F1rL7vUrxHHLM/MFNICfiYtY+sevgw0
EAxwxz3WcBREo/HqAyl3+SZRpEM0XklxzBUavQ+ASuRqQPYN9XegtRpspsuxcojI
2lIneYYonwe1/+EzreuPcCOGHf9ZnxVSJvHUZirmuuJ7p3opYmSIHqpUYsZdhXiv
HWdXfkDqMgXzRHf2BiBX0qkwDrGShZ4ssVyOErxDH9wLNIkGv0K0VZJ+DvLz1F+6
auOKgmouF4mZy4S8WhGrOIRS8tBkc9sfZ/peiplzkNCill+/LlTH3UllZffuVTDh
xcViFu3o0jmZyo1m5tBJrccd647Rf8706Y8rRzcKBl6RGbPW7WYyRBYSrtQlq0u+
a24EsATRelLTRkFHdHPGRgMn3dCzY46VvPExSJjwtyquIOlwnkOBGHWCkeGelTNd
26uLzORhADoR/E9CixRGQUzr3HwT/64B2qJkhhH0pIDoLjceMtaLZy0bIcs4bD9L
9oA8++RqLpp47UnqJCyUU8LdDMV7fvS0dhcgz44ANXgKIm25tuJ8XGOdbfs5qgQ8
Pi0YvygwnOK43JO9EVJ9s2gL1i+1uQPGGGcl5pATboF2BRigIsnMz6M6Ob8P3v53
nkxIVvZrW2nQ89KA07+wLN5J22PYaOvbHBqS4ADvLXz1cnh96p87c4xVYp4hW2hh
Uw24qzjy+JedE2mW3mzzg536KEreOPlGnduL8yiWk7DMr0pM+09hcccq1OAJlgql
AYdkzhC4mXKEShbYuFE0XiX2NfxVyjnRweEdh2pCpqKdNU5oAgcrkvQkla4sclWW
MfnoXzT+fiAwmwngnRlX9Vb58iJbqUnltwxK3B6a7RGEJ7J7nkWCB0m8z9OG5DF+
MFnbBBc4wwNFlljlX3WL6QEO10PK0tEA+w7LZymhbybHSeFj2WtMoJsRe3Rqc5Uq
LOjkD+8/RjNxrPg4XK9UWVw+lMlhqmm5O8y4esk/yHROl4B44FGYFHQ7RqjqsoVl
oqaDLz0Z55YX3YYeTtRLjeTCbpqtjjdKSOx8l5eB310nIASO4aF/UUMBAzgHeRsv
tGkgXLMBbAIJB1liFuSNbiaIMeLC37uHec3ZVa6yqq+t8EMyTaRxKWXZJxZlSxJ7
vh2AsO/07B7qnhW7BJBnvIciADf6v3Nr9B2Tq+r9zHEYBgoUIf4ljTyWN2Ig7XiJ
gga1t5xnPC5sbVkyUPCXdHubTh9t0JYiVwEdQdARM7PnaSv2be5bGP4uoRDTKxaS
fGs2BpG/uIGUG5g3/ASiuSCVvYEkzbTNpuO4R1Gv3//TUay84z5aFQd7u0MxpVgO
RKcxPfXA+ULCmmmZ79A+4UYnobEi0i2AqAopy/2uRXnrHBQs/3ckrtHLLyuxh14V
FOrtZUTSwdgZ7m6g3rb64K4tBFQobO+OU16tmDWT1xoMRAqHi7V1oGSzTAGysFAF
p/wIGSWRD+Hg53hapIskv1oFYyc82uEbIaLC1U7xmKc2jFa0ZNguKRxbaxOlNu1g
c3IHfzFozXR0QYi07L4+iDLZuu/BfFCY5IO7K35c1sznCM8lsDwmS4/BzKpd8FCR
bpqJbV9RkcKFoiGfiiNLcthNc8N2vrREggRE8JIpbZyvBzx1SVVT2Bhp4zd47kl3
sIqxD5y3UNdbrS6AMinSI7IYzPRoLKkFXkcbB6+Q6Ntpipia4JjF8mCuSKcfyA6y
jLx8JuAOsR/GAYWdUCkY+M/0HOmk7LvdNN62uzoJLkpY6Ylb7blDhOje414Svdnu
kMKiOysRXNbu3DL3/oAXf+XyKmCU4surw3ILC+dgkcn5kkt30LqaMBVqOm/z8LIA
NomTdcrZfMSGDBykQUgqIlvpfzA1HlPEhjOC0aUnDJCBertaPJndgwBfBUXWCxM2
NQtKrypZqS2U0It6jm9liQOCHPhzVwa+/a96wiRY7KsxlNgTEGpJKbTaZbkkvxsQ
uC5gLI/UKstRAnmuW/jYc0e2rrXXxdV4UQoQq8eetvXAtJZgfbLv6b94R0/IiHkm
aI8VMLSMr1pb4qf8Ik7ejagRLor2BbPcOdiE2yomlg0hKrJW6NBLcr8Lo/8XCdut
PgRtQnPPh7dHvg+T4yTJY87XBj57wHjd16Rxsz08bus36f5PlvWXtxBBVaChrcMb
UGxx1vo234nNlGAxdV9ttSrzqpLJKMJUWPl3SbQoWKKjFYm4Z635SGSdnpI8WphN
XN+k40hYr4bs5d0F9MA1x13oDV3jYUKQIoIjiTHngX9V02m9PYMz3vPQ2Ve6rfhg
ZhEG/tJwiX+mG5qZfvkgrkybQzUO+D4RKAqTSYN8gMMtS5cQHZzor+z3Gc8NWWUG
5VYbh6zmM9sMRWebjLFvKq7hoR7r/pu9CSD+TNgIQC+VD1IzJ42PRNN8Nh85XbwQ
bIyfUB8YRMLLvET2NfFx1yvcXO6jAxe1/LsQUZ6A+72/2XE/R+7OT02Um+rGwFS0
RpGm2No1nmR89h/rFhjYBPXdpO0zTTbAXTdpYuCoyOYtQdSNEp4QRaNfBBSUo5GW
vGuDxJx4uM53SuI6cv9dwgdbwj2S6ihvnYBbmvSdIXxxPr6hCGomB7RQiu09aNc3
0eHAduTVKf7NWhANgn5v22MFJcxjszH0lrFI8xuW7vUTWK1eRcT/WPlUKMpLDBKG
huz4L5sJyiGR34k/WREBX8OnE8b87xspge2CAgJC6fYZ1m7zufpg8lrySPl9fYvA
xIflC3vUsYCm6lWWYNH6X4jrylZ7lzjNG/WTgLvUakxtf0nKmbkocWdvEl5q9B43
aNwHiCgifC6KrLQmWP9VD9hFPChe7cUlBO34O5v73/v9XPXWy/DGBaTbAhmJEKXs
1gom0pAiz+M32Sgd5nOcPuMpybktN/rSKSKWzCGjsgAKX+AAaUZFoGIVuaIdSBOF
YVHphKGVMI9Fyy5P3slZvsK4NEsriXF4gxBHIAUA3PNH1WE2xXTfW/k8Ho5YDClk
E66uXk+RuCIrQIpPEx/pTmNsXullmRlgwNQ5xif2PnIj+Wc5HmxgsF5/l0pahL15
Dk84g6XyjAu0tYO3j7NrpLi7PtyTHqVoMpmX+xZZ0xpahU1afdIDdnONPJmGF9em
xDjbUBIswuyldzWwzIaud2RiTnczbYD29BVqribL24U2tgsgQR5mhCh1l7iv1u7K
fXKQ/OUb1tDlfZmcgn/1TwIPRkX8MrqTlE9Jtfqs9TaIZtp5IXwplEkFiE67mrzC
IdOGJVXUAgqVhOMPuo06yEgEjLz+R/uLsiHWlCO8npacqPuRTrV0zpKHHXYq4Wli
VeG1L64pFU8EJMBAQeYb4XAUC+Nf8xxcm8S1rRc06tE+ha32S9MZolqDlsV4wVHL
43Ih3l8ch8H/O3QbBc/5/BYp/5Sy5bG5JSszi6EF371M6lC6RSlUbKyr7cSQ4p+r
RXZuswWsBCITg/z2af8ww3iC2sx0LRLN7ApxFaSDy2Er/owhY+pf/+SJf1dZqY4K
PSeanVJwFf8gFPXBmNlarmoCSI3sNyV/66QGyEoPddjdr2wznG2nwlBY6v+Q8HIr
GjU/iXRitxoPLStD0enPCUz4D2vCGHRKuaeosxpISdm9XGn0tgj+yVSpvzNnhC4w
JmOFhVun4rGxyJSo3Bd4Pt3adPLuKdoOGXc/gXFv9xPdaIQZrjBnIP7K99lHhli6
M08CAU9WuPUnIgMl5CbmqYmewem2EMixxo4H4w7K0jehARG61Vcz2LsraxO+iorD
Rw/0xQvlC6OOF+rHl8KxZGgA6c0SHLhKmxNIt9ifuygv+ZJlnaRnnbGXO/6zksqx
09raK19DfuED6R1Bd81/UgLz+eiYgG0sgNp80FHslUNJ/DzY8lF162gw+lZqZKUs
eXrJFFjvhyEvxcsYx2XZDGs90QjCE3r14L4ea7QW2HtQ0HiOqP+J++8u6RA0r3ip
alW/ZSLGAP0LSfhDudy0DbLWvHMgbQor7ZWrbK7WELL/hwnDu7C1KoZbh18/yLAO
1lj1f8hCHuv5Fo9z9lB33Syv6Nodu0XlgaBHB0wXJti5acQS7SQwhy/3imut/OGI
P/P7/UGWFllN9yMisvc7EAh8rOXFBjTjxjjTMmRC4HtWtnabSFxtRUgyhWBBdI38
Bq87HeT5YXyvtNC5Qei6N8Y528mzKlzVt3GmNKC7kQTdW9pBkqlagna9o0gnEPal
Dxc6ci2QS5EvPalSHs4fa8utJbA+neUsKIyfcDLQ6vDMhjTTjJUyNnn8LgZyK/pc
ScovdtoKkhwXbi1ca73Px4qcWa+VHWGYKkI0ogzyh4C3aU7e2lIdATcxjGSY4F+A
Z9n25fJVqnSVUdcmTfGYrpxi5nD8TJLhUqk4VBagr3RBHbJJi/MUHpBHRR99AZ14
QITncCbq69V6FgJl9ZnSPwnlt79Q9YxXWT80DolUdFEb5jqWpO5nIW95uC3tATJq
v9MudcFeVlDc9PKtCLltG4b41mQ2zZtrFRo1+OwVjfNzlLBuGj7SE/L90LQ/nqqJ
O84ET5pQJDcuD35kvs8EXixYZjqnXHjWbuX9HMELq0D8P8nbr5n347QUr9mirit5
8Ui8OpWb9zT4uaTKNXylvYJgoTfzSwH4gP5Jrgl8oWCWLdmOt6IfGfj0ZVbjOOpV
B6us8jqjFVD2Xp+GoHevXNQFDlRAAOp1vym3xRU8RvccDHI+JZBsLztt748A82aX
yqcYoFvzDyahMuLaBV+Ut6tznZcBb+iI0TlgWhMsbn2GBXVMyqa0HKbGOfmya6q+
k+CnphXv85+hbjDnDb7KT8WEGmt84xonZcSlIuuPa/3v4CvWPz7iVpZ7SvAGrOd+
qNhqszL68tbBdMbBZw+wqpfU+1AbteTsyjuIAFNNiJR4jRZO8I8Be89+7l2N2tT8
Fbyw5Mzd+vksO6H28c9BM6FBTC+zTuYfmfaNW1gaWQImBdV01ELEvGyT79eGHxBQ
AyNcSqsw/bwuba1covmqt1fGrUro/FZrGG9JTvc6IqQla7Jl8LZMqS1pOWd/mIyz
quzdKpI2WcluSAwJCtcnh5XzS6CTn6sMzwDheSX1Z2QhMzMrMp4srY6eF9cAAuKO
zT944UNU2s7XW42hv+edyYfX8kiDBIDUKZChl1kq+WB13y0jNxU0HDSdr1SmG02H
OHEwh1kGOD2+MYPsQuTygceP5R9xIWYig5xTQUNmRFo+rKuUvnj95Crh2rDruRRz
MKtdanBn5OGcOfQpnOQTQymtULXrZanK67l8SOKWr7yMIzeD01bcVP6pYNhkBty9
8pfh1pMBX3cqrzQX/0+OC7ZgBRHLI8ovgGbUPyfmssb0y8Ia6qWLNU08zybSm0hL
EOsxGD8rIj1uJAiQaX+CEb/+yTjkh3nFitNKqoOSru6xcwbjlz47OEZQnVGU3LdX
gA4bcJFVWaDgjGesF94iL637ywvD/3i9tJNkACH72kOlY8mKs2BxZYjGtpa48r69
T1Fsog/kiVkmBGNlQS7Kg4Oyj4wLPeDt/2ZXZrPab1rGdOJPhc3sK4s7nRuPKCT7
cORJNKsiHBeuk4PBPxDrljMvPQ3DpptTOVbMVv+ii9b96EoawibmdFJBNwDQlmDy
gV+/nO/FPjAUXQxmpPVmL6FYYlZgcm0mYb7IcVBfxZzIE4Z5iKBtT15NKGr64xa7
df82S8OX9bmMPtNhHpl4gbtsc+0vCn718yB8nEpr7n+WGn/qzYaXzsgKcM5o/bSB
1BcWI9crPW4FOmD8RAMuxgtznrv1JmPV9m1ZAHcZdo6JKuijUQEUIubpvJgLrRXS
OokjY3FU2ujaQ6iIyoZA3rBKJMoAQJfIueOK9Y6DmczTRvrtFBobpGN74biimVF5
FvRj71cKa76cgn+q8bMJiPcCNmTE00l92eTJZ4cWtVK1NoW16aBlQM0LgnNbR1Ko
G5LOgX1cb0dlVdrpOiH5f2UnSCA39C83RVWzat0vDTECg5Jmroui5QeQeVe18i6v
FPzd2COCRTe+3H4hbWFhiB5D11Bzhd86p7h8GCbGIc1rCnrpYXGMNmWy4cZHetET
XXYu2CasbBeZYWZjasns9rTdktFCKfc1XtCP5RIyPCdoK5RallKoBML6kYFPUQX6
S21wiHhhMNdjYSMQmD8CJSSoV6RYuHvJsCtmTmejie8CPnRUUuLMgSlDGBDgyB8G
HENZWY1xGqInc5lDXw09CQN/GBWWDqltqnfa85jug/zmVmVQdRjQ7oUSssjInT/g
0ReH78NCQhjtrZpToFOME/0+0LDLxkbB+w14ojhtRHdfd8knwGm4+BFjzxd4YFb0
eYJrVYXb4Kgrv/Aym2bNUApR2ajyNc7e9gE+n1xICdlHIC1VaCa7/M/o0m6CUl0w
wmINjgWL7b7LbdcUk/xQOp14UE9qdb5XutGT5JSOC0Ox8z/uqCkiEaTV0xRDZF6T
6YthRUaxc6ao6HxvCNQsxsrvEgTaApWWX9d6SnIAomTZGaWBAQVOLA0gK5M+5o+b
zLGt/ar7JqXlMsh/shzCse5hd4xhwijfMI5MoB5F6S7GIcG4UIeEpcP7VQzXs1OW
wQ2SWpvYTBjot/vmBku+2jKgDB7rJP6wJqoCTuM7jEBE4Y2/aw/ZtFcimn+WRnTK
HixFnRpXBJwwg0jTVMvhi1s7h2FRuAYX2SlRGZsBPADu+eXBAmd1x9OX2AGq0wmO
A6kQwyNxUgtlTe82l/Corckc4OL5j2KUkISbfYAF2+x22Ep2q2Zehe+cIauMib9p
Pp6KmZwAY9UT9UhIynXyz68+Db9TlsvxmRCNaD1tELTC7aO8vEDyaqDRHKHq9q6p
uiO/46L9ARKKHVXeoo//FHSL9ZGAiITUHYnP3/zn6AX1hHHHGzR4J97oW/G7eJeO
yKKYkp0KxiUOHkGQCGa8orwYbAzFP+6c6AUOD8zb7hRcJKw5uJOhxpfbJVxtPCxj
jw8rm766uEQFCesA4sxaUeMiPkS8TCKA0AlmhdRE4v/zNLtPmWWoh6BcualRtpDG
sYlSAbDFLkBjd4UZlJqEwQOlYBkwV+rKeTCxROSwo0qu1TqZnktAUH/3486k1Zt8
qy3/gnWpcQP8d4mJfSlGykkfIrZP/IzLFEiY72Q7CGIJhBN9PsHx+bN9WgTlAiwg
fRa/ShZxBC5bREfzJmatG9i8wqB5iUMLQc6U+IkhRLzPrLPX79nxCXcpsyicUdxE
g532KSfTp3PKNBJTcFIeuNEbMjBXcRUnkeRQWlrmMu+EIf4gO8PU3xvDkpVpRxDD
mle40+1yTlc15yu4biq5OlxlaJmLrtyCFW6YP6+9V0sMtI28Ir9wijs+Pl8ABeMY
vRBB/eZ8Qh3lreY5VcKDP3hfneSsaRuB6LKJTW2faOTHTG2hsRWixoICyFe/CGgt
D2d5vHG/W0gM4j+U3rPVhUQmMZG5zzOOZnIfMRvitnhzDDZ441rpJ58xMFKbeKVj
IbBv4EfBMXh8ccCtLv9mEymrNLu+EgM4vKG68GT5ipc7xxxqMbgugaxamIKi+Fcj
7P01Fhn6Pnsq+Nbrhkk1BMQe336vPnKgliQ/QK3cCBf3/cJdiA1M760TkdSS+W6R
ZmvtPn8JTdAzwY/kiLzz5X6ocsVPjBQuhsQzCSQMOZHZ8TBPZlkpwzPCPJRILFOC
SyzmeZf8AFo+oPmzvZI7hz8jGLtP8UY/Zj51tWbNH2nvV+P2mc+tTpb+N6tY5LTn
MJ7f3rlDkvIkiHWRcFRmvYTXXAoFsLpOhF6fspNmfzxQzJ8+6hk4+88Q8IpRbY7/
ejdomJV6YZpwXFFAJoQbIZ6mGx5hPlIjF7wYt9t0OxqP6HhEZAeOrLsW5dMHXU1B
8E1ay0KGUQbFAmrNxvCctinSiYfok2jELmWa/YECt1+MpUP2k7jpgfEwOxrJ9/gP
L43hTx6dtP5ViHFMtdUsQeASPLosJFaE1rT0WJ4R4/Sg8AJ0gJC/DDKsulOlu3ce
XACdfxxl0YlfYbnW8GTL6NiNnaLjrV6I4rihyRg28Pp5mWBpo6cJnmL8PudbBMoU
fd70KHGvDGFsr52T8V/rAyk7REhdoVhH/afM0qgXEMg0MFSS87vdi+LS//G6nP3m
VMQzQEtbOrtQ4oCVeDQi+WxvIg0JTOg1vIW/6J/YwkLhWE+2O1g9T/mmmluQgg2Y
d96LD5hewFGXaFzaiknVvOMawBCJ9xw1Qq4U7sYl/j81wTP6uiy/LwKLrOgNdXnO
FEEyeCAY5caInXSW4ruvXx3zbShxVtrd5XowWx2xJ3yAu75LBuwLHF+MIhKyDful
ewjSatimGYOH6FwF39hMpQhlsPrnfrYpKd3AizBEQ2ivbql1FsVITc1gSuzniZnw
hLU0s/FRJ0vxVFZCbNT1z0Qu1rZAT5SUmnIelhTdWtJVd61S3m+xGmUtDKJdsfU2
MpfMe1YWdKECs7ToRe7v7yFDtJMO/fHkjHu92RmlRHQ9yJVjGmvoEyfCtdzelBM5
6pT1SNIaTz+CXtCy2hLZX2dHqMJ7QVVI2/nl3EGb86a8h5XgBjfHgZMOxGUziefZ
cb9OfnaTOoIxJnjJUHGilv/i48M8HgYqfWxiCW9isO7/xpIDYTIZXuL687sUPIlS
XN1fbnM51U4lGU7+jS9kfmy9fzjwT9+ZoEdfd0NROplNAFCEBsKHF0gM7nCMV+IM
c0HoybU40pmIIqkWQds4sdWap8AcgvtL8qJygTqn6Y/+IYs4WPMtlEHfxZAq8YtE
CtecggR2gThot8LWATNqCBV37AJmi0h1fRTt7Yz5bcK8os2QmECymRfs8/D6NOPK
1thzC+6k44kez4KL8n7127yRTYypdbOP46rKE/ItNhlni3VskwYx0Wl1zTZYUuaS
II78xWguETQkXx1iN3FmamYGh5YsR0x1+N4KnaElmD1QkuEBpQ3C3ET+TB2aHyrp
UhJLJwKumLYs/QfnxNqfyIKLi83xDwbIEOV5CiY4jezqpyvwO1RUeqkIOkWRG4Xv
IArPwxVvPYeLAdekU7KQ9LCyyQGJ5ES/lSMP6VV6CEs3Aay2NA0A8a9tKCa8nmR2
oXK5wbY0u4ERpGdeczUF9VUtUUTpWYUNaIIlGO5r7AtbRTkli3LiEH4P88vJd7fi
a1bGwHfgqb2G9w5GYT2Uc3QpZrb2iiBRRGcxZrNOKH3wLRziapYMQaSnu+7JpUhz
rd39u+8AeHgLXytE1iOS0ZzpXJui28dvMmz0WsnXno7kARdMBaHtivux8Qvl6unU
Imow2GrrrDSLYDvZB8fAWa8P3sXChzOgRX/OIinc3lAxnhIU52g585nE9JcBWgl5
72bnXol5cDzdzxTSKml0tEHIW1sstSKd3rhNskG+PIO0BN0ZEreB2085RNl26WLn
jqFOSort0i2Rx0tqKnDAi6sc12ExLGkqokEd/veBcwPrmhnElj0KuVGTcypEwjVl
o3x0oOApHj3CTXTFn08LNCCuK+3Ovm/kaDIK0gUAc16H2s1ZFrGvkPt4Ni+P7S+H
Wze4ds0zL3k9mT6rTH9g5Cron0/PgvEbTV4Im4lbylfDzPsd4RUI0kuwRNmmjL+G
PDNlcCTU7DSXxmgjg0EaTSRC+4w7KuYlG2iIxby4FNKBczLNERewGbcFgWlByTNn
2mY6syEo13iT3qvbqFByKqxr8drecVsKe9i2dLUBxfTigGqRmqoeBvN1bI5WjVEN
x6I8qCYRjnE2P1Liu1SlPSqogIgKy3O+ryKEO82zzWRupw0m3Ibw4yKSps/SEE5R
QTJCHXw/E3he7qXRO4joGHOeNQIFF4qRTAiDn9xGaLbXK96TALMXf/W+spcl5bzo
tZLmd6aLhgL0CPCN3huGh8Rdp/YLM9pPla/3qAANGbuXvsfIR0ZGSoqTxHBnrxSd
RE7WUr6Upp49u8pi4p/9bkIg05DC05DrJPdmHALVYk8n/X92WJs6d36zG34K0qSL
lAUHpCTCkdKorTx+tqWot6OHMrymBhISVmUAPVLsARcCQzPnTj2vEVMwM2VLuEvC
69UyAOQs/ngQZpCuGhh7p8go6K57ADFqfusi9wvjuMncZlMdhh9qJxefDW0rFM68
VdVWvXHCdNhRA76cBPHh+oG88XoQFfExnOT0s7Mbjj9Cg79B4fGgwVGC55RTMD43
xwScGQHvdylu1TU9OaU8mKJXeICFIJGxfv64iFBxmWtpLxnUUM/QiwoPhqWcORfK
kEawrnFmz2KkQ2aHQoYMJNsNtZ35sGsxC/ESF4Q4AB3YlvBUCdFD7ji9pFoLWvTU
yOCHxH09PHp2MWuGf5AWX5nGsISSHdWyh7GUqo0SfpXEE6W3x68x7AL5pmeyff7W
7/reJnvDztU01VQkF/ikxzleWdDCt7VA41hjonX63lJ/HaaHYVrevB8ruyzNMLF1
C1crmdBrkBE71YN/pSX0whEEgxbzNy0HRm6MUMAzIbRXVCO6+C01IXUZWkksfqzY
jWAgLz6aKZ76WlTCHYwDj+1Kt4s+KM2WYLCdb5oM/RX6Xx/YpdkJGNi6LzxXLreQ
JkJeb0JTTQdaaR1ir12svtJYl7ik17fl+0XFvG6MRSG0l/xyOmWFhHdhGEObjnI2
rRYDlB6uHn0lfZ+AyeYn3ohT5TCBFNTwFVnC1vWbuciHtXWWIw1EH9QNPuyQQsfI
5jpTEKZNvn7qcyONVskvROHFYPCe5nt0j89VFyZu6vkCpj0GbhZmuu7S7GebRtJj
sIAdxCPUbf3R1CwV47i+bOxvoDzlu4H0rU+w0wV5i3zE8d3w6VkQHPQQGls5UDcO
zrWFmSD35fB2mBcjB0opMgy1c2zz0xQ3zDAtE5qA3mDe3+4SHeWA/8qTfMMS1iUM
iGGa2BSFjSYa52BVDoc8L94DX8shYh7gQTxbGapUjGHnRz27v883BEoZJzoGZWXR
eeJZ6quOt41EGh881zE1wz/Krqta1zXU7lEn1mB1K3h18xgFL97b43WoAlj2aoK1
7Px1ZQ6l52Fjv/gDpXlIM1OQXQOE/OvFhWrSSIpl1/oKiBk4QsgTkLs/FZl1tEO8
HjvJainRomhk5UVSdvEvOCSd8PynPlH+XMMMMZi4frvWlEzqGkqw0T7L4HsTUNHa
KHXVCzqNGLSd0hm7O+bfDg3z9GoGLo6oFox/TEkvF/KCtmrIHq45jxJZAzwA9EGO
Yrh39uF/5FHJRWEf5XARCQ/Njwv82NuIayTWJ49YyTB5fxytKhQ2auFyyQR7IJa3
BEWE466GMT4fZ4sycOThH4A81Empybv5tn1cJhyelPtQQtNqXpp786MPEijKU85c
DZM0ar3WcxIYxs5w5XPMHK2QzD+jBQQ6ZKb3FqjzjdYv3t1You2Ajqa7cqkiB116
MPDQAb6MJ8ltchpaoKZhs+xbeFK52d3uj8szsiwUltng4vjR1H/z3R6JedNXh3nO
q+zw+/N31kGqGwKcZdd9znwmacE7+Lw0loG5chxvHnKSLqnluyfs9fLur2vcU7m+
x0omqFDZh9/bY7Hrbenv3bu0DHtG6zMoxbLdcUAAZYf0eFtBbmejjGlhI+ofmlcU
tdoeqSMKFxjwzq14r9LJIr4FxEhxGPprhplcI4ms1xHy5KleTFLt9R2grkPXq7bd
O5176kMpOdQ8eVMyexqKWBydZsQa9BQoWPDG68hW0LwkIiQrOLw6KZNLQDtZH1Kj
1rwvwZs3AoqxeDmDoDWxEtgLIn10DvCHim0iSCVcbxwAR2ut8zpqvxnf6Bq9Z1De
I19WCpaZWkIHU0L8AIxV2My6Y+Och4T70s03PL/NkPEFP0dSWIA1t+6W6+C1wL2e
t2b47HoVcPUq9j+Q32jdU+qohM399iPzekSJexy2+hlutOB9LRyaglhWVo7Hq/v3
ELhFUxAtpel+nztKxWwUfAp30PaOd4QshDmqCfKWPcJWqoe9+DGHKHYjJQGtEtXX
HX1DRhxmXOUK1HoQOvieSM0QL193YDNWI8sqkEHqrj+cA3FUzzSvsPGDVWdsnVf+
6M/nrUqdi6WrSUAeI6Oqa8s1YxLNrGZYWF3xKgPfVFGarUloodyeULpNr/Sih4gg
xA+nKcAWb33+UBkW9LFsNCmn4pXEls9DIbAcVd58RaJHsq7iduWyNkZWNfgw8KQf
e9g2Pdsmw9QReoJCfzCrGj/s+qTUZJp8Sw7NLIgtSWlJs1AxGPZc2K9jnxC6LlFk
ZBOc1iXMVynq2TZCVP8injkgpYT+SdpaPTPGF0gowB0eIXJIcBLZ9d7AwPaFtdcP
684HZbHjOI6mo10ufPNSodmqZWo3rQBzMuveBKy4+J0YuV57Yr4R0sybzOgTTWuD
frzZ+RXwPUQC17z4fGyXMJ7YRaZN3l4xkZLQJEQVKicnRT+cs4BvX8KCNhu9cgsE
n+EE243flgqzz/N6ntJkKddftYYF8TJFCqSpEtPFfguAxq0vpOeJypyJHFLrIeK+
L1COteePT/m2fG3qvMgfYmbO64oGgfbTNdk28rm/kk7jPYer2/IwQtjuijIF/khb
vS42n0jCuBDOOW/C4OBb1vBniV1UhdOMD5YJzCCK0QnZlE3nnVQUVgc6RkHaUMQc
4c5udJHFdUjLUb4DXDpaKkejDplLcMLXGqrkR/q3OY0+OpNNaxmJwucF9xEabv5N
rlQMG/fpIfW54/8DUT0qeqyJqFIy98ab8ge4S7EljO3iRMfsUKkIhKstRPSLS98+
4LdG45I+uXLratEiTnzkYaxA9s3RN1/q0cqxebLwtQ+Sd3rYjZt8woHA3W1W3K7f
F71qs6cj2u+uGkIYLcpXgV1JvmTMD+8Z5IjOedEIl+IcDFKoBqoePY13XwrdPaou
DU7UB5MHDBA4YDqlSShh0daRu67bb0ukvVZNjwqlCRF8OuK6YCI/20L7QCKy9bNI
HL9DET0zUa6CTuRAVK8kbyuc1VlVuvTFjvHfFeq9aA39ACFVa6a87Am0KpBN5lnI
CcHznvzNkXUyXYxfc7psPsoWgwP4V+noUBzeb+JENUvD3Bq47uytQbKZw2jG9Zbn
JPA4fHU4OHn9GaaJkr/FLNAqqku9F+5nWcNuoVTgdQukLGgKc3V4yoR9E1uYqP6S
FA5gBCEI1fWQmcFhfnbWIhVorxYrnU3iCs1co3kSF1x1mi06Z0LULsqKJBY1YJPa
/ujMqJf3Pg+VdPUXbjIDJGzaKtdd58o4X00P4+r71sTxDEOxDiJqG06w7s2AJhcY
DVsclWRt0zCQ1vq/coB40/uucA/+RMNKz9VeM4hyaQBXx46L+nXNN/shP9969Wtc
P9laUmqEhJaaBaEmQEIqabOYlf8UUZK7fW5nvc+t06dl+36Kps/aSzdAu///SJz5
A8TysfavM/YA6+DGWmak2m8h5V3JPZ9l76jqpX/7df5yjuUlwj9+BNOPPBSgdSW/
BeBhECfDg5tIMbftAGnS4zU8n7DWQAabZdzchn0EWz/bF8QQyIQMWNSVEEc5rzjX
X2lO8YJUPFOtgyVfZyVPVk/2CxyuJTayCaejcTrbIVns5BaJ0c+l860J8wfUx0Lc
gT2bsYs5P2Ca/1OWeSsdiBQu1qFAIO+uwdd0JV64oA4OgasbZCOwNWPQdHRwpGNC
LWLaE//TuVuB+cLY06pyMEv+8VacQMD8c417HWULpq6VJEgnt+1jPTXk4+cAMJgW
4nLSYwbYJYotRYeJXjtEVy2szKmd8jz1GBP2S0LzBNbj8i+v10OTgoWccjX7eusH
EYq2I7onKmeOg/AXILGFh9a0Boi8TPLbuKLJ+jLcY8fq6jDxBZW/98aheWXoMgOO
E16sqUT4slk6ZXHDTcpEh+lBDI/+gr4IdvLRFGV4iks/lEgUTN+9njHH/m+iwa74
WUAAle5ZEzt7IUCHwHKRQ/5WKByfiBErtvwcYf+M73Sif3kfgJpuXM8tMc8S3D0Y
YkfQ5qwxqAGxJ71+AXSDJkaeKGVR5KFBAmWxHU/d1gjCdpbBJECHrFOpCQnW2OjP
6rMvHNzR/VDtXO91TgUVm2SO7aC6pk+XFVYJxV5ajltk5ck7brFXNhadYj+3AdMy
2NSRm4ugXRXKQNRQHe7I+s/B3hTYK7xz1pgRlaaQTTBSYGo7OI68Vih77R4U+j7K
bmVosed+yzJgyY6z/ABonB7zqHOqyYnBDbNaFYybxMx0S7XmxgzlwhlG4vGpQUwI
Pt9/0TR3eFcmzPhqG5C15GOFLkNv92w/bar8erGvf6LGnH6CtmlTHxm2kM1wRmft
HSbQ4iUTjA4KH3itOxl69gqpgK4FUJuIZMOASqnhSoaECbAmzoigUdLGD3gkn7GY
hBdlf5MW/iz+l1gLqEiwMhLWQmLfvbPKfXX4JOEuYiZr6lF69AXF32vaOgUOCQLO
RGg0DZ0/ioemuFyoOhx9CJmqbgk3Am+KARNpw20xzptnDf3NIajffcZo3reEGYic
zwqt1gGi9Ur2CVxXvDg+F/jgZ9wuP8bXi7LyHIf1MNuYbmVOgAiJILXB6iF8k10s
qYPOIOPRdX/v2AL0LKt+5vcFWiG2mlzQA/WA3g7yQqmluZN4A+/ZSzcqTjrtkN2P
3jybhargIhxbHHOWh58hDrIGS3x/Xg4ZhvB0RifEMSamNOixwjJra046xboK9tTY
/Vm5rnR+r2kBgYraDc3ROO4IYL2WBpyZxu/azWV2CLLjSRAXXZ4MU0VRUXRW/Z36
8fiWmdJyLC25OCLrxU9S1XC51+B1EJy4GLNRD3chWao9LN13J+uxdT+H2G7QA8bD
Kv9/c8E274Sd5MtofDnr8RwQfzmNyAxD9CIf35LPLhdxd5LXjWI5EY7gOcErwu8E
buvUzxDwS7vnbabBRusDh9g1VVIy8ugzXQKgXgJEkxC0ROuK9wPQDS97kGVM/BfI
Deb14rcJwL6iiKVcR2G6v80SZermAcpVUPhLxJ0K6/zRXoI3edk7/XPI7/d8f8F/
2peT70lOb3TdBlCRA2pUU6F6+ibeEomvcsmAMxla7GzgbKwJAV5wc8oVhP6ARFHt
tUyqSMPlq+IZeJV2M56FOWT3eYuw2JkEXubE//rIp19Pav8bvBOkb1TcT9TTeUFA
0KpsVE54/ET5NQD0Bo6RsrDCutV1DtuL63BqtXfAXkDdTc3Oi2CWFOB8Zk0trEao
vVk6jHJ0e6TznuAnZFq6YV63rADMzCFWfpBsLsDRRFk0gScaqW0qrWFlf6ALpYh9
GPJveWnweKuO1ydAWVG1VohtnHmqZ96eN9P/BGTCModIykwRrIiN4GFk7dmzpGPK
WHb4GFPVBfd2GqG8+vizR4NAPNllz8TeQ9sdaZqQ8SCxGazTPQSZ4V0nvBd3eSxk
nh0qBZl3yV5fRFGk7ODOblogXIP99tGBh9FnVmfGqo+jS+AGj/Q9AstgDzJJu7B9
gQbPWhiWphvVDk24jjpqswHohFK0HQP//tW7ZQRq4GVwjujt3s3tuN5zDCAm+geV
8JM+IYJWQ3A0urDeC7ZVEF7GtQr/97XDbB91WXtc5sQlaZpd1mcfHJxKsrwqDLir
Fni52+DD5GVRHqPA6rlE2xNhRyL6DHNbvRYUVj466pn5T6dvP6NgAy9ZeqIcmkkJ
CkSFE9ZGMwUYdwFY/yJ0ayID/jx+mtyeGRu/TK4E9WmRw94IkR3wzw0pmWmLocw/
ktUyJlOZqOAgZsW+VsP/0UfSnyM7Cvt4AyFZ+A5+I9Hu9xnvteBZlNFgVAn80HWA
ExiUN/pMyBwLVnaCBkCjPZwkPmutb2lVL3X2pZyj96vZpJ+aJEpUIc1MDSEtYejH
9yakcO5emLy5tXvqo45crrJu73B8szx6Ur83paMJpYh6/NRylFYOZMb+Leeg8X8Q
YlmRAvHs/3/8PdrN8dp6yUiInpwYA7EmA81CyTr/oF+om/p3Sh35adyb+e2c2oZo
tNuUhUyPXceBnESRiL2HVStAXTCvjLp9XfP6Ty9rfn1GZ+GyBlmZR7weGAF65pYj
EvErNQEy7y2mq8uPpsNezdFVxUunekBJP7JrUDMO9FniPrZCZ8fiP6Mo5ktYrlXU
a+rECYHflzK91g5txjL62Txyp4eHmmkB4F7OVrRPdUe0orV7v9uwACCl7dc22/Rt
4tNW2nsDVIryZ68Yuz9B/tk6A5A+GesNGw+c1xA7HOPrvfm7tM3W2uHb6bgg1idh
8a/9UtFrThUnnNCqs5SwjewbrGFJ7LdbK0ysNEBwWKqrqpK6TWoTRsFRpQa5JAdx
l5W0E3ExFAGfF1Isjh5Gihm5dNABC9Y7vZKVCVCve0+lnVytpMA1chWeA/GkdHrJ
B42n3jYIGDmH14JgRMr/g7TcTxm4jWlfgJVZE7/723V7my9s+m1eQwXRaYE5k6CX
mOC2cxhY+Eg97jxp7Gr6JLUggzDgQnjrtfZd2Oxa8wF7aGTVeEhsM0+yirlbKnby
6E1t4CpXOY08NRLCb3OVlDsNK0A/lo83+OdVHS2IQ1+FWJOAXGJFubAuUe0HyzQ4
kRsPhdgvsokQtEKo6X2d/giKZZC8rWm7vTZFUPt1Pd8w3WGawVNbh9q7fOen145+
zSFA10Hq+C6oPKfvX8xEva3pdYobq1QW64esGh4cDy3dYbCRYq+lQ9uY/MbC5w9L
56ZJsN2ubtXcmmQFiwhiC3ciJwMUgyAR+lrpoWqSdXIQJSQ189yKlN8b8dwtdK4w
naShEd+O3GD3ApMNzAh+/UjFHnA1iaAUd0oBX7Jl8TLPHf4/lBHjd0W7i38i569q
xLZWPJ9CLo6i06O08TgdbRIjnHXpx9nfo+v7IPhMTF8mw8oMW1l8u/0qQvbULHsj
ZwfZd7JZrX5BgavFVkwNwkuAERo7Xps7sfoqYCEvbDUXNEZWX6dZKFmCGHttQnw3
Y5TgwPSRqQqPdBxAF3Rr10JOsDTEr5gZP7Ag82Zmhy+vLkKjem3p0a8BJpq3/u03
TM3VaYjbvTqlOP65E0QlmFON8P5xsrkNlyZBj6x3Xwny+PE8WctGShPJBVar80dm
KDIYA2FS5iUhXoah9B6aqKFMTgWOc8jAPMcAgN9Jx/ihkoYeGFzu5bMTHfH7PfpE
mmhlKv0N0ZObKX7PzJJrdFp5bfNZEEn3pSKtTwcxyCCW6CHEWWPlrSPUn27qCRI3
JRvOiPtCOLvyPMSdckPPoa67x4TS4YN2Hb+N5zzQ6x9jYgqKZBOFH4iQTipenyxg
+5wqJTYXwzGL5uPmBWw3UL5Ipwed5N1uTKluhhGZqctUrrSZi3XfQzOTiqtvlz0v
MzIqhgWMpTssKNLPBGKXiUmKg+49wTBW5bg1ApL+CpIBOPaegdoQyD5q9kLN/JoY
WVqQztOZVNy8CxrRKkkthNiQXzPDuQjw87mQYCaj2Se5byjzc8NA10yI+dzVlHuZ
NZYogxa4YWQpbWVmn5Rj8766J9eBS/y+MNnIvStUgu0TGtDDbQCtqpcpRGAk3/SU
lPAsRG6Qbfmc04bQINS0mawBt5wkdzuQI2PEu/J8t0K7k14GLjUO33sKwwbiilc/
TeY0BXl1Fy9Qx+Qp7UNFV4PsJ+XwtH3coKhsCpUcgvnuejMFHKYYYQ1G0uKK5fw7
dEo88Oo/Wb0c2pDL3p+ZVd8M2Fo2FSNyn8CpwCRVPPWEvnsuxooXKmJkRJKyh8TO
cN33Btqfy3FTOUV3jsmpRAbUcJD8rwLUdQ2jYjrRj2WTpvCXY3YlG+2ysUpwYTIm
+bhM2SqF0jbX50qDhfohqrJdIXDapd+rTHEf1gPmq3Ys+1keP9NKzUR2w6MqsYGs
rNhM30q2be72e6nwo9LfDsXu4fzsoqPtqcWjGeQfSSP0tvvPcMXee120NViBR9RP
NrIvoQVUeP0pZS4IwWKi2lXIDIcS/suSkSsRA5TaTveoUkpwf9VaYFxnwf1Rdj0e
7WDeezBHE2XQ8WNdTT+q8Py2Zb5aCxvmLFYdGrIwtn88tR/dC+HDXXV3fIu9YKDB
CJdPCcK9bAvq4fMd2jbhYmgY8GAgwZwct1JrAUb77vt9bvprygovwYYSVkzj95YG
wLpu/jdh15uJsAI4mVCoTTrFLg5XTcT42W3wS5C8tNE1iFD1tRkGU0av+H4Kk/4a
QHUXTwWSaY0cqmnlB/wFffZeo1ZFAMlJTE51hpp+WgnggRRqUa4vthSPWd2AosME
Yr0dwat1GC4pMK8sDORIQz/YvzAGS1gxn2BS6YQZh7Xk14m3BV2vookzn5DVo+r6
9ZiIoQrLQw0vbeNEuI+M83/ICfqZOIblo3HJHzk1iGU0HQn3i2qfbS5hH7Szs3Y0
aRjsk1L7lnJmXE54H/Vp09Gh8K6JtLb+f264ATG4VjdPh8M1lDCnAwN4hJ/1uJl2
qYWi/BeqC6hWkH6iSnVwQfhulzkBm7nnMxfNr+ed9DYGi5qSZWy+XcnMA+YuzXnQ
41OaWWDVLDcVRmSRCGgvZ2mWvB+320zhSVqa/WNIcACaqn+wOQpFxGzRloTN6PXX
O8UF+oiNl9hmJKAFtyfRV9e3xpESu/jNhlikJLfmt+LQARjovf7A3KL7jEo4Jbut
NDrjxDOGpb+qU+iYLkaKgj9sA+aA0rS38N0Ehel+pOvpNU9MTsXBxrEBVV0Pr2sB
sFTY8p41f20n3VV0BwudvjJZP4/MrFk7Bwm9Lf5YMYiYxW9+4tmtgWjEDprPBAZb
8nmqGhF76dGVATQFmCpfJF2Nez0g8yH78B/D32XfDVrBcVC56TBdRAjIKODj4hze
0k6A3S8B7cmgogmhnCSzFKfpvDOtWseOa0rr3KMcn3HGd9VhyjLnuPHJCg/eL82r
0DhV9+0mMxh52xzH7IZp+izYzK9/wxPieenGwcG3Kp9nSs90iMwgADG7Ioqn8OtF
j3n68M3QzLKu9ZfYj9IcNNePrysIbaWvDZ+AEkN3KzgmK1ikqDEMh5NxRllyvtRT
A9T+VDIF3qZOr4T5Ub+vb42vMvh6NrMKFpDkJQT3Ao3ef46t+/CzTe/3zsW1c/rP
BDrJlGOA+VkeWCPqj2Yb55hRmw0HfvfMN6O6gfL/8+NKWqaRT1HQ8B8s0addJ1SZ
GeoDYJ1h3r12wfWanaNU2mwcGia3HvoklJYrvHh+BLcFdBnxhZ3RcsQHaXBiuGhS
01kKYHt9qQsrN8REzBeTevVKnuuYQrRidu8AoVThtU30IS5LPnojOZ8rZ3mOwiHy
oXwBjkN3cyay4NKW93o5giryNQJMPaAZtg0RN9DYB1+FIrZF8DyfcCFWnFE8qtho
5LnHk5GT8CKQKbd1YxwqfVcBwpeGBjZ4pB/ecOzK1Txn7NQ2e2+wq9Fa94iSaknA
rw3W1p/Cb5TEgCv7TVHCgWpBoAGDJF2ljOPpSzMEMlogF25Z4h0ZvwGWzmAqeSTK
ogHqa3VzJ/FoqwHausdWR2ZCA4Th/6vqVuC15PqpCzr5OSAn7xqFu6g1/1B8GNaj
fgtUOW4hQoDd0RDG9ZA0Mllxbf12YXlZ+JXtrk2i/fRSpPL+4fBK60TlJqPC0lLP
Ldc52bPCJR94l1V4wJZ5O5oe9Ns9qW/x3wSNpGnv4eVLAbKOuT028GgsP01KjZix
Y/16B5PESabYYqR+WjgpYDZCgFln3we857WQzEVFPdYYgcSH0djtqhiXrr5b+qcD
oYhe1RJUluF2lshjXpvVdkYru1DCmhRvV6727Ynw9z2bWPtd/fbXVSwuvSsdcEt1
upZsRVvqeOCASQOmj6oqEj9SfXNRFK+QYtTi4Ctp2SncS2x36AEca1QbFc3zsdjU
/tyMm8S1zk+x4lefHZQP5W50MZjW47ztApETunbu3PnzhWYN8O60oeO3+hUuX9Kr
Tt6uIfC0Jtasqqx9vqM3H99ITlMUGxsx+cqCmL0xzIR1wDSVaDVRhAPHq18uPEjE
VfzbDM3djBBEd7GDYJCikTwyX6fa95FKw4r0QxOUa9cTrQFGSEarD5wZUUZXI8JT
m3PJh8WnuHLkpdspP06TuxOJ68M/al/oCmritspS8P6d3ERlXjhu/iUt+JjAVRKa
6J4Yys2kdXrVFlCIuQh+fsh3ggGNTtaRlbBVCRn1M35uTmUKnju3GAUWYb7RN7wJ
ZxW5PG3XrgckM2Rd+pzRnB0/83JxFdoKUzfrnN7Wdagtc1Ner5SM316WIkZb/szs
mjjQUGw+XVe+V3Qx+5DbDSChzBPu8ETTZDnvMOPNuAfVgYX4EcGXucbVwLK5dSij
vp7kiQr4pDTcsv4x7+Z5FIcZF9WhS1CJdJvTLc8utnbKKNng5zUYK74sy79lkxvY
BuwyPkTsi/uHBOoG31l2OSAZl1C8eJpTuhRi0F0IRAy2Ppnbyl9NkutkN/yd36vP
1M877Pfn5Dzen6MNNWB0/lD5eeLmrfP6NrqnEXunN2cHgXdGUfA1HtTgoEkepj3C
i9xe1TZH21j5vGQIjhHKOQ4Q3MpRyYbaDcomMGGvDKogdXyBuWznVxEktd6rIGOG
/dH1/eJfrjbxxtwpwpgymzWMJI0rtJeaBDzgHHF8vdBqy3brv4kG4Ka0BJHmmLzS
6JG28iKsowIyb+cFzRgSyO+TR5imAcFFJPbgJF32OVFWp164it3qKkQomYvtfG6z
JCVNF3gdMKXpP7nPltNu1DG5t2SGbYt3qm//6rVGmXVx4Aqj4dWPo5LwXI+7M/uH
RUL9EN6V/9xkq6iRnk+XU9dwYkE+V6EtrP1lSHEGIeW1496t8YUDE9Mcy5adSYXC
U692acCNYJKR5hHBA3TKYZEv8f1bdvFqLla3YfYHWoDTCZiRa7SG47c3RQN0jUwY
jTpMzLRxY1V0/89FLD4CtKatsp76ZXPcHFTaZnJ7qRH7GSIxH2yVhy0CcqjLsJuh
6OZuNOr6nQoYifN7JZhMeJ4qxlfemoS2kJpNz7olvPSJgmZJ8wUkA5XR7OjxcD7L
d5kHIrSOdZME4WuJOllMOm2nXSZmGmg0ak4SumTFENEJKCD6TUZSX4w+/4DA0qEs
L8xsbkLoTnONmFBGTfII1lOMAca3EkervYiUBoKGz1hR1TCGvy94HLjORPq+d85p
jtTqMxARyrECLrzKJRFVpA6gyDGEmN49T/IJUBSGHVL6Rk03UcLHYzeiWnJkEek5
PWDgHsitB/tAyKnaO2a8hZd7SImZJkxdpnDgHIBM0wcqCTjPYpfd0aAwc8yxR/6F
z5XL3OMoEDnqvF1VPbqHA2eorF4nAM5z34H1ykVZ5ZLxavJdZIOz/lqaDfu6cB0a
tvDSHycwCaoNHMBeXKEHAuIpfRd2razVgN4IWVxVlNY0TnUNmi/6L+R5aaD6D16Y
PgobSbBizJ/o7ENZLFKSKovKBGbspfhl8LA0gpQSk0bCZvR04YRdr0nG6ZcrQV6K
UGZxWGy3juDCgRL3YCyrkUFj5DuVAe1g1JYc728fztf8SUGW7nY2wJzWa+yraWT7
UyKRvC6voqtH1Km42OeTEvgFUWefxHd3Gjas7lp7BfQFvTxFEC2YhjmIOYSQxDbI
F68J485IffNEwub10rvQj4G0tNnaVgw+wn4EPrsdKKoBhSZFFbyV3WgltCb8p5SV
xtJA9XHBBfoz7R7rvWFEOK75c7ymgSIKjE1cjZTdLnFxueqrnIYBTbvlA00YPbg1
njjCHteHxl9cZVzuNInQrq+iqQ4URi1pYzzYWkAi+X+RYiE5dlzys0npmLqfzBR2
AQp/NV6phihD1sE2jb1kv/m1pCcVQbIm+6F+8xbM3obuHQj3eCNQYWK0TaGdw8Fn
1EhM4Q+uM35Hn40PErxoCMqwacxw1q1nuda9JBoCL9SH4dt2/MFcEP0aEe5tF7nC
lGW7txgn8bKL+8hjG64w6VJ7eOXMjgiyIb9726UDPaG/vGm+4DlswfRY3dv0iOiK
r40Im/9RPXe3eKwKa71f805UW8JjOdclNTOOamEgcwszfBryhV/B75e0/lc61+tB
K9JjTbragyWTqApLo7NmwdYS4FN8t/2s/M1/zPzmUsja6gqkxCVderIuQR5MK/c8
z43+x1VD4yBg4T+deln8VMedA5+Fg3hqqmzvfqDqyeToN8IPYykNtPJbrDadzDw/
QJG35TRfKsh/roR20EnkfDJ+5O7Q/n/g8L/5PFkjX7QhCAlhMQ/nH1buxu0VvFlT
YrwB9SE9mro3vKkllN8jfinVdf5vxhIFm4byebXg7VMUJJcB5Rt8zT1CNzX3WMig
vig0DZjd56JA7K5B6kUNFLXas/NIIACAQMWJyR68xInKJeDV1zEylGEYzLUcAzDZ
Zf+S6/X+ZtlPaJ8VW8sR4s41RjbE5n+svWQ0gMCeKkp399tD5W+4xYSDreCuZWcv
RzeSAA8LBbjIAkRfLj8T27iHH0oTDpwXOhp+kkPL4oHneIJ+cP98/0DjU2W8S8hm
EGl5F4bCMLwInpXlGxoS9EkA7SCyLqcoy171Sgc55ZAd/s+hOdLtvzSRxTn1fMsd
jmQ4Es2swopQ8o9otX9AlkkrrwreHNlCuxCD9AAcCSQ7HPe2nAanRRRQC9BYSb8G
a8OUi0B4RGiNe2TYnmaGtsPZxmeWs1OQVvaA2F/YtVmkyDFi0Kmeq8CtM5342X/M
o4nBfXy/2a1YiQKIeGOq8WhfBidrxHH5owuRFeFWb9qR9PgRtVWS4Xy16MdJZH69
zxYuZWyM0USXFBUucXsWXTxE0hC5beNqOpgiJqLK4q1wTWiHFgISSXOpYyWNdqLg
XPhG2q3YuiZsM1L4zBZ1AKIAz3KuwEAWif+5v8qWEcx1mvm4t6NHHKwByUI71Cqb
dKrhQGv6gYszSCHOSn45Z0lU4r/hCahlDnkPxr/BXjrymr7Nle4ko7/wSyJxijib
ItFD9yLxbsG8IUMWf4pDaw1zhX2JmPIuLZonNwIRzE/PeCPOPyi8z2e/SpXrzDCO
R0uNGtrkqIKxmwAW2JgASgQPGfDvnUBAkJVYOc+iD9K2v/B6X7lp4/w1ylh8UiJf
bSZh0H1PXo3WqxKlNUowrE13Z9oyj51S89pCL+25QEuzyKvIzKlsFtdwOJ6kjEpQ
BWKtHGB1EykcdCJVWBNTyP9D4OTKv+b9X8th79dFKBXlsx0np2nrRopjzqy7A4qn
mVU7tyTdBmguSLVheO9HSMGhGmp8hFaJ7+LTM7OP8TN19gh5NdNxpDgPrp2F5cFp
a8vXUygB/bqAbjW3HniGsiE8xI7kJOrPU/wXfTmuurUDmEpoyWIAqmb6u2BeC33n
STLhYpYn6HyTZImIJ8ABbWvnCYNKeDZeJox14enmsg+SFDDbhdsMMw41ashqHY65
8adwxiOGAR3j3ZK3T4uiczgh+Yi+SbOXXS2Xex95ovoiVCWfb5wRKFsPIoEKzoGo
CtAxqhoMWwlGCrW4lmjTZWKeTnDiPDXA4FVf0ehLX8HoBx2qro/GZthRFja77Bjr
mS/3aTMIbQClzKqkWBnHpYIRYSiavSDEJDJW37DaED/vg/40aH8NDlXRXiW04er6
tcJbOd7yxAoY+6xEXjHoDkoAUfaX/f6zXTeUYSfWstnyJFB+Vp6HALZd9kcxrxRx
7JLUK9cllJ+e+eG8fhLFBnV12ZVlDFuuLYqgoGqSghKJKeqHsVUyEns6jXrG5a5T
l+pyz9RloQ1TYW8p3tVpu+EE+NxA3mgBU90LfLXcKz8KXi6w6PH/i3f8D8F0/tet
kTtCS2B4DbE+cBXHM9qTbgcN00P6ZzxFNf2nyfAlQy0rAJ6NEYO03pR7WfhhPB3W
5FioP8BPs5qp7qnoe5vsuwB146ggue4DSFMj6Yi3+2umFYQK3fi5FMFt19785E2R
zPbul/xx/JhTZMX0Ev+5s0BKa3XcpeNL0aXNAXQqIG9a14+X4f9pZneyEsBHY9Uf
1imE0IUceKb1P4Zqs2Yyg7AFCBfMdAkny5cfQ/j6Nyn+HGn4NsPCX3IS3MuSIBAN
yFEn+CDU8hvwULnQBeF2silrHPVnimnK6zACaE4EXRdZQtqsiJSJBVd7/W4CX5NY
JPoqUsmSp1/ENjizzA74utpijaWTdhUrk8hlePPLKMyd85pKp1O8cKnem59aCfcy
5+GUwtkwhFFBJyIStYTHsCo90oIX2U8R+4RSjhd7wB9ulOG3kSlEdNLkdXhtVBTd
S9UBgSALMzpeyEJo17IEFPQS3FbVe8y5m6xQ0Fk7gZKs/FXSROkElphlV62ysdgG
5ZVeBhn0IcGpWRWnsKDrVkAsksck9fLbhnqYiL4hhLHuZzSjqh37uF9QsCwkYsif
Cc37reILT4SQ/FgrlJGrL2idrxgwjn588OJNtvR+stnP1iLXK5E5PiZKhITtwLsv
gXhaNNfbjo5BwpQBI5FZryg12w6bTpfnYiDVsScLHxXLKhrDmkstgz5mrttfW0r7
dDjEZYrLZuc5d68SFPCY3wkUzcuk6h1/qOyQy+hDcs/KKNlPWqxWQF8L3udyJOKZ
9Tgdv/KSbQg/crwVVrx/mZG1GCN1UV8RKbLYaiyWciQUjmIXF/Qs7ZAc5yhHKbR7
Cw1a1HYt/3DTay2ZGRg9YYr5pK4gavIDPvvGbfASi74ffMomOKxrMk8vHKZaEjdJ
HtkrvfPh6qUnfCR7bWjF+T8aFWIaWzaqmX8rTSiDkpjJ86ojQEGS0vrfJR2UMKF+
cTErVbBERMfSTmVYNsdrK11R/4NZ0QA96n2DV8FZfZqtP+8i7ppKphFq4qzeIxiC
Nra6eEYHyCQQkLwH76cxy0x7jsjsHP+hjyhPwa6h3Je7NTzFYKHeB+/XKcoAu90Q
SuaVQANAaOmoLDaDXwk7UVMAM6SNlyRMYUoU1bqu/8wmngxgsA6vcC9aftOjyDjz
S/BrsOFQ0OhQQHtIHHzg80wWFxEun7eo3b09gSN8CIOb8wdgvr4ABwLktnJebeX3
U9v9E6tcXqIbcM/Zkh6wxvyWmD1Aqnty9T+OYJ0gyajp/s8AojKErV0jdA5CysKq
i1pUBMs+HzbqDxHcFvYdkuQMJNdkbxfmLsnqAXWFhn/bDeuy+/iDjVUI6zvBc7Xy
i2WZJQbGsnn+ficntB0nQa64iimB+TDah/FBpQCFOHIwSZken2qU+C/X0vRuganq
nkO/9Me6V1mmG2kCNitm5glH9d5HvG9sGvnuS5TbJJhnkERQTu60iR4QVpEDBqW2
KiQRjIGuiPhG5l6Qe1NiHs8hoDXHp/u/7IRFAgQuTAf36EklsIWR/4m9olC2iYhg
+N6b2c3/Tlc7bZeaNjzsyE5W4spoQnEF72WmiW524GyqlBMN9L0bHbnrpl3rY0JA
8XWeNnkbiHnToU61VQazJitoTde9r/xQSRGLdmyAs6tPUVAp2H9ja7nhVwAXLNjX
4V+YnLSN5wVD8rn8FQFt18R+Uf92A4RTD6kE6SaARHMd0J4D8Q0qe9gB7xQrGhTF
/vuSFAaWRuLwfVy7GNfitrZxJFCea2mP2RrKOVqNmGQZ9Z9sJTgn0DhBca4eohr6
xDpWO3vbIRNrDW0nn4tIRZNnye/xd2IP3n2Yv4n7sN4rpNwUpp3khhcTmHzmNNP1
n3TeFRncXE84WXMe2ZLsQP8iauQ0Ytpt+af/ImfnDMxt6qiL9yQ4NeGuqjK2QNdq
G9u+mclMvLPK0V8nR2DhUBR1fNo4bWG9vTYV8tZfGkb18SmrfWj396/Eagb4iylS
jwEMtILvWbfuD8tT3TFofG9XiptJiw+yCA0+WB8XIl44OTBJduh892GaOT5muZAQ
5q81xB3XKpCTqI0ElWA/H7RrMVWSEhfACithVdhahfJ3ttIh30LnSkJzS7npXT/g
zEp3smy26CrOT7LzXojTaOSh+QehdZcApv3sU6iL9ctbE0hoKucigbEExZZX8jep
VDGmWcFaJQAu8cKn2dDYr6KJYrpesS2IacmVx6BP4usnTI8dScJF+ZqqxKFgjtAz
4eyz4zpstwu+CgLq9Np3sOv1+HjPHqVBiqGXBGHRSKnc7vFIw7adPbZjMYUCFaQ3
Iamkv26t2jLBvR3abFhckzXYI3CsmtsNqHFFhUdQYKWhIymk96YGMO1+LZ6YwK7a
0cGpBj6kKnPDjObcwVz/POe+Sa03NWifMyJicSJNsWyQgNVT9V6D8+czkkLoN4nn
XrRfsAVvLOtAkJky423sqnFITQNtINnj6TrGbprHlOqZA9+0dPSN4zxjU1dnokP0
7dG0BFt1fND5PpmxsyCm792AbQpgNRhizr7460ZTuYkZBiPYLDwbXQwthtRYVbzU
CmzFFxWtGX3fUdFmsHwxD1Jonnzo9rVdjCTlIqWP3Q79jCQaxwzJIvQlwo3WZ6qk
Y2HiPiLzARk5IacntaDSo25Y6cPPhAUsqRuWTOekgcbAdZNK57i/R7GdW/I05V8Y
qJfRQ2zDV7qJ/4F5g1TrvVCDlm+lOGjWglaYtQsSSgC26zCeJaJd3BZtaMt/ZqzM
CZ5OJvWc9SpA4fN9mO3gP6J6eZf2PJ9BXfwMRoZn15DCofe+LOiRlbyE5qycdeWY
V0AVze4MlkrTZrPWKXtGGqL4vIEUcYEn7aHT8bPHb227aQwSkI7qY+VhVASHS2If
lRomxGWDLlJgwdt/A3cmtJuaRelFq4a/Xm8yGIQKCSHROnirVv0+n8PXibFzaZYE
Rcp4k1LSYjSqI/vLE3W4S8TwH26dfqJhNOnsAQYwLHVrN9qn0j57jxWQYj1abMpF
zPb342b3PBeUeM16PuRXIYO7WzpZ3WlGVzgyI4Kd4qvExJY7OaAuKUjsayR1u9Js
7Acn0m5jXTWEq4OfFsaxAr4xhIEvXm9HgOYzMQk9Cw+foXSFdheqmnz0gmHUbSui
r3TF7ajk4gyYIoQuBUPvAdjVmOqsodVvV2X7wIfOl5ggThQU/X+iKgssK01kr+MO
C7I+1y/DJs0+/HsXztVauBo/gHchob5sTKz2ZwuOvCvBL4pfqAFomXiKYxAdI0eC
8EywznMP0HHXHhScyPVLcrVJmLHn1hzy/56nc29RewYpPyZFMQbanwQkyMJkQu+c
bidNV0XGHSohrvV8y6zuK2ui7wEtq190Zlaxk5755f5M/DjdYmsZHJrdWRcEDWbz
7URwffan/O4kqYKFWuEfGG+4M+L1sF+l0DrnV4KuUkB+ufpx/P8d+PNBJ6+7zrg/
Qd7feq1qw0RB4G9iEgWcpmlR2QalwkI4Djp+e4hAfE87tUfxJszb7DEjlUzw1TmW
uRymozgi+Z4Tt5t0q4prgZZJDJxSCunNryQkdFFQwHwX/TE3gl/69VvPC08rYM/0
+oxafjk/T/qSW/We2dDXH04rv0xhGwV1ocA3b+jzRJe3mmmE8kmsTLo77RdT3pON
nPKNbUjnH+GKvrIaF3d1p1fFSkaqjBsC0MRv5uqkoueZJttFRLZJNAdO1o0GDoXV
Mnd9M3OqpybO4t5CMPErLoToQ9TKz9M8rX2rnMIrfffG0y+gXrQ0DFqOmHA/hrlL
X9te5d/sc55YthATTwEodyrB4r2DMid95uy58Hk1v38Qct9VRoIpynrv6qV7eKHe
tL3VLhj/alr0YZAP+9v3ZZEz+bf0yLOxCvcMKC1nYBHonpbLRT2Qoh2JBeRa2Tcf
jUzVxuDOT/D0kRxLpVGHOxfXNDx2ygMHm5Ao5fxCHiCrHmWnlkC1anYm1jPxr4B1
vrd9u07zqw9sWEpkff9c9/Hyqv+II5pzUgJHw7NZItzOReFchIDOxuca7dTTWzyN
GMXmzOFtCeKcmHChujm0mn+A25hp8DeRE1bvzzv0lnlmTePEvpG9EuT4Nh0W0nUi
J/QQyu4RAvnvYOjxvNdUvD0HICGA+f7livogF3oa7z1fP809BDswoZUajeS73Rj9
mmyc3Rzu7RqG6dMpxqJBiywZzuGEgGhNz6T6DQCZcXEsY+NE/QfSvKGSWB0lJyNz
v7hkaBGfV0HhXK3osQZY/wT9X2R0Ra3mKkaQRN4ov5avo8EECXn8alPq0h3SOU3v
b4+2W1msVWMQlqb2je5BDPElzzGJTINiRHQ9UbYe4wdA+mDy2k0P4m08lV4/AZX/
8lziQi+H/CDfC0hdEFI1ZrMAnuBxH2EJilNUHa+ICwf5Nd717Iva0t+lHeeB35WK
veIDDyR4FWUVkTX965lwuh7T+VBAHT4o6dN2qDr4p/EfRKLIKl7dF5X/m3Xi2a7e
r6DGL8bDZKQa42ign01J3fFncHWGWZlWEcThXQhFSGEvrCP/i2D0L1xdG6o8byIN
psMGXGkrpb9AvZjYgNQnypfRy08QlFyQEW70Md2g2VCsfYVQncLBmq7uC9GG+bLr
ZvVBFM7bBvx5vYf4b+bQmtbC5zpVfYicm2HNKvhs/TheBfbGVFqouCkRxJ4fCpbL
pzV0kxnhH+JKrArw1IcZUyDda/nIWNxDW3mqV9I/LhziU4iNJW1ck4H24pL3uuKC
3WoSnJVrHdz8SyHNNxvnyDOy6CVOY05bhBs7EQ+JigPk5CHrPF2Bmh93rHzMGOWs
MUD/fdpJ+acS5fSfKZ+NKw6OdBjachppf9USYQ8CppcEq3b0jDc47WQwtv3rrzTj
EKXjWCcVkYQGXPqFkiGVQHFBUtYZdXEgwdCeShP6/45GK3htoG1D+41kDmAFqLl1
AsvpMfIqSs1DdKBNGmP7WrxCwSGd87AHqdnSW/IoiZFtad/ZvF71par3d6ed6gUQ
xoxxPELqr0Ev54WeWsmbRtSitZ50/BlbQPjd9NNwfCBUHmoGq/0SGgHztNvlWjBK
1WuI7QOD/fRoLckeEdQja2+zxKKunegQ+lGepiReUmIcZHPbHHZP+3bieUZ7opIH
BSiJy3MnwpHfX/Q2HxXQvcQqK/JPOv1hp+7m/SAjk/B4PugP6AU0O6cBGG4OOI66
y6GrX6YoklGam0k7UMQGmZAxXBZWD209SWJo+TZQUwnygu+g5Q1T508/XZV2X+xy
bfbfc4kp352Nf7KQZqvzdllxmJLplqKC/+WqNDg2Xnn37Pl3bbX/VeZyW/4+rRQl
1jFWsF+tMqholsr+k2QAT7QaNjvO3J0MjASB6YxhtBHyYxIIVGrHa+zSEmSrMcD/
4Eho+wwc26gptFWA9zOgMmevLh3pjZkx5+lHHKQxrqA2ZgI275Dz1A1bcAgZH7/Q
xLB6GYY0ylN4K6BUVUGCTvLpTGCxLXSVuZb+zwLEnc+EtnPfrpC+nD0znZeks34R
PUqKcpB8T1fIVoW7ZMIuh2Pf2rU+RXPj19VCWjCPMbhl72IY9epjy04cGZ87pvfO
sem9m2nQUwLoNXKjDl053KlqgySSPAgCCnczwjJuRzSJ4xVcWvoKFq6N/i0UY7Gp
hDyvVypW8MmElawrCFiVskcwj96pphUXYZ6H28mowTR42+YpX64EJzZXxvjCGaon
oeMuuWSIPMJBaTyFjPu9zb5Pc0gCcgtNjS8o8/OzK0SoVcg+BT3Nyz2yCXi9h/dm
oDkXK6LKrKb94R88/FLSNuRo7JfmIbDa79izWIrtc09nQyB5NLJtZNbftThcWe0x
QaxlRKPqbJS4pzb+C5a8bsFI0qf3H9D1Viu9aBUstU/QUdjRPTc+GoIBNnydH6pu
NH+I0YN3lHnyzYYnxrLZnKdTi1ZLGdnwIejWYFh05cehi50BlyaYfAvKsOVlBWHI
2SRjJmliLBQhMU5mOY3qLobbvJp0p9wvCr628xFqjF3oEdcRqA2JMn4MvIR7+GBB
L0SVb8Ma78xAtFbl9C8SbaVFoUPHzdH2DESAp5pxmt+HNKXCqurvhnMn/Y/WRPvF
hcp2ivgh5dsyjxg6yzO/3b3YpAQnIT7PDGxo3Uu+Sor5airXSAqzLzEHutwpxNjb
IWIHGVGasEWM96ibgDtPgIMjBLpFLAsJpt+G+RIZGN312aGmn44zvdx7t42o4gcZ
QquYvHq+YX27mQUgwQ1gneWnbu8a369XJ4YAnexP6Bx0cd3L8+atNZ2KBV8ou1oK
+PYyxD9mGB1Rjsb+u2l1Fyz/nYr1Rau7YHV9sop53O4gWRxRYA49xTF5LkVnrMQK
JmybpAb0W4sKERVJ3WxvUQBvEsO7x4cSc2aJImK7qvDDC/23xiKLGAlSKZBdnwuX
pdq1M2BAQX+Q0vngshwLZr2uP3cCPwHVvC+xYDR3Yn4sTYeEntazJVczLS38O5ge
7d9Z70HKEkI3pVcj/BfjRKej9klljdz3VSr7wxpDhQSbH4rdhLRuotxdVzCM6YZv
TlALr6s7WuEqFw4A+p4TUhIYj4VjPElFnCwUJxvxOSE8L/sVVads6Xk+s9mjOzGr
QoM84ylhFTByuNtl9wlMINcKzqyn7cDhBMMMtgXcPViTWPIjiAQNEJQbV8lPGC5n
W82K2pZ07DINEXSTXah5db04cf4bn6UTgefyhluyC6Gu0FQ8gHexxG3MYiL/VJmr
qI6ZAxUL4MRuj2676o9ggj0ydLCsBt4PFIhBjgsYl66enIaZcjQQdVefRpXWj/+W
BwSDUczyifitD+nAaiFca9OZp892QATG7eXAmnB7a4BMrE8oGdMf1m93gRbcWXjd
RgL2nrzvmdlSpvN0nvOqaeczlYG/Vf9PY+WrPCo9K59wfxczrOIcoFHKiQ0dAOVL
ZI47kdzbzT5ZytpfXNKOo/6rKDLcjqVD1SnsFUCYwFUIb/6rCRyAnHRgaNLEXrfe
IYCr3v1OcKw8rwaCIhENWqO+u0tQdZLi+CGni7+u14QXFQILTkIwobQJd9pRtzhp
yc90rsaqPYkgcNNm2Ny5GFjv7hEtJOFF7tMKIfnNGNsXg9WuxMAYjXRrKBL27QM7
UtRRtD0u/arG5dAX+yM+C4JB5iFHn4pYuwoELai6qxv8jSYxpfCZ7/4w04g2vl5I
cubba/tNFpInMzL1a87OcZVNNnAL0jxhtE7XicyfkWRy8RklKoawkZ15cKggmjgE
ljfVDKsVpRxQBR/tdURaAQFMoBxJEwossQesEPwY4blxVBiPAcnOlpDb/HRW7KrD
qzHEtc2CXi0p7qL6BMTRkzCK4YaZSUHpVoEJ0Zat23qmWccwx4hgznFCNTZEGAZK
FcbvrL7UpMDSdLNRLw+ME7FeZxiD8EcpMjtkGJ4us5OxDhrE8k/IZF6FihdTcTgq
e65gPuhZWcGCZ6b8/U6MNx0aavx+evYeXxDpSe8niysszXrZ72a1bxZAzZFRem23
Y7ziNQFhqf59dhLh3NLy1+BSw+jk9N27hqNzCRvXHfA4lb43UxpumPV7pLBNv3Xv
gYt1ndtJzF8HVFmOsaOGcUQEkDQdrlWuI29zQ01wBmpndZHsTwYz9Csyf8/XQtGM
EnFtBkHXnA72atSevPei6hlWNo8hfS9TG0JU73ayoYzvsiFVZ465ZJwLXbMM4l9N
aWWmgKVv3ZQ1JMSS5XKcP2a6N9/SrTZA3WJdEWM04WZqtT99anLt0VvnRfKfoyGr
V84NxVO42+BEX1MBxoiQv7wZU5kQ9KaW/FpAc2d0JNG/SWj9s9tnarkgK8CmBVNE
lYAUjSUlylxwfwU+yMZjB+gTSFsa6Uqg6s0ZA/26EFF38eiAE8LWMf9tmhfO7m9f
urdErJiymSignv2sP0EUEWPoWOvtmGOnMslfq68/QUuL8kadEmT8AhSFnkFolIWk
6gtjKpOc8Q0IJJ0yRIChxZKuFAtPzBA0VzYyO+34EBnr1i5BU/iHNPStiv9/rhEU
iAjdaq/UEluZXPd2iZFhaYE199fzvNxnlDEI0Us22ZXPsgmFXUcMqX5vruKkZdUf
IthZT6QIlpbhxFxKOs2JcwpoH6wrtdt7+ljMq1pzm72oo8TmRefY5HZgLXE9yLcU
o/0ekURTY7NVGN9UC9O7DVPWK3cuZiDDmpBJnAWDWtuSUmxgMXHBZtdJIeFe4zvx
1VyJ/L5Bs+vPhyLia/jxC+KUZOB3/mP/gJs41f15smh7hy/ovDNEZU+07EMcW2Qp
hkXa0LArHDKFi7EQSyRWjeUwk2+LrpqKAPII/L23caeNsK3CHlAibDLnOHjbYl/L
LRmQFP/oII6ZZz5VVPj53iFbPv2c09TFcUW9V9/JFFCrcU/swf5jzICwHTAwI5cC
gb+Gyjc3b3nFtjCMHgH/HWXeB1R4i71LMJmu5Xdk9UKY4lXTn/+lWNMEn8kmsFHZ
PsPuK8nlKdN3BXoEznqVaWOPAz8VFf7nUQb6ID43378x7BOIjSc1liqIk5BcUjuq
NE7zfw3p67Zn0oeEu28PHhBWpWaBBQfqam0ErgK4jnOTYoGKmGpeyI7/ZQ4yk7Wd
XTRCtUZ4GwhmeOK58D6y6xEYzXlvBMxC0R6XjjC1ZIf47/YLqQR0wCORFdD/ACSN
FuG2NvPNxBVRwQJvBU57t0JhxRxmore/xmwSHnlCUyvgQcII5mj+SP7sERMljWxU
rM1zpsQ0u9nJ2f3Ids/X5071Sk+i/uZC5qNVXF1MwWGfU9wDc2PbWh4Zye9UrwyB
XNrpRcDxKXxpTNYBkffcLUYlX8svjYhkq88EcmceLeYLMvCPVKzJbquOTY/bm1GP
0HUT8LEAFw+jMSNkTj2xRrtKZM2Yg1FBZC2EklVmlxrzXQojD35ZXmmLuPtugQcU
FL2pZJcJRV2XCFupA9fn4cKd2c4ia6WaNMdsMxJBwbcf2AfGTsNIk27A9BaUH7+U
xnmXCLvB03Yi7PTdrtss9VBQRtHItcSWjctQP3zOhCyk0oXNJv2RJJMLIo5nay3N
mK70B9oXOKIZFiOA3KhV0+6Mw23APxmCOsCocR8XMfmoReB4PhBdfBosaKnBSI9G
7p2Qr05sF80k7SxkVQkQEAecrfgF7Ih1TW60Qvi8cgmARZbk71TxVcrTxpRoRWNi
xNkwAKcDUn/AWYJiQUSwpeR1OoDyw25s40hfca4AdXXQgIURyPBAxpkHQEy1GE2N
RKmcIVXq2Sa9Yp378rrGjN2w8jHKvfmLTH1jzkdP2G3sMghhzq3p94HN+RyObnQb
vcUM2y3KCyHHdYzAGOMWImeYCQfa8B4tHUtR3/XYi4SGo4SnpTlLiJocvEE3xDso
Dvwlay0yXV1jSCJRWw6Z5GhPUlg8P6dbONER60dMyK3hp1gj19U/DTqNM3Mlz8J8
zjMVSdKqOBEGUbGogw2d+HPWYzEjo2t+JmG+bq35/1XJ6jxXY7KdE4+5/g9Fl1eF
UZ2r2gELN1VibnihYXKu9qFoOOv1bkw+oP0CwRJ89iKhgs/Ib9qd/uF5Xvw9hUu8
CP4sM6I1aB1g0sZcbNoNMd2TG647c5N6voiTX3nCf7NmVjyedwH1h6mfDprjtjNH
d1XbUhz3JoFsDxRfeDamgfXZeiFrUR/C7D0DkMcnsybFT3m9sNXkDUDuc+ouOzdC
rCTac8b0lcw49xbU3xjfQihRsqw5EQagDdVvNqMd1Ev9bsCLS9G83QQHqQtrBgs1
9SdfJNxkWKaf4CB9ltJ7tuWiPMtoq2VDY1iw8zRUR0RbHpcl6k12cMWSxIwaxA3K
4vBu/e/p5rcjjJvaK/rDEg7vLUHJzIIMS1zTFQSI1eBYgIlG6buCmPy76KsSncsl
RBu7IqARGykHx1a5RLI9htYH9OYWPBxNZlCdv2c9/H5/ZteHdrZKFGfWszD+wDEW
dyttaHoH2SpBP6yv0tvi/Xqmj1fAyuRtfa/8LsvdiAW0SNdgp79thjnkrLe+KbNf
iT96b3z+Zdvennmj5k0BK7wg/pkGBFzyzVqqCxn+jfq16xFegx620rgT5m2P9cGc
7xYFrqCN+kZP22FNLvO1M/7JhaeUCtj4cdTiZ+WWhlOJieNd453XVMNVK3GVfMnj
aIMiSpdb+lAeffA6NDEWRdliuZPQjeSSf0c9/s2DGFHddeOapKSieza/6QwTWBSr
CESrHko00eGg2aaztRfFR+QBq8S/RiI2pZQ8vwJjJWuaEb5b0O74M3jmhOFkKjPH
McEp+vlKjKaM3Uf6AuUxG9gwS8isOqnJpG4Xq+MTr0CkZJOxGvoeGTUOs+nE4tEw
IPDdAXgHtbM3LDNV/Izj0G1p8R7MB039Xj/HdoNtlkfD+nneh3tCwqUFRtx155Ev
Jxr0sHavjQT2mf09XTarvPjq1/MNZFM10uWHSAOmbkHKaFXgmVsMv3h1ziS36CkD
bLkuNm+t7y+vNjVfEna71RSsWGPBZgFuulo2EnA5zDX3etVhOxXYZz6Xi7ovHAhh
ZVr3wsGeNm7OFMuGaKRXDjDP4n1TaCrkzEGQ31bGhhFSjM+167roUdM4oX4K5LfH
ADIksEFgZ4HLVw8+Z1SDMON6nwcpgdDdTkN/UCtpKEnTbdaYZtAXF7wF47OOzohz
U8qbv65GF+GN0RGF7N5vmzKSwIimwHtpVMeDIJ2cNm/lO4vuLzGw40h7Z2WA+1d0
nO1UEApqZGrJkW6VQ/GW1WHIf1ZXd+b+cTZBtPw8tNu989VkJA9Gjbdoq8ccC3Kp
qJKGy0xqEwC+iNabRYafaIU3ZbEjqwFa8oAD1yttyscWELxJsOI6fkR7G8Zmsn4g
mlwQKonoXfCU98PGRO25v5xEAod06W36n4YVBkXtGUs5RgNz50k02Lh95ZV69jx/
LGw1DVBQi31qIc48DtWeWbznqrR1CNBM1FvwizezjEDPm9nLM7u71w7y9IBJEZVn
G36uiI918ruZX2pmBy7AZpZlYURJJ6/QZoTTDXEfs8hLgUg57XUo+G62/zvIz8gN
S0M4Y6H9cXXi6rw00MI900tXnxUsIddB6Lh0hIYvJDjMdpfjaIdaF6Tg9qFqZfhd
Q0VYuOLkMTqx8MubvOUqDtMI/MC12DDZd4ZCUMe0iUmZH4oCOwKskpoO2+1wdZPl
rMbVqgd9VLMi2OQxAACWfPHQo7tCA7xfcF43dM8uZRm1idZi66BHcagSzTnTEFpg
0pVkCcu2p0bvh37VTneU3PhJrENgPqhK2WU3FK2GTSvUsS6+iO8w1NC/zemUNi92
UfkFysFtPL+q8OLqB1UgfVpujwpcfWyp1HaWF/glbAK8XceDKTH6pAPt36KNu5Dt
YNnneRzSrBLbE7iDwJlKwAm/9EaMv0OLn+MOxOl2Ky7hEGk5a9blivZ1qZ7TjklP
2wtxlVJNHrOzj2j42EsmOfvwzAXK3qbVG/UcGXGmbDawLsTPWbFtvn/kozimkvcn
L2tmODx/xgJ82g3MVFwu1qkPIE838BFAk1cHTbF/J4jwApQkF69LwxdtUeHfxXEM
bLHZH92Es7mEsMqy8VECtyD6PY8UUzlzrbUGQAlYteoRIAHt365a2MIQdOV8tuFq
9hs7YvsA7PXY/hvdZDb9aW2mOqDvxlBsqTmIzw+lumN6hgO6d26MAkmwU92ss2/V
C4AELFOj4o/oKQglKXzNPNr3auroM4aqNfcGAtAq69ooteSbcQSZ8qQRvO6NF78o
K4Ef8aQQCizm1+9DTMpe93Cfdz9Xux7CrrItrj+PVwGyJ1KRgKB9QQRZURSZ2DM4
WiDBw5JdFn7HIh9IrQFPoWIE92btNXM8pJHEqXrvEAmd12lWSCv48srTGwe9emHa
9ymngj+yUoOXC0YHJLk+VUjWZJbLGUIF48uPSPZgrj860L3vACIq0CDe0Q8ykDG9
KIPv89FGGSm+BO1cuztf9K1Paq36R4whn2RiLwLytjAS8+K9fIxYjsAY5v6nAx8C
FNDvEUqrcXXga4gCwNepANhp2FAb2v6nf2jWkceX/j9ln+OJmm+fyp2TNJnGgHtO
He6Uov021cXZ14JZQvq2N2tOxYxEDs8LL4RSy1PvfcBJiRCZSjct1OAYhs7bOG/A
9TombCvegJq9FPcdZwyNRViBPqRqqYE507OWpGpcsjHVouDTT4yi8TY1abcKczo6
o2GInZX8s9kqrunJ9gdygfIS9JE68MYyqRfaCRGyOD0L9Vrg7NqgpV16LSYH4oXc
C0auHK1dlPZNAskv6ctAjlNLj1S3DeBbRX2FhNIhr1YJ7Lhm8Z8o5u4mq5U1JeCz
8oMWvn4nWGVk2WsNqYOInwpP9uHqtKF0CmmzDCOBETcFYlOZXl5a3k1LnUjupFht
HKg36ToMD9aH8cjtpKVGlYnx8grFM6KRZUlHIhEqxaldaL8w9aV0U4T8wOh4IrKb
gQ+VAtp1sG3jHasfMiZzb6tmXzfvKZQjQ5RYC/VdgMacpWNPA6jABL26W5rOrPhf
5R6I+WWL1xpVADZ0OsA2vO5lX7FZMMv5OYAlltBpx8OddGmy7i9zOFfCFisTRTOi
9Gvau0SDcBdZV/tHJcwoL8YhSpSHt5lFYmwEXcuN5R1rAGI9+rCNkafvhdLuMeHC
5r5aPRASg0pGfSoTlAs09f2t4Hqag2cQzxnEXyRARRsco311OCXQmNNF5PkmrMw+
g504KYeM+eoDd1fzcmvwZ286rUf6AoR1ZLOTVY2XsSZPzT1onXvWxZM0Vcp7gLMW
WurF4olDkH8J8T8wd6QSVpg4eJtmZ9H4mm2J68hHD3GJYVoF7iIEs97JmhdrOxC7
HBd6+f/X9GqaXzd2QJmuqrVzINP8Fc7BnkihCx3vIwEdJh80kXwSLYovaMEcrWZG
x6M0RG7ZcX+Rr4Df8W++yF2/h5itBA3s4NiiODkzMHXJzbPJd0+E1XZdrQV7Syo3
8dDvOvR69+F0NOt+ZIWRs+ZWXxcEkvoS2dP5WYlHQeeoKEg6jPHE406e1SREUthZ
iaIFG/8iPy2U5+oQK1PRAZ48Cyu+e7j0vCkVyvr5n0OF+GtYI+DpkqgIQsSIGrAR
KvxpQYtkcOwcWiKdbL9tQLlmpPFHt0HSmmVpOVLKkDXoC7wrMgXqxgAH5iPpL/n8
19tlAjE6G+JxsT6jMq5LtR2MpVKo4GVz9usxGOmpbQh0K0evQWzrxr7LmYAuIpnN
qqCnIXx3p1OoSN2gaXOazT+k+fYQ8WyclASNAOAQgn+KjxaN6Dwecf7w79OYC3Ct
YEbllIpmVeTzb1Gg3kzTCfshHqT+PAco9X+K9lCPrUtDwAwn8P1nK/wsg7xUe+uW
IcG6VDO+5DJ4tlEXT6IPkL2IMlmnsk8tYeeiUFDq9lAQ8fdIV6KhSZj8EBuBC623
uRFJMmdCQTL2J+szwIp2uTDusjnmmXyRhsSJBYk6QTlYJP54HxAfMzQvCV9cAixQ
13czv2U/2B9FKb8COB2UD8/piVtKfWE2Oi6NN37C/DxZEJM2JuQekzQUuzPcHgea
hzDLxAtAMwajjBZuNyxijeBpKRbreDpxayptSCqf7WvPqOzN+5dCGneMJTIwSLUU
h0kDAW0jRnaZL1afPTH1E8EMAbh8z3vhuVEzqZjrMzTWC3ly+ho+WtQA3bUxQtg4
vnH0WK81GJOg2a574QQ4wn0rWsXTQYheP3Y1AN2zJz313b+slVGWiNAlEhcsGPPF
TZNCqLOgpST7HGBAiuD9lNHAOA1H2I2RuOtvZWZXA4yEOk0V+KF4yjJrk+csbRFH
Mt+QloTxerdvwnD4Ms+NKmLlDQOcdrwMf4LVbVnWwiNgvsKXn8cEWEtus2DsfXLJ
c96URVvF8l2enHIncgbM1T62E2d9ijIXH3YuWJJ5zLDX9sB0xxneuNFoipK7wDCM
yihECfvBBL7dlQjwC/Q0SSKk3tg0rn2OliN7GlW1DBV450ZsVXq2Lipt3xAN3HL/
9Ms8E49M7g8/fYQENUQnmHMjEqOHNJ31aCJAjL6BVDu6u58xIjzMnmdGumrb+OzI
xH9PeUOMpwaIbE8ZKf5/5KBSH8tjQP0voDazNA+jU8DGX2oUWAsT9Y/Iu4mA14Wi
u/QcmDGqZV2ZhactPs0W/sS3Yml1XwV1RrOuTx0ZrtS+kR56xbkBWRMiIFXhNBkO
tnGSJGysIRb0QJwftJr/RAqdPn0b6zz+XlYs4lqt0klOIawMCE2zkUGtm1V/iycK
lL1J+rPm1t6coVfCmV1M3nNMuL/5mStw/L7Trt2qXRlExu7TmmZNHh5lLpRVlqdF
y7mPcEQnMrpNd7vxIQkux0FiOkpGTqfjj/N2YIW7L2OwWo0Ok4bcneomfEFcfXnx
KQS4Ae5FOmqg3EUWt2Ui/WfYDgTFuv6dbSz7A4FZRJWzavfcvUY9sl2rlD9qM67r
2BD+nSBw24RLQF/z4tkzfhN93Yi5G6k1tn/r7yYYPX5NrIwUdEEwTdsdurtSg71v
Q/fZzVntOA9a1zKQt/o2IuPljX99bP9J6uCSlvPCQ71dxfok1LBpStsm9zWcYFmd
+/IV57NvpmmFUEuqLF4Wz0ApxuRGGge91p5iEJFzz6h9IroKVkzLprCYAuqt9zIt
+Am6HZBB9Xx3X02MWUUpL7wSuIKCynOYInM8go0ij/L8UNam3J9qsgTKSp8UvlF3
Ji6YT6wwSrf9SbRXIFKHmNzdjFKah29gz+YixNKMFs3/NqGhJL8F5kEynGnhORoM
3JP/fExSJ/09hMXAd8wvCNzs7UktdUImy62A3MYhO0QQHG8wuv6a5OOpg4CdU9eX
7C/gdAxKKgPlJ+ifKrN5yCsGEnyfSCC6WJ3xgsmEE2W6ZA1/ALmkJFcxtVJ6R3ME
XfjLEdLvVH3Rjq8fac6ZtjJcs0V6SRR1nCxcxN9wPvqF6uQIn6W2ttznjIPOUAlg
snlYAUvqIxxGgpb5T8QAzTmws+n1kYx5VqrEe4nlw/Uq9M37Cc6736K/IXx+VwAw
UsxwKZn+dW7aTOk1pFxhfH6SiS3tfLYnnEm37aNEQj/YjIXAuBLjsSeSf4KiN6or
wOmbk6zeiv52yxhOhCY1mbUUDy9iZuD6+10PC5W9Xqt+Wk/hkQj1dHijpvlpo189
bEgJqEaslPcR7Mr7mLWIWRlmP5uxpRx/Y7wiSVvsmjmTOYCfOm2VEV3n8M/imrqs
LWjmvBqaDdV60NZ1109gH37m62v4CrndShoKIYcPw7OrS1PUNQ3Ud3Wi0IiOYulA
8iq6Ss63sNxPfDxczd0jMZ+OtJbO7K1TrYJywmBqusUhcNV1sJuH+W3t+rdXfQi3
QFfgrmHT+33KQ4dWcUmxWNe3/FknP1gQ4cjd9aSfjKfl71unHyZYlNwSP9l1ueH6
qPZR41BGIyV3Ff9eWq8elVpZ0yJqseyhb8JOSmQX2IRfbc2CnTiUWDKU1UCZIKAy
9hvdJuQOUmc7LzkUth40LztZjMgvX11eK4lRPDDHYkHhviFOO+e2O1ncGQC5/KPN
WsQSrtspZCZxEdJQDgMODO0VXj+H1w98BEYmghGfq4sgcDl1QWYGFOqaCnuYd1K+
RZNpbmV3cOQVjC7q9nH97y/2zbUTtLZGq5RpsjvqECzf893q5Urkq3xvmUss/vmE
slihm2tU/u01owSI8vBGt1YXMjJ2vflRXPqyktpnU6u+cWPCVLqvXiXPns/DDdyx
509IGiHyTBiNoAmbEanlN1xK1UQopQWMHmALj/QLiCVGDCjppiXml5/oXK2XMMvC
U2Q0AsEWG5NtWpAVTFA4VkgiTNDj6ifqKiQ4V43frgfeHN+IDkav+n5kQacFri0/
FD8paWOFVNp4kxl+7UTlDIsYeaHwjt/vtpXwiTeXWog89wutS/Q45Dru+QCW5Eqo
9RbqrDhm7bn63X4vy6OfpTstik6E4DuHdbnxGaDgLpghsqNN2KTAFSNpdWDbBjqf
BVr9YZwC+JIWU5xPJJK6JMfpDNNw9xxI111CY1+4BOqGeXIIfTF0DsqTBKgSFSuy
vLNYOdw7DvjQxGLNxgIfGD1odN2otBS+C8yGZAJdFXHAj9FkoeXZRMMPt7kTd+kZ
ELVAWa3fZ2qscgQfOH3zkBxFJGpGoOg67XJHpF5Hpi+R3N4PRDs1pevAdu62O9RT
J9VD3jBi11FpUJ3M2s6aZ8i/pD07Bi2YQa2bp2WB814A9ZSgbN7M/pikGj9flr65
cA0XZoDPXwnY48C7AylPAXfN5xtEaRajJ5J7Y6s152sC3dEimNIcwvx/HiKWDxSt
z8wQu9Pn6B7aKp/Jx1RZx4kOOV5nefGMc8lmsgjI9oByHF6w9CCbVx4kmBUSnKdF
WIl9JToBchNVgifrXEllRKkZhVBvkP/Ir564d2368l1Iscy9/YbCP90dPnDG/EKN
p5fMTBo1B/c7O/Ljk3jqHFvaNVLcb8SIGGWElZ38MzLsTle95H5dwJaetGjGL5o3
dQRs7ChkQi2C43kTXdPlpHqowI6S+q7MF2Oo0lxK2C6aahtAParwKfsCGemed6ec
S9dsPsqceufoINKFqALdEaHWr4Y8bCamFD6lWlndfS820hFTm3zLv3gBAqyHy5i9
GLjlhC8onKMXmcxiYa2TjOVVemSdekc9J27cEdoGgiL/uE39hQqwxZuH0x0JM35d
yYPoZdBkMaJuPSX4nDpbab1WWZHW0P2ypD56SMfdGVvTbC73ZQhNiGlqdQ/j4BkO
zfncyG0YfOJO13sArH5MkKjWrRARSkqXmHY/wNelMVsmq00wCTrZefd26RNwZHE1
foDzS+jk4WYPlajTPpt8a26c7Pwom95WfeOGbT+ItIbUlKodHBW9MD45x7cpgaUp
A+noZeyrvl9AlhcKTot1rDIvSA7uJrRxkmyBxLF4Fx4I6qRta/eQ6kWud8ahPczA
Ieb74lBrOzxPnloSOSflQrk1wYVJSlSEcC57X7i+/gwDnomSj4MX5SwLHyppg3rW
WdOeEowNISQiDRcBqjVdN5OK+cs9N8DJ7Ehk/1StTgOWUoJn1N/Ez8toSXQJ2aVA
2Yc1xdcw/OBaVm0FpcaQxzjQqfqrMGf/wfAUGP5RCmsKM60xwzZJ2RpTeRoe7hSm
uK2MshkHxL5+oqq5w60YdjnPGe1Rq8xx4/0d95Uts0eyKslba85sLEqGdVKujjVq
F68/mUqX6O1NO9MQvxy1MwFOhm+f2G2Q6dgWnhVPDrOltzKHn/PZV9JhqhmBvEa1
kXHTVNTFFN8VQUmFwIs40E7fSqa29L8yqGH9zqAf5fmtBHg9A1eeX6DFk6eIo/cy
OcJ9dL2zQVpCLMWY03TSbzHtUuKImsszDw9pabhYofXRUUQtqxxSQtcXMK1fclhT
Namqs5ru95dsK/nafWy/UOP+0mMRWJgCk/tFkuFa6q+xKTttgBLdaYppPyg4IMgt
Bvt2oVWBhEE2vqzHDUvxIrxhakEGOguIUM8VPv3jxxGexdy52cjvwwzH1fBKw3yh
GaUHWHfC2+Kocx4YqYjcu/Y6bnM29m45RP0/qjNcJSm404SNG/opcZizkZDV4Rs6
1D/GXG0qCF/qMImAiNqXjQDs0Dbnhllj3qatE8OZOV64ePKWM7XmVwilOyj4gOWQ
WVAqmjw66cBJV55LWdSXx8eoFnmpXGwII3wamGWU78su9rQssJ1MYhj6L6x/davH
XS5ypjvKLvPRagsdHK9mZMDCuBd8eaMKiOvxaQEdb9YlKSJHte2f+CDyyriL/XhJ
OwXqnoslzdTTJBLhz5qEeigFgGmnqxASUP/fzkpQkiwQbeWmP85KddW59EBCmEc9
Rwzl08gmnd38u0mAzSQoknKm5FFpHFoJYn7y+PFXjnGzzWlA8GlMR+ROr4jIT23h
CcA/o1XzaBEP0ycE4Z0MGoF3tnm0LEOoMzJgB0r7R2UkpjNI576oNyRcw4fsJr5V
5SENgFYRiUzIXJiatFPSeYfxy3xxma4BfnGiuDDS39QQWP0oj/XvYniIW7o7LKq+
NWUGmFBCItigeoXjY2Ij5hhaL6DViDd350rt6Dunzrn055utEUkkNijl9QJ3OE+W
2uLXkQEq4Nxpw6VGE89kgmBkzvxYA29F95UNJkNUsPYskiR7fpwoXJpoYG7wPYIZ
qZS5ntgckmx+FKKjpfkCzGys58ebtz3LYmII5T3IVRNlT+OlnBEa29HuSZj0YFZe
+b6I6y77ZnQt5dImB8MKtqxsTKeFSkK0rowTlUdsRbOp/fqDM5g6e7EASt7sbJwL
ZsfqGYPWQDdHVj39XHsOzMI8c2WRjG0bN12Hx8/2FpiArvrDJIAmwr+KT0KZYFe8
TMRzS9w/xH+leX48PbDzmuVqB+wmaQWoKGa2j3m7OioVKYFSDKQF/G9xqTPHnDYV
PiP9FYauzL1lrPAgll2mMhU7b6QD2OYJHsHmU60/GDOvXC34esHO+QltbYB8RZw6
WPfRd+ZMgVrJ2azEO7L7EscY11IEO8R1ogvkah25tXk7wxSDSHIfFiezPBPW2NCu
8jvCSJOcLypZgfVV89xd1bn7L+gJa8GGPTnAGOg95GfGAKvqusjzNnX6Y6n8NHHY
afoJttnSpZK4dq9IKvDeQ4p5X1U2GK8xU7NmJN19zvs2GwCJxYIqxKsylcqn4l0Q
3dT+hd1yyw1RwdaHt7sjISgjqbNB5B+LJz8ZGfALRMzm3d9YgocFzbqODUSH5Tfc
bJose2oJt62FsuObbo1o+Uq0HiaGGdPbktrad7/sjduhsddMeQgVWaU1F0rL7Osx
VaPlBuNihwfMWZcLTFb8JWPaU4hl6HqjfE1dXpZHUA/OlIvkG7VfkY0NicNwY+pl
dXsRi8jtNOKWBUnnZUO2SlkXA4G5cKneMgAXI/Z74Wi22u/uvHYS2VpvabW50Dgy
BEArkpcaVkfkgRLcTV2lcXwn7x69cUb3RDKfV9KB/2/VqaLV3N1cPtilZnUZ56WJ
NYDAEdKot+AhvZ4AyYklFiz9vL4TZu926fKAE8922UBcsqEZkk5xscw2nmdap2bD
Xydgsthm6OaA0Uj07ULRI3pkCvuj/dndrkH118NUiNEsNHZetD9lZUR7UCqQarw9
wh/G6TG+A7LY3+A3HFjhFlrWfBM2df84sPoDrZ1BKj45NViz/wOcJn8y72BNvKkO
r2maLnetti4qzptotrstTqrXY38/fvD1Ye6GVVe5Jmpri15fViCqeZ9EUT1I2DM7
N5NqIVzhx439SyxYglgf93Ow3S/WupwPGmLK1dPa97oITnqlyGUSMzMooZ92cH2M
6y73TiXb2HDbYT6UPTI8V3Nttbdj3CXKjwWj0KD87DUE0kDOaegcR1vLvAMLwDCM
qJr8PiMtVHTSf6DEnfcT0mAcYi24wTNuUCrt605as2pMRHuUHKEtDK/QNc8yLRyw
x01qz0kO+J+uiOHcCxDgjzKJAhk3VezmXWy0LTumof/Amv/XWaWfflQy6hBoCaxo
YOOZ/A2J8vV/Cpwjptv1pxvD8ghpjVlGppPgi8+Bot3bbxjlyaeCgPNu17s8EF5S
OraHNVb9L26GHhq3h+FGJv5fvXRLWh+2igCrS+TV237beEzHYGdksfuRdbq/ZQEi
49OHlmoDKqAvzG8OtXl+6p5+Xsr6pkn9+k/e2BeWsSbIlbgxld3UNxX6/tCWEHWa
K9U79FpCaCmm7ldDCGs5Iv58oTxKKvNBEf99DjNS/7KOn1Gzi+MluhfejxOFWoSw
RnCMcQWR6rqMXzSBc8VVGZ+jasQHzoRjhAateOEa4tM4cUd6TU5TyNckZgGGJZIh
drhFnL7659xMC9EbMyCQIRsR+hfLxjdumujtfo4wZPAQnjEE7EqRZ/5tDLEsL7UV
sqMGKWNau4PnDQ+O5gt/wKxhjuUtXk1qeCznJUhde1MZXFTmA5beRq9BG8wu/wfY
wtl6DEdTlnQlQz/Im4Dg9616jjlDF1zCVPGaXMonLaaB7Q8MNEt8yjXzWzwoJCyr
y+HsWQYzsTM6ItqPTBf8n25XLYcpYO2K0zlCvqhwKucK8E2OK6ZcQ76k4svx2pS8
3EV9hG9KytbmMK8VYW3B+VDIGyImDQ6cNOeh6iQEeQC58GG+FfLCdRPR6s2xTjnQ
TVC9i26/6VNQNJm/apP0rUIJ9dVl60bNtY7Q28oosaOUguk+2VDpQvsqBlKse8u8
qF0H1y8/qvSDx6jqy4HDpSbE6iKfRh8F/D3t0oX5tTq5X04ilJwQASJznzWiEWGc
PqOa30jzQq+zfglcZdJwalOUtH27axijG+snOjXqW5029b0c0RdMeRzfCDeXAWLV
HMfltn/2FYsht5VCbNTPeyTxCKkjKucgvsvlqU7++2Do3Ipdg6jo//kAlwxSZsIY
GtNeGBiYQn+/PzuGT+jGqXc8avxW/D24b87aFFyMa6dpgHQ9IqZP6FWJsCqLPxq8
XwGBRPwhjxl3Lx7d1wq0m5GxNmXUu2RiPmpdyqNNCR0a200oQ2JIeddJ4v5GB9On
JiLcg8/0txjcYlWDglhkVDYXOKFSlgevEpBNf/MbBbXnUETvRqZrDUIAYwx535F2
VnPzV3O0V74E7/m1flSAssdOHXfjMRI3iA3qhmw3+hKIQdM/yZYATBi/LTlwPIIT
yNwWCu+xxZzyGSjl8800OsZDRz+L6f5k0aWSym9uUzT8WiAwFzYrlgBPT8GDSgDp
8/GULQ6BuZ+elpd0k6rj39/54umtjcbHTpFyX24alr7qytN/uRklBEvfB3dAl/ZL
Zdu+m7ii8PXbAkMNUKNOcFyKj7q1AmL3pnUXnR8Tu/nEWhRygnTEhnjIwFj9UnuR
Wc2WhVfTa2+OZDUIb39YpTXsgOkcYYvvOoIDhyWkuT4PThxyjv6ND+sf3Vs887Q0
xElij43TDVZrhmo+tV1DyYXDP9QyY/SnuGAD15P8BB3pJwpmEjjkmfNlDZsAz/of
Wopz4P2nXB9mIw/2oD2YAQuBmJnLXV2iOGkWNQAtvOj5i20Os1ETGedvvC9yS90K
926Oe0y3MBRDuTCyN4WZ4jdbZPovFNAVbp/E6VNJDLevzUKqtIm16I8O5rdHoh3s
N03zhnJ5QOsM8fee74Dt/U0d9GWyi7Gyqc6wqG8RVVWBsg1b5jJyduiVX7NjS8ZL
afOXqjCaJ6JtT9cH92TYuTbdB8nckZP9KEUFaI96tlafkdSjmvzQW+Nhsy+7hK4i
IzZuVm7KbXLm80ml5KGZNR8rZs21+KjWBRw2Djba4w7U2OE4KuN4yeiH9vddxS+M
92yLpnwuenLeKMCI6qr8SJ6DNhyNhtoXC+UMbTdDiWY35cPaPqb6u7d0tqr4VwR4
glUa6HHVhNDaKT34hn/PLVIekX0gos4jPJiVA7fHtFXGd48whllwOpop+5gvCLlS
f+i6eBnAxW0fCs2y1mLnkerW0pBE+OPyhW5ZeBq9qoDo0fdXDH930sDO2cfvyGwQ
zUD6ehNk+wX2aJAhv/g760Nh8hZnhy7Lj7U+p6KsiRO69+a2TVIsGezusYh+wyfe
voCQoUKrkZpGree/yuwc03JG33y5osKsIDYVyLJItFoHFtkKebK987USSzDMzAE4
gXjkV2qsA0r63VvOstvi5IZq0LSh7QBMV9atvuh1SZcCCVnB8Wyx0ibOZxypYIrb
YV1qKXollYKlaxQG+J3wW9O2vqhwCjjMF7CHk2w0sgea5XylmBuo0qne2I50jS5F
hkg094EKeDp0qyJw9WnDerez0zs9pREoD3w6ks3trCQHTQHA6rM8Jfa03ly2Gv4K
WNPUzsByBjd6VCVlIX2UF2u10uuztOjWgEQR/fumJdk9lk1kEynWBYFHpl9sdsTU
Pqx0uLQOqWUkpM2OZ2QwN5XzEkGr2gxzDOZvLQYOj4bR7oTDOoZfDX+/RgQUmDF9
SkZ/6GieEFXyYcaZ2LF90Rw3aNitHhtUglSvw0P3m6qQKT9NrLBEIlFD7liu61Ir
jlfnrJL6VwoDpkw+I1lKrg11cSkYsp/cmailqQb62gB0ot6NeKNwkFDEf/stPvp0
2xXDgULd18kfptHf46ZPop1TutVbG/KkLVOZT48tCiN9UVPPgmk2xvhVp4RLHcam
4hxNW4EC8B5D9+CWgEo6j83YPniPNRwLf9AmQSqdf0T38hPov6zmwZP0tp3fAutR
Dp/UXpNXpyjJv8GdBOQoLoHTJBonOlDmniVP0A1MxC+rWJ9o+N6Fz3pSQRwN32uh
MtnMnhJ5dS3E2NzbkmJPMZ7FLkeF0VyWmT8bslKWiI0F/Iue6uvAcLkATWCpE5pL
hZYV0rMQHANq7TBXzujhNt9bJwhYxEByB7sB4muSxFD6gmnby1G+WwvUfJ3yNiLg
AbG6gTqr45wQsCltIYwbAZpI2nbatxJYCaOngYJGJYxysQAwgggTfflPIFf8rJqQ
7VpnS5dHz7Uf78kO1BP42WsoWljLLAgrmrglUCrac3+GqjVND0sUDc/HIwkr6s3E
rUqXFSDRfSEtLG5lBcM4dPg+kB8wVR38Po8YghCkpiEW5QSUpTCcuRDE/82mRpK8
JI+E9KnVI1TYMveaQv5EjI5Dy3c0NUyHW0nIFsMt547BQPmbsGHNlRnv/RI+7+Iu
g+LGAVkv2kRQiF9z/N/kg7XhcmSHltGyaWZSCdJQNSH3qPxrw4cOUIqDqOamklZv
lpe+YA2HQIY6qQKZotIZx9dn78AgboaQkXaxAm9oPM0abOXfMByHGV5sXQBwztiW
B/HeyAsk07E5GHuoxq0vGaVTjwS9QVP9D8cSL0xnXNE/UNNJLFToJyjLkvyKyxPQ
5EGOaFtA/MbT5bx0TFFRehD4KE2l3KIzlmjxf1UrXwWJFNC+JdrrdeGYLA4G0Kx8
C9X1LnrB+hfOyN9XZoixr1vvda4Yx1v9353ukOqTPjJIvBKV969NlA6yLYY52WMY
BMLhegfvFw4/lvZi6QU5fT5JNIzluSIcvT5VE308KY1dey1LJB8qFPnELm3yjqP7
YH9TxXt0ZOGsCQvqtCq2mcg73TLGLmo0OZcimlWaAtIvJQTkSl/FJ0goqHJmH8Vn
3KSQxXbi3twfUE+MojmKtwSarNnsghC59V5YxUKenl2Wn7nGmmEYbsKEM23ebuim
pgIT6t+JtWpPRyKsY4e+ARckS+hkxMbpQjucyO4nzgoYv3LXV7qySI4+jYDmWBNH
rlkR6gNJL0TB8eLErpOrLshOvOp20TywvI4LtnSvrS0e2ska3IFB9r/DQzvfELgB
3dvFsbyjLjMK92eGQgNVsOyKgVHSH3eyqcPeOy0n572a2JVBiwbMRRkaAF9s/Miq
xYlrALD0MSAzBZ9GKUQUkNLuNcco3cETPv5HNuL2W6eMYe3Ga4ve7Mx+KhyjCPDc
8N2ezcyzo1xA1SJjfhq7i7fAFnsSWcBOeSvOnMDb4NR8fMkGqpEQOOTOi6jhGiBD
8gVMABNWKQkpJBJ3lN5A8G+Je6qjHAxub5GzLYeiadToMG12bGA5/JuxZPKuHpTu
zex8Cvs4LDbpFkWe9X9lH5eeC8kMHhhxNBs/fA7NOLRFSaoJqzgohoHHMUZ0ZdYt
5ddCRv7Whu2SBjrr+Nwj3QSSRw+Vuvvru24GqGTK0TwRBOYX53eSddLqXmoDFvpI
o9bSFleplYkcEs+SBB2izSU0Iy/AikLMHyssQxh1nI1LFov1aKF4Q4f5VAmIbOzk
Ga++3rFNP0my387oZ7BXdXJqIJG8q8iZzJmltauD4SNpuRJ0OK9VY/C+3+Fgw0kl
4vpRlJXQuH0NhifDmudbeSLLMAp10tEYBwvPCH+rUsTZGD2C2oaah1V6q2uWS24D
L3NWy509KWz2GLVaX1hEVG9sMrryFyWjEwp0vt46EOLfLjvZAE9g7YSxQU4PIZAG
JEYQSr8ZhPiTBhI0ozx309JoH2roIgejwbZbnT78iVbKcNzoI/skE4oH7mlCx9dN
Q3prfgB83HjrTsmxiqGLWoSEwI5JGUCeDsir9HbOzwFvwx66YWv5dURVNJjoFzNA
yMe/bNBpXpSddiqfDPXXPs91Q4C+5WXnj0eq9NV/1ktJ3LUnvTaLj9itDVlWZm4I
jEfo7xPFBbI3b6UXIKJkTytAy+Vjd7Q5fn2Z4/1n0btdf7v7mi8rXF5O6EKNr2dY
tgIBh6k2aZcqtAGqIwI8bn+xQHi0+uriecppZzY2/pFipUR9mcKJl8FgMK/CA+w/
TfiKb8r67B4Xeaux6g5Y/gAh0nJc01fXzU/NsE23oBHP+qC4P4PkIQnZRbQDLgx7
q6CAE7LjyJ2i9JmSObd5nxlA5bFeq3aJtAo4+m/oquS+KyX4+4kwwaEzAPrSzQ4c
WVqsIDQR/7HplmmGm6G9pCQTPszRJER/k8A2Z3KmA4igxslgxmiqRGSGDccxidWN
djZbE3/Veiv0xwxtoRWA8HgN6m8g4N4F9rh9Iy4nntJn41nSXwzP8J+u4609rpoj
axLzAbXxiU6zjCzk5UCQ6ySjTCa9XD5E++Mnv8/nPro6Vgv3/Xp7dixfmbE0KKH+
QCZ4gDFbTc3fLexrJUm6Gv7TeSXbVTn4DNonTTbpCj6j9aXW3ZrAqujjZQ5QtNnu
j07fnJPCLjSXcq/uZrgrTTJJQSK8Lq+w/ZXQOQM9jL/b3mbS7vdlbDPrZhZNyU5J
3ltIS5l4k7cyWKS++Zrl/iYe6hyH8jNzXDbZxJHa11HMzUN9NOVnlRYK0joUPUbj
IimiakdttTI2TRTzFr0dhszHbrMi/hcfdZTyrUyI15+BpD4JaQEw/NdiGSS79xWC
QYNl7UUmD49ejPTiZj156SPfiiPC7rY9PAWOGjge5sykmTpj2Oplng5J42bpVeQK
2GwvPphgSwYk2yMUNx2Lw1rvV7owhPSvawu3f4UZvOHTJmY3BVseofDeaIh0mwNK
VNPxAEa0VouJ/9fwGnAz3MdugBDww+XX+9T4ZmblEfiHKLYs0G7V44EztJbOfPyt
dNVGYgg9Ql1qlMO6BO0AoZlZsv1EPwCWxKtPtU890ZISSHRLQdoAafdbr3SagaOA
9aEAy5crCZl5Zc1iySr6EpjQEUk63U+qU+22ViIq4YNhIFwzg9Umu8E+Ya+/fgtP
Iyh4hUdJ60shqfVQmobtB/coaPe02gOY5cUoD65CmuMkhNSXGlyKfw8rp345FbPK
zP1Mi3ZKc8qHJ60LnlK364fBZU+cePsfD/WNsPHBHKhrrCH1FHPMPooPO18jyBt+
6BoktRD0KFNUKw35VsqwtpYEMfFcyt1zSse0xh/biAbz8l2K/X4+IF6fNhbrvnp7
zwjHCbGu+OIqS8mxu/f/jJxtxfLLzQoSAHoJXgZP3ysxK3bXvzsSYMIyNy4fQpvv
79eDrw9T5BBx+4p44l4nvl7nFdCx6WPCZ6ED/QuvGWhRoXWxfom5o5GosPdubOEN
GdL1SSs6gSF6A4U4nmLRUOscC25fRwn2hksjlN3WVT+bdF5ohEerVeaBHM0B/J77
ergmao2ty2dEbmqExy/twhCcDcikXgMZqRl5R70IA5puQ6YM3H7/IeZ8+gHXjeOw
g2WkYvz8H7F86VFAFmrTt0hHc2Br0S+ry/M1RyVfQ0zdqLrrRRjPlK+KyI0uLKco
E0mxML+8D+i1AiZGw8nUBAxOUQVx1HP7IEe1AqPPjK5tj9NSbwDv7d2P61A3UapZ
oHldfUjPNJDux503ReUxA8SOTU1DHCmXTtE4pZpCi7TuHlhg4G/gNtZSu31f8RnE
IRR//ShDDfSxyfkYCfKmzFZTWZoi+n/J7F6q9NmCxHE7ninHQdyG9Lq7FTfBuhuS
IYyQbJjgFSN8nRmJspNord/7WRKBbvAmCar43zex6sh2Xw0S4X+Mk20V1FyOMmLN
Mkjn6eHXtpsUeHhmfyrC444nDhtnxlld+4OPNPJlhVw/EM9Ly4X4IBxkIDsTGywR
aFTc9hx1eFsYA33ToP7/K64ItJLL/YTsbvDeStG/vYdWUV6Q4RFPe05xNg54YeG6
p2jmZ4Wnu6Tu0gL0R3y5Y5682kbGo1kNetY4Nsw+80wBtJJGgqy26/ODPkACvMOs
K/IDi5K1Wxj3eOKJq8WmLUTUTKu/xVERaPh514l3xeuM682s49q1A5kG8m2+vAys
PBMtkAKKtZToNpLEpQB3XuBJJsCCpch2y7Lyr/sGBJnhO1oOTncpn3pHupc0TKCh
s6JSMK5/2M1H2hbMLdlJp7A4yE9YlzyXJYdURKRnCdMDTjTUMs+4oZe8SfM+ZnYO
AtmyXzHp+rvG+zWVq90He/7O7fxZRcueOtQFYq1TKjbi7327zbrLZt7uMH/eR89f
7mifzcU5PcKHelB8es9qgUZ+tpxdGSdu88IqzR58NtL9ZdXstWUCLyUqsA4Hbmfc
DZvymuJgGxftJexw7t2kC79uQf/8kErBrbvwCsr++lOO81f2qv1NT/ew/hdyoUTA
OTuN5yoApCwhZhufzBL9fWgmUQaTbBmA3Mq9GX2SXOzUm2gz33y7Ur9m1lBj0zH1
NDr2oI6dMouqidd+7JXV7NmoRxBBSF+pfCLSXeHuIhd/i55/xK2BifRhuZYM0y/x
CN6qX+fJwQpoChvcTOXU31Unzx0gShNWUg3WLzzFP3t14jUarEtHkj5LSi0SuSSJ
by4YKHhc1Bc6puRr6vRmsnMlsdYhMIjjggjaE2oG2MLvZxE3pz1r1VNkcNL9PtrN
fyajqJZcbnaLkwMbb2jgnDUz6TAC3kaCMDFCU7p5+fdcSfiqtrwnqXMVf3orsmdB
ZA9RmEOoErVNLkcnsNzxGWNZhS2R9OX5FU+Yrxebg/w9zWNMogRiJzaMJ7hFJUuq
DzbHNqCkeVjRC7qQgcde/OO315kekxO5ImhaQJ47d7nA9g9yiOTYQoCcoXjr9QRW
h4G+qy02CeaDGaBMwwdaNattCNWUcTtCM7Frt9maNkVEfWh0hpSFkL/g4NgerpXJ
/43yP3k7S2gwIuBjNJXG7UsGX89LDY0j4ydDKiyN6rMlQ+qcaE3E2iF+7V+s+ECu
HLTpS8C6O/AiPxKDMkWD0im+6ok6OBfH7aa/dYrskGBKSf5/hWkarbaKc0kkmN/g
wDTTg0p+lyXkO5GhGpfIMU+Facm0Rg9dEFt+YamKkr9ILdZ69ghD6yLdccq8+dDK
ma1AOuE8AP4PBeIH+dvsVmTKNXusnhWmgZ4EaUqRBgRUmYQL8plFdi95ymDNEVOy
8rUeqgcpZTlNFOwA3Q93QU/XqF39d9G0xOhbRHT8tAK22Utwii1DsFCmov9imYac
h2MtKi1/IiVjej4ZjscBJOwekU73Q8TBaLQAYGUxVhLyvgGf5TAHueNrKl+o5OmV
grZfxr2G5houBVj3Cx/MN8uCCBE2hXLEqOEM60jsFrysYDpK2rFEYFPACWu7yecw
MkA7+pfkSdEQBHjBk1qSO84IcTOnf4X6x3Djee+kkTdhfV+6cHXNrK6B80JC4LRs
ej++9L1YmzMrOavTSHZedx5fpufZr2ZnATZfcchT65lelQgKJJ6W93IDAwIbqe1+
6ILlwh5ZZOvGXKmBIsVBklmDGiXYNxZVZWnMUYTW+YndJbjptQ85RjapAdlSb66V
nAgcmOffCwxa2Iz7pqSMC3TolQXvIpS8tuOZVcRF+WH5qCfOrAI1/zOz8Hv/UuxV
ECS5JJKbMuQGairciuqjdAOVAiC/IunNCpeP3pdhJqCn7n6xqiY3G8Wp7Z+J8eOs
Z+d3a39LxwYCZBubPcy02O/dP11lIr8nEqF/c22n/zEsHLAdgkoQhcgmxpbkBaik
NgbKKNz5YA5KbGj7/v+fSiC4egFcEcLdx+2ZMaJJ2SKz+MQcm7TWA0gEmfTm7Mf8
LV5WyfpPeUUvYS3rMZQ8/qoFb07Mz87E6ChQMEG7b4IUlKAQcf2wxp34A3flcqJa
/eFrzuVQN2ObOxfzIottLPXVbtar/ntbFahN2tGHqQqqEKqas/rahWtEg5EZirEv
d3QX4Lph8DSXVM7y5dmSqw/SIihrg7/DAZH1WZIIE0iga9NGEWB7KRC6Xgxzs2Bg
6H12p89/qezZAu4tEyYiJqRko34T2AOuWtJBrzLs2BY568segpN9WPjnkoFc1mNO
y+KGlOFzPENDm/YiG1helWJ+b+V5r65CM+Ka/TlMVrjeLmKsQTSVK852+yM9LJdj
2J6t7b3WYaahEu6zQ0Pak00N4EfCdczDFJbRSNgekNFJ3o3PuX/hGYsf1sIq6fgK
WYmT4oFTVrX7L4lBkoXAgbdEN2gQ0U7ijCK4mNYKAlKnCJSBYtVLQghQtj9mgQf9
aGesJMndDjVHI+3EyaUmZD9BZAav8DB3PJ7YOOu/DmtdgAj/7W61Cyd4885Qu3Cs
PdG2ypf3bpovy2COe92sLLu7t7aqssgsR1LDHgAjVEUS7dAwwsDAL0uWTp56shQg
v1/sKn+nuab1KgOb2yq2jsKp7DbOt7/Ocvuwkm2v1xkoRk1GYWX22sUybN5Pia3J
qLAj5x9plCkFgUubgw2dYjnbFsYZBepXieVKjmqOGeaARfSBDTZmu6UEPwM9ox/P
JDW+fifc9vQqD/SbVQ8R6peGIgSVVjx3uPyKXAr1+v7YM/+sEQMuV70R53DyuUWH
RDuUBTrlo/QHES9npE27aljEu7IDSLQRtudDWdxZC6Rs3KwevWE1z7OH2GIAu4xR
36Z9vInuuP0pSA0YPLQUPy6cvsTl89wSXSXw9RT0XxF/lKBykJKTp/CC9Jy4TIrO
Wa40ah1My2qZrrmwS92bN294cIbSEZ596SSww2dv713PL9T0owt/IQ0P8JIUQjDV
8Qvtwsx0Q4l1HxxP2MIthfMpzUY0HbQQz7QpE8Atu9oSFa0sTLOyFssfnLCWCB4Z
CYxqDiknW/c+QI9M0zmzsOHeTGsdQg6ZAFw/exMFI1Eu1R1i5k77Bj7lAiHQCl5R
T9Ls3z//r2qWay1PvAR6o2lHuGGbdl9LtcSYhC8U1bBORmZVyE3b3dyURmF53szZ
vAnXx98IxhjMaf3vtxzIQEvl4srJ3sYPUb4GmEXM2GrTR7di2Gyolz+U+jmYnC7R
g8E5bW6OLPsMUBJSLKNyV5g4+3qgilozOA5n9HQy0/NruNkoUZTObHL9HIyhZdPC
AEwYeSNPvw6ofjugQB/2mBf8x6JoP6+ILn0x7SENdnwAKuvW3a2jzFp1CJQma1vT
SXUPq3npFB4XcUMWdzhfgkeu6g9tQ47BXneheozGgae9bH+27eH2WevMtUSlTP8b
hxG04NvsGjUqmtXEEiDSZGK6fWRNu0jpuaQE2FP1YjWducIbgqDeuMP4qu7JFscE
l5ko5GMEtZ5a9vUc3G4oP/EoLYFvkZnAppQyNl9y5bGpNXkaPKtFi1gq+hqbCxxU
6hn6+NXg5M00gzZ1z+UoruAEriKBOXqR/HRriZmmDE5KpuPVbdN6io152yHoToKm
aT9mpMCB3sJC93mTiEBVmgaAhZ8DStzHsU5o/oKr/+VpnIytzH6fKevOH2A2LnO1
1bFSQ2h0kT2vKAWdrBLuKynvEZr9q3so0Wws0XaH3Y1JEl2qD64CbnlhNLSGPnwz
GcRdP8InL6Fz5mv3N9+4Px9hZiYNKvscjYsDDEYtdIFpPN34+C3iK7S7+hMdkDyd
MzKZGdXLYYeQ5ss/cVlUfxGVs7sz1t8NMZKxNwIgQoqizvRpvsapiZifiBIjSIUx
KCRWvWUfcN3avs+2EBSwYjyTv9ujFRuLT/X2MslLp/DRUhmj8ez3JSLcb2f0Tawk
DeSNmXd/siLWK1xue30ujg3wtpWICFks6TxyewGFYJmy28sWVHFfeZEWVAzbGj2k
/VD/MHQtUhTi9BU4XbLuKBq+FYgjytcI2cxa8nuhPqUEBiZRWdkxUXuX2jXwNZRL
IxlakprIZ/lTQpmRVWS7YZD+eUFaCxjgrOxlKfAChRYEWbVdx0QC/EDkdx3yveKG
Odgs8+PaD++thBbCxGl8vs+WYy+ppNhk27IvKKfisX7W2K4wfyfmJoIDLf0ADg/y
7KF8twyd+ImcuFI2+iOQ3iyeE/ERSDD74clLR4Mj/aeFY8PmiO0WvoqpmED5GIS8
CPWKg4CFjrPGIGQk+gKXE1ceQpU0tUM7BAHDD47QcP8kjBEPTeY1uinPmVbHx50f
RdY+iCk2biQOj9zzcVpuTUOMqthn6w8g6lcssvL9kJ+bUrUEPfOJT1/tZYlhNRBh
andwl4WgKRH5qn0VRAl2xzalImge9PM6vNcARC+hulyLMNyxJVPrZaeEOBNk8pfS
jfDGJIpp87tefe+ErtpWXT6PmPmTzVXStaJNe1kQIGqrywhMJXoZyhVclhSfpiFC
BZnT8O2Ik4CIo2OAUWqtD/qRl1zQRuEi5Mc5biQO0OFwvtakWXdNUhH2Svh+6BwC
BiE7koEVFBPIo2naFG7C3Kz4dYfcUvlJMWjdq/R4FeLKcWKuaOh/QRMAUGZ38JD1
8Dm8mX6jf4LfhV0hTZnNMCca51c/D7N/jYZMgNLGYxKIVHZtHeCmZV7WDAgeLQZQ
Nf9j9JmwP1zw+rx7r/KG8VcCPEUcxceq328Wg3ApuUW5Bu4D13QI/V3pi4nOwnyJ
OjPitQ/Oy35AIEsbAKXa7Tw6EiSYJviqwrZrw4FIuC+dpCOxrGc2teMjDUCZauP2
1muBpvcdwW1NKQn3O4Nd1+mf7733KnADBwcgasMwkhc2Okb1ka+uO3Jt+JIJfPYy
HvKak7GX13+BVHCbeHnu08N5pn8XczbnA3jq/ZAgZRdlyFqhYdySzWC4QWzgJn7C
v40rvARuYXofd10xUZKmFbjeE4Jas29A2zw7o7+YLuRufliH0k90fEK1UUtr0hi3
K/h1A6xeR0whB60fDl6qj10EGknZAOaj0iMLvB6Vo1p5/UpKJrANk3dlKc8IhvxT
6YDo5cmXYf50/bqGgF0ElFHZYC5zUlX1a9K4brwz1XN+FEHeOCflim6/iMEFx76P
j9dfAajrjmLQgM1cBv1pdJt51rCu4SRRj2yR+o044OxrYan7NA+aMdw1j4pqMri4
gTQ2OSMFWN+bUUhRiGvFTUQVSHfaHsTa8KznEwJRtQboKWvrX9LVw3iHxFeAgZ26
wptw3tVOUaSDPAzejNcHr1px0GYYYkVEhIi6786j2zMTqP7cdbFmne2gpeYEnZCa
WCvLXY5dsbkLtpsvk5TwhD5H+ZDIx1+974Q6S/pzu+NO1TAJSFSRH8jbqMs14jt2
DSYMQ2dkwWaeUCG1y8LhKnLgCsguYrp96pTGMvUxSVk7m3fQx5uF1t41uFti2xZP
+JffQFyN9tBSOHbE7KMwJR8GHDzDUOfdbzzQbxTFyZjBkH0rvWGnld5PcMAW+iIH
3G8aBzg7MXy/MZNTo55RGs29FXav5xug0y1ngpdAJvolS906UHg4x/btx77o25D+
7flKTKyfI6STaOQmIr1J8UdXbAKEANKjZZl2Yr+xQIt5YbqcNBs51G8wrkLLGFVU
khnFV9cfCGejWJJu0lmqfn6k9oU3jhT9Ob1BVXd52yeqTkNj1XYkLH5gKSe1aUzK
u3wGqLJnaJGvsN4qZXWUZKHRhNft269WHGIb2lr6YhT63LlMdXtcrgSeCXXRRdsZ
CCROGtciw5ckX891fwB9OjxCythghq85Et8S6Lfg2lkNsdgzYPJd06aWM46Q14Po
yQSjncPcNe1tt2sRdbwjrg1fXpHhP49BLNJEXgA4WyPjyl7Ei42qJ11JkvaPRV9Q
Q0sGwNl0HGNJdwd6WmZGdgSn3ofW+4ftCdcYFomcn2wcndh8UZV9xhdnFCuhV7HS
flBbok2cwFKAJezbYXNZLyTFyJKKL2+DK/gv8UoL7Rvm+S2M95mEGvQ9oRl2VVGn
yzG+tGYor7Z7hLTeiuh/jpRf62bIxm+qy4ISkp0RKiAVSPsXVjp2ijBVBJyRO0Ay
NH1Ftr7L6G4jZEToMse4y47OdTnqRoystfP4cqQgbEhgwd5Jh8gpdspVTdExPSh4
m2tWFTZLF5htVIQuiOBYm5lTzGKOV5BRdu/a1h4jb/btX61kHYohHN2QOnR0B2cq
vppNo0IFs5c2qWP8CRT+7+Bmys8MuJgbyxFeBY0uH4mCDipcCJaBQNCuMBRzfv6R
LwmsKnEkVQE2rzWqNn2GfcNJPWVXOzgX3945R8VYkRFyovDDEoT1h2XjtrbHElRz
j0Xg+WHFe4pyWZ3u3xgvuw2Mg0LmWCphrGDLRuRwFyVsROisPLn/Pbu3Ssmq/H4r
lEWd67sEMFBl/iIRJu72wS4Wna6tHEtmO25GmnMDPXPoNPbU3/jP4S9kYgt8ZzvC
FcqMgzkP/LozbR2akt4tX78PMkwEMX98Hoj7Z6oriqU0Upln1/1O06a4A/Cx76tX
PiBuUwc/07giiA6NSZSaKdHBHEmaDsJvvMJ/WCdbzcnPfTdIlnEQgD5qlrhQ5afm
gCC10EEQ0aKRgAnMFiQanWOUAaNG8rCMxl2Yoch2YPMpZ7f36zbDM4Ojmr/7+U8d
ATaNnLwbxZGWcBppdGKsgP1Rk37W0Ewj4xrBt1o72yFCnSUBEX+O9bAa26egpzob
G7SEXOROcOO6BVx2QMl+OLIxDLRB+YjTGKypUdX80mSFuO0tz311K8afaYobdx4O
a9g96GSzdiVIOvurHus3MvlNo6JjS7wM2O100ckYkHFJJrZS7u7q83XwKzcViHqw
w09qr7cB9xQWfbc2hU7lUC2JtH6Dmgev2TgIMA3Tv0ZOt7/3RZAL747JEGAyJ+Mc
ybxiOdw9QU9H+K05ddx407dAtNE/vTgrPPJhTXt42HE0J7yU9Z6GwJN7EskI6WCA
ikz8E9nZiNThJAI7sr7A8u0ielu2W8PppsgJhcbzAIGz9hI2o/uI9P8LVGhJwqdG
o+PgRlI1nSIuyG5+64sX0wv7tK8kW7zmbKlD7e+KaD18cUtgYC5zCXJnfwelt+r4
8S+0z0w3UjhnmZe75nxpYfXuizuc890ZdglQ/6TtpFuz+VX7rhSfIlV4ao2ByBfE
R6TN1604ZopXllwdPY5JFBbNVrKHne2HGusAJq5SPAl4UygGmLooYZYy6QcgTRqd
UjXafsKUiFG1ggdae0I+E6aFb0aVmHgMf43XxNyqEjFUiRyOmKulF7sN0D8cCRx5
osHcJchsuP1vxYoImZKvctlGHVkSqC+7xM2gHjSGcU+MVzHLckAayomnfN+U733i
C/HeJNr4q4sQwVLdDD0zW+KfBSKMfBa8Ky9pMC426Rot9Qd+9Y+sN4Z+nLdE7GbI
jD63zNVSxN0xhoOw7P+XBi3BTNEYmhtqWk+sqWmSIGXEaTQUp7TFK9zeZci4XeE/
MoyIaRWdb33Sta3iB56FNuDXU7eopXsWHvlkxXDTuwvyZDHVtWKShFraupdgcXvn
SLLbaScu7s+CnAulNnV5yrCOlSYHeHxU73Mx598WdtOjmzPJYWwk/9eIU6QpVVxO
Tk/CSjVcLSf3O9ESAfTPhZBSf9WtOw124m5RQRXEEyn62rL5WT3R8ANDeH8n9SOF
s/6XIFvGdPuGtVD4cHonw44m9Phyiu4El6//ssedc2HBC/XLiDIW979MleCr293R
3ajAq/jDmBg0iMIaS5BGrLAXzcAMkvWvs271JMDlK2iDyaGwtEqFJZu1w+6utO3S
X3NeEPqEBUhBBQqtnUW+yWAPwl46BlpuubDnAXRrH+z5kPDATDabOZKR2r0Rm4GN
MkyW5bgqxqa7io67CMiHwcVEMyBUz9Afg3Y44aZcZN2NFp2MBWzA0GmInbCFgadU
Xysjhwbgcs97d6eRAvy3EE2ALypEzeqnhaZE0w5ViwmdkJAOv980Xb//rhjX48ZC
RWwYxN+4DbX0fyKTYhs22wowHIA4rwKk/NPIEd/ss8IZLqSZbglWkqcLeF1rKVHI
MUIM0OLmG+/6ijKqqfz9/UrktQBOBTgxL7wzoThcJYgk//dhH378IIR5ia2DPkE4
6vef/BnfLyHonBXGkQAzoola2/1ohXlGt4HeoJQ9zdLKliR4dwnvV4/hjJ0JZRMp
DC4IZYhQFQWye2f4yziT4yGyZznBvfL6wZPxu+FiUnwLRDQbGHrbo8AoVAJqVKEj
cOl9uzLS5Dbl3WlaSCf7AwWzuOPVahdfLu35vpCa75bg6qguNU5+P0QiPL0D9tI+
ptFIDGmIEKKNtgNcETkB/IEYPIx1reb8LwgCvMRbGjWiG6TUp3NY1vljSUFqNgJX
wX1gDkgK8Da9akPR17KccvbBclQh/d2Re1XBOWFuzHgzNUNm5yjT20KmUYABNSVt
xG4wD1ZI3qosLCyamnsmBet6o+BmSGlu03gSRgKsPpsOkSrQEpXEJBS8PaZKa92R
/lMwmo1NyjCTNt4D18lV4AZFI0dZUolvB5Vit2v/7cKtd5P97JeOSQpwYdVzUmbP
j7gU8cikY4XLKV/ZbtfsFUzEJ/rWQ+NfXsCKhHXb/lLbEdq94Ho4BoCzWmjwnANG
OD5F5Gm1GxKEGjrnrbDg10qpNZPqlp8SH4OJg7MutYgiTD2aeoZ3vlR7GNkFF9sP
Q7OyzhXytzAtm33Ngxyr2O3rRXL/grYExULhxmDSbJKCeP8HKO+0vVvS20+sqgwX
oFexEvUnEk5TUgafpOqDnvEkztAo3EDP3u13ZPsB9cpvbf9FIkMc6eA/CIwCM3y3
/O9JeYNdbt8sbGAKgGp73SRzgxY6VfDin/WvGWfGhUgj3HxP5UlI5jc4GTVZDXDA
SNos/VfkG+D8l0zV5yjPUOia22KcWcfxzvynITo1dTfeJBQY48LlAlCRqWoMDynp
YbnwqmduwYHCD7xHGUQpHDdeqda/yENlD0VJ/oHL116OrIA4eT4M4sS47GEwKbY6
lSJ80Hrh6X6vQFwo3inbGLV1MAhCwbo6XrIWFjE+oqWupbxY35ToXSG3LsObF06Y
iNfVYVIuBuAlrq9TyiaVCuz0ESVAVDrrC6fwwjzRxFQRpnxOtb3gSqetzAinlf//
/sX05wLCn2dM7GMWOPZsC/shLfRr/vcBjVqajBvZin9iMbow2lVvWPBH2kM/6KNd
h0ncz1EPpWDAlU59eNy+JbFjSkGsT/DKPecR0Xk/udbRB62hgd6cYDpVb1N9jXCH
Eqtlp+cIIWe9qIyVIOuQWk76Yynb1iz6CLbBlkjMvQNjuiCHpC0TTA/z5Y5bvMtY
lb4bc3YyE7VsoDBgnxU5QPHine1+ZRF/yuks76uu4+MFN8M6DAaS6NZyZcvgaBjN
bltBdqNN9YrQLIqxBMTLeZPY1y8aCdWIMCsPSFp88CBN6016tyFJ/35RTcKrI3WD
1sgm1V5i7Lj8IbaVyyS3AydNMMnoE8OffLScLYg2AGW5Wt+zdlqBMaNsooGfWnB/
VjGoohKODl5oqExjj4d8eHG304rCGIF3rFHWN2+T0d6VJAj9K4mm2ziKT2fmpI8G
ZZnj8KezvEw3WiDznLrnZjDmTEI68+mJ8P2gvSC9oIO2YlWDYX+gzm5SJpJG3OkJ
NFDFmQQNjJDMyME432PBJMctv5TQdk1F0eEYL1YDIhcTqh4XU8KCEujYI3xNU19H
V83kEnXfycUNktWS8m0SV36pigDyxk3KEvGBBKiR62NbL2rHMRMgj01otVOtSHEy
y8zanqik8/lfsz8Z7/mICP0Sj8B30Cs1sYw0uV40ICbx/9yXm2dGaMkEEXfg6pBz
UFQipI+bkNQweIt8RG18Mk6SjR/6l76BlVK6SEVh/zG9LtDwQLnKFT3Hbqgk51nc
mem35OYi3JWkVjLzcZoyWbBUJIqDHvx2k0ofN8k5ccoHprwPxOX5aStYLPbPTk5n
aonBBDapnt0MBbwFRGpJcWq3oKSxIq4IUP1ZbokS/CiF7MFwhbd6mL/sO9Kb/7/t
A14io5VTDV5G38GApoaCvwzcnTHHxc8VlQuKpVqPWmC0LwYHMW4Dznw/+9RyA3bC
fGdj5KJqyE2E1PykV9eWkroI++PIznMkMLtUcFxBzAHFjUnfESSHz9ctpBduV3+y
Y5koI11w4xT3MelHbGSOn6DUPRm5fs8YRNfQulk6QzbDEs/c2fF43xazuvwhOplq
ZffukP6qPajOJDbDonQtsddN+zXnc+ZoCC0S8FRndQcdPx6P5kLxyd0f1aLU9+EV
GoPgi2/yjlEdqcgGn93YL7ThI7dp9kQDIldRje+udDwcGwL08KACudhXfLewE8GV
wWYgFK0DfYLufTcb4n9XrL8RvTFXKvU12WZdBdaeKhGSXv9oY9Vpqmm/GVoowmiB
13gaeupHxYJntePfD0OdjfnKPUqxH9uw8fQhDYnwCkddElUwsTUqwBzqmu14ksVF
rMqtlt3dfEx9stNB8j+zy1nbfZWVTdOnryaPQuLEjffd7+PP0Hl9fp9PaCgusdRY
o5RFh2VwTqd3dT8ko7VR5qZIhr+WnQ5VvhwOe2aTWAAB4OBFmPFd5zH15p0AZnXR
pTQgegeauGS8nsXq6lH1aQ+Jf5P+6oFcq6lx9DXUSKwZlVL+HKdZACwMIl0YrrXG
GNFqGJKzxcwidK2QN0W06EwXt0bK16lprS+8Jp7Y5aatGG1beH+Ypum2/8h4ZgwN
PVNEveYiMNvqPx6BKXBlXlMhahsOMdge/ZpOh8Xldo+dSD1R9m59tPvxh+psNsap
MOvgF3qswjFPp0M6XcpiYY/Mo9UDuSfFMfJyQrBW48UUkJZGzAHmDVixX6M1Gwwg
lG0xoiWUAJ4ygJ7y7xUAkCJZIcGP7ybfj2hX1gicroajvE8fPVyKPQquxBJhVoTv
y4OzDKUbVYicgERJ53QG0wVt9P21px9DCJSOiYG9O0wmCvjCasnl1lajNQE3aUPl
jnPJApSkHRB+ktR0CuhtzVUHu1teZtaNxRGPTa92ZBBY6WDddltFMcBXwKHrqt1h
VJFkphoUgL4JPJvHjr8IAdAR5rqqjnZ0yd4af94XtJhCNT/YI/T4grOf9aG6ZhLr
N8voQjGQLTrQlT5n31icBr3rPkdkX2u6zTjX0OkWKAbvJxtPWB04oLRKxpAO1hQm
RQoF2kPCLk9+iPOXPd0NUsWTfixjNNg4x+x3npwYNltB54rgG5lX+iBKFI8FRtpt
SUzbkeG23lxOjrtew9DjUcIuFCjFPAUnPvW47AZWskpN9sqFSSQajYfHAhXOPcrU
ue3OYDZoDTXm+4OGC1LgZh0gePHxWvj9Ms9wMRe74CaigIH4xFX9CaOnIiGwwAZg
c+6HULpM5HL88LZvvGvwbH54dSe75brKJ8BFA+UkBshNU+B063EgqIYi7Tc6Kt41
kO3X63siOKzFu8eYqt9MRg92VEmevtvVvO2+EsPnGFIWOBipBbAntmN9sKRPclc4
xgCUDEeWFuMtRz6XTGr7+ECWzLuULROJnKEtykZ1GjVbK0ocplW8I1K9cm0wHSqB
um2HiNORwPM+c6jz5Q2FgspCwcU0Jq/J29U0/qGbXehc3K8uyJm9wQU7m3PxSjpM
YRShJxo6a0WlJH7bYhgIaiCrDZrvcZkE/hzeoAeCOLkp4UNNjm8DzN5E37294Lxi
63MUbZu3UMeSmW1G1oi2kAwHqg1SHsa92fdqRAiHbdm1vt7S54PVw+VNYCPiVvpb
aAJJEx5GtQsYBs/uKesGWKQFpjgfKNc6+hdM/UF93RB9pbW1gQpvwhgX6qLUjvdO
rtHUSj+quTOSnTVP6MLuVWE8Rywz0AKCdFKKc770Uu1UjLqkHyGhP2zowAWugf1z
y8pMjSBYqhmvXydilL2gvFb39SCqy4VarNm77s4cCkQ5ENH88I+KcT3czAnb878N
xji+agIG9XDEg2UTrP9Fe7O8Uz+iw8p+2oD+ns+BYgkmN9C36LegFp4SKhH7W9Q1
jvqSbIlg6Iwl1HhpV6hU1Xp63hfXhAgZ7Yf0eG/wgK/bIpalv/lgGAtMrqtJynQg
e6pxOd7CefE/25Xt13EhHbskqihwlDAzIftQB30ujMNJd7uh+eECEzDxq8LSglCP
2fZKbrxUeultNQi9YkCsqWPNjDwPNtvYc2vbOJCvzxoktgYhoEHDblpvprrdxAFb
TZzQdBnqgwOkqPaFHQ06966QpNJvLFnHz6d//y4FYCSTlWN5KBfX0VcCrYqyGXHr
z2UwTksFmAFVDgkWNnY8A8UNOG/9flZirXKaTJlkTX3X4/5U2hJMEM75Z1z9h9WG
kpG6eMNdCelcywQiGVZFdT/tG7aslJXE9LUKwMrtwbLBQwVOW1zOG2VtM7Zl1vA5
Al3Y2VbXRxAaR9dFmU+/LLUF9EI8YvYIRxzzOGHlmpoA9yFW3gWB+t4X2G5IM54k
DrAGtEP5E2yWIVEFErjME59U7BOlAdqnmKk411d4z3yFIDm66lGgscuZ4YXwGMpb
ue+HYj1/YBQdrc6AJgR0ctJSx2Z23WVyegbNxl9uP26r9mVksNx60yKVCjkX4kCJ
OpwkDSyVKH8KQnfiPyy7bWAafiUCHrvzZvIHr4TVRNlAeoqnsJHfuUT64T6IN/um
at3KfTYaRtxRvOr/k4zwoHLdNozCcuDPWnZ0zOX3O/fWlqA+0VQ+4S58l9TJscGr
H51ELZIDYEkbfL7/UU4Hg/KQfWQBxBsd57b5cAlrHt1ogbn+3ZmsbvMh224TYLQI
NeBdWvrAta8DvbGB34tEXgtd2zy0yq2D27v8cgmvLiKLq5MitkB+gmDEKtmI63BG
aiOTh0rqzo1bUY2vDhHYsadVX1Hs+zVSm37aq46o6wRJfSuspMj/ULF8omnl17pI
FiN2iDqzoKzZC6TSEVN5n6Dt3zLMQKQzLAZ662xWUjHPKM+bsmqst3TcA4pokZEO
HieAxHGyBrp83hGm0Mf+eNY+o21gRtpLFdg+/XsD//oz4tResh0jhaAQE5ZVV6mr
VZ7toM1sLu69n5DhxZFspr8QyAytkHlsXIIlDM8hwKqtuGVU+cF6zhoUhP5d0x1p
kug4lGJwLRU9MKYNzoAjceF3TItCSu9MpNbBQ/GxuGWtIyXCe7nKZ7xgikDaJw8E
bumF4bOrCQXrXnkvXnuBZ70wQFjfDIqYZlLuoASmXN6+zItjQd851mUKvDKgYvV7
9oTDh2xmwqB4ki6Dr2VEYuvDxsppQsoJxLuAsoVlbUu2zKKO6P7WTLj6G3zergEh
VOa/IKr8UPeJmbBBQOGC0RiXMSVeRB05VWjU2fepIFpNRG2leIDlhIqPtQNyY7zN
dcBRely8erw6K73dpUBjcdy+VjLxzjpaQMrqBwXQULH429RilpBEug6G4te0axhO
PWk2IvbcsR6ngLct2MDIBxoTOolKKL9Yl+6R4NLefFQGOCqG+o2SONovg9R1WyyW
zY3Q9lKiAKbB+n74Sb/tGoCRc72yKsUMPZF7lQsjAFwuZgBJf4Gte7g094ntfyQj
x3MxCGkd+HR2+4fuWZkFm/hLY6KNXeoS8uNabVqKVXBLofY6vvO1/QuCejN/Tf0G
QQdzv3gnOVv/2CqcOzksHGo4YxGz+YUPUPCj+YpcTy3zukigWxvyO/Ye5vtXKSiF
IxUlwJEnjxXwIMntPq9gWUVlpWza1lpkTmrrXii6XhW9FCnmDVP78SYcALDaskFB
n+x97PTjkl6Sbthf8j0jmvyZNvWWj5ZldjsfTYx6k2pPt5s8MlDmB738xOoIFrNP
bLJma2YMWuvlcEuHH6OAyhDEyOpTwfrcBgn5L2VHyPLFlNZ5vUocMJ6v1t4IJOUj
VfonxZCAWP5Tz+KHZXbA7olCfC8Hc3w74C/BA+gxdgIS869wodnpDbznQPD+9Bhl
PF5n8Z0mG8vo6MoSoOZ/lETtK/cAJciMdMoTIW9BXTNPh3DTe9x2nCabD+JeF4x1
7F5SZDn2wbjRFp4lBA5Gt4PZSSosOqNqkFKbSfVMyJThTNT4cXHrkuxpjo7lLasm
CM+4vrew3YUsHvFucFifBKK+K8haCQz5kXuVQNVqGpTX9iEiL7E+3FY4tGnaEudc
3tPqdT1wG9J9PDK36Cb9kneyAwrZG2dVYVDRSg+VxgBmf6MgarqqpO0lizxZfajF
hRtE3cXjDP6epSPQsfhD9djWx0h7iqQSYNUeRw8Cc7obffBmTui4k9iEznoNa/EE
TI8yqcnndstFtGuCXQuiff92Fot6v/opYQQeWwvvfnNtAmdujc7DewW0e0UNurkk
i5230vVzpzJmZt+G+m7wGpRfAsiN7WdnPWKdVu/ekRKeymUm7Vmr1DlwZ2Tj4euL
etqjcYb8+LkXxwoq5odxG/PzGteNX2vX+hWtuzkfkoYsJHab3wg6JhemiH8MpHq5
omHQynbb/fa5FC5tqWh37A9/spRdki3RKuHhizEe/c5YSwcbPjXAFxp5k3gVSLuj
6JfHfWbzby0hm+eOIilxaM0C3i4oPyFsAK2OaBE7Arbum3ImELVOywcZsvkFAvAj
vlEzdhheGKIfOofjs8Yuw6ZT3YIG3y+XdOeJad8LElJnyu1s+qWq0wuZJ3DMgweZ
7ZeDDWcL7OxbPx6lVekUcrh896/IIIQC9qnNk0PFFS9VPHAaZousAfUl8H1hY3yS
bwO7Ac3n5+sE3WnKNOWFifDJh64/2Ep+g+O8bqnDpr8MRaT7jEy3/GmUzb24oGwo
91z9tz2RF44G9Tsw8Gjvajw5oZzHfwMfPsX+q1hRlTvvDPKzEErSjbsV8Y7qDq+t
pkyQyE6Bw52F5Ex2zBcOzV6dsvYdMLNrD9VyiiJWVIEIzuqu5MMr3YkMxqT3x9Gp
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ThzlSugganamSS6uSeYlZO5iOydsIOiF6Jz/jpYHIzlJBfHpgf+p+fpaYJTF+LqO
5uEywUXSVgcYG80HmhcExw3NgoTRIvthCuHLbenkFXY+YjmCkGG3ME0/4H8h7xAu
ePmZxLH2MwidiYFb92crlbR1CBzuoBbOToqfnzMf8eE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 25440)
qGYsyUlu5wqpQH5zu8Kh6pNRynSQiTJnqBaeB4+/RQTuhh9K70rtEFuyj9/gnzse
XDyAseMLNTZCdLCYfWEuOE8ksPuelRt3saTuxLd/SgfWoRHrfokD7jkM+eddDaxm
V8j0YxIhcH42GNPy4QEtWYaVfWI4zwcFsl1x0KznhXZ+wE1H+bbFlnughvoOL/vW
65Sp2+1lklczE31xubEMCcgM0poChCturu6/CyjrHMFw9pk6TcsRoHN84v8PLR3V
F8nWpnYjqsE+pG+1rvhEz1WvLj5mS0L9vF7NeAql5FSTPbc3VzQz5gWX504hhNT0
LSXMd4ZTwa0tmSfs1RM4ipBSteYWsqVdPuWnjFcldJcv+77LGqoeN+2fHMheDVe7
vIAWlkU25WLIYY6HnVjTjWdOWfRZdSQtrHRGiqmPX0l+gjwm0CME2ZtBx1i3L1Zq
Rdypn6hDbI5KMYxS+i6X2y4FtZo77ig6diMfuh3IykPBhZF+OV5k3jQd5fWzNvvh
bW0wavjz86yu3w/6V3FlDmNBJulULnhoOC7Aa+opWrsuc24CuqipRzILUSms5Oa6
9PThStSRlfNeCcMe0l+GF9aZJj3IYJw41A2taSGUkcVdcoS0P1VGJa+CwO+XW+wg
rpuoF9qcOo9QiAjKJFS3AQilpSrXohHn3bHH+SJKsA3opBluWUKVS274Z5Wx6LNT
L4d9edcIxWBryweShy0vLGxBkOPJoTWrGqEtxl5HV+Tgmhps1w0MLBHJYZsU8EIF
9FNp3f5c+k6g8g30SEX23b3V77NENcdsDIBkn6+Kb5WiIBr4FFj7t/386S++IF9k
UZKiBCocnyxJ/Xd66g7QJPWPIUgfeBx6y7y8moAxpeQtGUt1qgELWbvGBSsnmDTM
Kfqno8MiFRjyA6BlDCrTjAXPGXsjBvtOB6zODuYdVmpMP8vL+nzJB0E9Yg9mg1gx
jckhqaCoYtsn+M+xl2LbaDFfVU45xLxznd87ZKHArZmSBqJfsen/FrOA8FxgCle9
vjVDlWlFLHBLjJvvmfY47Ez7oFKDVjgZRExF+Mur+VHqyDWwwwAffZ/XiAKZSAo9
miWLnO0VW3xkX5Cd/Z7J5LT+ixooF9bKPTizzDpdlVp67p1g0BdMqzPmMUjkSjDk
1F7UoKk1O7ztA7OoP/sg8arYcGqh1uzHrFI/CneGjrh3fEMGTJ/nfVRLaQsasAMM
ttAIywiFMvIPVBLzrG0MPzkyGNdVK/J4QERHWFXlKdC7elsaEHF+Ydiaaxsxc9yk
Uj/HfT/q9LAEMyddBXWgo2g/XXkeZyBmQDS7LtDbDlhKziXI771HjNztY8LMX1gO
FHm2r1gNvSICwh+xqO0oxh5yaCBF0i/CjHhjwhTxX1Znovq4vp5x7WZ11pC+X5Uf
TMyp/ZN3dTkdVXQ+wNTmy6ADGdu9cZFx/ijLrTsg0VWjlASfFCWqxgwcMIUwO8W7
wA6+aiqHWmgCm2A+RwN+apTWZ0mhykg4Yva3R0cfMWAQ2PHNt7c9A6sS+gQOUUcB
2AZaBw0G8+ipDY+aFFyVn2gvxCgFtGF5zqkBVGr72N7RRbpaPAo6H5hU7B7tnK5X
iWoJqvPnWhvzc0XLib9S/tx/ohIJJo8ZuFNSqhu/+d174JfCH0jmygQPCVPuI3ne
457Pu2Td8SwbAtaETi9SN1c4/XfIbv9dmzTus9ppS3d28W37Cpt777fcXayJGPRd
4NEvzc1nRnNl5nL0YW3wz0b2OIg5HRVsyNO9Uo5YwGP2Ecrc50fpRtCxPj5UsZdO
knlEsHmytwijj20FaZhAVViarkp3Z8mSbVQvbOvbOoTN6CaC5HC7HAp8t2WeJoLw
nY9/LNxUBAwQDWU9y9eiVD53CoBklTVpH2KAUgG3IdnVH3JUilkeZ4iMLrhqucwg
zSrvHSZZGl75jCMz1u8eVCa+hs3r6RAyk5Xkmb9MN8ohjSmxqbNlrQLz6drftTeb
ZEUEtKti1cOESN1vSrq15dB0fhFcjyqtzWkLw50ne6g2IlRZwVAe4PHlHD69zvmq
Pfc9RVvWRWQAUDoRGPjWMJRDOtMOGypeWYKYYA+9a22kg69X0lC+0/Rv9zmeIL9d
XcRR4HIZ/T+5RP0WFJes97d5DHtW4V+VGAT0z8JyjTpErdL4lY/rKc52SFrGBFTG
GjEM2NLOMb3xBZSfxHPQnfDKrbdtU9dzBCsCjnAk42MzbH7rra5uheQ2jcyoVWCQ
adfkD5sMO09zO2QI0CJ1CuD4LGlPLKt7sLTwnPmaxXFPZRLYSA6L8y18pX9Ciace
dtU31ayMc5g+6WbrdtWUznso+BF0E5e0KuzgK6iIoxHMuww4vyJ78OMLccc+1uu2
JdL0aYx4aHQ6pE7cP2Y9VuZXhE8JuOGG5YJ5oFf82hg0iJhdQ4Fa+3P12Y6j0Ihi
8rUewDLi/DA47IU211bVl04QS3pNfghpShrca4CRn5eDDMQG544XEY0OgH3To1EJ
XDZmIDwZUpRBXzfT389xm/NxPSZRjRw+t4r3XOW/t5DYopjZIfKii1XRzWSK6ffD
H8gEPbwjcY/629WuqKPAkBdipMKlZ4hxjieEylMzQkmjq2I06wcCRPIenOr9w+K+
QXmOhgq/F51gQFVX7EA45GJugqu6TjDOMkdc9Y5a8sLECGRhX5/fOzfJCJC29A3Y
br0wjg//KZ/qvzVs44zCsZumlML9qU9QnO4CvV6vF5zXBii9ws+4A27MorV01tH4
Ke/5NBnGslI9B4SKeorYWXzoHoQ0koNWeG6HpS+1YAQx6JbS/c7fWRXD7CJcV0LM
w80w9hDCrJj/OlnmH9M1KBOFeed0IruNKqSW5tC2VviGfXrLz+FiP81ec7OxNLh/
iryKipg5t3Z28oLDol7hrJLdjJW3DDZ8lAoCKL0oQ1lU5OFxBdfkFbUtYk9jJYmS
CqgNsF7ZAQ0Q1mE0AVtNIUVj+nKeofyjFaMJsq2K0OxCXmo7wyqjRVaIs4KTTwrG
p5GMXm5hdUiws8/2aadYpMAL2QUZxhvf9DjHoz+4SX4XX5NJU6/GEbYT68CoIvGr
tKIi8bLStGq42czrFYGEFZ+SBSZL6Pgu32bwUKGLczpHspeHbr+UxX/RudDnDxRh
xkrPRL0yk7/mXjCldH3AMreZ/UTrIEW6CcbHXdYZHFtEzisvA4PFk0/VVWNM1BOh
1luLL7SudisZIZUIHGupWaua0+UFd+NLn6mntsgUDATJn9c7I1xRPkJ1dTwlNYWm
XVIupP1G2W0Gh3LIivvhc0U860XwvY69qhdMRHlUEMzrVYzvmU2h4FO2pSC/1PYM
y99+TEL2HGwn4K2WMkNFYa6hRKm0UL7tEF5zfaFxm4U3zGg77goj+1bcocSJ0wBF
fncFKrLKLLyJeRzzxdmvOLLZhOod1kqck8Vrk5M+lbz92bwx7OsRXEzS5XKwSS5Q
pEOdlhxYMnL9eW4tyIvvFb9q8uPfiHvCy8KSnlviHufyiwLHlisqkShPhJi16mq4
k4zBMVDr1ykiaypQzwkDaw3Rx37WK8cPBr36pvy2G0Zc6JNFxINenGuiCX4CayL6
gSXHCmzZts3sdkh2OXd9taQGQF6Ybqi/rHBmpLFbK3igi1waslYzbYPoRfqE0YdP
sD4SbZNlNu4xbw2lQUtMHUyBr7i4ecWlNr247lto5bkBPb/tWPaSOYVSosqhlw9V
rs21IymHQ3/kVpW3w9rndrvMbI14j6iw6J3/AuZjoc2RwIFV5nLGYD99CLM6dnD7
8+CI9H3yFe7/2aJ4sXFEEj1rPHZEmayvy/meIzd2DvVMsBTqcnc2aoBnTityq1iv
KOra5BYyH6jWkjUwwvB4uVJOJwUkwX+58TvbyprqJlNQDQ8pD1VBBmxfDya71yAo
tCONc8+VxiKuFM2l0V+lT/MoWd6Kv7pNY+hXBwyQesA0k2SGTAQZF/wxYC5/aA8H
QpVR5aYD86lSLrH6CwoPYog3+6jKm6C9EbHCoWKO2YPjINZkm/DalMygCP34zCMR
xnKa16ypqQF+99tSqAwJOVoPPWJlfdxeQ4CfH8Vvacu/dWiKysQ984UagjnVMlv6
waSAeGosJjEInFH3LxzxossWJgIs4mYEtO280Td3raDzMJ458VAMohRki7SaQByx
1qKZ6n3H8MozYbb6M5aazqKfycbqTIIgothbMVMk8bFvijKhN4GQkpEBMey8eB1L
LCM7BvIecX557n6UorGOdIAkhhCrjricPgEX6pmMvskiEsbXY/ViR8alJyqG5MXY
HpFoKklCQr1bc+5f1qLUuFuJRkOiXiRKjnhCKfwO6KL2KpFIDkOqFICgCsvUN40Z
k/V5hRqX7mW7qFSGFP1zvpYQbT/6jdDK64cmoG0CkaGKSgiyRoXD61ebUgnlZ+F8
dCxy5gswmu2uqqXJnC2UbGCPL5cgaNaXi0Ot5lHPzO9+roPMgqDR1AMJzBws3iLx
+687pV3ANOT3JCcBlom2NeAASHAb6VGBZgJWRLiWl7QLoF5kUdnOY3XpjPsBxogz
Oft89pCB0qGvLLFAz+ETm/1i4CKqHEvrvWBqCdFDLWUWHmWjgkVk3fcopw2mfMY6
1Yhw5Jug0mztNhyP30ORLPWnGNwHQKB/sTzgXQw0Y6aEtth53yTexpjG1/NJZ7a6
v295vu4//mwDrzc1wvgY6UBS+Cj81KX13apXGIFYkDi7A94df2jRxYZ8WqFJh0UG
Y5yfThdMi+XlEO2Tw6YAV9nzZfWZMLLub6F+2fMz/gDXLUEY7fDBlCk+5+3dCz38
lTBKo/7ppOoBulrdihHx7RD+Gpfq5x9VxqCjrgUWT0WNf2rvNyPt56KMYBk2d7Bf
tAg3vEH5BXRMhmsa/dZnn5Yxf3CJTFvfjdH5UOsklkNc+oMizhrcJsEY7jsZRuvM
czSSlq+zIa8EOJl+o93UoS3CSv0P1AzPbXvhjSkSZLiv0n/yJnRSdtWOsyFojeUK
GATayq6cu6L2TK8MEWBqIjyL8y+L8uC33HGUPuU5DI6Zh8dLxGHvQPYfYyZ1KTn9
pt7pUyteRa3su25UPqlJKQMu4xO7Ezl2rIPItXWDEWu11/WuZYTkDOZU2KDOQr5c
9oYlYfcB/3Pz9vH2qSkeP1jdPcDFCuo9gv/ZmASlHc5FZZZCKZzAuGzdYUzlpccb
S4u6aUZv66E107ZN4D3vFz6nMVZHVuqJrbN9RW5o/B9Clme3oOF2F5Qr14jzd88g
tqKbIt9n8s1Fw/nM2cpCelpee51HXRKQexIP8rywnBL16pFZdFPeNr9mKllAWTa3
sc2PnUGR5qiLJ/yluYNYnH+Ti30cuL7kEaMGkVXnxVqZDcTRqidm2fgWZxZjmTp8
yZoU+0gVGszt8/3E+PThmZfGBPSKkVwRqO+GPWhQbLZjL6dzplq+PW7WOKMuaB/y
50EVu5firUOqnLoHAYO3dNk7zjakikH0S2jIo91/xwdaZvIDvbebO87uZ7bzaGcH
LxnzQIByTP4FmEnEMpOxrEfvvyMhehw/6YTUnocl829FfxIEgi3jaRXhRFyEi2WX
/1qMJS8JswqYEaRdYJS0H214VH6drtodnyvFK+D5DU+OBvCPRQ2E1EdGyTf1CQof
R1vxjbWVnYU4U0JZ31r/Bi21oUI50rQ4bNoTnl/FZEJ50mTegF1CnBKzq94a0d3Z
8J5C8AMQY486lwQMounZDuxhczEhqFeFAUOftYtygpoZ6D2QyrCNFft7nU2A5AZL
Ht2X3xJhBkiFKN829g5wzUsN5OaKneoiLKG0Kl1KzSmmqFLebyNlsxTGDHqL/ju0
S4HOlOce5LK40ai73/bSIZPFr6kSGIDZivQf45tygprd6RpbeWkpHMjwWI3uegqn
dkXeS4hox0VVadQAmzVQ9N4ZRL6nMVALf259AdSDvX8DHDjbFpByB4wmDRo/y+rE
akHCbo8PXTtmgCQ9gt5T/lG2G7pI2TArnR/nra35s+fosCHV/VMjWa+Ab4PhyST7
Iix6s3ebssFEBaJKjKu9nvUfOXMNzoOe0aS+aQI8k24DL/BB8AhtNc631/ixBfdf
jcIdF4HNu8ppUq+PKXOpa0t47UNKzY++TEzsCS/qz/UjvZSS5uk60I0nczUo0Cy2
JdbZV1Xvnlk28dxOAZnHxdbkov/UHcznXuJCMofJ1Vjq/JBwRfcEOtYD+g7xnfIv
ASv5JAGhiIrqdyycKnOrnHuYmfYhFKxeSAuFScWB11JUc9TsmsE0xZe4/XSaH7GH
VeF1eaNdAZqlS9Pidl8cyOUUIfQHu+WyHELW7iqXWCfJXkz3gFgi6WSTnlb7W1mY
qoNcnmCSNO5DMGsUMKZFE4Q10lUwGu5T1zrAzjr529KEGlAQk6+1oCgO4LGbGTc8
qDoJ/ko/xlaVqiyK+ApKanmuJozacl0OxerJF1cFrTWS2uGQ523UjibSRuSfK1OM
4YOvGGDu3j3jK8FVczwCGr/8229FrFD1oitnVyTtlyqy6VOGVgZwSYZlou/VwGmN
/ZTudYqtc3ZmXjFI9HwSB6rttPUfGJC5iBKFAdvZ6Cx3qU0hVisokyOeQrl/Tp8H
QJcWvf2XJzVXU/tifMrDh0KA6o7MJ+hc9AO5UGjmGes5n9jv3DF4xlzj7SnUBL9l
/JGXGg5G7mPnBAD0ya1m+sdZieX5dY2gJ/nrkmXVAacb6BwFcShnVlp6Tyn39Ff4
kGnovr/TlYjsJV+dnmc8vRecCz7uNUzhKdrxEh3jzNWDVXhlaaJnFjyvItWPxvtz
GyQG+QIlr6k6eHI+c/oJGa+3Rpz3jlnQF0ADjQlNvyIDVF7ud4/EZEmd0aminHPE
7E65Dp994G4O+jJk7NPSZ9skxXnzzXaAE5TIckT3JF6uFzPn+tosFkZjJ592OiIz
NpgmTwSw4/g/E0VbZV00aYXqlPfpU9CMPSnU/K0m/1GNk/DNcVKCytOZRCrPAO7B
Br+t5rnhHrJKByaliWHX0KIXgnEjs/H7u7US1Mx0FSaxcsbCdqDawqOARNi0QL6a
mp72LTzMSdblxDwhQSxldHeXKNYGAFVG/BW4Gn4wS5P+c+79mmEO0Dlj1pC3pVVq
LoHCM5i+i0FA2Ob+XhQQVH306etRKkQJLiQb08smwyTYSn3op5kaTu5igrQ6KoOe
CQrnuiJvRtkO8E8VXhgSfQFJ7ggSInYPtSqR+V6wu2E3zXn3wOaXCstmz9V2Mw6E
paRDjLCtkRDqC8OrmEcX2/CwNVWAXZOViEUBWY5fDiLFicJKz3+qsJyi78in1Yct
zxehfw9eMfolnSLyiddg5+GQ+e0MISZubAXXSFahTWQPeXf9w9jbfJG+V8fFYKos
/YiQcBe1C60xlNRn1erCmlkBL2bCsENsUaX154lg5DRWNE2Onq6DQOANbq/5FOic
FVxzdZTVij8YCaGynsafL5yVSj9T9IvYeH/9HQqmKsZuN8JjO36xolIdE1lnXwNf
KLVzjw6UuOkCIiOOfkrKWiy07dnh9zdNxcBgem3evrHmsBLde5ubyO09NX7hUta3
lDx6pKCTeIjEAiwDvf36bSL6/tA/lv5oGX2r534Y5TFjGw2RoL7V+YezZYmeRApr
NywgMo196FOimc61otXVmt7m4GkS4XKfZgRGe0wsKb7cQ33yHaIv900dvnAnND6N
0LFUBLPfypil9juB4MMTvy8YOY7mS7LSmyfyZVHBZco7YzCLtg/lsq+rxztgWtuS
kZswBjf00y5+kQg+SPszOFqv6Uz1vVY8+d2P69ZlQQ4nP7+Hp3fSqzt3pS5H/zT3
B1V3MOZLjz5rSN4/Qr+qxA9PhSxCene7I3gMqD9fxx174PBV7gQ95JNYwtsOtkyL
LuQ7IdmqVg4Dr+iaDS2OUBetHPtN9ZHubzW8ruvIjsMcOSY8QYoq/P0yiGjtAdt8
rGBrOlL8V1ATFwQ7ELvXTvBtsTZqfxOB3c9uUONXZgXbINqUOvZRGU8VfxuWJ0mc
iNYdVExOWhki9RPIDHssOqftO7nwfmdkn9FbYAF/uB1WjTVjyB8/BwxReWKtQpg0
fN3TSvZ1orxn4T/KBntpDbCV+OVK/1kwljGlKUjq9fvr1DzGEteXP1Pzlakdp1oX
gH+f6H3/kGr1qTw/C7lKqeXCkfF/sIBrddbEAl+g+am99wg+Hvt/QrNSoF+5ybuk
w+q5FxOpzHoKPYYkV4w6cNb5+bXLZ5XuUSey5zixQcReEVWwcJBAwAWACLT7Ws6t
RyRpQoWOpJLbtcHoKa3cRlPPJL1imjrVyhvvwlqo8py3TRpLi7NG3dAKxlFqt8xy
X6444icC8Im27I7Xkv8YauFYw/58/EX4kfukbOKuKy9/eqne8tp7Udp+bkifnN7h
rVDzpCB4oczOskdGgSzYq19VFDoidNa50lTIDqTiduQP9+C03sB09Dp1swkfIDYf
FG5iO9SymhHl0Miy2BV46qbaJm6r1MFAb4Pl/4bBgdIMoeZoBAHMBPCB3Dh8CmxY
Mk3DbRamhD1n9W4DHc1VSDb3kUZyFtf+QVFi5UH3zJ808VfiT8D9IYb7O5tfLKUa
9eUSD0BElOXDHpVj6z7WllC2bfjV7PUBaerGG1BznJZ5SKrjkzGC8Ot9BE3a9Sf6
fyhhC6jToHYMobkBmddcU74dL45rcNTFemFuQWaDy3vK+v3FiemjPXJ1/pToXfyZ
WMKMnY7DkPUHj06z6lGmz66/U5tJui1SFii0mm0DoEJQju/OQJyJ7EZ7b3CHJo0S
X2sACO1vJPXyuQxbqNLMXm+mM42qm6SDWGXwQ47mWMy2h/2s3sG6Ylo/dLZbsUaA
EIWWD/D2nIT6DRl5YRi8pVvDmGz4rOgNCGsZTtCVI5MHZtzbh+sU4t56cv4YQlY5
TD5RuIdbfl4u58W8LslaOoUD1BmNIEzIeGwE1Ebvf1B1QlhfyrMxJNnM1EKxxBI4
Mdba4zfZTbg3GHFrfsQBog8iNjvLpb6ph/u9QiTZGXX8h2FdjylucviLOWkbWGc6
G8e0IYv/xmqw4ooDEfTTFoY5IVPDQ8mEs6edmdpjEmZbDXIREZTlAXaIisAKe8FY
McBNll80NLrGwFb8rwdSxBUEcXPJOnfY5febsr6Z3yTvm34oV3zLUY0l06qauG4g
oFjcTFwa/jkqnxbqno1TU6/GNWLyRwG5QqK3wYD4u3U/TtYJwFoGf8Rfs/0gSMAy
GY11TeY5PVpM5NG2jar8R5d8SXGvEYbfQix7kxtrzlHLNgQj9oHQcrDvT6/mDm/z
V8PVR/XMCn4L6sHM51jT5otPaagjEiZkEGofafZPveLHonRX1k59S7V7u7wvppNh
DVXECa7vo71wYYfGQG8+1h+XCgJKB9fpxya85SUOhAMeFqXLqmXrLd0tSpu8y+hv
lJTWJ1+Y5sd/F2ggqs2m2CvltM2KKFYd/XlpVP6BkjdNDUtF/SYb5tEIoQzcidSj
pjcMwGlpvxYEu+9HgzBvuoEFrax+ua4sAj29X4kl6WeAc8kyfKePTapY6+5+QX0V
4h8SZX1U6nZtzfyhgUdeF9Snt3u9McCnpN3Kxbnt6ecacs8Ok3T4O1lRxEq3hFAe
orameL4v1S9fOoC5xgXzCQ7QjrCxj50RcY/Yw1uL26Fdvwu+vZwknI0yNQIbf3gB
26mRcWTmGdhNzhVq6npoGd4M52gR271hjwRdVthD6rFq0I4pjiR0bSzVXYP6TUUZ
pxCIBNKV4G9posqvdFG1hoePMIjfVycYIaPW0Efr/bQ9YopvZZZs2j7CAzBtUSe5
x/GyYnsVAfCSLEGdTbiABVDp9DBg40axDpsv0/pWvxIbwm+7g7+GSIYfWy7Xb2Og
RJ+RRvXVauzLmk8UZhO7bFoDtNkzBRfI1VjGXOkuyJ45P9dJIvVFIycm37gObPNy
9bmbnWBzSWAkkZdLMeCYytsvEs8wJFmCO2mTaImn/b2eE1TyQGGKOzdEk3n9yu1K
H62pn9WbjWjKIqOcq9EpTO045Cn34t+sJe/hFWMNDtj1jOQo204gw9i6iDi92Fnq
OoAMVEJmuRqtlCn44QzUqL10uPBin3qpAgBw9snO8aNe6TeTSHHlUIDSLuwRsUTE
3/AG/Yv0wx0Pz9w6kFYE5RP7FJHqPx5Vb+7mWdo3kVh6GvlgPtJGYfKshGYGvOa2
kR8e3BOH5hhMaxRMrVGGwW8fmA/kCsjOhgpx2ogY1uatI8D/3XL0rTMp3xcbzlCZ
rUknLsSCXbeZRri6bowuccOAGP8jXe2zwnQDuNxfuTWardLimkoNK95n9ANb72fJ
pkX7JdsdTrBWq8kfPVYHrpgJ98ub+O7NxadcVF6oIPq0r2dgzXGD5RsSjwIwG0sf
o+F9Rz7ly4he9DDFKV2XnUHfs3Hw091LHNV/vJQELH9enjgSiPtyD6aDnPSbi5Pc
LmZFKuUtpKaA0KjwneNFEXS0zWvG/hOuNLdZZzfKLhE+LZsuKMz3S7S6HVcnf2fn
OWA8noa/jVit+qkboAyI62h7390uemRQJdML/ONk0pBA2PvQOSMRCdmAFCsfn8kB
0ZHJ/CTLRIHIqMCE9a9VTzEYd2y8hyE5CnKYztIwpJ306AWceY4obklxnBw1/IQI
JplDBI+Z60hCNdFqVFrmjJ8XVQSh3Hwv5ABK0ktYZUyK1Q2XHrte1QPrK4OXD5fy
RbZZ31/USy/8E46Al8Q7CltwdbCju8s6AHDj5lLI86wxVxFPEfnwug8SMu6Znbb6
Kc8ZUGRkm35tC/uu7snUwhX7UZbO9BGyR2G9wL+8W92VG96JBDmiAGDQp6BEX45R
moKXcx50cQ9Qc2ZCe5MolTam4Ta6pTwiZVExeBgZkZ1II6X+qyArMw0usTcGuCkB
qHck2CKBeG9qVQxJuxbus/n0GQwctA54lF5Ngm522fTjpOmW4G8Dh4j1I3S0ujTi
Vin3I6fTRCO0Enxn+tdLSivQ2w7cR4s1A9GZc2FiVA30EQBqSGSppsGAU4Ujzt2E
/9GzXcOM66u1Hi14MExZTutuKTwytKkS8+msiRGrLCUOwR4Ht6TGZy9zdDCSPyU7
0wOoQj2Z4vK9tKmfbhHFaoJ54CG04oCP1sq5fLHDUSrPvv3bObL08k9/2+j/ZUNJ
haY7Swm/MK/tAiN4IcgaeJpJo9KVmk8MCW52ncdi79SecNyv69Nalnxy5xKK95s0
qgA2i8XItdCBKHW+fB73buII5wNWJPf/URr4fdH5pN2dCHMnZVlr/wArN6L17LCV
2dEnIJyrHtUNEKcnd91Gj5M1IwCQVUz04yiRDdW+nuCBXNPFIE16wFE+Jxu2b1e7
8LqL1DDMLwEJ5Itt5A32f/kmT1A3xbBoE6vIdfB5HT9dojtH5tfZpLJ8UgGsDW9Q
RSi4BTZ29nTAzvOzgxINKlkGigDrEBj4xjAbp0cS+nxKXGy6hc2xRtKEg/c1O0WP
A1RjfqxHoT1e/vZtZRtvR6OkFe7z7+gWPzaYc0TcJFaiHwDJlirs8IMz4lIvzvWM
bM63j5TN2VVIU+1FabfvPyJF28kYRtbsPwzegLqEzXs49aDNBn7DYN7aPg1/oUev
11KFNIUsL+gP5WsKp5DcAw4gzD2zDoLx89EAM2jqxapU2ZZdwOA4Q6je7rXgfg8U
wVbjLTBXD+o7vFQ9CHI5qXfhj/F+sdvf6cDJJ3fC2ECa6QlLVD2U7kLc1bFdvVdY
y/C/4x20jlnLS49PuPvThXdiYh8AqURwhgsJQEmx10wV+5T1nUrlR3s00xIGKN6o
WyZeJ/DmAUGNKKOuO42IlpUDQxIqxod+k3EntBXrR6DRdflsIUjnymk+dGvC3y47
koyr6+JsT6asUDPW+7c5uXpalpIdFn4Y1DTr0ntykhjU2hDW8xSx9ClRzi0+U0g0
4XjyYXScDqg934lnczdcm+gKDOXFNAmEOZed9KjU8Do78qgDi1kdpmyhY092tjUN
dNHXdGo+wzxZrUXSjl4QMy4rSvC1fFCSC3huecK6803bQaYOG15CXoBwlraW40Ly
TZ9QXFznLPEXVGv6ZboxgFsoTn6FhGGRYnXWhkd773CBJHogS8iSUlFHUHz9OH8D
oUwudpkUogbSY4TA09gIwtASEMhjLT4sW1erORufGCx3K7WAWm5DHy35WMDK+XbQ
I9ty5BT8mXk2Wn6HJMlyKNgNinhtp/lKGwPRYtSIv+m0zKC8A9R614RAZOONii/G
IELWifF2XYPHbqb+toThTHFAQizcpwD0pZtIOtADIL1MUmiWYicsan7oPP6TucPo
w86ycI4lsQUQF5onbnenIJNaqbw1GJ1Xc8kUf8etvalOlFuYK5RKexXkod0uOVVs
QsqSL3lgf8LZ5R+j36DWfh7j/ZWc8+jbVbKIGIRf9NzXN4QaJq2OyLMo9du0YvRa
ddSjhSEWTwF0scrGC7N9mEF/fJdlHf48t8mR41vegMGbmDLvqKtKDXlWjJqQTo/O
dOLFF4ThLQyXVBn11uxD3GPzqlygVyW4JrIKubrHh+dO9Nnq34FpdpCiuURM/1Ao
47vpVhPt4zdcRI2449Xge2FKdxnwkrM58v9sqtgGaKZG/nvRe8FyUys2PMV/GJqJ
O+qcfDZdMqiGWeRfkoGT9T1PDUdoMNMM+8osadyrDMmfyEZH6usKC5o6NswF8Yro
uo3AOkzhyUT801wv4Y3mijaLu758WHKVsAzbV4LCRZBrugvZT0SraHymI9J7m3BG
75OL+7qupKZBSW9Kkp3e78STZ3NCKS0nOJam6pkWVNxK0y7aMcWnUv6aXHG/TQ1R
Y4+EQ5wWWQs4Va7wGp+FFEVuhuUN5moccDR0c6NqW0bEEYPlDnGGTBdxhdOyoHPd
r8Vi9dZaLvNLkVBXS03NeUI+fBYUJoWIP7+xMmab+oHpC+JAnvG50sqfSwiiJuqr
9ShjxiT76rYi9HlpKxrV+/1f+EKWx2ZV2uXCu2MtlYUyur7E5hLPV3bL2xDS8GTP
HnlmBs9r4XYFPh2fqlxZKuzTBFuedonrNUEEs8F73pf/D3Q8XourV4buh2TXtkNc
SKFn0Hksl0q7b0G2bN2fos8BEkNAJMarv70AloSRvtAydcgD7zYCQ1E+sTPzqeiw
E5aJGMSVzRGU1leg8coQxDIqbj7Zc3czxcRBe9wCDOu9UvEZQXhrcTPBARmj6GZA
PbKsRxhdh6QpdCZPn05s9ZS84TjPRcGFPbMpqf9eOEyU1h2yJBATvk5rOIS0i9jD
TDtA/XwAI2Z6Nq7VUBTbx+fo34Vr2DWj/7d4e87C+Pd2k9S5D64Donno04IOx739
krEaXv4PU5tOQwNI52ZqHa+DdnNd11DCdsiLJlAbEzK1DXSfIo/CaYi3DN51uRnQ
65+On7OFCXoVAZJhsfNFmzECLHW7JKKhJkAW9Qb4EM1PbuWaOQrQ98qr9wjPnMrd
nJuKw8RsxWjnbamv0/Etfj61LyKfUTco4o299UqumC/OeVTzK+mYS+4rF4t+f4QW
SowrVhdKAWCgF6M3JbLlNGl1qa33h5RwhbtmwpQezhomPrfELQnpsW5dXkA2U7g9
hKsoSA9fcCQS+WjQaf+zDcoRMJh8X75ElJJQbLYzUAMTV5EWx6tlI7XXiz/4NkYF
iI62UZBCSv1dn9/R/qcaFSZ+f7TVmpefPA78t+q6e48KJYRloUtg8TSuyWM1pWVO
PjPgc9netP+92RSajxkdJDz7GC6JkLse1icwHG4DOIiMP02tsdeqe6XGC5omh0ch
LyVbwFlm6Guge92TiwGlOJRVPs4ygZtJF1XIzgxlCsrSs1IBtVCwQEnzezYi8zVB
F9FbuXyAVfD0dzB7MI9kAu9R75L0dsGTz4nKPbEB06+o18HnlKOAvbjpMrE4HlXW
gbvxoyRe4xUS4X5G8SROg6Jpnnamc2mDgxzwsOmfhy0ieI4FloRtdoKLMu/r9FhF
5AF3cC5KqVI7JAPH+d2DMhTSInV3EAP7nUb2mTjbikUMlphAn2T3UxL2wQD67T+1
QQGFd986APkV0T2mOIOqcCxnIbH/d9/ugVafiq54JVZGwy3tImW1UH9QuAlD7Jce
Wy/SDgU/OiLuT02vI6n697rFXUnuyJfkrDd1+D+DYP0SpaAB6ozZQy/XnDy5qTGs
mMIf678AfACzkuGhk18Nb1AFdMLt8/paZC7ZUApfa8q9JefJ55vSh+5HstF1bqk1
tViMDpe7E/sJQJy1SxfYD4FMuFG0IeepU57BXK5bIkiAbXzT608l4DLK66oPSRiw
/AOtRfBGT5ol88Em62kf8g0mCwLEtDk9JEU77LRT2GprYotS0qrKAF+ScywmsHKu
yUoh0K5OH9q7iqB34ArUiMOJHXid1AITBbx+6OQYZKtwZ9njH2TE+r5C+wRVnR3M
jAGI6BJ5Lx3QM7YbxhgtkhEUZbGsDwMD6hl8S4h+mMAddsKD32I31JOGMILLPKt6
lK7hNw7lKoAV/udd2i31VGuTWN8hpQXQHzFo+E3ehP/3nisEUdDHMCdDLAOfiWzj
uaMB+ZHPkuRd0dXqsoEh00Dfe5EcH+rDl/ThlQdAIs5MgbWB4M+EQKt4PHQFluiw
E/iLq1vsM1Yryak3h0N71pdEXEhaRT09kDAiMaAKFgDVTQzDgFWJYEfyRWqYvbhL
9hK18FG4wKygVeqiZsqHUrdTIfwINir5WpLM4zZBG6FdW9Qi+16YX3Jf9HD9VmJ2
kaUHdJKbDov2C9ir0jO5ScQKVhd4P5/AILOF9X+bjqvcU0Jg3LPwrZGqn7dTSiHe
KviA2B2eWT2mjqdspAp4q7jzkg2AKESCPfk5mTi9auMrJeuKheZmshTohkk7twwO
08GpbUYVo4cnughL066y1wFzx39qij7UP8bPEfYylUfwksml22fQHpg1lqPrh+Xq
uqpIrf0xlGSI4zYdOW2ktld/2Y7SbV5VEORQP4ZEXjMHB4YVscwIpMKizItSYgSU
XVjFXAxpu+XtydVhgMpZH7Zr6v+Y0Tv82lfDq0ItLYlVeYvdIAyn/5JQG6e50lPA
iMp0l7Sz4HQNseo2AY/Y0xBkrMVa3PFt26Ucgn7NyNkUrU8R+bTDllMM/ix3rH6B
ha8Ypn/yBA3G57eREFM2WCcETJ4A3ReRMV8LINpVJh+zCgPG1gHITWn6vSgdrNNW
az0Urv6RP3S5b/2RX8883BYAUklIUeyRFimHDKpeRtf3pI72oyWv+tneuUFMw7dl
9spUFPVPQTs+Tj4Ewz/RnXlJO+zd3Jos8SPV49+0mjuQ/l8oN1FNn4aLFg8tQoQL
vkcjjX6FHghT1BG25lFK8necfnFC6udnnBj09FMszON9dWDL7R5Ptvg+3+ndr8fr
A/HSNemfPHTwf4/qMDIXrpGOXtRR0ZGyGPcnexe7oOnyifkzgzxecA7qTcsBbCfE
312fTJL9JiFE+XLbDcW+4p5SpTZQb/C/vOR4JvYekrM1OPR6gXrK9WrHIAl5mguQ
uxmfT/c85fV+o+S+pQtg9oAu0h8NAVc2xdrmiJSC7cDpjJho0iQCFoEzeUf2GyBA
YasEruQ64KL2fe5fgqvvonxnW+ShPbcl/biSePvsONigp/zh9vf0xdlWnHs2oJSq
hwvvKT+6QuM4gmonMfb0qIdc45ZUO7jx0W8ri26Z2urtFxVqLmVRdI6ze7alPsBS
eJAaBeMe+cukIeF7Dn1vzYci6goc3MlzggAkhvTwmGoyMVAhzJZmJLRsQp2iCSp6
jOj+IBAqC82ZGFAzBr8NjWmiRrt/6i+Z3aW0x9EUYSgb3NPmLAjFOgvPHRmEmrlf
1p53jnWgfwSyOb5x8WQVOJYEgtAiLIYnxbwb0nwuZa7oyQ5lHr9x10O1V967AYE5
hXQ7W7xZOAhmIfGAlUkC3T53znf+tqm2JJoeMkwWxxwb2VPU1Evi4fY6fqJmUj2p
/BtRlXx1WJvhOyd/BmpXNfl0Y9DnlPsDVIzRstmTxzk9ulZoebKys91LFXEUMlwA
RZx1lVTaXCCAHYHZ9QsT24exLchjfAhyjxBfpKHK1scqsB/0tuYAN3XTj/k/OU4T
gQxmZGE5Bu42mE1uhW8NlMagy3PS46bJkxYeseFIFfWFM6gwGDn8JlXd/qSteqZ8
RcpipR9LcORLuwE9O4DreRtZvUfPMudNUoNqMaj4v+sMCIn5OS1Q2RySoM8xdbZl
ktUYtoMON3rP3edDx8kmJk6x4bc9w9wQaJV90R/sFF/B3f5f4nEIgTyW1tnY8r+j
KxF0AEZpXf4INvKfWCfnj/vqJB5C8FeMugQoyyURr65p2snNduyiHmhu/t5pdKpx
3wMjsD6qNHuPO8dbVWU8H5i9qMfeNhgosGmXbK/S7ghjcXAN31RC4L1wdYtJE0Im
PN6FaJbmKUQxkPDaYNh/BCishl3hfA0f2JFKF24L3et7FjKLvgLWRUZRLJmJZGR0
CPHNupCO24y0e2/amHuF+L2ubmkRMG2b3AFSzdPSOxB36xEAMg6ulMHLucTCR/22
S/kH/VCBzCGd1kXL3eGAy67HFpL/IFYQ7XjTkx6SZQZC3XYye00wDgEL20inUslp
SDjLp6pAMwngaIJ6wb4ui7L9m13wsnP0iD5X35PkCtb8TRR4Fw1yCoFDAUX+J7Hm
Ywqc7fi/JhLM5APOwbduQXqbyV4+uAXFvqakbPp+6ZlQCDVHrR9kZqbVE57fM79G
pWfsQaThmH4I8T/rFQ7E6nKmvrtasykSP7qPj7h+9HeYZc+SqHo0wIgLU9A4+n5w
RYCRRnwSEKGFLr1uBnLSyw4i8Yd7JiNsL30tt2gO0IH01GrpCVEGKCtlO8QhPXZM
7cpy2KGmcqeZdKxZMx1x4vAMVXFVBcHV62bXVITZG6powpI6b52o51H5iSOEyB5U
eXZdMZ7XQr8qac7IagulwXOZRhtJP/3+kCfc7ArXwC4EnN+yMApE5mnlqDkPNX/3
NvR4SOZ72DD+q1h23Ra4QoS9DcEUJqPWpGe1vBba9b4oWE/FELIFDyPrfflH8WPB
WaJWS9uPcFJV9k5CmlH4VZsiPgOcayNcWo+ScFe8BCQQbpIWLVkPfvgK++zNf98I
rPQdHzmJxfLsfzzdL8hxbgGqAyhQTqF3k2BmSD5lfxPcf1+0wDfKa4kbJO4ZF/UW
VBDH/mcHi9Ze1iXryag+2gSFcLBu5TkMdFCSYUXU+Cy4zopGlCnzxmYzr83pJ8OU
dJHESrF7QBEsU4fAghtyCGWybpmufGRpKI2ukLg31/0sxXjcfT9VV6dsAc6Lr5pT
ugxCXxcz7CXe4Xowgd40clCw4LhMgwlbs6Z8fcrOarkBcLV8dZfF5k6X2BewfULv
NzGU+dGBLN78XPzJ3JOpxMfTCXm7JyNbUb9b2F+vEfap7tvs3B30ne9bHLuAFfIM
FB1xrjiu6hNQOaLRnxlP+I9hIe7pGFZF+d1Wt8NbL02EfV4ggKCwU7XCNONNJo7c
Kb00JQWPZSCH9n0ahqyzctEPCH8Rb8+0WsL6PgkQo1kv3/AtB3AUMt+QAK+/j7gT
8ZkMiBzaYHQSHk/CIDjzLdTrKBKpyV27UGt0UKylaT3yYVJ1fgyxVnv2p6RGx6Ru
Jr3/G/FqSZsFcWoVi8lpQo7YaYyo6wBgqsANFho/Rc5ZpiJClfax0iV3V5DxzJh/
Q0405k/C47DUApzrZmXrqi11sS0iwD89Vu6TkkQitUEkTal2Tl2a1tD5BPvaCWCu
BJxKyj8Sf4BmkPFHyF7bQZaqhA0qCSiR71FewNUMFIHpBrBywpjZ0gCzNV8abegy
CdOZCqEwaxi6F1mpQZnsMYElNfK2D76F4fw+zac2cvt0dX3XNMf7+9NeX6zfNTxw
hZ1zCoup0lvFlfYb++PaRgmuGjdHmyx5SGv2MzovIWJ2ZvEdSHo72hZmgtPidMp9
0WGk2lGiUAvncjcHd5Ryf1G2x69IRP9v2/++z9SgeQDoleVKS6hU0Yhi6ML/58hy
7yIEZ1HoCTc6ei+wezx63EXu/5qU6KkQCcTxhNsVD02U2B6uAJtKQ0YJm35qEgYQ
MEnq39ukWbSpVhewOaDMwwqIt+HpyEfGsauVXcpqNBThvFpjAC8nhfE1BvdEwsQ6
iwss4yhwkJgNOTT/wopcJrazfL4YD86Y24Q0Qtm1HDEvcr3aAQOATsAoPbwpG9ho
XpzoZktovpAVCZR7Qm+I++J0BL71NUvwGohvLwMIwLJRTnNdTJgjmn86UhgpOxAo
/103MScomQhh8omSSnbZmhez+keDeSORbfAfxyh9NHzg3bosIFRfthmxATq7/PZ9
WXk1ua8iCFwY9KgJsi68t5mtbk8KmQi0sQmJt+/bnXn6YMvA5b6HnV3MVzED6zwp
NPe9w3NcwfPHsgZTOznbT8GOLW4HKsQhEb0iAm5d/crQrPLvpNe+VMj45rfwRqSS
05NmZcFvUa1X2BrKrgLoCzfNL2NxSk7BocRZAXPU8U4lXnWcCCj0HomAkz0wd60n
nbu6hEXMZrzpERNwSC0/DucPzDVB9Rq3ON5LJJwSc069HkQjtVKr5q+RgJuyofaK
fpprfcA7aMcVnpBpmYPYr26sy0elqiNK8E1tAUdY48QKKWCIN5XzP3inGnommC9k
KyQR7MMh+zKcwSzy0Av9KXoLSEpriw7hF/Waas/RCHiPtINzu2k6FUq4MXLcXURq
zJo99fwyO4lxrykmRi7NNmbFhiMzKELRuAYpz7b9DtvvY9rMQiVAnn5tcujD72wd
M/YlOWvV35RBsaqNXsPUIwkIR6/ojR92HrqQwap74ZQyF4n5ZnY2nrFn6zVyCXKZ
vXe8XOsnf6xNtG9vgKQc5c8h9rqq7tD7lK7DNZbebLdPXPEzaUtFCLHbpbzLmm7i
exkl/6Ilt8H0P+s+R8rAnXujDTR88/JkpCkTu9rSlDLEvGqkp+Tx3qOYNZHB2w0F
YoRrY57oBquQkzdV+s/v42lniUGVXcaIgsZhWCdHkz4U5/gJxHRuETm1ekAXG4ey
QLWvpgcotvnzpth0wIgyBWpy50vP1bUml2rG4kDgH6XwwyMkx/VAE5Ti6DHCwAEc
QaKLKJdNeA1KfH+xf4o6VS9uZnhnMYyY1Srwau9uqVis4SO3wulIPOeU/uxP/K50
kA0UkD4DYFuGSqErfKdzh+1SkP9jTO9JgMdcDKSaG9Qq58MKNo2QJe0EN8BuPPrV
XSbCGBldakZCxL1bycJC3Vog9NWc6JYx6dpglhwEqSEFyhjvW5YPx286MibJxRgw
9FNgQQKT+x5GK3QrZbzb6LROb7byaNyZoZzq2TGPN6fWDU5nnuRGRZcRCeiMlqfj
Jgc8eXJYPQn6BVMmtLJW1gcVD5kcg9k/ibCChC0f7w7e8o8B860Nj9nAn6bzQlr/
A8vkTceLzd8HPDmbCFCi9Ql8o/2VIpNmWX+8/5vQqiz/kBRLOfqI8NLgrwveBlbj
ooGLnEr7LRHk354/xPQfVDXz4y2qZeNSP32Wlo7Ox9RAK7HSdXzG6IhVU5lCQO53
P4DRO1WBx9GT3WNPp3Tm1gK7FygN//bUiPnpV3k1RhknW+ZkAAKJm+BUSh37JL7s
75g9jPI5TMGVf9kQ9v16dfy6R/JYETFY3U9Ruy+No8/ZLnhpHpYXCOXXCsMcG6nI
Et3ZbTqDwwZRT5QYbqsE0gaBQQCAyLh6bsccDRFc66EF13mLRAS09KHU/Hb/kDx3
3ftuJ3yYRZJTQZaDSAcjOJhbkN9WdyQXUS5sHS6GtijuNLVMyV4OBNwEwq6Aqn/9
Ft59LqXe+t3uGPUSGv/vcIiuc123EtH9G2nvMraJZLhN9nWyUoEUMbyefQisMCo7
F+7lzWj7ZAC6TYkKVK4oHHBuwWgDM66Ow1wiga2XwI06Gpvzub219uVq3ca9xsxu
GF839Z1NQ3PrbW5waQQkuHNIFmiBgX8E+c7LC4hbDBtvOXUvH58eMfZhXuIxumTM
ePK0WAWP0H61vXJuMGlfAwFLeQUEO3eZ+ANXdeeWcyv7apwh0cjuM1I6eO0SNg8m
d7nZ3bq2FYSaJwk3PLx1bzgNZVob8YnWLmx66dwCw9156mm/DQG9fPJUO2d9AlhH
9zHcpAtXur94y0ibZBFbjI11DfSUe/Z29RysUv014gDURY8ubsOvjHntFis8hw8W
1VjRUkIz5TQ2CCclMGYLfvarreCYl+j7zOyCEQ+ReJXk3nd/5EAqNgundfnBJhgg
z+1pz4Aoci0NiqLjkghyR3nnp+xX6uzrofy1Q/Kc2PYpW7M1MITNlsm45kzoxmXI
idC8CwLnLUxUkmUbkmjxdZxQlTSwyAL8DvLrGHzTxxJzFXHxQD49bwBFYvmXqygE
cM6UBZdnByA8HbnjTo6c+jwibr7j3dtV9o1Nh8LPuNrSCZz+bWNFSV1X4Zm7roy2
KjAQ1dnpwSsZuFzvvB4qT1GR0V5M2TT/+Ps67VB3v/SuncAkpKHxxGc+quDa6HzL
B0rIHmsZtRFfOYHqLCjir9cw+xJaoP5S2wHEQxqn/8enZkkNfMTJFpBIbaye1vf6
JmoysznK1qCVl+0WSCSkG2Tnw/zQOhps1wNlQ81LwG/eBh3ptlKPHY6ZPycrKNtB
1xPDy9WkGYe/6hzbx3672G7+NC9tI18PV34cWKHbqAcw50moTQGrgoaNw/IzILOi
/1E4+FkfkaU4QCB7qjsLcR7wssYEnMEVd9cKPJPL/T+Ig4KYhjSSesAaMHiifmjF
hlJljwiQQ55lK/m7WDKLEG5OfQg81Hrjc0OlmWoKSuBTKhxaZD1Ws2nEVeMEjoul
4NtC+HYPymsYjy39Cd6AMwN5svIcsltmP4o0neuiVrCusLP/LsItuVE4iNayGmVs
/PBQPDkHH+6uShKw/69O5JelcgQQRxZ9NRCm9I+FJExC/DU72tKFtIGQPR7940qr
memiDrbL8AXS4Uz0UkE3wFq5erMt+FLroBXNcNsGNix4jnGuAhqkotZwdthTKeSM
hAzm3RZZ1hNltASFLoVFIGEpMQ4HGNeA+832ls56CwLvj/jRkM45VIvHmmjPXDKf
CGbxE9cchJfoqvPs1PAq/D3RR7aZpS1G+SaXzV6BoRzOpBj1jSNS0mgRtmqEIHWB
bT95cOPaGhLEQZooNmIRp2+SDBHyTfxd62CYHZgNb7N3tdZzH+OqHfDVMy7XoK02
155rcab6pYFAeQnzqNWuDhoxCz5W21EkalgLcGi5mkK5N3zHBotK0++dhOfwp0Y6
duFhZ03tcd9CMPDPQdxiPvS79EGeV5RMY6y1mZv3H3rzgwGGyeqiOVgqcLXui14C
APEH8m09+2OsdXLjvGhd2LyjCudjw1PfBJZOthfj1hgS1FNJS34kgnW5iuBDsfcL
g54/WEbpll2gb527tnn7+H1PnzufBeWsAB20Px6jYvyTxp6GJhKf3nfdfYRjzmul
xggsmnT8mZtFRXxnZkVDWjYi/DE8GShyEL5L6nQydXJCu1jOUVOOgrs2pvJbOK37
y2E572PukUaM223kiCJWiiVK2CJmTAa25Nfds2z45gLkE51eNIeKEcqJC/RHcw0/
2m7xUgUjb9cFfjVYvCxK2pmbokKhzE6jgw/OtdCJClOMpkFUd7WX8gWiSSTwHAbT
1eDs5VZHUvypaq8vZXfOp9I3O7/wz1FF9Jpxle0B/M5UBMe1th6r+EZzQhD1/Ekg
rHuETQe7+li/RJkk4nEcxuY07uB2m8/h+XtFlDMgimZyFC2lkwe3OCBzGx86/eX+
Vqyubyo9Ni4dnaMGtNPDGRxsM2r4f6obYDXjYpRluYOdN/lyk1eB3Z2Q0GPP284w
2+BJ/2jKrv1qm+mpJYF4+V1wrTZKF7uSeI14kFu0OVD8nFcZf+6b1ZnHZK0F3ubu
THvlQafIqLVDX69hXhkVQm+tLnVE5FNvzZgiefUHJUMF2ATb7lfeTYzRoxc5um8a
BLRzW+nGawk/D8YxrCJ8Sap88mLIaZQRt7suaSeHmf5mC691f9FkvyfRO/8jOb/W
dyInA7BivAooVKjXAcYNK+tIKVTjXY441Ng/2dL97pBOGpgZ3JVODC1SXyi2hQUf
Mh41JjVpuLOEMGOMdq1ky0ewB/UDj+dmU712rC8Np0eUnRdivkHdbWHB3HA6H6vb
nDX7D8E04DDxWRwX3yFK9uYldD2gXFAggf+xCujOcP65LnmWj41vuPixTPYw430J
YknmUmbU4a8SEleghu2P+C7Urv6aXPAfV0JFxWoMdI2m6PTNnhXiYqnFsm1jILiE
rju2NyZGn3FkGhVj4DWnMUeSHHCzNxoRgRnRBc9odN/7S9YevrXaip5ElZK+0BXl
uouUIlubmLCuFVjHVje5hRKDag6x2Y8wuljuaVZHythjm85WAnkALXfKV6lQ4idF
3l67NqUwKI1pf5k781LTRA0+9eVJjxfWGutYFEJQQuFswKtUokUdtRMHWSOXpC1m
kVPF/baUp6kfO0Tb05aC7qYgPgDz21SmPMHPAo9/GKTylz0riXBVm3qBQ2VsSFeL
JDH9IzQhVTfZMtoFX5a2s0trFNbECb7p2WPexXM1kd7S5riiSZ1wg3K5UlbWMV+H
/Riw5AaqhXV6snIsGmqzfYP3wPHCAM9AGaczy5FAnCbGq/yYgYcf7PkyFYuZoTRp
DBPYUHm+4c0NSs3YeX+GPeLN4eFpXRnvzasHqS2x2HU6gmzWS5alZY54ifDkW1dv
cKtkDHJ6ciE5Z/tUiK8nMGNDwKWHddq4S4IcVM+SXugTqZv+YKV1yVQWzxRaaswj
6RHvEfqGKSqbO215eHmNXjnt74LeH23r3b9YFfYpFJZOjxpDWTdc9eO+2evaHP9R
1qjFcOngtOYh1Y+DE5FQc1SvyH0tU2l6ZlLJuCK4To/qENbm14+z/Z6qhGhxbl02
eyc2zytssIsT4GvkzAQjBnKStp/XjY6Fe2N99ErovbCpXMl8/05ckW+sgN+G0PWn
0APOyefNKqRAXQgHZoQ4cBltFbCFk5mRAj7jum8/Y4ndWhqj6fSp+r9sQ1uIGuOz
/GRRTHtio9Tv2l9nmPY0IT7L+Qx+SFP6wMUz7aIt5TAd9eaYi/MwTbpYFchBGGbO
qk4xRb5dANrsEtBTPSE+sky2d65hWFbU3VEJFEyFfw/JPWrfLEeFyvzyTOLrCwE6
xacstSo7dEs+PRv0l+PLys4iwJ3VlR/iDkwVq5gT3r2f1mXfIZ+BAaO7Gn2LQFov
eaZY3tVMfoFUrHlMEDSiqqNPMErH9vwef0vWBG49FARo/aiwoqC1doTS9hFQEH9v
+LJB68vol1qo1leNb75gQdTJBoqLQmssh9zw7Lyu6MihnCqUd+u7fFYxUcf9p3KN
vtiaCPWT3l7FmWR3YLnwHjyjPGrlBkH4co1bDlCE+PYsxK/ju9B+gwUCIhaW9BV8
SBf1X9Q58zOwuw6D9HmCxazvU/ghRtcOuupom3uyNsylx6jYAN3waWvdzPZY67eT
9RDIRISri3KV8PDJmNDuB3ags1vewzasdjqKv/xH2GX/HkEEFv9KUqpaGdrPmYXm
iOZbSvVUnlw2Xrm4YfPQ3UlEoFL4xfade2nPHtIoA18QNcFYR9LQ6ukI+/7mOwxv
j0k9h00MR0cMLc0XXRymTgUeeV6LZN4XkAmrlDWkfNn+qLhysLYjb37yfffFAMMY
ObF35+iFPWKCEEPikjI5zMQDIqWFFKYI2AjMqhKJMoIxuoygAVQh4pbdt6QVHkQZ
hINlUEAhZeE2y3um44uVjXTR7vtlQbPkC8e9moWz3kNIyja5P7mX1aN5h1mFoubL
BDLZweDThwDA5PcEkDMFWdKMG5k0guJhK0+KL1zbaj224dt8H9rIT2lGzq6Jdi7l
mF50nKz0ayJPD+kR0CKUQCKoCuLbByDgmfvJFXDtubK6D1A7R3dvb3V2Vb2wHj2u
ejYRDefO9mvT+fNKERRQw7Jlb7YAJBjMgWm21iUnMcCZn4u5yYp0fr9EtZ+91q3T
fknhbtwEx6yyEb7Yo6voULFQn9zti+mou3lQjjf2rfLzO2Gh7OHxNOgsOwoxi9MO
C0rn6t3fGyNRWCloC9ZFJ7+3JmK4TV9gCb6ezMrMYb0JF/Z6aKUufFU/CbaeHZD1
+pdzoi3QmNJJru6ISacSZk5AyFCy19+QVxDNRbS2w4HEb3uxjhWpuE0IkWVwXrTQ
9DRVqec220wz4UtheoFmdKjEymHSpkoHaOLIO9ktVTZLKBz85U8if4OjmXh1FrAP
0vgLJ4VKBkwW2MLQNH3RVpaWNggjdPgl09CoTqdGzdmn5H6Bf4cEkkJYDe1P4s1w
Xg/HQPRvRzvqtD+s7T03HRSyyVzDgeBc4uy5miMi6Jo1ueSyHRDFp/CBch8fzPl3
rf9c7I7ZF2kzjj0i9U6FRH30fInwFdPK/0d+KeQCWbi2GBS1a1DSuTyO4QngM0SF
Ntcd1kPKYr2gp1qOXupxX6zb/xy5LJSLKRBvBzYD6AFQF8nUxEn0APeeoff+vRU6
K1gpwHd6ArKzQmDy2Yx/T6N0GuQdR8Ne44YTfrJp+75+v7kyGoegl5lBDiahJW8Y
EtP1HY+XAZ4774jkOT5CT70tX4h1b1d4fKt9jnBpGxDac8/d43+KVwS3gOntveql
cvLmj92Zp7M59iY7mgCcKiGTiKNrVWhGOGSfOEIvHeZKu1vkKIQaEjDa7iybJKL4
/PDBIABbrbKFOAeV7P2+UujBhuUjOznfDhWN/NOdux1hVL0Dquj/QqlwGwgvd9He
2flPm+xopOcL6y+ue7yQg9+3lfQvltTa0QkXAOkQNRWK2L6cJjzwMIaA7guzgYiy
V0//z/Szvf0ZFN/6mb1L4S9F2ET9jIJJLtvrWO9SQbux0OTI6LOjlfx5BX13h6pQ
2WzQwwQr6tDmG6NJ7wmj4erWeM11KJT9GfE0encaQjyD6dnwFNi4PEkmphGmLxnc
MUVD9l4jl18HCyS5ahPlIotGIvrMazezpdWgsfoejSFYslQBoE+CXRnGvMR85Uk3
9n5t/KAmi1oEmXe6TL9K+4q2ujGKb6nGa+Y90jn2TF4zgTPB+yqvx23xDCLudE2f
QfBkdTS8Pea325WSOVcFHH/ZH6Fl/4mvxxU00DgZRTGXxqzXUY5L6bzzhKj5M9Hq
y+LYhBrDBV2mUQKwuRFUCWIFV+ndLrULqaif5xI9VvlHhKB69gnGCEJzj0pvBH0x
NNwnIOwx/YqJtsQ3ag0AhcxEi7o63tXKvkMd4nuvshEY172xDy3gal8mrBn51H6f
jGFPCCnt9dw/Cxqcvtqlerp0Sf1AIUVIpH1PNulXL/3JT4iY3NeyMd6iTs1+Gc9k
eIQMxv0TaWDIZJ3RBRw9ujI+lBPkwhoNQ8y+aL1BbqOfA1vMLCKPgD+aojR5KPBy
mFaneRCUinofQqSkWvt8ZgN2S37WP9j8uetorYrWctzoJcp1Ly8xAsqcScvGHSdT
t5z2VQuSbxg++TWpsz+OSY8/iYXYgTlFkbE/RpBDDsQE7oVC2gIow4imH1R8ahaX
gGKR7OvfzFHy5XaYUCyuTeN+HFijVMlpfGXUm7P3Osi3DL+JpmF+6S3/pURVa+Vm
KsZBjN5X82VVP9X+sn0vyCQ5y79rYomxvsrashCO6sMkWUkW0BMLSFxhMl5UhR6Q
AeHKx7EKuLpWQMtkVXv+ReBQxL/qcYuLmus9MBjIOn20hnm1ERhH2le7doq9Ly99
8BKVWAD1ojDUe/H2qJC2oTTpnIIwPic6ef4CxwWZSNb2NIukPa1NVype8VHxiuP/
877dg/PZarStYBMGj5+BiqH3Oops2/HBa1rCVrWq4jEdrzMKRn2GTxurVAdq9JLp
1BKtCd97LIpFDucvGpqsRPW+KclGeKa14lYqfxxu/9Q45norCxAWmX3fNihbN57t
DT0zaIhVtndwaLKq1BpA7L5cwEjiBXQlloE5EdgW8pGHVtEpqzjShnqfLvTiLrLM
r/sDFCy4AjE/HwFUS4GqEtdw6qMMYeMvubOEiedmSGzL2vDGeejElIELUel3/vLR
68v/UgzFp8fc5rN7pmfbRzc0JXeVNo6AI0jF7SucSHx7Lfw9/u6rX8uedTatLtlE
CbCyuThy3TSwdg+sVYjjQPzcu8k+FEI1z9y/tKELSHPOqUwrW08cxua71o+BHUqz
BlSkTixOePTCKyVFdpF3xe2ek52GVqCSv14oKJXj9fjfSKDegEw+GMkaRzpqa1he
AByLwUEMY2OS/VisiH0sAYvpIc4b1ygy0z/wpPkbUNrreOt0yxVj/myPmjkUilk2
TRRnj5Stb+WA+CPx6+ddZ5rtoq+77hWoSo2qBiOy2st8o6MySkDMRJKEp2Aeh32n
ML+eUy70nt9dDaVHmAfp1jsYLnBud2z4YmW16Sh1A4/aRxpr6ZwFKUjDTcg60x9L
yiwFxpE0QVYLY2Gll94xenJqMOaqxZkj0J1euEgZXiil8GyiuosSitIhIAt7TsQT
oVxfQiam28LUBLoYNJ/Ge8Z3FTeclj0N+B54GdCnaIXQ59+FfofA1wQVib1JtkSB
5yzpk8tSomNwXc9GRZ5iO7RPyskygTxmt5DG40gmevV9BrikvuA6Lx0JvJhu1RsP
V+yRjgNMQYOHQkcs7dxRK9YORvuKFagbFKM1dJ/rlcynXs+fKXh3WayGQb82RjIU
1rJiqu6d4hudZ5Btkygkw4L6v3GhAFnNaAsDgb2g1cQTKR0LRpeqr2jWBnVjx1BA
F4ZoICS86eTW4jPK3Vsk7bk4BBg9Aawxsh54GBZrpmXy38NVqOuccmdfBj5X+yxP
c/7v4bmpgeJY9ikgtyrRvsY4V8t3KTHXUmqhg3YI9Sx1FvP5sbY/RZWENBEvW3+7
NBfEyF2JisY+S4jnmtnDFNysZ2Jz3LKmVEhC0X1XV0K3Pn1CrcDhfKJMZCTo6Qgu
Bxul/nsQVW7T+34fYW2Rpry/Nz3tdNQ5pluYGQ1Du0aEaU8cPz0pPdE3ijnphH4P
JArdm/SWKxQtex5aZOE7ck1PGG6A00A8G7xhbZocP8B1n9RWDSgLoZQlgtiQoASc
f8Sq2lZbR8p7fQ/265ujY6GgHildd8s/l01M3OLxTb+JzXfZanp88uAWo52ZqJHc
D8QJUuRYTAqMJZVcTpN3BylzwyP5ez+u8mteA+n4PtseaVwEaCsBbC5AzRTK0cIE
Z4EYH5mPHtJpbmS+xJr/6zSE9p3qmd+oDPhEe5mK49mjC0g3QGFbBNWVdpLCH2Ld
9kbV02qAEXv5wWwcSaW3BlFBhbBhPCP7oqGwrhAECmbhbvH/NRYsFk9H5AnL5ve+
kbp1nlw1AIVNz2nnolAPpwPBJmKknMFOKQnYGbm+xg5vP2xhQ6Ge+C22a4RwZwR7
Di3ZiY7+3TOow1VhAvWR0ds7NdyXfcWXXww8EnFpIYIs4iG0DURJVuMzWh03kuci
xhgnkmhhTDTwZL66IiryPwwEcxQvoa51OtpVzinRWISPq5pTs51A63euHzEqNNnC
N/wQl5owmn3bL2lUxqtSq/8l13LMnCogM9mnPrZR9d4uv67mi4cDU0Ja3n7Zq4A7
xHRcUxDs49xHOJGccn/VgOu6B4csfer8uRwWncFinq4aFa6Xzaxq1DUOEAsqTVPs
+18DuG2EpAFRHMZcrpvqNjg7BcAIImQdIDDUNwbOTbqRNF8gzYiJI/XkywfoliAS
gIte8cU1rY1cWDND0zDvtmRe9kNrYKj0a/O410zNK/HZnaw6XK+yqKOQjPwGz+HL
pJ26A71arf3EQKH3etsMOaezeKAtDS8mg523OBQPiYzePXYB9IqiG4MGE81cEcrk
WmyNs9qeOuj7urE9b+rWESwG41lnOAtJd4nOmgsa0lv4dubenffRtcYipA0ik8So
cwRlWQYmfRCKd4MdaGcSbWmaaYVVXPxyqgvk6J66XZKLv2wisaRx33lQa/7/qeUu
ZFwbUBOXbU/upzDne6fuTx9lt7XodmN/81BUJZUtcc1DivcgmTG5J+jO+7ICV63R
Qo9+Vn4I1r61gfF5yjKbanaT32m5GNEBZYFB2dv2PK9kWPKzCC+dChn/8UdOkbl3
60MzWZ6DnEP5CSGhmlhFrIa0vH9LYcbfW1k8DsQ5uwLmusX7G/et3vogSns+nf/B
sbB9Z2kXAwaxuUJ7cHgnLtGgS7Fh3X5RTKh6CvjsbJd8o9rvfoOrcHmYOdg9Mn1Q
F8AsBXwKIoXras8txo+kkcTL+/bYNVaabMkFZddxjAb7y8H1t9NjsEWgBgVy3UK8
9EjuzoEk1QEsjQtWJgap6v9n7bkRPh/zIDO+z4aHpmyGZMZIDHn/C2QQN4pkWgSE
Xp22ufiFVfOd8Wrr0DU4ggaZZq/v3nHXCfSTaxNU8W5p0QTvHyHtyy3WtUHBf5v6
whK+DSOHP6PLQJ0n6IGWAcK2jCrSIJgmMPjir0H9IPZ1Emc2NvtC/RIPQ83mo8ns
tmh8kv6VYlRWpYUoIVeDChl6WEq+TtAKv9Wwfw/cMOJ4IlPkSfJY4S7/Ujjp3i4r
j2BmqT4i/KsYVTpUCocJEJQtMd8F4wsl+NbzjsCn0spVfRzDvN/2RmTdhN2HU347
W2o79qD61RjjuHL7Zj8usNHZ8lNrS1RpS1ptNjUaRA2bDDU6DVuIguMnm4IjJUsG
AL6JN7ycHLL3dPV2LfaGKroD54hLQgVbaD9OhWWdUfYS29nAIN5R0Iu8Fgc3qblq
zzmlEA9M+lbW+Jh8baJgIOkxx3bAg6JCq8HqsuH3yKMvPSyi5wt4p3up03HF6eAd
HlVf+fJP+b3lOYXAXtpJbC98IeoEHsuN0g89yHql9PXuWEm8ITC6mWb9gIeKSmpm
4NuQhjnlrTSKknU8LVr0lYKqyH2HxI5FHxiki+od6IAVEyxaXQVdmIyZODxl1QK2
JmW+r/R4CIvcEiuNo3FMXS0WxPHnDEB816qiuARiFYTgoVwnH4dtuxCmScJVNRMD
j95gOr/jx2j+DtykhhcFjZPvCREJo0rYZZMi6+O3YIVbiMG2g28Y/AW2+BgBb8ls
2OafVTc8b99eG7yFBGqxa6f0qmLYn4KZbUJz9AUVM2gkU2oUFDjpVCe97CcGejz8
DZbG+J9VWhYxvl8m4jl9hFk1iNm6F5l+7QwmNF4fxXv73PuKKjoBYzQp9Set9drE
xAevxciLAwB2xrhHXFXQmsSBSZSvanjIsEEoZDMHcQ3MpSal44ckbeOJL6F6FEVP
rH5i653o/cc/2NPO3XxVM0PCs1i397EcYaX8jwMNfOH+wn2C43lVraYhZiFSqvrP
rh8Y91w9KoUG0sSF8S4RVzq1kuuodeWbXVEEyiWbPfEMEFz88TOJt1Ey2fjf2Vmk
7gFNzukXjPDg00+Qp1M9D7HMKvpMajDh1p+ETsQZEzSfaFjUbCXCXQ0d4AHxAtpZ
z33P4LEE6RGvVhkShbyyVxoM/M+8x67+zR9QRIRMYLBzk5620N+/vv9JBEnOvgc/
QL7MF+zMErrnwNX32E6N3KQjqK9MMIRsE/zR9PX+aYp0c4n96uf3KuX7Byc5NwAo
Yu0MDDOckfTmm3P0MkvUi3UYN5q8YCOKMNr8a8jSRHDvkACbb4C5VR5DJVy7IhXu
Rm5sFBZf80jACTNJphrNmj8whrKbt7qy//EPoi2rblh03hUy+sittjkq0BiZ8zIu
AKNY/aVATtf2FNeqx7TtU4dIKxZpDihekBrRoebqXta6ggf7pcsVQHX7eAKfVeAL
7r65hxAHhkq16wFOan1uVaDO34B+w1mgb02MevRJY3dU/TXe1Q8O2+G5Yc1/4QCv
G2oWbVUl/X1HOm2gyjV5mjyVi4ls19TyyhNgKZWiHSHOqUeqsURGF1gK4EOSIgCE
L+zKaAPxIap8NIvmI6Bo1YtNNqNNTEbuyJMWUwPZ8UZMwHsrO4hvmFFCPVS8ABLL
IHmqlmxTYZyeswkxc+WRw2xKNpii3YKdt9q8MwONO6BX74i6YpDJRIT15Wx3xCMB
e4WhFmBRHOXsYHraE25NJwFMVxR57iHSPUMTO0vIryNDdhGK296pjscDKI4598oq
keONLrSuaNXrkX9muJkjP90C4It3mEgq9YazLwMCO2IGieXXAZubqbMfLCvRx7bW
NDje/jIidvrVbXhQsvgjyd1xOlX6qAZjPUktvkPr04yHB7qufCo1zLxmQfmf7z3P
5PQ3nLhCf7O/b0vK/I/x1k2RtfPyZUJn7J4/3xAJaSiHvmyP/RRhIFOVlc7ljHvB
gSOHoYLcVCEa3WadpTbOnNHOOYOepTeB3FuypodpnhaNjsyS2pW+xdsN62qkiRhk
ozISh21evjRALAZKfPe9+j/47s2j/C+QZvbAhp0EIFSORbLSjRRvVUg6rcXDn1a3
f3qz0ETjrZITwNQ6d2gonZPMRgIxeE9gAo25zx3n7NeVXnl7sMQLC9Awk5j6ijnT
NRJaLYLjbyr7aXUWDx9CwSF4pz34a6qPQqYLHWk//Zd6sm/PoZ+SUWGt4ZRIi7bM
0RGASWL/O0EvSAorEkX/aN4o6LFIetETgnqm+mbgJ0WjEd/YFANgT9LyfvZAomDI
j6KcKFfvCT4kLAY7G+ql67Ij30aBWJ3YuVyL1AFfCpHoAeXImqLvxXpH/lWvekdZ
DTRHmVnjAkGk0vpqJ4gRqmguv3RQO2HCPfImU1XiE0+7i3kaTlbLBgZt9jQQcwTA
QlBnYxdz+pI4WA+YiHFJ/TPR3UYaBgqgFlwk088iwk1yhD2RSjJq2x3DoquK5VGP
iFflDd/TB1Pf4W/mCLPX5APYdf9HM7L+yTb+M1g6yZPJk69/q1u3OoBcZyGGecY1
8SRnJ4MCZPjQKlVQXLLFZM28wf8oBHUZP4Da9I0IG7g9t5/EcmtTkEQr05CajTaH
RxZQemibRRE1dDH5G7J3UVhLjdbq+KpCyE4CeZ7qec5U78ni0JsAv8LxB0Gx/5Gw
FX92S4ThR8JFOqNL6fnXgjF95tNaIE7VgoQsqpJma3796wcssqvCCNWiLKLaYLgt
B/ddsiWv2Mn3uiTgou5LhUSjcTQsXai8yeD8tJ2p6uelCD7Au2bbjPXaMuxmkzLU
HHNT+HJT5irmzDID5hy/NoKzmhXf6bx263I7DTPeGNxxwc7cT9i+wYjL/DY5Rz1m
jMOkoOgGB7MwTl2V/l3wXx33BHLNAYuHNPqPV7+RICA6NdVNPb/mKib7Osj7NgE1
prvl6V4pCuKJBSUG4JH0AP0aeVwEDQbHbs3mCWrq66aEs+G//JXZgJyBib8/vxIa
AM4LrgNVrP48b320LhB5Xy/db5qgMd3kMSmwBlvmLOhI3fOPY4pz5yYTGil0loAM
4jP6oxmL+y/TGGfi92ryE9OehVUHwMaA8yk58Muaiag/CcJFKzRbEMEbK8qwY7Bz
pEQPl96MZUl66IMwN/yVgYc57L4LceiKxVNd6zU0FkQg1kYy+pUDHmz5tpdQ5qrL
kmiPxd5IZGhcNFX0IDwsiWEafko9TmLtJkibTIaRFVgILLYswlkE+76Ix09z/fOx
S/UxukCdVxRLmKIVuelu+wGfpIvZaT7Wf95GQjp9bYppE4W+6P/Vc1aNUsdJ/Izy
PNpmoGk+jPPHSSrIb8ufmqMDNJaOnvPgJaXVgNVX6xcHGgYf6M+JiwGd8txN4i0v
q4Sx5yQp8Bgakx0vzl49r1gZebtBUhfmAinPxrTifwhNdoo2b9LIgloP9dWWCFRk
MzGhSmTmgT+VuPH8nPSGvG1YutyWTLpxgDWyvMw9PoGGOiI4hFtweo30yVeuU9Jn
MqZfB8fp2efBSkHxpz669bNnxCkmKcYeSm4BcydIKeB6RBAKo1rn/sTREeoAJDuc
I2Ywpe+kzWSBRjQbCn3SR95z5Lj0q9r+tiskjpCt14+cTXbnS63xI5AclRUE9L0R
rK16eV606bQNz4Xv58smJFe3/snqG59WxDJJcOhTmrWHo5YKJiK8hE1eMI4PKYPT
SweELCyw77RYTmxt6NzEBThf3cjjOMmPddMPJtcU6uecGqMEl3sl2ITk7xovum5e
nM9IdPZwGgVK3+Np7nK1IGzgPF2bpUNjYvMjn46rsZMAVmg8Xd/0AARaagYwSnQT
rx1pi1TnJoj8x4zHg2qyP7+894eV/VRqjd8ou2hj5V61S11L2N1WkD7Eugietqbq
/8mMIGbHiu6vtD8fBRO8cymhVTVn88FqT7q1k3J1JOiDi53MsrP/0gul+ZV27qiV
QknWk8WZnyzROaixxGzZhFklilqxEjwgOH4CeFdPHsNuDn5R5dZq3KnXwyrInewD
JX59RrbhLFn4voknGAjncDPxkfMwE9PqZatIN33GC50RNl4FRIRrdHXG34t6+0GU
42g9a5PzY0QYj3YoEBXBpX1SZltQbWxx5ZgOay0UwYxYjKUhA6V4IxdZbstgdrZ2
nCGDxGCURWDRhMjYhdhKxgYoDjBg+ZncOXSKbsEPqUt/p2m2BxAlLWRpvFPUbJOE
FVI2sqsa9q4yk/mqnNNAskvT2i6nB7Na48m3xngSLmt8uIywpRArRloaTnU7OjLn
82Fdy7BvHqxdz16GLIoJjJQ9h7A3vdmRSltWpkd58KYDWponS6zTg1MQd7zfJzD/
N6CZy7JPOK4JfqTqH0DlCi70t+McJ1mS/7M9lwGnu3RbLSVhAWdNIeN1Q3URy1u3
8X/eNoNmk//1zHPFRnBuU6SZ2rjfOn7K/cYJ0Rdr+ynHeH48ZWSXlB+ZcUyBweg1
ggLfT7Ne0h9O+qJ68R4v9Z7YtOdGfNXRrZDMNNmKCmshgFqeLcNwkpWB/bKAoHl3
PmCBSvRxuTi2Cancr+YtJU79u0RQgc6jC9CqipFcNokBwB+rYvZCZFbRTe4DwJGX
63V/QGI21p2GAmnTl2TvVNIvaMc8bYxqKantshqegHQZjy3GEuLv8rDF0LODw6dH
AIFqSlhrOwXB6VDRYxROaTpNhb5NlEHZwpHMKxNC++hY+KevAWqKEezQOeE63/Fz
y9mudbXMYu7jGgAWVDzqe0jEtJmCYF+H0hq98QeRk7R/w842hBzuGnrDH7n57lxE
+Rp8vQpgyET6SHXKfZbBTGGE2tKSmnBafx98B1dfXXPeZy82iRkdtr21XCKntAP9
GmSULWQO0S1+vNMDppouJDBzxyXf/gj440uitC8HFR9hhiR2lCw4xe2ClgJDHicl
X6SlWhmvt8zplqA/4Mfiw7jCc+VeG6sIaESLC3s6IRRkK0uF5IDJ0Vw2dHWllRDB
5XHz0qjQKduXWVnXiFZxAo78R38Xl9sXRUQxPM1izij7B6O5QaseDsojtxwbDSl9
VqH4Y+9mRjDsxpBj3gm6nbVlvXXnbD1jtTs/FuYMsp5+U08oakI9YwZinyZa6Ru4
2DOZv2Z+bmoxMKAroLNuUaiu4xrACM0+S8As2JrjZa/xsqUGgBTt+J0OSDdUQiGR
uhLBMjMLKxbZG5KwJyqdbS06/2mLqrlxMRqBW3/on65vokjjgqIz6YVa+nzvslnS
as5EY7TqWbfJcKuwur0sNzyuIuJIFzlsM7XlyKstTlFoa/NWwG1JcJSC8cuUdFEb
cKeyfwix/8NErn/wEyUHMShIOxsRHc1Z+OfPIwTRhIOTQTIFeI8nW58jBpfPhbRb
iMlwGtuy4q2uqmIrbNla8M8g3JYiEsZi6+wpwC1WSQV1mo3/cIqkNT434HUvIZGQ
J3iR61l5WYKuiBCWJdtKZwFvvVwLktXrQID3eu2QgtnVVB4plguura5A843cVllt
p9HEkyYQjCHGII79xsbSDNohvcfNIaFyUw9S5uh3uBMsLFpMdqJPApShCpt9doGw
EkIAkybOCzXv+k1IjSHaQXhT2O+zUaH3aLIrn1RrznK+r5K+LN3W7Mz/g5brmhsS
`pragma protect end_protected

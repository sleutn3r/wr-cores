-------------------------------------------------------------------------------
-- Title      : Read 64-bits timestamp as 2 32-bits words
-- Project    : White Rabbit generator
-------------------------------------------------------------------------------
-- File       : readTimestampModule.vhd
-- Author     : Peter Schakel
-- Company    : KVI
-- Created    : 2012-09-10
-- Last update: 2012-09-10
-- Platform   : FPGA-generic
-- Standard   : VHDL'93
-------------------------------------------------------------------------------
-- Description:
--
-- Read 64-bits timestamp as 2 32-bits words with the Wishbone Bus.
-- During reading a disable bit must be set to prevent data corruption.
-- The Whishbone Bus addresses are described in the wb_readTimestamp documentation.
-- 
-- 
-- Generics
--     g_timestampbytes : number of bytes for timestamp, should be 64 for 2*32
--
-- Inputs
--     clk_sys_i : 125MHz Whishbone bus clock
--     rst_n_i : reset: low active
--     gpio_slave_i : Record with Whishbone Bus signals
--     BuTis_C2_i : BuTiS C2 clock : 200MHz
--     timestamp_i : Timestamp from Timestamp Decoder Module
--     timestamp_write_i : Write signal for Timestamp from Timestamp Decoder Module
--     timestamp_corrected_i : Indicates if Timestamp has been succesfully corrected for errors
--     timestamp_error_i : Indicates that errors could not have been corrected
--
-- Outputs
--     gpio_slave_o : Record with Whishbone Bus signals
--
-- Components
--     wb_readTimestamp : module with interface to Wishbone bus, generated by wbgen2
--
-------------------------------------------------------------------------------
-- Copyright (c) 2012 KVI / Peter Schakel
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author          Description
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
--use ieee.numeric_std.all;
USE ieee.std_logic_unsigned.all ;
USE ieee.std_logic_arith.all ;

library work;
use work.genram_pkg.all;
use work.wishbone_pkg.all;

entity readTimestampModule is
	generic(
		g_timestampbytes                       : integer := 8
	);
	port(
		clk_sys_i                              : in std_logic;
		rst_n_i                                : in std_logic;
		gpio_slave_i                           : in t_wishbone_slave_in;
		gpio_slave_o                           : out t_wishbone_slave_out;
		BuTis_C2_i                             : in std_logic;
		timestamp_i                            : in std_logic_vector(g_timestampbytes*8-1 downto 0);
		timestamp_write_i                      : in std_logic;
		timestamp_corrected_i                  : in std_logic;
		timestamp_error_i                      : in std_logic
    );
end readTimestampModule;

architecture struct of readTimestampModule is

component wb_readTimestamp is
  port (
-- 
    rst_n_i                                  : in     std_logic;
-- 
    wb_clk_i                                 : in     std_logic;
-- 
    wb_addr_i                                : in     std_logic_vector(2 downto 0);
-- 
    wb_data_i                                : in     std_logic_vector(31 downto 0);
-- 
    wb_data_o                                : out    std_logic_vector(31 downto 0);
-- 
    wb_cyc_i                                 : in     std_logic;
-- 
    wb_sel_i                                 : in     std_logic_vector(3 downto 0);
-- 
    wb_stb_i                                 : in     std_logic;
-- 
    wb_we_i                                  : in     std_logic;
-- 
    wb_ack_o                                 : out    std_logic;
-- Port for std_logic_vector field: 'timestamp' in reg: 'Timestamp High Word'
    wbrdtime_high_timestamp_i                : in     std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'timestamp' in reg: 'Timestamp Low Word'
    wbrdtime_low_timestamp_i                 : in     std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'error_counter' in reg: 'Timestamp error counter'
    wbrdtime_errors_nr_i                     : in     std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'correction_counter' in reg: 'Timestamp correction counter'
    wbrdtime_corrections_nr_i                : in     std_logic_vector(31 downto 0);
-- Port for std_logic_vector field: 'disable' in reg: 'Read Timestamp control'
    wbrdtime_control_disable_o               : out    std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Error' in reg: 'Read Timestamp control'
    wbrdtime_control_error_i                 : in     std_logic_vector(0 downto 0);
-- Port for std_logic_vector field: 'Correction' in reg: 'Read Timestamp control'
    wbrdtime_control_correction_i            : in     std_logic_vector(0 downto 0);
-- Ports for PASS_THROUGH field: 'Clear' in reg: 'Read Timestamp control'
    wbrdtime_control_clear_o                 : out    std_logic_vector(0 downto 0);
    wbrdtime_control_clear_wr_o              : out    std_logic
	 );
end component;

signal wbrdtime_high_timestamp_s           : std_logic_vector(31 downto 0);
signal wbrdtime_low_timestamp_s            : std_logic_vector(31 downto 0);
signal timestamp_s                         : std_logic_vector(g_timestampbytes*8-1 downto 0) := (others => '0');
signal wbrdtime_errors_nr_s                : std_logic_vector(31 downto 0);
signal wbrdtime_corrections_nr_s           : std_logic_vector(31 downto 0);
signal wbrdtime_control_disable_s          : std_logic_vector(0 downto 0);
signal wbrdtime_control_error_s            : std_logic_vector(0 downto 0);
signal wbrdtime_control_correction_s       : std_logic_vector(0 downto 0);
signal wbrdtime_control_clear_s            : std_logic_vector(0 downto 0);
signal wbrdtime_control_clear_wr_s         : std_logic := '0';
signal wbrdtime_control_disable_sync_s     : std_logic := '0';

signal timestamp_error_s                   : std_logic := '0';
signal timestamp_error_sync0_s             : std_logic := '0';
signal timestamp_error_sync1_s             : std_logic := '0';
signal timestamp_corrected_s               : std_logic := '0';
signal timestamp_corrected_sync0_s         : std_logic := '0';
signal timestamp_corrected_sync1_s         : std_logic := '0';
	
begin

		

wb_readTimestamp1: wb_readTimestamp port map(
	rst_n_i => rst_n_i,
	wb_clk_i => clk_sys_i,
	wb_addr_i => gpio_slave_i.adr(4 downto 2),
	wb_data_i => gpio_slave_i.dat,
	wb_data_o => gpio_slave_o.dat,
	wb_cyc_i => gpio_slave_i.cyc,
	wb_sel_i => gpio_slave_i.sel,
	wb_stb_i => gpio_slave_i.stb,
	wb_we_i => gpio_slave_i.we,
	wb_ack_o => gpio_slave_o.ack ,
	wbrdtime_high_timestamp_i => wbrdtime_high_timestamp_s,
	wbrdtime_low_timestamp_i => wbrdtime_low_timestamp_s,
	wbrdtime_errors_nr_i => wbrdtime_errors_nr_s,
	wbrdtime_corrections_nr_i => wbrdtime_corrections_nr_s,
	wbrdtime_control_disable_o => wbrdtime_control_disable_s,
	wbrdtime_control_error_i => wbrdtime_control_error_s,
	wbrdtime_control_correction_i => wbrdtime_control_correction_s,
	wbrdtime_control_clear_o => wbrdtime_control_clear_s,
	wbrdtime_control_clear_wr_o => wbrdtime_control_clear_wr_s
	);

	 
	 
process (BuTis_C2_i)
variable extendcounter_v : integer range 0 to 7;
	begin
		if rising_edge(BuTis_C2_i) then
			if wbrdtime_control_disable_sync_s='0' then
				if timestamp_write_i='1' then
					timestamp_s <= timestamp_i;
					wbrdtime_control_error_s(0) <= timestamp_error_i;
					wbrdtime_control_correction_s(0) <= timestamp_corrected_i;
				end if;
			end if;
			if timestamp_write_i='1' then
				timestamp_corrected_s <= timestamp_corrected_i;
				timestamp_error_s <= timestamp_error_i;
				extendcounter_v := 0;
			elsif extendcounter_v<7 then
				extendcounter_v := extendcounter_v+1;
			else
				timestamp_corrected_s <= '0';
				timestamp_error_s <= '0';
			end if;
			wbrdtime_control_disable_sync_s <= wbrdtime_control_disable_s(0);
		end if;
end process;	
wbrdtime_high_timestamp_s <= timestamp_s(g_timestampbytes*8-1 downto 32);
wbrdtime_low_timestamp_s <= timestamp_s(31 downto 0);

process (clk_sys_i)
	begin
		if rising_edge(clk_sys_i) then
			if (rst_n_i = '0') or ((wbrdtime_control_clear_wr_s='1') and (wbrdtime_control_clear_s(0)='1')) then
				wbrdtime_errors_nr_s <= (others => '0');
				wbrdtime_corrections_nr_s <= (others => '0');
			else
				if timestamp_error_sync0_s='1' and timestamp_error_sync1_s='0' then
					wbrdtime_errors_nr_s <= wbrdtime_errors_nr_s+1;
				end if;
				if timestamp_corrected_sync0_s='1' and timestamp_corrected_sync1_s='0' then
					wbrdtime_corrections_nr_s <= wbrdtime_corrections_nr_s+1;
				end if;
				timestamp_corrected_sync1_s <= timestamp_corrected_sync0_s;
				timestamp_error_sync1_s <= timestamp_error_sync0_s;
				timestamp_corrected_sync0_s <= timestamp_corrected_s;
				timestamp_error_sync0_s <= timestamp_error_s;
			end if;
		end if;
end process;	


    
end struct;


// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DvVI8N4SI5EAoQ2LFA9mAAVSZB5vBJMci/9ldd5h619IhXRZC6913ASfDgIoW4ft
xjUyZLzx+pTwLDKjZH6wKsBw2i8zIgt3a+HseBxpPBSxKtnb1jZXcMhe3uMGRdUk
76nkeHxCYBlWVt36xir4haoD2a59gm4Dei/bddkWV84=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 19616)
YOVFEL/alS165n+YgG+OIV8caS3R7lXYqePw8TXRfUZGX1uUvHQOqQuoK28jut4r
yDEz230Kd4AgH62TcufRtQ0YultPJAsbtzJ4975cX3xzg2aJhFjrms9yqff4Cqag
uWVzqnaDFk/UnM0qSTKUUg9K8QUxvXQoAGp7fvOWXg1BeSSyZ0c7WIuXIe5ziCvM
Hx4Q9Yyty2bqlnSyblVcXU6fBrcdiN0YpbAVi2A1WO3j4jXqrdoxGBe0xYMfLtXx
MELNO2lqlp4sg31Do45Bw1EwiiachW2h/KWb0plJUFaurFkYqeaxERgJObGUnJfA
H+qOTGFgaM9Rb7/fuDYtarmQzoifD6C6axfhZIKj6ysbHUUrkfPNWgnU/OP0NgFW
RSoVtXvRnCdtrH669eMdqeVaK0UfQcmo6gvvfTY8kzOkssVd2oieCvs05Kz7p+L+
csHR4yp4bBxVR/06dc7acK/lpO7k2MGPxe7GiMKJq9BYeRhKkRGKO9V7+PRoKxtc
QzloCFwp30RrCEq81f9HV02yWbR1lF2xkxZ+60f8GCP1xz2/KAkaMXKLKL0K4YI0
HnfM69XhzoJWKDO5Lw6gE9Ehma/OcwzU6yaLM5q9nCQXmx4gK4pKHjPtZXUZlKOB
i6BCaC63+SpfxN/ykP8sPChFdZrJGanwbDuRy003vSn1vNCB+1Db8IGSv9PDc1or
hGcPL4XhzyLn0Ml7F4rypvG2x2j73U1N8MVQluO18Gt0ZIsYsN01cKcjcn5iV49V
oZk1BSaANU/OeYhSWDwxH43ukJraaIU3/QBea04Bu5gjxjOKucjfeaimMbgD4lnK
S8GnoRVCVzSj+gziIQhr9wI47mbnExiUYnkoJkfrq5Han7e/DBuHsSX9hg3LT4sF
sWF4YzHbYXMGHzbSdj36K1kNrMxErXtm/8u4jAVbwgs4rMWGVy+tLAjxj+W8+grH
IOpuR8PIErLAyezOjUllcckPzHCbWo77zr9nst2DKEYALwoq2/0yXSviKZwgqYFJ
KmgOyXHmJq8Tn/qho+mDaF4lvHT1sqsMV34v23FxaDhJ2AzLNSiHcaJXxpazHx/a
2SOmKl4WyWhXV/SAqELgSWmwxlvNf3dggRd3qI7DaqH5eWFNYZjUJxhgWWBvc3xK
/uNjxw0Bxss/qWfo6PA543mPOtPKbuhJxjmOEB4xohO1ygvYPp8XxL6zYQel0hVv
U6pMHNQhgV9mn2oqkfIx6BElytJj29TJA7pY0rJxwsoaSqc2IF8WDNiaoVzRZ9n3
TvG9vc1rvRpwMgo9AFlLz82Z+IIvmC7rDuXWSzY4PGo5AmhnDRv6zZX+MzIEO9io
SwOFmkglnoA4b2fmPI3lHNAA5xw8R+LAWwa1TMLtJFs6YIcqSFNc1eqCyOKXF2mT
dAvIw9T3CUIDsA+DU0KryRUMNq5Tp4J8OFNnXqKj4LC2OPSu/14K4awfVE6E62io
AkYXuWECRmcUwIodSUhEgGPiFeFH58FSiKPVJsIOBv6ScpnFPpoia2Tu242sSMuq
LnhySLtQi+1CF0lGVQEqu6T/Wl+9cC0VER6Q8WRmL4WbdvVAf31+2/ZwF7ANxpeN
yK3R2mz5IBg75ukmkF7C3rlhwxMVmZ+UuSu2rRgIWlvFao6Qa4XZ2IKDRIfMFY3e
oLUqVuOvleZWapo+cGnrcbrdkT7ThOP3UzqbrEP+qBxI2T7gV2JP4Fg7FC1BccG1
7O1X6mNx8MMPbIm6YwSHndeWMHSZgMPiLPDFcrGS5p+S1H2faJhWoHdvsISLmDZY
XoR8j8kbm27WFya9RnMPraoW+p1TQqkB0a344FlwsvKkwqHJgQ3OzTz/sPaNCscW
mLUkMWcALIv+PJnNc6BlYHSvMckr5xGwuUbh0+10r5AVRZL778qlZt4ZHJNBX703
dFTRvzX+tXI4M+kh9F0R2mPzFBwdl4mZMV/u2qVEUaJT4XBaGxvM7cIg3XCHdk81
5IxSQjuKrbYPb2j1C+hLSlM24vGI0phP5jXqt03aMzEPZz3rL2K9IohWMpPyu4e8
Nx2NpkPepcQdIT7cxEtJRD5wonGWpSvxdPaWX+cfxz7nby8DJBEe3vHGa36MsjkN
YicGYTl5ET0KFVESmlgbNMW7hefBSx5N7sowrd07roDcfjGd7csEhUuuQMUm4S+B
FwsXhs9MxAUpE4FzV+Qr63klyCYqKN80o6I/ykiTh2GzAOGPvtwTuXM7I7vW5uiq
gXjbDOG9YiTuIW+L8j9d05NOG4uo8y/LjoZU+1JhntGgdj61OMBGX+w81DIYclSu
WniX1IAsaXxLgeonCUIhVG5qWrMXLbj3Ar43+gHMyti/5Srz66pG7bP2Lnz3D5Lh
iYSEd6zeMpf7FBkqH1ytnUYjwpN7GU427sPDX/bCdhWUtqjDM6ie7Y4+IdFrXwPS
6Um3EL+36ItP0kHsm/jRQQb/N9IDkMvbeicBgKG6qRWYRJoVYA8/1EBZLwUjYVjU
01Y4/yagD9VrrhYiP5mHnEnIcoCaqyXYi7dGm1vFVEYcIFW89pVKfeA2F9ZMM7cn
rgmRjheL0pNjCM26GWo/xQRq1aRp6O9hRAmOt3ZRdVZmtK7Inn/fpPiKLmdG/wLe
vsGGR7GBLzdDSASACieNnk+mYMNi3WSCKe1IKhis9xgtueQ+UO1bKlTGXzG7wVv3
qqs8R9babxRL8GSpSuxGnOWeil/7omHI1XNhrr666Nv30Oekb5+xu4QlDQFfxp/G
IPScXOXwRRal3t3vc3FxR6XR3OfA4XPQOS6o05nsLhiNzzrWQw0yzIRQIY8z4Nq9
sziujVJ8lagqe6roX0goEOfKp+basSQlaOcuVgQ5O6J1N0kzA+DC2TMcVblhA3M3
7vkfHDbQklqy6dhDWbw4tTvNW/66rVAvEK+wDPhek/sZ9LLFlG7cD9vKctTYPd7T
ATJxtCGkOOBBkVnePfhmOCQi1wneM8S75ks0jDf3eqO4furBs6xb3ZDzNl8DXhfy
YpSyQ2d7Xx+XONtqv9oNssIZ/NNJ+fTRM02gyQ2pT/2aujcjWWkyN6KE4SO0cX7w
9VTn9AZSyy9nwHryTw71fRc0m7e51w90DAkCvOcZL3w/bBdj3Y2fWMwIaiCoLpJQ
GHNBXDk+k/FaPqAjPIyVKSjAF5s9bD3xCPy8D90Oj66dkjc1hu/3pUkmWt2BriBk
29mZM47Ttk+slqX6t3Q+iLaFZ3hepNgKW6TN3R8bIji4W3BkXIzpOEoZu2BRK2UN
4payEDwCNu32XfAPPTiTOSmAgMuPcCjvDMwp26EOchpqUXA2gF59gYZFOsKjNVpu
zBAakVxPqmzxC/rdC6f43IhAf1eLL1D6LljToDbQ6eadHPZAJ+CiUFnn8t6pFeed
W9owXmG3RPEHllOhI4AbqdvZxdsbOcMjXsBQF/ktI8QtqnmCU22T3J0D6sVKQKxJ
iVxf/Mfmg1zgYxNSiT48MrcRwUFdM2GgQ41ZkliUt4STiArEebzd3cIBfbyiDgEn
jTd978PaI12U91kEWKALiV4Bng7ZiyBnvQDFPGhFDmTw90Wl8poW0xkhTjjRuJ46
osWQZ20ORulyl4AT1VVY7FHdzMh+hkQcJSXEOiakOghoc4dyR3f4ENGbxo6O3zjz
G6f4VYBvGOl3udvvBblf/5z01EUcs/+tnEHMUY9iIeyFJaNlBj/42s/j1L6kL2TK
AZ5aXcxGzV7xESj7u7TZ1hDA4Vk8/0IE/Osyd8Wul9f02obAefj7ZckP3TmQx0dz
QRUPEYRbhCj1bBsy27m//XVFzVWotTO8OMzuA6cHWJ4ZhuPer1Font6eUX54JBnG
hDCPRYtVlhMfxri7X+/0WkB9NH5muuLFrur9bgjfsjd/SiWqlRD3oBXrQQ71eoao
iHzWcnofaVLtKjIb5pF2TYw3GUXZ36VIGv1ZnlYzl0mwzecHOcZ/35hYshOwpFas
5/3dF3ZP3XbD/Pj0Tl3tiuggBSjjAT+fd8qc8M4TtkfH7Ix1Sh8iuTmjOcBKmjyt
3Qaexc/1McGILFfkd89o5V2MApoc1h20xKej6saqtTou8VJ5j/0iTkWLFJcPsqJ3
zZx3+u+V8RJ5QcNqTMzUyB0WkYJOQHYpYlJY8vSN7rwgpZkaBAlkI2GwicSf8/Pz
lZItPrzYHQkqUtV33rdQj/j38u/O7BauD1wAnQ3dLPJhAnNYKAcLlAy17nqS9PLH
xrmu2Awg7WEwUUcF2p9gIEAFKqFQmk5rLk50j4Eri8c2Cw6LhAhbMM4jEmIfngeY
QqUUdw1EktdAuXiTzPZrR7W5Cbq2IzBy2ksal6xd8VDuPfB137sPTnNAL8LPTgsC
wqT4ta4/zLxwLOwKe3sn4QoDxweiPP4AVhH/gj3NfBteoWsj8CvNEnwN5M435US/
NbhLbBLx2xAXsPlS5t1DFKextrWBuqeohMS0Wp/lEZWzbc4nbpKFn/VS+Wh0Cg/X
prZ7uZKSEDZiw6meV/aGzkT8/Q4GHQCH3H0ZQQvOO6jN39neVVCdG8MzzFTSXk1J
zpQdFdEN+bEhWDgJv/F0MM72z5LDmzrRqg/kG87yOEpfiZGymGdJas9dYkzWzHhD
WWvY8oOb6LdnBZbiRbgDUtJOPbE+L7gDeFOxVETk7074oo34opVs+BweffSjFHSO
bWeY3UtzR1oLfAl9yEgKdYOaNxH0b+Jg+FbjZNafUPnk8pYyhiLbaaNGmWKWpkMR
0se7whpdm7P0le+mgBvJFQpeTfUhaxlVHR+YaIAeD9VwdnboDHv4hXJmeerrQOGY
9WvDWt/zYGM802VsQ825uxF57LvkJaw9cynhhiOPYcuGHUqvnzB/CNZFPWV0QaIn
4HxbyaE0EvBqCr4RTY09hKoW2QsQBzjIz8Zo0WJB0q3YbIvpazfRNpOQJzez21sh
qTTFoJIJBm4Off1LOKA5LUQdtTaH+4ODuah+O1hNAysZGEvzaUAvaPD+0M1E6aTV
Jsu5viNG7xVmEXrgv7fRh0p7TtHdXwb6ugcaO2p8H8Q76zKdKihK/FmIzjPEw6Hc
oN/JV+T384z4QatM6Yh7nVT8iPkIN959bEJ224BE+DTCXEUdE3PsIznXxcwwXKSO
hAVUbyLZvNmayes4XIhbaIloq2yYHwg9R+DuexQ2UPPOdWRXo+++ZDFWBzt+Uwby
JhjbYNdIwa5ec8HlX/NQJyETI1K0/xhea75yLozinuAoH6BPBuefbMwELQycZ36o
nHMYMrZA5QYs2jvU6hpjleyWyeeBVDKQfwlkLhRhd1suTxCzYGR3rCcputlO56ys
ioIHVqXWFDfffOIlWkRzbKyhpIGhoJTI+pQ8ucqQb9meD3oMlN9My+sewNlPtkhM
6lAxBTuUilPTHgUVmHhuXu6AXQGoMqUvBHtKPEveQHCdo3WJCWNJvhpelNcI+TWj
9kuFgQfuuPHzNl5hClwmfy2uHVybxpBvsZyThscRGy6v0s1ZVW/h2NlqZTVa7HNs
OapTBKNTmufCCYromljjGtPTfm0uMQwroJguEUbvfU+8mrQHou9FKWc55Tx9eZgE
Zk510H8Of3brr1uINhu2uVaUQ2pvLOzkFuAykzWL37COqseNT55KfvoPa4ifPBXe
24eatKD51/NDPsLtXNoOKHaNovxaM6s5v2mhE8KbYSpPg6J7KuqpiPiDc86bYtnj
FI2fsH6HZxTGZK+kwoWGatTGScgvgnP+eIK129YAL6H4Dm4diaFU1WbZxvJCJ+KR
AOcxExnQf3gPftMJjK/VC+RbvwGbPoCHHUX1SH2Jt2LN1rv4ouoPO3riuzLdvyHQ
3lF0VsFK7970WqhOWh//QVFEMrZV9UsSl7B2bJsB6hb7lUSZGQ8+ACqeCuzRMlpP
8nIYUIAMh8Ev2dusODaPh7mgsq3aavoRM2+sDBfft/HsKCuhWdw6u6KBLzKCteaj
Tz6vWbK4krwD40SNyVYL172dxNJ4VaqCGKbwNmGUXL5FAGRP5bWsFET9Qtv6Lh/D
yJEk2y4IGxpKHSFgu5T/xqyfcN7WHkSPWtNN+QWG5hIRJDkFLUb5p479SRywzyEk
mrkv76lka+KzrgJ9pwtHV+w9b/MJ6PrnJHN9qeJB5KccrtBiZUXe31XllEFqdgG7
PbRcNuOBt2UuvdUtenpFTv5oqeO+b6BN9DK2MIzgG3ajflnp13+oi+wdm0r8jx1A
fhFNxX/5hv66kY4Jf3YZ+aK7hTWMBwy+3VTxpeMbshMp5s2y1RLXZ3V6TaQmCGen
nrwLlhoGzYLy70I+rGQ0RPUj2UvwWRUZFfkMHCclZW72CeO7rLQjHLW/srSGJ3yU
cjRNuZUECtORMDgRdH2aU+ZxQEirMWsqxgoGEXQg2jlbyYTasHCkrN5aSfsnwtyJ
RC4WZauyHd+uWKBYvLVoZuUzGVc/wBT7yJ+SMqalbabXJpOJehlt5bEG9XJEaVo+
OdAEE152vmZtD5WizCiVCyjZtcUZLQJ+GLF/flhO87muOCK8n2ST7nkOavbixgVm
jOnUGSMy9URp1pYcBwAD+xV/XqJfQm91MCYGYisu4rDCS4JUkXTRxJgPGNXeT2ou
2c2ioLubx7WLk/nDOuj2KmUsuzXA8zVeAHXR93nHOW9yzdOHaNPFBaYNhyNoXroA
/um0BSS21BiMeTNKlCQ/nLVT3e1tBunPiATXdAqIjA/KfzPB1gcnCaUj39Cpgzl4
A08vgpuwho5dJgOIYQWkBOefmhWwoY2D7vwpNh244puoYjURHbseT5cgpRCraXkK
KTo29Wga+MwLYgyil/gKgxZjfQBNIhm/uhe8PImbVmI1V5Lk/v/jWD37d25Bjqpn
o1TJw2TUsO7efLOnN8gpf9HuDSf7p3E83Rj+zaKduOCfBSa+m/1pz9AMJCRol2uB
gDzdRp1dTSCIAiKjJMjskj6BY9RKfrhpsFWSl5a9iL9Cwi3HNYY9Ie7nKpVamsh/
ZarwwzvRhpX7VKZLSDiJj+PvPPZaMfkmG0T+oUCujN39B0+8QBs3obg/WCBiHK5w
LLX2YlYTicG/fDokLOcLDVYjOpKmCJvndtmgpEWEhTVehqEMYN3jzu3uUQqRew15
WkL5f3rJ0KVn8rCsOnpgPV9zLZJDAMub7F5kSx4oKSbcnaUBqMZSSzZ4PnKV/jlH
Y1T0rywkxashbtzmf4VZ1znv7y9WuxJmX7HjovCvAl+Mdfh5WJNEuSnvo/cZCD+z
zW+MVq6fWmPspM2ayuWp7a3sGDVFkVvGMOdCiVj4h7kWn0ekPYVW9VSyUack3zT3
BL+5ClmHSiT5RBQDQnBGlGHqRAQCpjjgxgEOh8NbwCVPg5xYInJDHRhhpSlSroYy
QOuxGh33idtJzf/kzbIRGQPvoxoqCSPks1fjMFeRBhEvK1hhmqC/B0qn0sn/HaNj
o+uEQNM7V4+kr3puagQcCbfCTBXqs9RKaUV+N1M6wEBnrLOmypNdLZ1whPZ0tDgK
XbEl4JJop8NgC8OOIi4PqRr9jJ/u/SRTOpIlYYF6pb8uBLStn1PdnT3kNuF2yZ1f
J7iXrGIQiohdM14ii4X7NnhsElGlsLs1HmfETLCJdM+TPnODggJuOpYtkZMtZU9L
JspCOLaqIWH0VMc81+ZuLpjNJpuBM8PrIoUY3cX/J6zw2L7cBT5BNUWaidAEvz+M
Mr9+53/BlxUy4rztjrOyQruR4PQUxJTLmKBefSHQ+OZ6ULdCzSldXZQ1jNcMNcry
dR9vtDZh9ZIWZxQCZggkIdYrrr89k5EU+eWbrjO8FiDcvim1LPhAvAftQbibggWg
C1RfEki32G6s0jObN4+IW2S8eSRq9iRycwkyBuYUj+aK+w9F1NcRzzJihLt0LVNp
aFWslh8/kr/VoS/beECvDt67oEllNIiSqnJp2t7WQ3YtxsdT50KNOqN8oMva+ChK
HjhL9ZqM2l1xvQYAwRmGf1LcyL/rOYEdl3dmoyVv8cBXN8Gla1Avcq6TAUOh+/li
J8zzfhJwzTm+VHW92lJ0Nz4q4IlW5U2QFoVVgDq6mZk/S5u2s+/Dv1EMTge6Hn3Y
Fk8VRD32lKmLg8h0dCE6V/Zjrmpr23WHX5m7eu/ZPdVo097ILpaLYVQik3JdCgiH
FU9c6y1Qzs1YX6eoTysPzn7kb8mtibX2m8WnRXkIfUnX0fnu/CjDI724y5hG+rN1
ZnxY1EGV9BREW3g+v4ICCXfERR2FhOnEpf7y84b3ZNEQME6HsYxtea2tTyPkcapq
OA/TEJ04fUfxonIZ/PiUQD4N4P6vP1KG3oI4yYvhiGaHQcU7nI52qoSfyAHmc/oF
LFx3FRn0fQMiwHaBLhCnVT0DagK1+lDLI5NnZVcCv5s7ttAM20tk5EZaZJhuK7WN
0lw+/Zb7Qhm+Jh9wpJmoLOLJuiHsixPnaaUY38JSJjjzBM6Jy3JyL5XxZZA8a7wC
a7Nk/tTjg5Bnu22mSQJCE+NSUEtlOkdpOzxgFWvlIbcZV/FlR3vxO5eoqLdJFd2u
BDpgh50bmn/JC0vuWWwIzAycqps0Ay1SHls844zEVI73Z5VLiB/VQIgjUJjgctQt
NE34elgnXDLpZz9NvyRKnXG+McqUnS0pE/hJpTHlM56ifJYone+tlF8kMssmBfjr
Pj5aqhK9lEzhPWId+bzSlAJKLwfczUG07jRFuABBEX3COO3zrkxQqaL/zZOx7GSl
LFXTMyaZVpdhlN2aTr67RIcuVmcigM8KHOkL0TUKpASaXWMA5XioIoRc/noiOQKF
g4kpQMwYILEqPA9oTjq5kNSpeVAt2kpD6jFAvBg/HaABLSYpRyEQaicBrF74CU8R
IxBe/C8Pi4gUv63FylIeE+8f2Zf3yM7RwHuK7mf7/LCMikUij+4GhBuW2yh0fYkv
LE3dul9QApoCcOIWeSrqiGFzzpWAfrK4EAd+DNBelfj9KH29jIOGmAjbw5thGQ6f
IqvpnnyEO/w5Tr5t7F5fiM2U28ncdnXJHEQleJvKjOGBFiUHac8QxqjSr7QOf7mq
/QLttBqyU93P/y6eIDpmOIwhm9Aft2qvHxeGrIHaXX4NCVv6gnlQrhmfPfM3mzPu
H4X4e5RTzRNSyZ5DDz8Fr6olhrVWYD6En6+Ibz4bfZlvYF7L2RLShauKmUkKkD7m
UZJfhFj9edRGm/C+65PW9IJkg1DIdPM+JQN6mW9PIPolbNU5RG88+nHJlR93swJ5
WDYHCzV6ogRQlmY2qQuyAlVGU9g41zTYouxtAqHJYrrx2ny07TpZ1SmFUC4Nvd0w
tvy5HVHmVSM8oHbF51nKY5XktDV7vQmHvg89QqODyTfdUCo1Zb56qJcy0L/Kv5He
o+XSGYhUcaKkngZY1nll/H/7AbAuSfH+kacOmhv3U41z8ZUd1Q5A0mdb5fVwCeS0
CLjb4y3uMO1PsycLjKFZ0oEvz6Mgcsrf6tMkgNcuymU/0M9umtKkuyt6u4bE2u07
HqNHWMYJJqmLeJsgDm7L4DC9+ep1U4K+1mqRxHqlBqPEqRr4UEoV18F9btqNAV0G
Jjp18nohlsB847yvBNQTsiK4Wass5qp9BxCZcFokd3U4SjgBFe1gshDH4yy6Bs9Y
+SdaSZevufKqUXMOgo1fiESane08+SA5aLpk1kscHO0x9dHEQ7/pxBkEw3KuywSP
TstVzA/tUOTf2KFf542D2EMAyZ8xKZb/PAmWYU0Y1ksLlArbgsugNnaMtcPQ7ONq
Io5lqEijuhte4xv7HC9stWS3MqTWGcph/cPJUGWpvg4GCjgAu9NoYNHrAnqdRyuN
ZLPzeP4BUsaOhpeY2hs/OH01Q2JxaKS0HurGEMQ+dwq5s9s/7WHhJEfwFHyfdR33
8yeav4id6BqJPxmZA3KEvWmDiB+39Do4eQRMVYg/rvkR6UiG/eNVuh+A+y6VF6Xh
hetjAeW1joSufghmuxuZgGoIPnkbEhisrt2hjqnQrdi+3DmJC9aqkad4q5JmpN62
Ck3DydkgZWTSZuj+fBqbpiFJ3EFFSFzRO4rKG5J6dpjOTEO7BDF4z0nQUxs28WSQ
YElOzcPnXhsPUT37d/Xe8LVNym2QEdG/Bqv4g4MbBmzqZYQIAoi/OwHBKfRMN7w/
yxbEDSiKyH8G64tvVxtapINkDP7bCc+Qo4cXqPuf7WqWo/l4SfOS5luQdCmdu/pT
+L+Z3lYQuNBmIQ3ORGYLenwrlmClfSVvd54vJMID7zcPoyn6dafX2iq6p69IyA8f
dtQ5+hF2zV0KY7EsP0G8zNcAhZZG7FWDEhFPRgjBnBofMurUhrViymlX4Wf16yc2
2WPq9n+6CV39/oULIN0gIqpZ6t2AXw/57pkb6ltqTulRX+fcTcaV5KshNGd14kiS
Vtu8SJzuUoWm0L/SWcaIKUqnm8bmi42Ok//+uLy+IiOh6ChGfSpKtAHELCMfAtdh
VrMgAWfvUPuTDEWCi/Ed7fNFgz+lViJH8RJ3FZCLwYglfL8Djr2K+GV7cs7z7jk6
BH7Rw/27sQhxaVKnBJ7nMockt8vwFvKM+uG16YkOa0ly8H4Pvzr/JfamtIZh99lR
AzeAgFFm0H9uck95nO0j1yqxs8mXjFhBNZsKCg4KolFt3EuaQxbRLShvJ5LvYnnp
C8ExxQT7QdnVsDnX/wO8iyEoNHxZq/K/mCpa057be6mC4WyembdqtB3JfE4n3i7X
Q8be5NEygOEXqcEYX9TKfxjhqF+uLJ8DFyv1/qOb9WbrPS7wQAmbM4d2MlPTCYUI
mfGj2DdYUw6qf6IIi/hdC6RIu54mIEmzxP2Gb/a0Z7S4LRC1G/CRZKB/WvZGZ/z5
iO3mmxbjV/iZROBzUn+CFmc69+yMSg5f6ZYaykdgO4qGH/cFUYv+/ftd+WgHVx46
JaiuZFzQAl+KGsNB242YZjFCAa5eQtDsk3uvAje+hmoTHHhlKcdA3NDnncrAq5yS
MFUroKYdfPx8vy3eu9LfF5nMGiQ5/DI9AIGVOnfyY8lB1djdEBQF1Z+fUZv2OTx9
nKHovyC4MQQqNcgZeaCr6+xTm6Bh0FN3s9kz+k6Xv0zqUbQoSHk74L/gtptZR1Jw
SsZgVYogeSSHjoETCZlfjp9clfQqGDt+lUPVK/+FpEqL2zs5gsGA41WPlojfgBcx
QKAkB01t6m92qI2enDa9pZjPUhp+6Z/O5SNYKtnYTNxgJIVNEEHFZ0bYekTIKD6Y
/R81TyHHk1k7j1SL91F071YJnfcQX8j9Mp7yaIgBCHkmdUnNF38gpUESys+UT9g3
cgqI1B+dRzVcMCeIqYO7BMGiFg/ge09/GOB4+JNr94bgIYKVAZVoiVHeRn8lDPj7
jI/wLdw5wYiujTj+E1Ya6JVsh/PT65WMyhrupQj5dDIT8XPqLsf25nt68xihaA+J
ddPE3KnqoQYmHGxmWYe8unRxIAOefhfwVW/QJo3xfEVe//UdgnzoNNyO6YvHwRrO
kxSH9anu+NN5J9Q+gqWKJm50IZ/xmechytxS1a7ibP+Z9+Mg2V2escaEHgXyGw1S
Mbwjeg8A1IcuVmSxz+M2xeNNPZI2DZ6nXF/m4FDoXXvO6p/XPoDuTKmkUs9b+O57
Hk6iU02s1nlqVDt8GWzNO3uKukn1rgNEKDoO6Hjw0tF5Jy05uHVwviLKeHwyClPM
x0wVG/2vzsfknCbU33eYxbib1rbp4/O4ik6q0I043B5v4LBzDaMCDFybvYYXKulT
WUpn1+y/+s06QKaXYfq30My8WF8ycYFuUrOnRQXftwEeLsiQPRuDT2RlncGSwqBp
ywc0QmNW8ceCcU8yICj6R3EBIUmIEfiWNhujb4e0wWE2fL4c9JmHL8Jaa2J7JLfs
HVk6hPwr1GeRUqwcOStsuOQ5m2+LV10OFsjQu9O+QkpLhDAhc8ZVUwWiD+agSd4F
kZWTuSldA9uM+tgSxFV6a/SbqwCHEJOO1VzTdU+Ma6wJf5i0cthSeL8lqQDr4z+N
bHfj+8/NjHR1KXo4mvi42dWHVFpQAFdPANBMicHYcGjuigE1jL4h49hP6KuSUrjV
L9wy8MkFdId/DbsbzqhKjlFcWoFbm/e5BoFc4NeKt86W8uUrqX2TbefN/RdFutuW
ycaRuGF3amtc6J3+wW7pYvjoyvpQ30QZoGCvlucytGErCEocdjvqSEbmDp7wtDdF
0PGT6DyQV0O5WSBnAej5WiEi9tlyp4ha3z1D868mVs9CopAVAxOUGpqB2M69s42i
WehBb2XYqtGKtuQ6vDAvah/3i+qPg8Q8hvE/r5zzeXTNwOW56f70xJizgR0lwXmd
BpYqat1+2w5gWb/0zF5LF21RQRSnq6SD5KLPFc7depN2GN71eCuHLY695Lb0IYWn
ah+RqXYcaXdTz4ym0Dv4SdJ9oKnWnaloknc9a99Mjt4UHntIt1QdwMdEOgsnI6cb
mNT0yYrJ1YNeFXoWG27U4nI+vNr5+1PGUU5m7At33NDf5lDkA+djMD/r3+5vMQQ4
+WG3xcOxhLjH5XT4tmcb13fADw+IqEpvEyUMtagUYh4ovobCZQV3qqhCDKZhZVpr
BztlWiaXMJnmGvRjyndszgGNeJ9T5sbGXBZ3z7XabsNbNrLP3Xe49OdK7tzdQ9Xh
gpcGmzOHYJO4r9PTyHN/taRcszAvuf1JUUbfvDQr4aklLU3J/LtEyNDg6mdEnTXy
czqUn/R+mT00/IUyIEAgT6nZBNMi5tU7h/AUH4xRimTTfjUUshol57w3TBs05Gqp
mPgzsyI4Z4JlWsJIwH0YMeXVxzXOenckQC+I9knxDYI3IFY7t1EtWPcgUKfeFNma
BMj5JbyeY+zybeu3BZLrL134zdw3MWVOBH/aTc91yVcQZiV/HJBIkNYbEPl6TJUA
p0i4j2b744rluqzl+/ZRm7No1lsGv5WaQ/LuEYgn8Kljy5Ey7d1SkSgIxVaXbYRX
8J1a98AVdvTG489BM7hDBkc9ZxCuoKXL6cluQK4DnQILFgxb9bu/3KuYgESbB5XR
j1KY3xqU16p5yk7ZLuy1mndqs8o42Lc+ODU0T1A0BGiQNeawymn0CmbjmfJp6YEX
suPfiM4GcG9CsUsjOTrse3KemQ5daWZ/dg64JhJgZZld386W4xKqeCBaquIzNps/
K1xJYiEvYcTqbIOmFR9qvdJHL7y7SEmYWi1ULekzm/cDtFLZOr5WWSc1XB0AbmHc
kCuw2Ik8PFR5ckUbNEz+6thI5xSPPX3c9HyD92MTfza3lXy4qUxSszbFG6T/EX+s
DSVzyapoIR6i5LTE2n4aw3ESskAg4GSyQOQ+2UGmXtbqFoi+5CraxyzKrNjpKgDu
S4nQzeAC97oGIO8QLFw0VSJ/Sxf6TGcGNKDn0VX5/RaJjTaBxOnotoZlvef/3prB
67QddFLOjiADGb3GLpN6JQSXR7TXE8Oy0CQ6QLt10l7F5evm8jkcBHYFlbFNKxxk
HD1Ew4Me+3HrDGEBnb3Syf+MuBCmsnarou19sLeXF+LorgNdLXYR1DQWlHVuvm4B
jsdbQWN2LFYyvxp6jpbIUvMBqTrxu/MSpRCc+jT1ajV1SKggGdqwoquO6ilhQe44
OBBDfVAV7kCHubeDG8mfVeUvRe5Jb9Ju41pIll+xgCb9mcdyisTGE0JOAqdIPXcd
hUiQ/dpp/20gEgbgAPrjuhnfd3y9gSs075jstvE7mmXu9wQAaZ/ipoh+cahiuK0i
S7For/hBfOeYdx9Gq9ORDoqDtNZlI8hDSFqTdGqb/56FMs4KrCT1P7iqBEexADW0
pYwBCVokI1zNN8mxTdHgYHj8yURur4FsZ7QYZt+ibfBfLo1addPl33JXb0yrEk1M
bYAK3BQekaOqPXCaf+JSbCBNWid8YNGWII8srLbjL3lcovWYeykEE9dw3LH3Bb8n
eXoo/uaJYfEkvuwMmSk3bzQl3HnyPxXUHeN6YTCVHfcLNzCaBumgUJIQc05e/M+K
jWTk97X74vJEYZozCChwM+HkKx4YLuPwISfffAvK3a0Cz6sWp6vlrAi/GKof5fCN
lkKuL7rZVlFtZceXpqZvo3fxSxuyf++z0BS+lbT4scEmZy4pE8si9AMmGikzE8yd
1xfWd68rxGLPzPsXyrev/fHNYjzwJtMng+BiC/3P6zApiAzkLlRyrrWTOsRVtgsF
ceMTFsZsAvirIHUHEUcuC/zulrmiBC2nvyUwY43yP8Hhq28KLJfQb5WwIHBshNuY
NrXmEKfOvnZq/caebllj1NU4h705ljomyEgazCap/MQAmo8HyrijCbM3OvFEMtPH
oXFsd181wXzT6mkRfoUbsblU5s3otca9PW36Z//uceXIUOTIuWqTQEHNxwQ8MT6l
S/24OSXNoCBMELxW7nGNMTrpzBUlIJAJWQQ+7wFpHxE3X29TKnqNovjsfErgj7XL
Y9BtnBvOTCRGcj58RrIRPYpCTHpNhAr54l86nj+m9tNpkGqGU0BOg3W8ztlvzgNN
kxGWzp2rzMgYllxO/pkqR6bwawmYz/KbHhxOtbQ2vZV0tF++uSGr7XoVJJKxa+fU
yOEHhaSfF551eQA4FQef4dycIDZsIpdUvXBPTP6GrI4ClE1owqMbbUUPDoDQZosG
2UBgBig2xrIWrniySjh2zdKIwkGxaLrFLJfS3mArUM81vhHKQ+ZS/scgBHxaIL9S
ZyiE2OTwmWxhE3Ew4Bn9kpjaJL7y7f0NVrgEkrFCmUb+2ipXMlxh6yEQfV+zKCt/
ZI9ezk6yphuHwpP/Qr9D6uH6al88UHhxyi5g75StV6Kr/teGz8LLVu7VHAZDWVS1
R6B1eBAZNdcf78fMkXtlSc6434HXHemtnm68uGgTXpl79xTDIh0h94Nf7+5XO2Mo
2aNRuc6n0r/Stxglra+fC86QGH950rSUXOuE3CQ2RbjHNO0TIJM+FQfOZRnXMnQx
QziWAHNw9pr906NXXXFKb2QZr2xlIWNH9HU14oJZZHvlxkkFeJD2lB//8+GzilDe
Sb3muIhjlpuk4em1aI4vAZzHSRA+dkAt9BJJUgLmaE7dPmQQsFXaf7TsCffzYIPs
CmdfXoNl11FLhGL9imzu+KWhgzfOGAEyYszfCuLphSwT7WYUXJzMFSv39Pfmfr7/
GzHAChEurwO4m13a5D87FJ7KkWPoUtArjrERD7R9ZjyGqlx/VyUomjpNTNd8KFod
1IN6gSXihBRL5THKOtC+jbOGfMpejEc7+RfRl3e9E1h4DQpyB9dyO6aeJU2SSq4A
+LBfvq2KhPR+AeROngM/ZrN6gAOui1avK4F0ad0o8B2+zx92GU5LD1KnGZ2wICOD
fGgdzkIUi9VDA6o8ZzHhoJKzGYae0nneXDUVMfd+0IukSolnI5+T2xPeUURGCsmi
HW7B37gdVvbDJt2KiCrpJd+buFXTbet9nGgeF65dnr+fez8siBj9/JkkGhe83jUm
VlEO1drAEAjUiZ0jv2XHmy2BolJUCTD9zTmE7nsbbRGXwPedWAACubGmeXRU2WSb
whGw/nQAh3y1SNp2ZVdaPJsj8iJ8IDYWzNbtc8iWiobwbBq23GCClGxzEsnJ3izV
wEZShoMgcKWR4wccjUMbTA6UpUzBfcTLdLTviHc37oPgqSL4Zs0cXtSLXGy0YoEc
OfUmFsYAMGHqTKAHibxdRcLDonoHY10YLb4AuYq2V6DX2wCGDAQxBsLJfW1pRW7b
g9ukxi/TtWmQuIBVnbI48oP2p+/2LABcEvqE/Mz/Aa0v2ZCgUxog5OpBCwG72GbY
MG6s7CCxS+npUIQrSw59p1sazyEPhA8gZEjAgcIqw+ZPlpohnyWBX/IV0KP23Y96
5sqv02iSCPqkVtPqFz17Z18ZiAnqEew9ICstxNAM1cAlw7NOBjSA/YtvpU8D3F/r
pIaBBEz6BD35ObUrNunCzvT/u9cCQnMm0L8xgw1kLEXy3wu5Y5Us0AkV/r+sN38U
vkf47MlqU+HpIBwMYX3I9/3Q51WvBdw5WcmBjLo+y5EPqgoRdT9nJZzHrzdbuhyW
6/rXRFN/JAq18AyPGXlg/bfa3qd0dSNDFFZXTWfBIvXVwJiL5CMMQVMvntJg/F8n
RX1bpm706mJ8AwhhOPZN4CoLbsXwzCZfXE3K6V/VSUUBmcM+i2hscqFTvAiir83E
mSznbtFr0dP1Qdhm0/euLpuIs//iwrKc3hN7S1eMkBVaKyfhkpi2s/+dBpNtu0pL
nuPHrdcSHlu8ceoKm7CtYV1mdWW+I9FqV/cL4PeKI5axTV+v1LGaDKpbEQQ2oWFa
SaCuECBeUZE78eMiqYUoXyq2hNG61qK6BSBin1AW3smGJnh0jN9A/CLhn1Bmw210
ZOvA/0lIe30jxbmg39U88VzQbfPLJX98vBKFFl2y7GLMCc7S730Qpxuudy4w48Dv
iL9SxAGZNEJfFfWJXTTkwazXaXz4k4zJBcwNkvlm7SjjRf3nCo12MiYjN8QaqQh2
Z7CK6YRGRqvGqxBQ/LeNbJ++r0NKwW8nyz/TPPhoT6NjinV9/UQLMFLIejG8+07C
gkAH2OVvpGgcKOuKwOoP7dYi8yzfXRxVOED1TjFqF0nszYXWCCF6cFCNXXk8ZjE3
IkKBAl+qvnKaiRPo0Vvf0FHNvaTZ5AhlmACh28CmE1CObO080HFHByFuFd7aTVif
6JzvC2KNrnSIUpdMkhqxBDpI8zHf5bHM/mSJNHxqxE4V3zIJq2Wq4AKJNCDlIhne
FCWKToCb8RaarsU3xH4FrpSl/w8heGSwm9ACDTS3It4a6F+krJZIlZ8fqHAr4OPS
Gi6g7C3gaygD2i94WoxtWAS5guFbLplaqyXB/Zssz4ncSWHw5rl/ouycpsOqjqDg
80ffm4cX0EUJiQrb+uyiddoo952ZA+Z1t0vm/J64nhYwmM84QsLfd/RRGJIqZRQg
KJQ6vgQJCLVlPgTqS23N15vBgfIxmcYSLMB5nQCTIyX6yir4pOGGhAV7eXgRwvbV
FpttQBkS/vB+AzHZuVsLzP85IvCljyNXu2CjPhl50AYkzFBtYt4wohiYJk0NUq0s
FGmr3oo8R8cIk7/G9kbsKWFtc51pKIYwPZKmjri0tLgnJOVI18Bj7lZWGjp9U7A4
7ek7X9et8ZscfAwUPl8dhXQRuXAy8jB49ChiLXO3gi6I2d+pn+Ig7sV1MCj33sby
oy25ASmlJUtfDq/fEmv119+9y8d+j9kbyVDz6SB8VK0gDy2GZd9kr+RnEkHlggqd
fLWxux9eThFQErpZJBZrRa0UjYKoI3POxO/w0WB1Q46h8ffctlIMCcHFt4xoq9GM
fZEWFq6DSzgPT/nKeyYwlx72c7Ln98y94Vb/APHpoO85KYmpxYv1OmLBeUePl3Vb
R9Z+Rhb0ShV4IIokR1n9zomq9VfN3GWB6q2tHVZq+DVj5p2m02vYJeREdIN25hAG
V7KUEjC1Nb74PNAEW0k4xMnCK2mbF3giPGFYxpKG4YFZkLddTQRHVv3CBf+KAEfA
isGaLvFHTTGErzjfwV7+xZLp5jVJYSXlb6IZGalqbw6qJqO2uXdT8D8sCGGy+3vX
Ss/Lcz8FY9htLNgL4WJ1aATTPh6eEmF2eGVgTt9Pcer4P3AcOXpcXT79ai1Fpjml
m5YyY5mtgiZh9cDFTeU8+r9QxizEPQ4RibXkeqagt9jvcSktRqCnKc6OYPi1NRe0
n4wEoonDDUiAkiwO01bvVtMCCRVbLe9be1XQt82DlN2U6sQScmZDRQ7Nt+WEtb6n
cFl5wuoG6sVsfHOJoYEAVzZ95q0WKsGTs3Pg34V0xKshbGsHh0wR3bFXzYtoA3As
T9mQPn/fhXvmCywIPPS82HVAao/YNA4tkqaf+O4Sx57P2iHMCN/2f7VyffLB3o41
NpG01jG++Ng4Fjo2/FBTFFJeuNeVixCm1FnCHmnfkl9gqhgZgucp/HBGd5kLE5+p
g8vCITFrky5INJalQBTuuBN0JivwVDrMmyt5K7ZP6nkDdGY+01FLO3ae5X7GT7SN
GcB4QDx18uTHZQIeqq7cfeGzhtRMtqdynSdysLLRLQo70NvA8FF01VAp3Rp8brQv
+NVwh+kAwaF/UXXoNXvhFiIUj4WSxlyybgfNK0T31ckxie5Xjgp8M2ePttW41nA7
UFBfbutXVNH3bxbB8H7DU1MHEbrQLvos1aJ+lDK6SLy7rJPhFLbAqvMMG8l/IpzC
Cvn09m26spbkr/A41+cFccjxTn4siLuZHOBSDT0cxk6hw4AIWS+fT5++wQr+q4tg
T+EA2yLNJWiP4/fVO/7uWtztG+d/IpcaR4ceu7jkyJVlb68vccnI3T4TO/5K8UTC
L85TVNewvdi4WwY6KTyTZW1ywE5GJ7vy1su4V2HFIqfewQQTjOFLvfPHWk/75CqG
p9TogvfzynpjnGsSt0egQeztaKwp+BLiZLNE0J7rz7ywUmbhS8QCr6vIeom1c969
lhb0AkC6AXKO+J+iaBf1Z3qFmu3tCI6TuFTz1how2FcMZaIfwcjinly9zmV4SWz/
zoRBgKfc/b2At8BoYk7u0owBWulVKB4x/mGNHyK5w4a2isqv3L395IAOmWcL/BOd
vBIg7zdgNeZnkH15JRdmfWMagL2OgAt5oLOjATfzwVaCyRcwhav4i4GwHyAOURjN
7rlJA6OCOLDNIIJgBd894zwKIP2+4GnTNuUOaXIwcsNfNBrAKYiatL/NzHFCbbFq
9uWFL3WZrUnyXAA4NzXPZ2jlATvjyrpb7TXy5tuko4Inoe1poi5fwdiwWLzrwm4g
wA0l+JKxvJ5eE6gZXsRlHsUoPif4oYUcxzIUN5SP0wM1HFDMqePqHk46zoC8+srh
xtns2gwpliGUFeDMxEU38JuugvFLs3wrURrAOGox6IvG/s4mrlussQ/EDiiu+hXj
9T2EK7GnC0pKWVLtBIERyAXHpXdg06r8OlF/HO3FhGuQT2BzuKVt1wmwRLshtYdq
1iCubvrd4RseAac1oO/EbLnHGzGL0jDNBy887KZsGFTjEwlrFL6tMIxPfFb0yhC3
mpQbtuL9sShr8IzobR/4zG64D6gSu2JAUEqN4KZvFk/Uig9bw9KgJBqgejCeaQuZ
zIeoEgz3ZDHKcM2X31i7l2wVC2kxCAfG16d2xxcHTY2ZNC69LoVezF6R+D1sAQBS
xuXaXbI4+NCOi3ECVOpsIp12vvI3wJi/V2HGt51kpkz0ovoRRxYhn1OtfH4WleCI
2kLu6nsTKAx+Z+pzgQ06o9clLE3VYsZAucbhLxVIPCsyps8T+7Sy2STyoPBPBv15
zQookdQ7jBAS8sJEylY2ivBH9tiTvgy0UR20+dMHx5c6pSIAvDRXUI+vTgjeDGdg
urRyQSusNgJlxRtpYJsa436/Rl+LU73UJPYacUZMan4Qi5iyozzED5KWh3G5k2NG
4tzNgN6/CUYvcmArzKR5ifvb73FPCOOJCwJ05TnMuyfC7/WL584MZnJl8KgK8Mam
9lq5jPsOxdySwkQ8Tql4RfUpI7UTEK91b1pZEUCG94gHSW3WVDMeV5e4hyRsZjmT
goG6bia6DOKhW3PEAqYld+1uOfJpEivQxdptKoST7O8Y75V8mk4D9MJA6gG3LcQ5
nsQP2HqFAv0IzxHrbQlE4PILJPQ95OevLFssVWklyV+SZgFAPJF81egM0R/tLEL1
8fu3d3++zyUkwh2quAp/E/KOf0hiv0o0ngskdEk14IWM54YP3e1RzT44NQNQdlq9
A7qi9n8o1Zu8JwZLhowbG/5mDSWUSRjGUrUbeQZvPAIsl3fmMx25aVMJ/6ucRs/U
Sguizj1sbND8kSExlgXkqnQgPK3sq5rjE+2JoO5aovLWCHOIK/IxxprdBQBdwQcX
WFQ4oX9HXrIEsgfvt36FSIckTZhAcuucCNxCR7n2bIn2kk2u4Il6JN+0I63kJhQu
wk99N7+0jzCh9y0r0evYEy3Okp81pjwbOxZsctxbNUZsxgsE+8tr0O/Cd5+r9CbQ
/kNYgI9LCYwahvwdurlj+GVcj2SFBG5cSGzgmI9n9zzHLrddD2gGcJnuzDINoGEI
AR+3ZyZlVVpiq5g7V5ola99PfuQphwkn0BwWW+dMi1a7eeYktUTXcaiMATSAnx5r
M4DGV6W62/LJIdb6jqv5kTATmxDRHtnSDDzuSl0LAoVlt2NRJbhOLookha9HWqzg
nmC9w5UTVT71/vtJMeInHkCMJomNGq8Dw1Crv1sbfe0xLSk1J/gEGarZiYLuHwKL
Wyr5TIaqfrAaUcsGI9Kaf8n3wKezV0kYAEjffzuPZC3RuSRvBq2Xvsta5t7woe8v
u3+f2Tfm/cYKMXzE1QJXZEgog6EYKpJnffAyNe+foZzUdIc03Fn8oPiowv5zArX9
QSibc8yMqrj0gBL5GrEmdd8EnuJyjnTcvrO0vgFBhFgv9JqJMQDjDeygoOi3o+Ei
CFtaDpS046lUSXFhE6f/8OrZLYmn+GV/RLB4yFbFT1GoETTdQExaI5WNU1YZjtvP
bXSUJLp3Sf5l1xiiFTajPhEuSOv3sPk2R2cqIDGHC1nyV2Ugaq1MPczmuCUNto6B
KNQj7zU0BNy8NUeB05IUUnT1be7iVIcxauYBZztiuY7QcrGQX/4t8A1katedDJKM
STReooVVzV/9MyuuzthFP1yJ0Hd0UiOpvy/aWzb9zG5sawUVjdFX6wvvjjPaFyiG
yHgOVm6WZaM8WeuudK8VXV449jPIIFw/ni7a8aP9im8JA8twXwhR7brUmqdlGSNm
aNoe1PQUunU0EBCsk9G9r1Nj3CaAIXMjIvTjiVuXCtyVlSe18AsiK3svd10fB6yi
D3x76peCwcJt0doFqQb/9fu6u58XRL/Tk2eQCnnGA3+6yTIqF+GWZDVIdvYu/TKw
4Qqjv8NyQEnYyjmZ/CZt8tKgwLBhW9/UowZXgCB0gUpi1Wl8bToAxOE/vsGmmED3
ZAvxSdDYShfNE6siHjWAgrFL7Z2XKJ0e1S6xB/ktEUx7TH+eXFj/Af6rgKBP+mlh
jfbyx3r6fXrKQxzQCnmx8nNOrNZ12i2BKAC27RQqDaslPJ0NKXgjH1mYQG6c3dVU
OaO955TdB0zHkX28/GuLrcBf961xzuk6lD1qe/gnpJE9Om91RfB4Kal+0zz1igYY
ONq5kfcrkh1fM6dvTcNAax2Q30BEvZljLVArD2jaBtSBkD/WYDMks1kDmzavcIr5
UUC6E2b5Ruc5gCfiwvyMdDxHFFMO5awt3W8lC/p0b+dtCPt3kXM+n71Tgfcqc2HJ
SA14tWTSLb9cTHTXpSCYZnryVgC1uGUrnk1eRJAgg3ojQhgA+E9gMPsLl+imhJoe
hjbxzlk5HwA5r9SrUUvrAazJlozEF5gidaj8JVQHJQ2g2x1YQtZo55Ez4z/LGAGk
zZYNGAkZa+7+4tF9hHjA+54K8bvkbm9BO6Eo0vLt+FTYHE8TxISjF1q5ZdPhnli4
09+64bATTIhP1mw7Wf3QWbOpQ/MTrMoHrn/IyXCnFf1yPvXPa3j9jpc8E8SCuANM
CosQ2ly2fHix/io7fIxoon1GRru9mpR8xQRLqvNW0ZSrsx1CJ5JpuVGgKBI34agH
TYESCIaIYitLJzdvM0Otg0729GVGY1C4f8EnDmoXQjw2BckjNHX64MqDTepTIMmA
Mm91evTtejbG8Ud5YWCCvhWmFnd+VegLvjfPYXZEfjEtut/IA6L3FLDXbZwJ+Xdh
f4UewwEvFCjF9fl2446ZQhmx0OgDOdDRZxLx1S9/fkKmk2oD3CBN1Et7MAz6/Crc
xuwIKotG1BVznOkYrV3Mp757t3Di5D4KgoC2K9hy+pBipDWTyCEXbrbb3DeFqg31
tUsFPZmJ7tehRi7K9fq+MIX8mUr+OQgEfBkDnO0p0avLy6NSWphUYU3kKizrCg2k
K5NkHxZpXIWogAahb4IO5g6mfiOfTG1FLFJzZCIKkGibAEc30EMs2H3Bw1mWM15u
FpAoRzdWRkiN5yTB0JNtFZ41Bc1EWBOEsyCEpDwpRHlSQDJGlOa5W7fAEhBOy5HK
S+iAqRhmaMjdB2zC8jXZ9DwMU3ETd/Fs1bjRRmBTAZ/lahQ4UC6WlPJ7qxneVAk8
QBnEhEMrX9GEqApNKgOofkJ47vB0srljekh2tv0q3J+Je5ofjLJTntzwVi/X3pp6
pUvCgovy+5W44zJxAij8MMwUYVJjhM5Zh0AnRVIyOymR8Se5kbOA53LAMoal8mdd
6BtKg5mOFGx3QTuW5nR7kh7YPIxb9QWJXEBq0yUrfvXaYUvTZ4ACYrEaJq8zBswn
+fBrlDVPnNbn8y/v9R28ZG/zZ302nR0TSakPSZcoj25e+oGd8Ioc2JtuvBCUrmAD
rosYg7pKAM7IOkN1RjTThWzC4JenNHEJdSGeYVpfpIL/1j29uIS7wl9IohOU+XZP
urNgtD2c/zvaix5Y4Z+MFhb51Mx4dQpVc6+9+i+aPYWZ7glmHRZuA3efdgIfo91k
Xo/CXp1EYjA+sXW6YyQzDFFsAJnOJUeBDNPzk3zw+6Y+Y95JP4R0DQj8yyBI4ZJG
6YcmOA8mWqGsvh1V4wIGNZ+asl/EDFU2tmxs/BPYAD8tGJhbhNfBADi0ioiCA2vQ
MrO1eimCgBkDH4nHbstsOTXFiTzGzVktbj+6IBKAzEYa3wV7/zRC4QhlRmYn2fVJ
G2gkQ2SEX8j9TkR18sRdaMuDUSan8bKLnfgEvMFu8C18RH+BckV635SJBShlvcf2
zjG7nE698HM/nh4z7+zNGrvY8bq3tPgMJkWSL7YBmINpwcef5Ach5ypRHLv7cDZJ
3wgzQB5dFeeJ+o/WhxPDAMroqV0U9GJ6stuAj8IC872+j8vlNbmBb2WIZZqoqG7y
yOz6K1WXVXi+sKfG18Uj6kLJ+jCb0zviBEYfTvyZNMYzHwaUZ/m7Ym6MMjkcJHL4
h4EYiwKSkbdo40boLIjDSk7BGC5gWCNj6hXIRjvLOjjofnY3dodhHv2SS+UMVx3l
tx7wC/3l74yCqpVALp1k+TxUH8XItWsOl2DUIdUCTBw7wXsM+KW3EkAJFzhfVlH9
eqivbwwk29lLijOQHBe5lu23mflCR3ngOK/74mu/VjIBx1Airk0edepT2f7wdNSw
LnSxexyrIYXYaAhh1j6Ns8jaF3me7ICQzRJ9tEHuEXyxCWY8rg7GW58q45IeCVNB
3ZniksUpObh+34IILhjYCEaTHLdul30LGKOi/wDQkjnRpSSNZg0j3uVixE90A4sC
gqn6ZZrlMI53QB663Dc6kznbTcGTQ0gvygifU1R+yOwkNWxfKwatPxCZY4syNjvp
DPMFkEiE8etVOe4tCX7gp3CGyTTkthEN+BH08SBnwKo57q+Z0bARiRkWKyRDIguo
Z5s7JdRapwgdMQW99Gr0niIGowowSBkoA6ojNiuLuzrkI5DAwiTcWUi/Jl3TdQZE
xVIGFe+NI29ENwfNzB38tf+OGgmUM6AOReWMQW2tnqfUOdvIm6bQbOlSWX293ONE
mErmtWH/cnvjS1XfqF/vv/yCAzwBUIGDVaSw0PQgKL8P7Ojn1xspg9pKYy45OR4r
TWk6AzF9x0GeccwiRKQ78wzlppTpLCKvjHNLXZU3SNa79IOwDVHygzwAQl7/YvOf
twjCUUaKa4qvThnaI5s1NJILoytztUWWqH8VtWaOuI8y4HB4YkJA/gx5XqIQQtKB
QmSS5gopAGBSaTS8ejdRfpPAJLV4fPmzrFuON0p1FtIXtzbNAY9IMn92R6EL7StE
ICSlUPXvQJ3IFFS53SrinaWN9TQhcDfl/SQ8BcjdxdqF1ryvGEImQ6lhUtnSDv2w
0jYjAL16U/6y18mIzRH+mOl791Uz4fgYApgq4boN4qmEPe+oVrzyWr/uXdeCbjgQ
XJZ7qBYk7s7+eutEJkSoTFKzyMSUK1U19H8uO62ZtsGcPqOL+CMcbNgQyq3/uAXe
LCEubLHTVoSElvF5QWm9d9KmcXJJM7ln+un3v8hcsUWnYJe5o2q+3zDVJ00zfuY1
b55qoK+PHFFgs4iwVvW37L9qniGuZ/jdE+3X66OIW3eT1myQtSTvV9cYDdI42uwZ
e3Jj45GUTQtENs020YwdqhJB8aQ1261FYYapIt328QirPdpEriAul36k4VjPWnqH
Lm99s6aFyLHxlLSztaNs2X3Xt42xsAzLljbXUZFZ0xPWAvWFodwF8HZVb+rMhLTY
yErVF8Bqww6q9Oqi368YehB2pXn9M/0gg+0LlR7HbQzNaFl3NlwfnL22p7LAVaVs
/bn3qVJdstq8YNvGRkcoYdCltsMy5bZjbzS7EpwOhf9Jf/wm3QycxOZLnQRMvHJW
YMyf4/vOKiYQbWlJOFIUdBnBSTLlNCnD/PQETky2mg5KfuaIRDDBeglvv4oGLa4P
MBRkfitoUPpLGpNvUVxUJSxFvog0HBUQZl6/WZxUkpksgKXqBNU6tl8//CpTF8mg
lF7K3r4chCNMVP8VRPZkREzXvFf/eGG+gDrVg+zkn4pbkMNnUHb/H49As+YRFtKN
pbP83uVXW+0QZqRiK/u97pChiPPghQ098HLVCjVbCH7wRt1vmYicg7sO980i38fK
9tX2z0CuO0YAxehY/c+E1fFR8cnqcCRVMxNrkRghTa499HbwFsTkueSPxCjo0Bbn
TiqFrTOjHM1i8Top2lBefxqMJO+3pvxaiZHQN1NfRURTr0pmZ018RRLBVQrSDGCN
kahJ8rqvY5WucRl9v3VlwdsdxHhEOTE/tPS6ZdHQqVWe+zKhVuhZCD5In+7QOHM0
wA0bx1evVqllII4zUAbIHW4E1evqDufSO9VAJrv+HljXh8gU3KNQfKuaIlkwjJzw
6ZU8cwzLXT7+r6DnJ2VxzCNLHTwK3JALJA1pTYK8ovxecUnq90IyYtLHs7PI1MMr
KMEyVvkHkPjy8yTKpl4RWLqIymx+XbM73XE5cn99VcFyumMqbUMVxpnnXuya74S0
3IPnXJEwoavVmZ4Ae7EF46xg9h3RWtfMV0baxHeO92QOxBgBfhCzGXBgQDsywbaj
5VPGBtesQi2kThOygqz9ZF1kKd67j0wHpW973XAoM8iZH2S/7EY7FFoUzUByqNt2
GovqvqNt31UtH3yv8e06UKR3Hf55aEKaYg3RC1tmZFpHnyo2ozSmyPZjYIXDM7sE
+tSEaKoQUWpji+cp2Kkd3OB6BkE1tWKf1UQN0gsmI3Oyg7aTWJvfJUEzsmPHc7sk
Bz8OqyUEEaL2qbNeyKDGwB1Qsjm6xT2VW8e3bW5SU8Qo6OZj1upEjbbXtpA6zlOB
XF3lWrYZFYPCwiSz/2EBwxpJTlP/kda+M62rP6r3mp3pB359TYuJkiMBH3/vrVAS
BbjKvWYVy78Xmhr17R62E3Bs1aDnzXP0ONAcmXUsJI8IadB4VxxqKaToSBoUyh0V
OJkViwjWlo//jKdS7FAKVYlMRl7gpe0o+ep9ZEfnHwC1REZqWmb0bL0G6goj8IgN
hSpSGXRUeVWERZ6LlATqo0GUBEeeQhPwtut66F5nC+Q2cjCAafxQnYPrm6OS0HwZ
A8idCbBLUE9bJyjNm9x6qWvog2hfDSw3D0/+jDiMnAZmYwycUy5vtZgANkWAW2sD
h8rc4szw/742mRiFD3rgp0yOLG2Wg2GoQv6AcNE9HdWZ3SEibDV6NtBGqFTpPGFo
xa0eK4h2EUwdbGCseeSIR7MD8ksi8NM3HTymSFQK29Wzb8MJUISAmVfWdT8ke2Wz
HOVpJ050QR3cBgOiK5FBRkRJwoNX/vVD4g1yUpuMhBgxLmN1SwPgh7s2uyUhoIph
RZ4fVHdq9eKp876qDgZLDXfS1N/1NYbP8SbsCaoA5YJxMiGVpQL9PyOi8VooV3Pb
mnFTpQPmhibazhe74e30Zt/vEV8LYAyfZmKKGX0+IBdFcCYeCGhEYb5kllayTnTI
hbz3331WspRknqvYgQgX5w/01c2k/M8D4QBe82koVE14h3qHG6lpcAMch9wyseCm
9Ime9S/FmP15RmaMKtB4JTII0bihxL6/Iv2iighJHxRHcEZbMbrbbPfUB1I3FZRM
iYM34LczRdChIi0SWdvX7NtUCTsasu4R9kPRhjxAAzeGziTMajD61L5S/XzUf1Zg
1/kS/qFbWwgu2N8mL/qqJOcLiu0DZIoniu2uFwZvHTE=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MQNgnhUtXDdbrHRm5rQiG9bX5bR8+W1K/RxOLI1CiXKwM6A4BUdougqKS2UteBLo
OtqN5ZTM+yeBrTMNWPcjDUESRC/+n3RQvXeskNmuUrTlrn9PmaBoBkTqn3utqV5Z
w5WKUI8dDa0yD3X0v1fdawHSaL32ymf87lN6dZob+K4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21680)
GVQE+UKRl/RNAcVQ93k+3SLfX0HgJeXIz7DR9qJBd/ZrynFonQ6hTeBr/0J2vVB6
c68Dlq0F9RGhn2A355/03DoGLOupm6o6eL2STZKt3leZjyplcYibIgVctKqEqL8s
LOMCL/dRUU47n4VX8h4smNBOh61+XVWIlFY8KgcnqGwvXW13iqjcdpKEaA7NTTbC
HAOKHyQ/RCbniNEck3wiY6qCcdK+A5DwsQqfr9KQMg/a5izBxws8qkcUKkKBeMLG
g8e6OV7Xe17GoUqufZccI4DcdQtLBYcQp6f2U2cGTTuuvxrmiDzHOTKdJp5xYC4r
wxY7qPPnKwGZg4g+/tXIQyglh1h0hUsCy7aMTdzfdAwXGCsqHci5ZX8cmZZONBSx
ehy4tE8v0OriGXeUZv3HcunEWJs2rsrP2HY9CKB0obiDLSDp1pGjEtq0aRXSxtbP
U5jDRT/d1e52dujyMggtuwB7tbDJ88n6+rm6Q/ZLQ2EWN4OnnJgENWeRknRpzsrJ
IO5lzpeoagTsE6274NLrk1DWIjV7IJHUyXjKHr2S2SIQutIs9ZOFd7GT9/VxttGC
ilbGobGzVqSJ4MyIwzLk6pkRcDHj6M2NAWZYb+4xSd750Ug+vD0HVnHCbmiMksvE
yOPDf/uNCattkwp8xHQ+55sY1+HLvABRiCjfaq2xC3tcnLUgfBEKaO9fTLjDEepm
rUtRxHCFkVH/QzraQ3NJ9IXItF9vDMeRStjr9LhqTylFbRq3tE42PJUO4zsNVLYn
kQHnM86CJ9O+dIygqB4K68WStjREB3PjmR5tzRPefS527VjUTFl1kAU0XTLc+hq0
AagNpsVCaxFWuQuw4s44SncZqX+lfTgZWDHphQxB/00SKrUGKE2lxCBUpAEfwh9/
frmFAqeyzcI2AR8qyk768kx64+q0JMfnh8eJ9eJez+xb7NFG893SROFE6mvkEidY
DxgDcviST77+KM/th7MOvzfYJuDw88mNCg1XLfCN5R6jR+RtyUVNS36Q7KesKqe0
BdGM5R+nrHa3w41QWvwMZT7IJhKjCHAJ/i+oPTbpiqG6LvA++zsod1i7YWmsZMmr
SZ/fxJOPqPGlcbvxqgFMRDFFECHl67NYeM4hfIzZNXnQ0S4MBB5y1avtdiVQGok4
rj9YMagGGoeFhasGZDAjngj5OM2Co4h+QqeSSSBsJk0xXC6GCLH8GrMjwKS4JBn6
7rj/Fw2vE5M4yAqKBIC7N4ekKrV++qKm2qmVwASDM++UVKCRK6kWchL1w69tldCB
7WDyhOelh/JgP0GQnlFuiDoGG+Y9hfou8G0IofAnG/dpK6esNzoNplkIrTOrRJzg
4fCQMsskXZV+oCUhuqmyXibIyn6rEaq40D9c9g111+GZ1DwDtHysccs0usfy3o7B
MY7GBSnOTtfVxQOxNjE0CzEcQjDhltsYnWPcaoYMjl7qHAR4BQmf7vH4NMvBJpn3
fkdTeQDhnG2mfDtOLNmhfOLaYVdHxA1IMNSjlPobTWoxPocur66eCE3Egtx+3X2N
EeunxS80p2ZldxTQ3DUHNjaqi86GMh5FOpEDXt5IwDXmGPsVFOT+wAgtnwVuIPtY
9CT0tDIIJ7T6ivQZHX8w8Dc4YHAZCYcVnqjUlIhFIP0gRWFK2hGcZGXbEKZuSuo9
APwRG9p0sVRGKMVQR4AH5l424/hynAt9K4e6zzK+KAvmuB5y4WAx7ITJ2tdzNWWI
6MgDmGPMpUcGMp1GUNv3o8rfK7O57/SpTKPCxHfcT1Oe2bdeMgCi0YbOk6+GXFyy
cerqF82gevUUS4crKnpKt+ksY7X15Jx3tLycVyTH6eLPBQcmTyDVjxoo/4ZQtZhe
ee+KXojhMBDthIcZWGqoTepLnDZy1K2lFOy2I7kaSKUBtxoa4bwnSGPajWRSKBr1
NNH2HIVwshPB67Wh23WsexifmgmBn5RgvOSKAqj0mzYJvnkXdjFNkYjJffMY5W1k
/fHazONAOhjdkGSDkObeDrgLjyAKP7uwQ/3fHDZBarYy8GkyWq/MbRD9PIM6Hg+x
iIGTEvYumVmAgUbSWp2sezYnktS9RjqOEsztE0Ea19CqCf/1KV9FtMAeoiMKLkaG
RjZzeCGxDVFOanAKVOcA+vfX50yag3l/MCCseuXXysg4WchPUSUBhbx4jkxmnAMT
MPU88JNDX9dpNA20XLbu7Uas88vRqcxJtXmE5qA1In+buzY/9XBJBu7e2Xw+gNOW
Wnoh9KXzGcd3/YQHXdWsxPG39r9FWrmqOoxGpr9aJ2zVDOwNSfv1/c93oHudsIBj
l+GORyp5VJoTwHrGRV+EzEk2xfXizPc3/T8A9dfGPKEy0EXU0Zr8WEsAQJ0ixcUl
Uu7TT4Dr2cHlKqsCHjf7uWNpEJepMGQSAOHoK+sVxz7kt/u/xz5xp0DKsKU2vQ4o
HksmrADOoU6ZF4NbgSdZhnzyVTX7z/jflDoOZxA1eDA2o4VW9lOBjdb1emD6qSvY
p78iMKgJtOT34QTFt9h8J6Mc3544iMmvxxeWI9/tf+ca82QM7otazGIDjRBkKXae
06CCPpezqzrVAiVPMbmIpqmvV0dfXpoi5XbHokR7VNtihVh1lb51vESawrRSrIjJ
s3DpVCZD+0wKe4yVuKt4n9O0swAk65Ew6ZxcGQu5eE1plAntKZdRohRZyJNSUsTQ
wOj1muUfOn1f77Mpf0kByzbBBsC7flJRDfQILNCA0oI8E7elx1szKIzY4UG/ZqIw
W0keZ5juRJiS09QpYeZ0WOvyoF14mmMzFQHMn238mf9/eAvUGFNElfkrVhmDawXo
2KNPkKi1dzO4QtEp0d6LrWzNASCalq4vf2phZh0EqOKXG7Im6PIpguXuCCXS/WZX
Ze5dINffyg5AUjbd3iSBT4pn817Mw92UfL3lXs8zTJHXF6xw6NXplEeVNC7H+3Zq
AL5UA00so0CYGJkRWlUH0EjLFUrxCZT/oo+f1AiboHP3eblW35La9/NAhuaFB2c+
1AUikbI1A3e0IMJmEhYItHJEn8bZ6vBoN6PKVaskf78g68sPqohFxQvMl1B3Y4g9
5ww2hirPb63Lvbcl3qVF70QMha8kyjiUOEvrX9q3QjbVT72jFJiMun4UqVTkyL2c
BYMML6GVTM8N/g9BzgGLbpgxKwNNsV5rXq49XicbHHo/9isFoVuh2XIvAcxGM39Y
lphHbFiI1lCw5y1c+qsFQbCOHssDSxnwQ5C4Y2iRoRcPPSEOdS8LA/4HQ0DqCUk/
5bA6NIy3IqVV07oxvTj0t7eJLHcNKUSgzu8fyavunlPaq1utUA3sertAMbZUC0cj
deewZgi2XdbeFbQCw53EPIlVCv5mDLXBlDnj7UMVYUSL/ylK0KhvvzQwU3+3cDxQ
m6HFVuvYdUxp89NB0PBp7eXi4Wl98NNb0y9h4m0Yr+MR4dgEeh/ob9GN1Bu/JXcT
qp9h/m9UyLA3qGOjyHhWVbMhY9GDSB0q2DzunXbKHnqJZ4breLD3Lm7Y3I1gCs7B
1Sl1AQqKsij5FKO17BdQxJXPlDAEBambWJarr2kAlRhrliU7mjXfafHNoJ8fVxok
cAKquFjJdgOAxSvpXMzHpG/yrpncTLXk5UNsVkbaB83KQgrWgru2q/Z4R3D6jEAJ
da0hrA3m2RRIykr3T8+SXnA2nUVMfVLYY4NhCoaPR3JXnQxd8BKvEbrvey0Jg3G0
/StQgIVZuddW50ifwWYkgPIJjWBwioMYW2niDUkeZsdM8oN+0bqMMidSmTva0f/t
e6XIQw4QD2bVPOElx8ZJ4f1TqPhb2bPbq3xesckN7zrgof+VxAUun8I+KKFTwVbl
v0F8f0gJcL1ip1sxT5hNE9NzTw09FgxupyDWZ56dDMSEkiLEX2xatW1AMe2nzxqW
hFH9lG0ZylDst/zOiAHehVcPaLhd/OxGMCXJGFEPJKj/mTbNrklzDNHAotHNEXcO
n8RT3hbyqyNK+yUiksUEyJtSYQmTs3Pqk0AR/ZYiOn5BCXXZqOBbJopSnGlAFNyf
fjZKfO2WROU6AYZ/OL9BVdJoSgvCO1U5Sgb0MwDNue4OAG44MfhboW7rLBLnlNHe
5vFvjW0UcP3x2Bj1pOeNlz1I6pAAtTRYAmfM5QE4RuPisnY+Gjpz7tfx8nUVJ3Db
xfEUttGZgCfPlin6Rc5c0hWIDn1e9CDMQMQsvZlMRZ4gzzkOGY+eusgsShK+isOj
YY0Q6TG4adppEBTU4bYHVYRIrjaia5ZzTxJa+A13kaLMfefwMyg963qDsDJ43OBC
4e/JEbMJmJxKHP9gNmgaY+6HVl2flR9k4r/dp3io8x5G4x4R5Krv6VITy3dTMj6L
1ad5+bAqSqKBeSBhXuCnYFehLF4RXt5oasiBG09mVgMD8Vej/rM7xWIFBzAy8+df
flNdpyagkO+GRoKWAOx3RwhKXjIGr8A15AdFlvKvAHsouyqAtwE87bVXvAL2nMgI
PZl+3O+9OwtKVbr48lPCnvlm8R6eJUt/i56ibW1hQdLM4yG0ftkkN4zaN2XEtsGg
tYQAoUb4EOt3VkplbcBEwiAMRDzFfCEj31lfWnDo0TIYhb46CcKQnVDNhKeODt+x
Z6Mj2XXHXYKAT3sELl5qs9OWm2yrQOcy7isfTMFQdPpLR7qmELnsHsUBExm3z5Rf
o99h8ZKvzLASiJ8wgkxB7fnhtJsVbobTBhH3FUDlu/qyl9q8qehzjE53wsefhWtm
BiLdfNCwCLzD1lU/dvDBrc6plbrVUFNYrb6O2RTvyfFgqB86/GGbH03MQbHzVIID
be4MH60iY7yO+5fB9KZ2zsmtnMpkwkceim4Dv3j3tQeVXZSvr1aYIh0yQzKklnLR
yrwHOhPCQpP03DQuIKvjKbnXCAJi5+VvVYcduxlkuWCzpcq57rzryhPyPiVmnFCE
soAbtBs9Lj2vKOrza99G68hu8ZJxonB65X1hfuucW85M6C6ySO1WQa+OqAcBmjL5
sILayy2dioyQW0xi3tQYaJ/dcmUHPbUflG5Suf34L2+mXXQbKgaaCrtUm2+nszq6
8l4ybBwijy+dRXN5Eg9EGy6E27UrfomcAYl1mJnvKfX6gJqM2pkJjsZxjGNsewVL
Az49vw/0Jn/NQbud88dw0Iks/nf+9h+6Ei/Pik9NKn3xuA+uU3qORUWzQOkKS3Yv
ovYsuLlzkeAz9AgV6wF0mhY7yYshN4Rob530ytl/eKFoNLEuTiCqjazs1mMeE9Kj
c9n6Zo6rI39N8EHj7+lLYiKZBEF4Bcu9hgE2sHHrvLT6eD2zlHp87Q6eZnwuzsAJ
+glc3kZuufbO3UR8sEYjkzWKjNXCROWokuFk7KP9e12R8MNN25sDjadlxN1cuNMc
AZWlpX4FMvGkt0DkLMgw1YAOJT6ooeuxD42tVA65WpAZDfV8oeAUbiqn/owBDJtR
Lz+ffcEaCr0AtSb8tc2DHiolcG79rBzeaOHI0VLfBS5/bQRDQKfgCOVUKt0fC14V
mJI6OxPgGSkhzEv6AgnHt0zYANS+jVC/3OTE4hD9NL0qP/0RDiM8cXQpAuTX29tV
8UITF2mzY248wzHt9aUgnP8Q6zDf9tdWz1Y8O5nxs1cD/ZDu35LrBMGRDyFexV0h
bVs8iuFt90cZEeYjkQMZnV3U/nOlw1EdyqE4VtHjlQ+Vx6f/yVrLTHfblqB9+6bK
Po6QkqWhYNbaziynO1s4ydzh3OMi7gNuBNdnFnYpBnn2XDR4JPcTBdVaQjLn1Ldm
oToAmuSWmz1aTBw80ha1y2YgJPUeJWLTbJBRhG7yv51RpM1hgzKs8gTPaFRBi4JX
s/Vjuiupkzc54P7hdQZY708foqX2NY4w6tPzV99hBe27XLDaAhgAh/eHw8x8us4g
t8JuCP4S5Yh7ia2NJ11plXuFolTZaZUaMORUywZ6s/Ja0pWtSrrbxcvgzx7ZaOgH
Nnslu5GFSW++8tNhgLWafaxISStxu41IRmjP6uWpCBmPll1h3BHLNG+MWu/M54Hq
YMQ/Pm8aCHjC62aeNXJiZTw/6A0j51lnaY0MTuIKcGJSsz14Dy24gc1m89i1E2yG
146779TCLlXfzbSICFkQujXGdV0Qn/2SkRYkzhqc4m7wQ5GmJf2V0CAVqCN5ROQ8
IowVtIBo1G6yjuvQWH1UWrAQaGpELkZ7JhDrit5JyAR91adiJajXb96YLuU1PzLd
wHULbK5ytr4RqSr6tv9uE8bvgz/0Z+Ix8rG7Y6wbOLezgxDsXHoN53JINboQ+fE+
goBbqA5L/rm0+MwUZ5vPsrL8a9iGJZgj4GFPKHc3nZ3JkV9g02QkhbWxqOvAvI31
t430pH33+IVSAohmoBjPCrUJEVlncNwvrdulthCq2kusn2bnVEuA2FJwFVLmfmJb
IuXp379NPt67nk/i0aSj7a2qOA0iLSVo0HcprF0GmqZeNWBZ22HviqKKJbAqvLpv
TeaCicFUjIp7dlPer2Qe3y5TuCCXakgVDH5BfwFY245w8cysHRZdxwvlv/CD9Iy6
erbZW/Qi8rrCYbbape12Jr51DQzGAXtNqmRhcKy03iKKxDqwjPU+W9gReZn2mULT
GNfc4e8lbvSKF60HnEA37bL8zPDraV1KE35LysGM2CryRvEuEVDi0xlauL88IKBg
Ad9SFq3nujghz6zfHqDTMTuW3kx8PUl3gQMvc+nig56j/8fF8J2bnUnZrIWiSnjZ
ckkNNoHGe2Icc3uvN7LTkHTLouOT+0Qvi90L9+PYiYTA6p75PukVflNEuLC976wr
Hm1/op37cs2sKgruByQ2gkiDTUU7L++g3ZGwa6wuUZJ/X050HpoD72iOhXWgSO55
LhqJ4KknauCKzYc1ay/FMTs9l5LNfWczmQ9+1Kl+CoDy3F8L52eNXHuO1jkEdw4X
QgKBYCxGTkok0/mC4UvPVDJuyC7K3HViVXWZ2mYTYlfXMSJREbZmlw1OTjmuDDwK
41J9Z04YoYl5sdGUK0Wmn/xm9corJoQ4CIjffNx60qwI8tCWrrRP8Hq7+3MpVnLc
Tn1+qh829mIpHhHnSsV9Aeig4Et/nyopnrtdbfExMra2QtjHKHkF9fMAtD3l1bMV
yNe5gOEm2858ZIKehpuICoa1OeaAXkFByMyQ883ujFCNJkBbXw6aXXf4BNxfktB5
N0ukf7Wd4pm/VjvQ+vIrxec20LN+kVkHmQn1ydmaBNmzkUUzbObOauay/hdUhhtc
mlTbAyTr0dWTi3p0a4uUSvrlFW3/2Ef05jplK2pxwFD8+PfxBNCv4KBuk/PT/GYa
fgOVRQ6aVbl6IhMN4epWbqNWFnkVIT2CuVyHptL21tYTuCSPqQSJ08z1JVxLOEyI
CCoWimeV+rfmYytcUjQhAb3AM6ruPeF8UP0bHybzD/8gfceMjkOPyZsAzkV4B/Zp
OvKgTl3cb2OMykLZ0eFfD2TKIsD4P3fZ2oGJXPt3YmDN/X/gGC+LF5vN0eWzdHWL
7rXGyRZrRiEZgx/k410mn1vzAF8D3kTU1G10o83AmsgHG32A1ynvWrOV8UEEm/59
mcBpRQBOsXHEefRZYDiRLxFLqeBn6uT/gHMHPLXjiMx98b0zm+R05IcrnrEJUElR
M9MhYlUrtbQq4JXxh39TW/AvHcbmRyEMbYaPo53B2TqDzKCSQtbNhj/vGuTqWWOv
NbZ21Bvdmmg8vY9gk1nlIVObpY9GSxFk3Fw4y0YdimrJss61mGZZgyVtsncuGKu7
CZrO8Kd0ypZT0N3cY7ybeRzzeF00NClZsHt0vg3VRKNItpakbhb3yTvRjGqKPaue
3g/KC6SxMFMqEp3mMOO6oOxZu91IXCPwaJtS2CRNOEfVKpxWm8LhuO9qlaWMtuwE
55cZ+tsL5LLJgA0Iawj53Zj1mTnuBWhS/iBEq/m9LIr7VxEgLL5sAzzREIhOEKtY
YHcgDCCK/IacI/muU8yLNoWBMMi/bwNXQqZAJ+oizriQ6Du8gJkSqA3Tmnk6mSgl
ZzohmlXIxQQX4oVndDxsQb/7v1aG3S9e2vonYgEzhVP8C2t0r6DBLk0X1/7OYRIR
JGBERwvjY2/OCjpaJZY3Cy4Bn0vlq9vXuxsF3JeH16DYCQBE+rE/yIjhf6I6hmhS
TcdyzDW+QuI4BSwQU3ZWJK386jkDdcYzQ7uYobgOTYqJ/SSJUlG6l3fZguksOPUg
fn4aKAxljVjfkLqeGUXo3txNPohv6ghp6VAb++3lIHDdC4+JuYw53GO3h+RkyOsF
lY+oNew3x8jFRfGnMZXPn51PnV9Y0aQB/FGl3OJVVfMsJLKXws2Yt5CMYXbFpUId
auhTWxE0HAyugfiEU8veptM7+yk7c9jaE6b2FC0wHxgbTWi++NPeImBu+qtp9Hll
7qEAhTrJ72kslV4U1+iS9zwapDR3yMGiol0/P4f5wbFheCz5eAlf2HEOLysrUI2m
83od7gbVBQvjaQdICeUM5gNwR1uVK+WIyfXEp79+obpnPiOTkdkv/DoIsbpDjUMn
vadlOeZsCgYEG5sAtGuL91yVotYS92s2LM3AV1NftcU1D/K1plSw5Tufn2kepSNt
H6eCouSwCaATbv4bol/mitEeQNDrXzJJK8edKAe7SMbzHXz0IZEYSmVHON34SLQr
b+PUP7thNgFpn6E7JjoaATrO/p1A55oD18RiecPX+gRJVGZDU3ipYkyq3WEHzf50
CwECJ2Z32htzyUmndoo6wLBftSCAsN+laTyCDb36BOPgtDW14mxf1EvZva4ne+72
XT2OFDJzoPVWj5jXQGO4utWXtfiVs05mFmxcC+ycKL0+tMDxUaWmGEMHaoiMrTcs
G6GJDlK0OmlgtND3zGwIaSe7yrBPVcNYauwSodP0WX2saHzStKEUMlChCbSu+Ues
sPr96iP2mUxsVMuNeU7nzaAVQhOYZExFUEvq5RogWb1mJjb+3WM/sUiDs4vMD8RJ
KBYLaH6gIdRyhR3A7NfsV24LUroJdtgb/+A2tDB18C9hR5SmJXF8P/YNQgbUKEIW
3WdIhUXOj1BDd59K0FL92KgidO1ZRwKgyyErJ5GctwaG3hmeBAZRTIX6/W//hdME
hR/DaoP2o9BFf9gXNbh4Jcs3tfXbq/gnwsiGj01aLXohkaZtkp3jG+VbT/nBk/dq
KrgMs9+l1zdIAGnGH2D+RmZN9tYB37omm+/OP3Dl8aekiTsO+M0viMQ935S/usu9
0J91d5b8GYT/yxIE7MruYPDDWghfecGXsgcXP4mL0n3l82PJK67DZbqTQxWLJec0
sRr+08dEQ44ED+Qk6FdOB1gCfFTkeegqzsQFaNeGAOscsrZDLnaW77GA6CaO7M4q
E6soCFAG37tSZOwCVjOFUYZjq//fyFFiPrh1a8or3ykUjn9FJ7lCd0KUTbRXq7xQ
YG32BZYrkUX+1M6/XiHlnMsi0meLHrytfdQfbGTiZGTCXGOL/yhosZudeyFI1urW
/FDpl6NcQL/3pVpPG50CVvKF4TgfD10nYpFA0Pi/Kq9FQb/eDK6gSp7hMNPGrSpA
6/dgPk5gIi6O3iHA/xTjvsEqqJ3ATd6SD0Oq+FOocwSd31kx5gQ3ZHvZWGRMtx2V
XXg3tfGbFoWwuJ69iuqTp0cmEsj+Vi8L6IrchNPph9XqOjI1MAq0ms/SoRsakIK7
tY4GWiA7aFnge5Ugme1kCa398U+9HoCRjboGd530sHwrXr7v55qdvhXTrBQ12pOs
qlBULsrWJcFDYw5cV0gemW3kQH/jB1oG+JD+a/LsJZnuEm4sIvj5nJswxgad6zl/
dfiz/tNjS20qo59v0lQoMCxC4ilQRk0XH1+6UmP+2+GoIrdHy6sRNvcKL9QbKC+h
cjBG8IyTgxHtCOkMyNIVDTiOkpV3DjLZG/oC6rKLmZ5LzDPwHcwcRM3koc03Mf8V
Yy8woVPLwr0oOQv46JHIA9p0ItGljxXMoEY4WzTBoRifWPuIMiQkIRkb7EDZExnW
xbRTyYwWh0HoBYEnUXt6jyY07+gu1S9dvPVLSTPo/avmvij/o37tnrlHZBbE4Xv1
WwF9dg+O59iZQazMQDOeZPT5hx+gh2lzF0Gjre2uupx+DR/bf2C68QiuWDYsnoph
eRKbpjx1fvw5ukkGIpHOya0jTwyV6nkUG1cRyxWfhfqAjf75zq+C6ViJejKT74iE
dFWV4DQ5mKHOnSkq/pzqVzsFD2aa7RVru+vXyHMJv7T76/sNayq8FWHpN2p2RA6R
jN5NiUEpkpgCNOBi6dNdYLNnOm9vRfMi05k66h/zKxKrmk1xb2yOKZcBL9BueBYS
PAOFpgppuOXU6pVEFkUTEDARum/tBKmwkxNWustjxDxxuCUsyXa042bjhAHpKTZS
Hwjw7yjmKYN/DcurEL9QlifeW8lAsezWw2d+AVGJf56SoRk8CGrazgTYTrlrZIwE
12PDxU5qMgmqNHjbP0JlaYfeP3Lv6SrnR0AWYZMFjqfSnftHqbXbRjh5T29vD/ii
EZUW7kkHXoiTbAJAIIOZgaPvKM75XQSq0IY/fsPnDooQ46G+Dv5SECba1VodonKp
7JQCiit8CUryNX2zDKkVCBspEna/2MMIn4/i0AOYFOLAMVef+5Pl1gbUmXM+x6R8
JP5hijiH3dJV+MK9jP2Jt24Kmx99YsxgsazURAGHz6H2moq2BYKjMmbAgocOFcOt
losIq2w7hfAnkPWrnGoWNprRdLcqLeYiBWU57HZez08FVwxZb0F707fn+yvw3s3C
2IaDvwDaL1I2NgMkwUxkiCpFteGRPjjP2psXrsUVdC0WlxIhSoJFc/YWq29scJdY
IqVAJTzcsIxVMjKL0AeIVt+IXeX2AwmXdZ72KQKnff40fahu+cA8ptQuId/JuvEF
lRKTfYfce2FtbXt8JCrxSpv13rKNcmJOpLMGdnZSgzgixS7j6DCLdQFbpzhxxbe1
Hs5ElPN88aHxgBRyx9bNhX6Nzw7gI1xKfs6vlOca80xWxgxAIN+tSso763cwhqfx
3jI8mOIM4eKh91gcKYdUvxttosj0VebH/YbehnkK8Na5wtyNbEQ1XG3AT5M3EbDD
lOHDG1t4qsABtt2i3MJy6S7Vmcs3vroS9uZtf+zdyIXIuW8/W6VRCuml1BAbhrJX
8rBHxUzL4YtA8TNcHH1d2q/ifGSOZ2wuRLGOo+TvJ4XyUN63UcObZ+8OF5ugroPL
aq7FtOnsXRAIJ2U+tU3Jv3Fql+dxHnbtuUcquAKkcD9Tlb2A8d0rYl8bqEhw3le5
CpZE5UklcJhznJvn07Xd3LVzZgXxZ75k0RBZ5LIsECK8kR7obrq4IDVVv69G1Gv/
F8mIfBPiquXYiUX1L+uYUJ0DuRHKpmIDpCqE4IdLcCIgmclhYd0YBwRsBez1+fX6
wmxCMY+TFcG9VGsY2HrKdfsXmDynm7xOMjUGYh7MGLPux+goiP2ycUq6v/N+vkre
c64MY02X7mjauRgx9UnYQGkbKh0o8HTXIRH4Hie6Lgobaq/BK6SOSd2W7GW7Jye5
bqvV/7+FlrdEQPCAuN8MHUu1s9/qmjRgILffc0iWdz3+vwMrxNyWSC7EINShp9Qj
DTVE2T85D64mIKIAbScyQSdnq1Y6St+05HwlldJH0OcicxqEZSG3fbUQLDDDwWRN
1CkeB+GdQIOzSH/RY5PdKJsPdYD5BKTnhxFQzZYHTTnIA+Wp67r81b7e8J8pskPP
SCUz/WdAwwI6RMePUgPNLsWfw5TMyJe7wbHhpsJtUCVQ8mtLZsX+ssMHjFkbZ3p9
dp6ezoHF3rCQGm7KLnjKgOc2EvT+I4e7EEJN29tg256LzBBeO7wE1/BeWGcWhGyz
DRwFDhThtJNC3t7uqSlIVQFEM3oR7gGbM8LrLo60vkw+em8mUKerL+g+tt4ap5+F
5JN6AFykGKXnfqrD1fZn7SNVsOoeuywnrSV7Sm/J9VmQKTZSu+EEzjr8mOIRFjYY
3/bJmLF/hKC1pda7FcOQPindlO9/+jQD8BntEucpWOusf9ClXHiRuAe3f6TNqxCy
S0X6uRUXUl48JKWTvqCagLpt8LSQOGB8byU6NsR5OH0kf6Sushd4PYSJ0BjIYUOh
2Ajx1AJpMvL8bX7axAyhH5tUqMMxw2RpxYwjLNdf6VM6NXuLblvt82nzH31PbRP3
t+gwbJxXEpCJk17DM7LDPnNcJtArF71qSQD/rh5RiPfcN94w4ddnVuNmq9bGCnEm
rkulhO/og3/lfvttQJEURNElxQMGTOV5f21OGsnielQJiDzKfofCJAIDS5kmPi21
95NUeDuY3q0i6KCzduNMPmP6DpiZCalA5llr0ZQpFeO8A+LSh7vR9u05kAPc1nla
N5iuys7OZ9tBHMo3+NBcskkwUvdrXgRHcaED/uRH1nmebOMyoLZMG2ZbbP3Tflxd
m5+uCHTSFolan2pbPeZvsO/qdWxS3FUiN9A77X6pkUnWAv5qdLdb15CfqdYubjh5
AJCA9BwSxrFyzJvQMtS8RW3Jq2GAmz5nSYNsnFBgN+voal2Vg/cDndHjv83PbU5t
+ujmYhIEVZ4K2ZK2JECvT8lrGqtOKyijjNrmjkHREqYrxpog0ITJrKPAvwMwZOeD
MiEd3cu2J1q/lyOImmTc7k+tbJN529vCuvu7RrofsSoXPBG3E97iVn4QCr88xJDL
7P+h2WDmq8Tmv1noIWCEoTSXtnZCJgkGzGyvS0p9hL6wj0HreMpHNDh6v++NRqbH
bfc8jZLG1/W9hnsGrze6dO2i9w21Fu8GtJeITa6LZZ1KM7cIx0mcAzmkq9nVFtDA
YwxC5c6BCMITKZ2I84q8th4zp5hIyFQ5ZnEKklqkK2Rg6dTWreFXptH0lnP14TlB
DyMhR4C3mcPP63nWhCJDzIsReR6DyaFfph146b3tSnxelNL6+mYUqEUpkdkvWU+W
xoA6sPASU4YPI99IBqyT7tmcXAOeGcg+DhGkKb4HUB3qsfRscXLJyTgXOjnji+KY
7kFemhQW5ZDvOHwh/trS18RTcWu7BbCCCEMbXTTFfSU5eerNToPEIZuSZhJxajyw
P9VgOckPVZ6ooNfouNmkXwdtOe+rxry2Ff9hAFJAVnAkcK33hY2TP0LpcQjn7htf
k9KiY+fHhQOS0XHQxpdlWDqhap1J41XyfNRJLdMFuz+nVWOrm+SrgrRLb4eyanBt
+zs+W+xrYDavrgGTnRBVTE2I9okuSYA9Bhpg1Y1mp25cic5rBHmtkkV/UQoktNqd
yz13f3B+oyP9c5OYeUICmf8ObWTmmgBAh0G6OHiJ7FRgpli89QwoswmsgG38Mxns
FGvLMS9fKAzwKGxlEaFeOl6HrgLaCaXTg1IOts/aghJ1d/dLSiDs4tpof37Cgbhu
zFnwGPMS8zGK3xbyrNp92q/3NCvPXV9QI1Mxu9ppzj0bPj7uQVpCjB4ivBdobuiF
3jHpQM+7P8EppI/hpYcpyB2t5ltASUQdvAm1QGk1OZK+J1yNa7gZ57KnCkVpS+KL
IXwvTPbqENG+JUDsTQZoBpb5k3ieI4gwYzkU/eJHUVhstRBfQeYmTEgFkdzjlmHR
ECXw4d032IzBGiDGzcGkWfzx8cToAoJ02zYnFJLREUPDAuan5xlViqcnlq+lu0Ao
pECuguIGET6Rn+q07ajF5pXNXpyX1CWwRRLdWkYHRc/ZKj6RjqWT6doTRKzyO4Ki
+W2/2dNiQusjYSMoMyLlzfr6X7suGvIJDpLwNCW8WpSS9D27A4sBFJEJwT1nnogz
iH1FUQc5noe+qvwSJFZ6kOQy95/0RDVjfDWr+NsquuwZ1DF1E0j0UoVNx8cPzJ2Y
F7FH8/y7fh6eQQitcmeJc0iewhtlVFW8Gthvp/zlNOix6UVGVvVX+xhdncsJGAk1
gb97VPTGGHD7aVmaWmfvKQgvLWP4RUw8rnNueXdWYAmpFDZTaUiTVWiDltlyDJSW
IXYancQ2LGbJLwGT0qRdfZomzrbpiZz+RJrcKUOCesHKFOizkiDStNSty4HddFRk
IEP981tQAi26Bl+azrvq01Kn9/MA8ZBk1Kfint8KdJGzw1lyUS1RCAO7JWIOcqs0
Bha07BHwlbGRmP/wQRRlx/GL4qUqT+EdazifLxD6LJgRhjAJnjI+O8L46AlZTkCE
dKy+zm1t4skrlL2SHVsdG9KPwFktei+LoFbS/eEyy2C55ACcvRuC77jIQIbsk1yL
l5ac7JBfbcM3iAJHHdEeh3fKmOK1SqUfETDsEz51616zcDthlsuI1Gd5eA8jbBcZ
9bnEJlWsCUXnt1T1CBRM0lgR+skVX2LV4WujEG7Zm7IkvtVuGkOvghLYnC40lo1t
yuKuiwh1ifoxEeCvssjH1VXbooy1AjNgkkvf4rHEnCP0e2d+YE6IYyjKw14sOn/S
DtcN91cM+EaAw93Gk4BGBDFgMPFTHKB1ZHcatQoQ7F3zKN51CHgLcr2bcRFSv36w
mUoKIfQ9M7yOW7zcgg6hEO7rbkzs/BhAnFZoqt/6COZwdW0fFhyogkR91z05TlYX
yOSjONHbd6uvdJAbfoT4RbmB0obXSuNCMqCVZTkTcsPTxWiymtauqqFqJ5BRiSXQ
fnlwk7HUYlMyPmiXa/6Q/ZTnmpJhaOMiP4T1KX0mBiDIq1rMGEyK+VppgBmfR2PO
GRi1XrusdPy2x3WarWplHZoi5UgYXhg37LSj0v9JfXawH7RBE8bMncRChofTkKoQ
AikCsgs2DK6poVi9cAmLrFncyX2UPJUBaU7tW1QEas3ZcsWjqJ0tX3CZQJ4tTmuI
i1lZ8YqUf8yEwaRKj2JZKy/0DY8GNz0wJ2eIFGGZ2Q5sRhATZdSsLUoYXMsxZWFh
4iJcJLhR+mMxUl6i0Ux7l9W0b1/B6Lg5wfzbw5NzTCd999MzYVLynfYJVAlQ3yD4
7yKXPUsjc5SL8vcxrD0Sjz4fXiSnDzEmfUnKylKlyqlc8fdBxdcHQw7xiEdXkT/g
X9xb7cXzuOXj6tVydkxnPAY5FthGhigcwTANqx0otzuMuloaLqUeZ2OLoC7wQDXG
IBH61o2+0tT5kA0zSg+uGxzK0eOkvhHp+9rUgQbyqgn51YlkquqM2aN84P/OrOIv
D5YC4CPAAIz1TNxRBFdyi0OA0mfwB1vtR43XETmUxwXS/X03ogQGwjakP/K1J4BZ
yDUfuOM74GCsN3t2gouqA1z4Qi3Kt0IudN/dkvXT0caV7WueiPB6Pko7obLzbDKJ
3dnhalt06wiNi78r3pUlHvWLRImcSwjCrBTpGH6hr22sAunwpe9LQf7x+w2hBg8A
uCsYAn7BqsyEmYQvQl6aRxvkonDZ9gZtxYrgktmAJLvtjRaYYSreubuTs6Hbv6D1
STc9JiyorgcJXo0lX4LRYWGXEVP3T+Z7NG6S5RLhpRtZSQVZYpwuyVxxYcNsCEMz
e8Rw7ex/M/Dijdu4zbdoWTiXwx+TDONqPTA5ePXeFgUvvuHEVlfW7y2MLuT3Pfqd
QK4RlZJTfwiO6xun8tpOa21juUkMtb+SsgSK3JZSEsXdrkf4W2DaDPqiscEd4NJt
T0/9IgLh6AzW2jO+7R/6YXW3DMkmgKSscy4glBzJdUgJ9NwAqcOR1P/TpNrIc82s
lhwikxvAwOfCQm0UEVxIWgOf5gCJVhnRNYsUqsFDGlJbBBi/mMe/mpt37VgBPgar
Ww5UinmplORfHbLfVBbRzozwFwBtvN8oqTPnPMQwhlkZkCphMORyeyZPGkAKhlNK
rOQ5a0HJpU2YcB1iaHStHbjLVV9gY2z3MJux/iASXtRYS0M1dSw/m/Jp42hkfpEP
C3kDeI6K8j1vSRdA8s08RsYxiI47tOWaXYGSrdPhoBlfQXLSjEBlqr+4y8x6a30g
IgU/PYq3HxVADkw3EM8sqLcrEkjni2dHFkxBWJ8MOupvxZNX5ssQ7Gsr42j0Kyac
TLmBQzr/P1jmHiwoENkcmEA2aDveb0llO1XuyXWXAMvKz9WaBqO+cuxtvuxwGCFQ
rjGyF42Y/8IDqUqNSmLahRil1wRm7vRjRtBEs9uykU6eBfcZf6tOjaoXMQdzTeV6
V9MTiPJgo8qsrjBhyq/+LYKeaaTvAVfTO8XrthtsZS8WQ1wrGc0k7t8uF8GYjA9+
K4O/weYDQBeuDcrynVWX5J6M5+Kbkt9B110rEMUrwAvQ16LprINbbueMGeh7rXnO
GS4bEPzRfVLf2s6LE+H6V+cZIVVzkW9Tqmx70sXCMCugYufHJgFOsj1+cWMrXeTK
W38wCA9yDBcG1UDwHojHtlz938IHAeTH9F6obeF6OVEfStxDxc1xh0JIb1c9LXt6
jWVA/XL+xxrEea/8j6YVsL9VIIyWH/shZrQmA4klfqnJZiUOQtYH1hXsR4srytjB
NM0KuqsjZiSF3Hx/YPOwB39+4OzenkGxC0JHyf94zPerwdxy8umS9SWVmlWu4QHZ
m/EQsIGww/f6+m76XJEssywQi/eKxQfP05LEqjbTFLKq+H/QTgfRrUlyh/EtK5tZ
NFjxxfc71oTc5zxdU8U6MhcAe+N4ZkgcK+PgKM7jW7KkSqYya86lqVznJ9HvTDWl
iWYb0f+OdRbLO6CmQ8wC4cCdaczI7XzhxrNwqE7s8JF4of6ndE/X7aViLmcStKzA
n2QdUEjEcvyQu3VgR0kTFepfDxh792qYUj97VAWTZCSyBcilnogNkFTxNSxOOwoP
8v8NcsLDwoMQd+0gX9L7+sn27raxJ+SKSiWuaimSUsEPJ8WvHYK7b+Z/yZfThFsx
uNfO8jNQIZBwxmaTPyhF5/IIJ6OkomZr3DTkNFchE0+puznF2hzzVezI5HqYWVIg
Np5iMUtlLhjFAIQj5hOs7NwXANaMINPSyZKIgz1ezhKoVzoMH460H8RXA2Q+G+AK
X3KSwMeCKBGrZWWOnfXBIs3clO65Zl55OfjNYOlTpbJH9YPCt7eUUMBjYx/IRwKJ
ML6oSnBGWcSWS3e40E9z/XRx3nGogOC06bwbN7zI0vKpWAM3mKzEhXt1FYgigF0R
+X1n/yi/lAMShKedoRmCrS+3DKKJ2JDhL9fO6M+Z/rnTYo1IErvZaj2Y1vNWTVgH
BfdGjBi/qFMLAo/oAm7Ub602gmxNLa9nnRHS0yL9Lm7lV1nbjRXyMPuo0rIkRkn9
aJZ+CMDcvPuLjus0v+BVFXh5CNRgnghGttEz/JtSt1RFkDIgKUR0pSlUlN3fYLa6
7YNVxPCkCaiMwQFqV8fhH0kZOovAdqvFvYRQVVs5hSdECxyd7AtzoyHLJ9zDhsmZ
GLGsu6HtYmmt227APlugEHlsqjYonlJuQC7wd6ItNDsRZ6R8cD9M7UCSbUPTHnKY
ZOSpBhMSLvwymJIXamHcaOrasVyIeStgEbzZWSswpTIDpa0na29K/OKOCoezg4LQ
ShluYXDlivT0hM0inbtYPYHLF3B5nQPcQFaln/4t2TVVqXV5gnUt9DjPqdeAmsx+
WoBR7nE8ekZuq8gUZ9391Y9ShmMEyoqmFi5FU3RCu8/vr9TKWYdOkc9eo8x28JXT
NZjMJZ9sDr2Bd0AWwaTLExVPVLb8mt5pLKdY5u7zPDWYE7BTfxQyaGREms5o25Zu
HBD8gpyXoJPuu1BsIEhQ/1WaSB47/QUInxUg90c2SpGph3PDUGUd/fIb4dkPx/vF
GPKYZXzH7fB3OC+cPmOqpgRWg9NCc9q1K/GwMNfMy9BOYlqHCHSUolrTSJmRrClg
kZdy+s3jR0ngCsvP/MXFQda4rmGkYUo/6EEkkHjGbbZOtrewxmQdZ39sb5ZZx30n
EYkoyL4YNjSpAElHT4LDJAI2ff2uYYhv8B3je1Li3pFXINE3OOqHD1Kp4CUFrkdq
Ur7mbfcCCrwmc1MtmV0tDZG8ZWQlDhL2D4tThmPq6UPb5gFIinsyQetr7cS/kWod
NCcC+zxewD2RTfo8bf2ek00tz2jbFHP5qEEruZmr/b9RC9hfcg/16EpnOtaVxjBe
oFhwvOqkmJBkaq43OmveOc1KqujlOhkrFlHt9DqOQVEhv+ivw7B/zHrrXq9es+VD
f8b/xozlfQcFyHmdtHdieJqejRPl2lrHn77/6oO7lunnEG+zMluTRPGb6PlGsodw
98ldDN3L3p6HRyXW02r326lglrykopX7GcZtA/wmwR2whHv7ITSm2MnqHAxgT+/l
PiE6cDfMKTHvJmbEu4pjq4/SLI+KnYweHr3AkttbiCza8+AR9E0mEGxN9Eh1nS/h
WEnPwpVQVqqn4eC9tLNqm7pR9NVL1rz4H/hOR+CUORsEwfhQiUmAGY/TL+JTEQiz
ehD/X8OaGGK6rKv5B6t9q4iztAVBfvW5biss63z6IvJdEfkmAdGNl9JEL8jHUvIz
Y25neidYNmqfp9Cf//hH8bz+d/tr6zbMgAcRlG6F1EFi01TnxMCgvZ7gNEoeKfvH
jp+hPAnYx5MHW+Y8Pinf1UsyX7wSLMqUEthJqYw64D8NLJHTkHFaTSOscuRNjIoK
tJKmEeOG1RVDPehO4TXEBXRrWjCwjV1fRhtG4BxsZ+3kDTj7w8x2OPbzVnqoj5n3
9NjF1jKI2QOqA8Gc2eiY+sZtuECQqJX5qdrgfql1VhZW5uNaPBnG5W2oXMZ/hvpO
3RdpzMV9fqYqrcY1vWxfEIsB4N/Fq6A35RA805EZYG4GhESB1d/a13NTyNMEYt9K
H0zkItlEow5z2rGAVgszOVPFrHotgxsxmPWQYtQx4ioDmdLpV/UhSf0VBbG5DW0A
Kov1IDF5d92nWgGqxJMzGhfsooUuiJJAdSij1/fL4onhLq3Nk5lZ7ap9XhhYVJmK
M1lg1Tv/l5BQbwWazElCYsmOSvIZ5xUE/yz86fqZOGVPmJrEVwoMRWqkIFplIO/s
aJ3dLnMexd4vn16ejCR/DjcQmZv4cHBDcMatLO1CAWHiT+PaKZmfAqQ4NUdrrzup
yk6s5GMMFp1qdgR8kbaRuWBZHY/shLqQp6T56PpyfX/lcbVuZ+y81ruphhoGh29S
uh5LDn/ja1EtgORikTFdwtErM9HRBjfnF8QFtQ3JwZS3A5Sh4IEv9z5ohhOB+nsT
eaEiNaeiXCJooxeKnWd9Vuu9+quEbMs9NnnNOEeLAOaKtmyZmmlcpL0AvrB/taNa
0trDx6+CU21lnSmvEmi1d7PEZvWjbcoO9xlfWOyXNAAutwUN0rlajkGunMk0TjrZ
KW3b6nUNeIFJHganH8nRVcT7oPwxptWHNWZ55DbNxfhtawY0b93/8HyKuW9Zs45t
vfJANtZ/1UrKrjAj64GEpiMUTdjAR/6t0bT9TVKPq6BIt6RZ5RoKAN8PZRy3XYwd
IBvzr1Z0WzH757BfIfgxQwogc7BdAhCVcVvGI1Z5lhKGbg5/XjqWnJilT3e2Ko54
PLGFovIa9AhMNpcul7qWXme9gcLA0AjQLmT8Pn/yzvn0Ll8XlzepYR2NeSebqmdw
TA8hC9dA/+VLhK7ErCBiPn/wqdl4iUDclT/RZEAm0USmcOo9SEb9xA+DlheQLApy
6itdqq6P3+ZMRzy7+GBUMhAZDk3ZBStG8nfhgmx03F0dAfHjeedIjwclJ8QYF8XY
9sYfa1FZ2GVoy4vF7BmHcWusHaRQb7T08+VhKH9UK2H6H9G5lfUhgy6K56SweCWI
SDdhRP0AynwOGjywFCHI5IyssoO2u7y4c+naYR1gyfIqppRwWHHvGl7ZYvG0As7y
Ib3IjDf/Qg8jKsgR92cCWwiKOrwzEaZ/qI8MCLSqndYEBNdoYvW3gCx8fVFcHgjm
8iVeMHb4RZDuthktDGoywOp1m64KQjf3r0B2tMOMXKCGFN06lqrNKIjbkCzpkZte
hfPIjXY/NC8hahhvl0dGgrnvuzB+RUd8XsHdUeGWmVJiozzidrSZAlUaOa2wGNLl
GIvlk6QxDkMMJdgAddlGANg62hpUaV4d+KKvOuayDt7IC2L7xMp07ecLvmIsvOPX
sk0yrFRU6l5mWGWLyx5zj1Tw7yhyUb2bFwWkC20pmSeqp+G5VKJCEyxUsrncp/sI
UoYYKIwXYi8e2BcIwQwBoa1gTnh2ijzTNr4K7SlGoBNPusJRHeeKwbkMA4cxlvh6
44PYZptLiMYeyaXojE5ic3EwuUhvkW2YS7I7Z4jpKqC63LehFwj+GFeiWga2tHdm
IXKV8kCCkT8dasaSobZ7pafhM2GMNi+8SKdK1g1Eq4qG+B+MP0Io/tW19TrCNMVo
6qqRPhcuFuPMucG6S35q78VXw5HrdZycjuAFrRnloDoXeVBAsWijZDXXKPouCU5T
RaAT63TcRzuUfIHeDRPnsXeD7stx5tZDVyglrEFiuXQpbODzmYQCrYWMy7HBZGGZ
liot2Z5BV+xhX/bDpHyFbSDWC1IEUvQZs745ujPVvE5qZsbRyK2eWY8Y6ZPUfljZ
v2tRvrsv4UT0FZZmkzwRLcxlZr2PtfA03DkLXDp5DZBTkidzWRsVzJ1H21fa62VH
12WuLbJ8VCIuLk8ZgLQ3IIr8hlA2rKbK81Gv42SRbShcd0u2r5LK6E85ef99/rVd
WgzODpexd/qWdMKtT78Zg5nvxpqs3DNUXI9TrMizcIlBnkU6BOeSB3dgYYxh29lj
J/GyBCEmloK43UlGVjGTy6PbxRVwM9uIhd3ibugjOlttmVicGncVE7/dlgycaHKo
CRojQupCNjjkoflLErZ1YjroJr0ATJTkCfMMDNoAf3ofGcJkSgkQhInqn/ViNZh2
UR1hOjOuEIkxpVYkS41GIA67Km4vg/3/Q/wT0NN8PGIKKMdsDv+P97sqEk5n5kHd
WS81f8RJjOL+ylVtpIzQSGtHV9pzTGTKCL1tDTs07crXj/XVwmDcy12WtcSRBIRW
Dxb4GQ/WS168PJe4JulZvQs6XLSc0viN0+LEbJ/Qq3BU9C2HpcrYxhS77AwfPoDU
Leew1A79BOoKrpxH0iWhJdiLytslHxm3crmiacYlz4DmzZEO8oshWZjW5ici1oDk
Vq6uu4fsDzziiROHTN7Hwj4zTq4IgBIZwzpwFtycIOACZu+sP7T9P8tvEG9+Vc1x
6KTcv8a73jJ1FJJEUPf0UPZmWCd9Dgbg+qxUxDcWR/eM5UHWBagVSn1JsSgFH5mD
XRSI9Lm5k3cTpmKRejFrTNPf1CllOOCgInYrT4jqSsrQThEYgeHvv1dewZJOcgdz
5Q2fha2ZcRnZXp7XjysZOiv2FBIGLneecAWvfSUB4Anh6sIH3PesWuxQx318qYzS
OGVYn7WaZJmMr8V48CoEW5H8bSliOeegMQQ10MY7qOBpFuYdVT4q4HI6bJsj6PhA
9HAYJnDbHKZR9eM3uuKzfmsmIh7naml5c7yJkYHQ7xKEuz4obcnUDPz2kinna74j
P+ssr57+6bbxDUZ4Fw4L0LoYQdRkmQTy/ZdWrsInL4U0SEbl1Z6yIkDk8GsfGVZO
2tn3zHjg/WdwGRxC7TSfib24ZZFjG+CnmEhdW9ONZnNmVgcwSIsVHMHxdaq2ExN+
z2mA9mKUOdGhLhy0wiOIwjxFTBZqczluZGFTpFgdmvYSfDtCswa2pQmO5TvDjpR5
dgMhEF1TRemODKiS+SMW6FmrKJW8ZHdhNRNa9RaAA33ZQiYFGqcw3kw1LrXACcDG
VGzHKzvYRx4eRYdiuUtRTgK2T/nLnF824U5niVK+onpU3KYj3Vo9ijwD++6QVn4h
kGP+prcdLg8Lsp3TMkaG+j3LPGs7ej/ysQgjHwJ9z7hes5VrElT7tNMLB+RutTpK
4XH+dUs6WWiKDsME31nS0bXCJ69JKIjY/XF7Wect75bp11ISP+lBG9aVK/5UH0Va
a7GirVOChel5ydzo0+4/k+ifXCX3oAOIjsbG6an+5PGvanOZ4RSeIQOlInJS/UbJ
OO3o+F1jcI4aX+Q29wdIQ5QjKa0Ws8hwtwniK872H7//Jr0VaR2Y+H9sqpzxFyLH
mzL9BAnj8Y6ELqceGkVdcNsGpwXFRjCtj5M43sbtEtCRK7qmZNEV3eC3RrAXkHT0
Du0k0ATAf9NcIqf4JT0wh8Ulp+ZAiA0SakbD1YpTYL4fQUWMzetFzoTu/MZIcwvM
XyNqSh9vzllOAgXMspOt8DTZPc2epZHGSmeaLJ4creIWjwJLP2HITVqHtoQ9CWB/
kUwNgl1iM/qACeuElbCWXQlZXTDFS3CW2wAJm46m9EsW0cXmqfkj289BgfAyJSzG
YlmlyWGzr0r8VWz13hEcux4uCn1p8g90VM8njfY+/olLd9rXwAG4f02we9J+L46X
0xZSJj+tis9sy1wK3MTEs4FxPPcRh/SWR6DdfBHwpES1I9Dc93RNeqbFBf/g5JZl
T6D3SCRWtIqgx/D5QETrSdZN8xIoOTYmoI9ry7TmWgz/FeK2YPmucgrIobA5Xf/v
I5cQy5jDbF4nCwxCKBoKLYvico/Kyy/wVlCeS8g6jYa5EARWHxrok4rSjkDGXooI
KYU3/h7wInFb4eZpsVeSWvUQHTEnWaUUgXoJAWPRUqsXT3XIKr/MrlWyFPyvrg0D
RsgKAtMa/mu6K00TKchH69ODP5JYfHaXuh+p1G7gBGRboNXttZcDLAnHTkdAm24b
ZKM/47cpqdKFbb53TT2s/FmqKb0oz2eLkAZ+WAHKKQbNCDoloRVV/nVptcCsVNte
OLuj0VoYjbTzNOG4qJCy7nuY6dWuxL4ovo1t9/WB/dKNmTqxTemt8ezwel9vc22b
7/jZnu3HtS3QZ182eL8QXbWL7saxlcQ2MHZYvrp2TZKpfm0p+ibkWfddTXBJKi2T
txO91/ngVYP6vD//H9om/sWBazElW9uny2OAg5t6DyGIzs14QSFuPSv6uRdRoYpP
YKgVaUOVpm21njJImD+4kKIvb3Ue3J0HI7L0tU2yZ2PMzxc3m53b1FfxxopB7Wyf
GGm4BWbFakF74aksp5H7tzEsRlqKYm8kv5uevQSF3EP8ZBr0BQEaKDbL+bq8B5CI
SRXW6JJ2R7jvPN2fYWU1i6zD8mQoEnkde75QbnHH7DdlkWPeGyshQtjy4ml5/p3y
/ZXgkUtNQrrDK/Q4whL3+7cUDumQTDeI2DnorIbLLdgvh2qKZV3J2KHKGN/ArsDy
AJ9m+p5StRRV2PAM/3EHvQHeWnbRM9MTBQ1LRQDLZnoo0Ps3ah9dqlTP8trAezXU
ME/X9j5Z3b/PUN7nyC5qzabm/LewJbE3we7Sh6yiGwuz/7pPpC46pPUHxC61p4HC
N4pLBpoewROoJpogppiH2xRb0muzcw0Szc4arP4LHBWewKs1Xe5ME4rLf3wNpgrH
bgzeI7km0fhw0gRMxwU1pN2UgBfyfDuzmCfakN4bDvMKLuf+iEWntKMEmhIrU98u
Bi8lV4wZN8r8wlmSFAxKpn41XK9JmwbOreeypSQ2iZOVJvAQBA6C6jbXH9zzjvO2
S52DrOYKLzvgteOQo6m9BXfErIszzN6X+e5JLpEm47d852krCy9BaGar6nVsYelJ
B90P+FDR1nze7djNn6S5RJIdmzJEaVqvaU4kD9VvpHTiAGoFD0ELdXa4ZQL6ja6T
j93UcG+9v4KCrIQdQ/a5oIGjJQX/i6ib/PBv5XFiapP8Q7dRfwGQ4Lz1UdmRVwsu
bAHasP8Zn9C2NjDLh6lhohqX8h2Td8ihyl6+NXdk4om8hf69TyD1vSiHAOW51gBY
HbYD69UxCdX7XIeAuV0z3h/paVnH4HSMTYuNsb3w7fqMZdi8dfNDkGeygMczQucT
tHq5aol3vD15hc5QSNu0NKMsDPQAzOXFuLNsWh7voj/7hTgqnJ8TcLrIaBi72ZDv
DUrdIJqEiavN/tEuj3cTNK8Zr0dl2a8WZ6A/CJVP0lcKiQ0qo22egOSxtTUGmz9u
+N0QaKTnENU8D7+1o89iyuxLy4thEX3KjmRM+f7XSXb5JbANdE3Fi/g7mQcKuLgf
xCzUZ8vpNKL3b4PkCEKn1eHZgn0hFtlihnz/6rhvWc/rH/h/IE6plTIEtxg9QoHI
GdHHB7gc/zMop1XuqospkfoIVSR71eIPhrYQGOcAAP0FQ6EKi2pUjgiJ4C7YiIuF
6leaxLyTl8KZE2i1Kx53/8KkiR5JZv853qwzLD5wUtpuyfstqq39xHp5mu9VUiAw
toVBtyucpkGWb8StdmkohFlTJ8BmLXhCz9Hd6w27M0Xzv2d01V1/FsWx/NW7gL5v
anqp7Bp8hMF8WlyrJU0Xj6TtXxObrcZ8jtk0CFEBJlBcB/vIFzXvI55HrnLknO41
Yd8KKK+ZEijZMO5ed2UibrnT2dn3HpeeP9QNByH7EL0JceWsl9h4WDqg44DJs6oY
3UQ9FsZ7c5jLLYuTDnghBzH3ieQDygKMRGthFRKY+v2OfCBJBd3EXEDtfvz8M0oE
QLWqkvBpqDQvrMP7ZH5YE6pbk5KEEUcSzNMWDeNhK+AFtSbbrIVQxOL9Cpb4nDwL
edaucfhMQgRrPWKj+xV7izZBriFLTqYHiOxYZF5chkY7kGgQfoy98UXbQ0BzSZEr
vZ/eTb5Pb1T6qEL6gMd1106tEZAZ1J6KPqBaCa4hW1JMzeqEtd+is6UEWJ6oa8Hy
4RtfPyHhxkXo0/GuC4cvvWA3rpbRJubAyQt8gUPP+JRdwoBwiKtSZInOB5wVvkT8
vusCo6MpQyLUtHYAOXR6NqmrYIykG/Bowux2yvpEJksoTEhVzCvZtXvX2LK8i67/
oxWLU1gs8Zm9IdvjHmSbR/nYQw4WLhUbgwnWgbxdU9TM8/dIOhWfhOlFDbwRzwOL
W/fH8QIRHX6gInG8QsMc/IRd9FInk9Fl03vAIzhrZ71nFJ9EabF9o3ucu6yWAm++
1KPE9lc6Gs5F6xVP97v6/S/0j22/+JTudHkHBwqpSBhUpITUsKAvQkFMgOWo9wh9
vowyDha+E7QqeHiBV2jy2V7JsoTymPH1WRfa7aEOoAEvu8K1tZvUPnZm3Mwi8Vgm
HMhNMnXveZg9/vLB2VsS/vBHWaLD7DU1PRMGfITRkCKpY4T0DlF6wU3q2irizQ9d
g6qyCmpwyccmbofconrPXYg81CvhrERV8PyAaqccdUILL9oDPOsf10HTSoUxNdNC
HLV7X3VP46/J/9HubgLjrVLo2b/6kpsWokQysyvbKWOl7+DVZtXU5dfFWKocTQ3U
JjtLOJc3qFHHtQpVgZV2U9FG5kLn/Q67sOAo3Mh3o1zGlWtWVAGWjCilPSdS82jP
wCCFaxPOkz1d3aZT8ocuL4Q0A6gb2FisBdfFXnIqVAf8qwnHDlym1ZvXtvOLLGuV
HK2e9XWW/9uTmTVyKrGzIJeXFBZkiMA8jH6wTc/lFSKEbhcVSRhw7uLY4S2J7+2A
farLphdDmZgm1Dq2EckML7SeEsuJeb0GXOBvXeLcKNwGLIpabHdaavsUoKo2Zcxj
bUZ2yXrxW8HZ8pd8yFcPWRpYvKRGAtlvUwj2XoobwmhjaOLloml/KBLTOPKboxbc
4mwhP1idP3HHwPAQ12jVrKkqCXU27/Fzc7RtzioYGKVqWDTihUGiGz6lZY5DCC+W
pbdUmyBC7ZKiNrVDX1PcNSNVPNzWr2+Ygo19CISnxP2AVDh2KpFYbkqp37w039BA
XbyZiEqxxid2iFyaTkvXHoMdTbg7IlenTME8k7+1LlODda5dMJ3zMNdjdck4QuzM
tgYi3Gwu25jbJGJdkJWGFg3pJMaRGKtxTY9ZrxtfxzMnJNjbuJWgNhult06dXvzg
9ZBjFzOeLYrHCyB7vtW99g5Z5EHi0a3zOGnpECOHx3rQygl+rqb7K51jNVO7xsbe
rpz+7QKrWbUa7ME6RtOGXbhJIMUNi/tNm/bA98bjOXxYrGf6EerhsifXBgPIOOes
BMnuw2hOMUx1oFIIUF3GnILDD2Mfr9TGNLAauSMBK1n7TnUxo2Fm5og6Gy5lFU1U
hGx+AQM1Sh301pQE25x3GXr+yXKP8kPrN8L6ovTdZjIUGDAgJgWIXgjFjc2wIeB8
2WAN1kPngKN5YxRz5uugsS5jcL5C5BwbvC+wmG7wQpkigrbdWPnf0XZF1kDHOALD
Uj10ziyNW6RaN/FezPzLhB5O8fkQD8/bRmL36rQ23LompTADcGs4tebrYT24DG1V
PQJuy9xgiWg24iXCrS+6ZkcZW5JhHTPRvuUc2/DFn1b3ypeZpndLNpfOhcftyOZt
KWXnqaH+6Q4qBsJjA8pb1r/ND2dMFaXtcGKfqNJxnW68Rw9l0GBoO4zWAR3q/GOL
gdM+/g4WU8xNbz3cQL+Y6QyvqpV0OVPZnLS3V+3vrTQQNZuhSCoQZ0kPyPER5m4c
BskYtdRB3No+FYVYBlCke8Llm+sqwGUCzk92HMzat8Cc7TNXtUvSEijowiRvDYuF
A2svA3K+AhOfoLhQ9DlRRuqDjzYCNIfQ/aZ3fV1JTfFWFlkK3k0XuLveJm/KRSYa
oCMEtnWQp/mlvMQWypoLPme37tDCuDIVkoODMroSqOVmtfdZrhXYtKdMY29BvMBs
sa6T4tAgaL2jSACiQIeXLDG+qlQ9EHHTF4MxtnY17u8bUfwMmiXwKsu4revyIdIo
y6GM8YAmRdM3wIfm6KBkYjugj/yYWnXxNx9mz2sTL8jZa36dti4qedJSk26p3nrT
+RsmIo0n94h0pdjuZWmk7LMaVNj7Gd7Q2RVdQ5ksoBTG2VwN+N4CVwJlFoXGGPAm
J+knvEhYz/2tTDQL/PjLuh1nba1psSz90iIiHeR1rHJ97Ay0cGBA/qhGlGw8V1FX
KdESeDFZm59RXxPpUhERlMENQ22lyOeUfRqUFthmmPWBAuNmzKZVOQbhP0R1J7i1
T/ZoKbdT9+oBUBWl9jqgMYuAjJp63/fXqc/E3n7P7C+1f4l1lBw84l3E91pKf4sR
wmzw+f3W0ck6qu5ygURrmJWEIv3SssnH8Rps3hSX71Dy2+vP+yA3YRIqMmuq2YG0
sKxUuCxxEOm6DccW8I49BjOjeb1h248qrSjNaJED4QF1V7ZRG7XyKf6VObrsyG3w
3S/Y/qTxyWQXKqVleIETNs9Kav/U6vmcCASBHbJU9B+Vp9VM1ezIPGNBOOGfq1mG
BvV+/4t2y3pQMUptBnHP/642RRgAmVKGnLmPGPa0IGsh7HYF4oW7x8KyHFIpAwjA
UdtkvdQR48G2Ldu6n0+AZZWhuPR8d4QQhByac8vP5TPQRN4cHOxirsex6qBHey42
E/OzUmPeCxPZsPhG+lwpR5YzKPRTxVaWKL1/XUjLE4Z/YK3pnNEFDU+mV7GY8tXi
X5F7a5E68Sp1mJED+KbVQL0Dbj5R9HMfZlvCzEA9Jt/TAHswAYQl1UHQj7dm9FYe
7w11ntcEvHvtSu1qV2uPGgw+/TIH2WYYN32+3uOxzvQ17ewAw4LEzFSmJxs9Fp55
GLCLTy+wdM1EI0hxMfRnXDGGuG0bJQh3XIWXBmA5ADoL/QmThS4Jprp0L13NKRvW
uj243p9NJq5FGdWJP0aJR6P5avBzgO2vytbFzQEkkp5VIw1peg0jiVcX1F6lDsUT
UAb9OLLgTd9oHHMiYvH4jODXrMvmngR0Y6sx9pR8Fv3l6aIVy2AFaSi9e7xYmm8u
JhsVN1IWgaFMfB345GSB2nxHFdcIxPlG7Uy92MJiE1wT1saDh5ZtY+Wy41XYgYG4
BrNNmQiglE7mwcvo6PuSn3AelYymSwnBsuuwWdCQbt/8Z5SFDRbDn84fhRIJgnj3
8UwmOwipy05t+lgr/pS9rkI5eLXNI/0wo3OjbZK5OfYu3dQHU2Gdvqxk4MN6Maql
deA0mltnXFP80BDC0EeUZctdNa5sKMPW2rDl8xtUqQYUaKvU8ZjjMjfDQbClswk/
R8oQhfMrznjoZExAEehUPPfzpqZQkkhRwFHGajF5OJlgs0gZ7+qBe7fVD8ripzCE
M4GiUKoZn2qTWSBloEadnWPlLJ+leIqbRxSXQItBR50C5W56yeM5GRlrJ3p+s4hX
TjUUw9X/rvmdKfB3kFbw/uPrqdYkcKbFZqxCpYRYenPu2ZQoNtxVldQXgMQ0+Jvj
A1cMTxUnXmT6SjOK3+j/2SvUBq35RxSIr2bYUfQTr8sAlbs61TONmhn6QFJUGEbl
Ilgodyo3TWbdM+GmG14w1hVDYFD0oZmVCmEwVhVlh92FDolNvqEmFJ6C1XKIUxsp
LoJ9TDBj8qHOs19POyz08HRoxv0sVxlOvuMFUbNk2xQZBsYFHCo1BwLKxoB2tcx7
RAskBzOUvivY7HkOEaJYsbrT290wPgfloSdnUrcfjyA9TEWRWA1Wk4Vh3LLw1Ut1
vtGa7wzo4SCvBAZiMtcYE1pQoFWzzKJAnsh6uwMOUV7+U8tXZzY6GxAvY/F/2JtW
IOQyxKjldTR4h2Jx8Cr6IrSZ8JOK5YVnkf/rh04/8y2Egd3m7Op3tc1mQ1bBOf32
mL9nxPiZ17snSh1abncFQQuHKFwmO5gfmKL6lGRGP0e4grWsXv05Vx2CERn6EABo
/DImvIKd2uHpClXMYbd60HDC9vOT/+4jCF9638gYwPk/gRs+MfRCFqrOh0EIcKeU
8ERzyBbbwVHN38Pg7yOtQGeVqTA0c0ciQjdjgR/LpKd7d3jwqU8fWOajdYd2dE43
gEHRW+zWUOscVujyloEDEb5YeLE6wUyiLadIg2NaPPH/85vOMqEd5e6e4DJXePyv
Q+OMdekJ88HKmsw8JOaEvMm2EXoibdjUxRRf9XztctHYXcdhRKxEA5GhRl9pA+iW
ON57bhbrCVRf1EBTpth9k5UB05FX0D06tpxjmyWB5yRJ+dLfzupIiUeL6t3W8zrn
TRJyvw4b6UXOYnTPxvZ/1+iX2CqtSq+U5ox3ZAbwd8hhVvRy026nsXhUKUgOp3mQ
1PoreEQ0YNuc7V16dyj0asuR3mqBBUpNTbdn6aZZqG0=
`pragma protect end_protected

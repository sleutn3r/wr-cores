// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
n1sgLVcQ3oCuHKK/JTrYEkT+39fYBut55RqEBZL1f7jxTSi4YuRzMKsrUIkq0mQv
etgHq1FQCD8TtfsRnqesGEjiBcz/artk9Z7MEiALMFZUN4AeyYU9r7GwEVakXe1q
00QmW4tYJpMTdU3EbINCeZ2W1najfBG/KLUSwtsNqzI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30160)
ParAuuhUYVLigLZt+rDYSaUZgzieqTRCT3W/ImUPCnhkCD4/wb5krxLuqZZgtwI4
Zs1yFIS23CTUZptAChTwP7TqzKxdAJbyf2ppx0tLKZOWGzywSGc9FxRkg0JXMb8p
N3w7tIPW5+c++NYKNi5LcIoEFwyWGO/NCWKvx6yQq5OHOSlOI1SmU7dylsvliVDx
Mv6JONcHNEAb380V+NaNs4Kw29Outv50wq0pSrPccpEwAiUL0Qwf1hOes4cUhlsP
+VMSGIUTLhE0fm4KI2Hvdxp42M4x/wrevum7dQlOlrA43Kit543VchnxfFocWHqw
6uE92E5h/e3a0Sc/AS6wOPdIXnOnzLk155x9ghnDena2YIsqenivZHvxYQrm5y3f
69Lg+oe3t9hoXA9EZ0qCW/DWVUoEPCbTUbDk4s3I37u3nDBhiJyb5cJRX6Pj/J4i
aU6nZ/Ai4BQOv1CyZyJ45VBe6dI/0npDZFaJD11DnosOV+d9xmE5pmXJWbxSwViP
+HaQPr8z2/meWhrgzHeku9LZZXww66NK1/ANahQhQF05ljTn7Wse2i01MbTHqN4U
CqyG8LxPvFglucsH/MXwCKIu5DkCjJPLWAU9refesjdT0bU4VgHInPtb1dX65r2x
Hrce5m8/Zd/RQ/wf2kk4QgIEnCScqzpR9mok1tiYCifhtPkNHNA0p1/Z5cfTMmnR
BHVFeBdy3HaN/3vEXXCuNtAPX241U0zhdjkNWotrMd1fXu920tvetM8N/12bsQW0
KpJD2N37MvaxIqunFyusx//YeJsNrx96DLeXWyocDte7Rd68pSfBYKKGZIo7jzWI
B1+vFOYPU0mauSf6WyjRCSvjYuIzKaisZ195g1NYXu9/i7K82lJ36ZlchCfsjRUd
pZeWWQmpPEf2xOoEldRBmufO/Si+gi/nMfU3n423vtRO+1cQfe8FmkWLonxaSif4
yH8DNbLBle74zAhaAsxU8GXNn8SjzDCpSf9Ajz+0MhLBqz5so5n8A+eu7cP7td5A
pyLoLC7DJ5nk+VZfBwsy8Nf+pVgM6YfClPojqFWyPcWjf56Ewhco/KYyW4/aQyE6
+VhySOI7lkLXyPQDpkkUaWNJk89cUFMX3EbY8DSvqWzq+rznHyhfeCUxqGU8wIqo
nVqYFrBfVWO2qiJ+YhU7uajdh8IK4leBLd8TUaufj7PpD9SziEOs1zcxndJmTZVL
mpmuJHZTErFNWc+L7irl8pmD38jOKs/yjgUBdk3VygjUkvUIokB+oncXYNeSfWom
F7JohdgrV9QZDiNKtU/tpvHlPf1gEQHjdqOiyEi3cMfm3KQ9QH3Yhi5jOIT1GDyP
KnrWQmi19Y2k/xFLVsIU6rYoSCMHi9J/Clc8HIb1JcJm4wjLZvBay0BQktTdITI8
Yk5nF+ty7fMFg+6ivGXcSW8Rlu6MSL8MZMLFvsfhk7JKNRHvOzlwI60Akv3Mcbjf
EQPOp+hSKOsClZ6yjrp+oghm/KBBtg54Plg+IQ+olNa9G3SLyQuwGNhD4eYj7G/d
tZS+go6TiAk79zw0rD8mA/7zESVkaY+YLAXglRUFDEGBsSYYSGzfIZ48inyoCEzJ
1ho2a6S9AGcV6+zODKK4DRGHz2Pl2tSwEs+ogGkMe5SM2WNS8DBiqKZrveugBNvd
T/7ac9GiWKyDFNBUGgnzL/xMvnYtr7iPPQHV4d0sxCVdn163ON/ObpBus02+Jdb3
eTNAzMsgaV0cyeuobnar7u49C5YSyX7oqpFLFjD7w1Kl+uBc6VStSg8ayKN8DqUQ
GeClN1a4iXznD2CkbfVdCM3jv/8EJfu9EB8RH5qGaw80mpAi/jkLj3YI2KeWFU20
A/2INIqtTXrIpvkyg2zZsomx7SLXhPo94nI+P3bIb8TnM9CC6Jpq5W8Zm6SUwkB2
J9P4jiSW7BEhX2hAtmlBvi6E95zyxmOCK9O1GteNWASNHfamnwt4R4SezrEdpKaf
nrNBq+HDdhcYkHxAHsaKUF+MPJhDTXICw+faX5hAr5i/Yc58kP17c0ICQhsDauTy
zetAXu54MAMgOnMlrfnt5QsgLjPJOwbHQEWK9bEAY4BKtiPBmgg06yKcO48lCzNo
YPk+SRBWMrx7v8BzVjHqaK7N3Hl4p0bNWn0cjl1maw5JzEok1tbCAiTsygOMoRKh
sl8KJx3BK7tL67p42s1vcGr+3QcrUi3h+jNMiQstLsHlqEQB57kwI1aHlFjPIjdr
3QeFHL0w+2cWM8pY8uaLTHcSfWr9Dc/MBHheMx8iO5SX0dm1EN8l+n3vKKqfzA0e
sQYFeErrYuZnvDObP5erjlY23J9dolnjk0g+gq9S30zsOzbEY2FkkX+07km7x2nt
1kP8bRuOmKH7iMevNtmv7NfMbnkT0ZduLdW6CR+UOsP5ZUVeftvmzm8O/zhxq/Vv
Rr+bfNiictswrL3qU+cotSVDLDQMUo4JMV3Hjjq363aj686bOJ13/Y/2C7ILNr/3
8U4RPMpaXWVnyO19QG0q0I/deu7tUtphmHrz7pIKR5HkQQARfnQ7XCGGzRenwkvh
UGRogSHJFXVYUpYwBgN4/qzEfMyBMZ06Y9FTjHoQWKblP1YE3XjvUj8okCBZuNA+
koHiD8HO1p6gNY9XoFmq8BbkpqW61HxFmMR2gQvNy4eKbmli34Vrf2h2tyhtKSTY
fBG1bf2JLMWeB12wT8hzxP/YDCsBO1IP/21A28DFu4+siPT3RajUFvvSLjEKOq7E
V+Wcw5wrbKA25xnzPlShen0NFTPT6seFLM28X40FyKMQegbRrl73XbKWBLcyB4XJ
KeFPXxtx0qRCG0F8i69+sG95zwGxO/rqlsRGZwYT9OGmTJxkk4fYS0RLVAi2TRgi
YL/MeEdD5NU8SvTxZCxqR9aYmw9Pl9rcVbQmYxckGHf9Hio9jbFC3pBGUb537hH8
D5BZGSxziAqyhhU2EfuSOjOmKfqn+AcHa4/TanyRvuvHgojKCvQfeK0b7UNMl2jr
KPIXkkRoRvKUw+MdNO2Mu2OO/MRL3q4lkx/DLay4qkq8TN2UNoGPE/vzF973WeR+
/BeaphnnYXm5Yr4Xiubpi0+xZa1ciew9dQxJjB09TZH/7BhGH9cAfF/qZnsfaPhc
vwpACEmrj1kVmjlSEmHQtFgc2SImRgHThqFxqEBT+TeDPLPy9uTN6QEUJXoGcBlN
/CfzVilSjfUNcGyFo/EyKt8dArYkJRVuzx0pN0c7dnft2gCHtBFYoji2tIcRXw7P
DFvx8I1ctK1wMqQXQJBlOvpdcoDGH+wZmcodJAd5hVyHr4pjpl2KSXMP2Vfwjgf9
PxFnfcV6tIk9iajTuhIXopHYUEVv+udmwhBJvuMLuFD2eaLD7T+YKql4R7gNdJuu
qwCQEZthUmTTUymlQ8vTcHNKQvmghQ5/1SZMzwqOLxnqReXKmHAm5BT49GPGV/MX
H0QI9c9gXOTBx7Fh9GZve82TOUbk+zbjz8mr5x/E6BG2AeNCQ8sAD2Y/9Wtk9T8+
OQb/lsF5yPr3s2FF28uI+k/v3pcrXpXd4qM33x23ySdk2RL5N8356IicE904IkgK
fbaUPM4f8A2jEeAdWqB0UwL9c/M6hnmGeMhnsB1TjKXtff4NgW73Z8T3wxu0fUc1
zGbSp9zAc8pzKU/PJnHtcSaXu/4dJuKmmFTW/TnOk0LUTHv2/nDeGijzYtf1Mga7
EyF+EXkguSRZ12UeksckyrbLj/h332osMJQ9ShveIHx16TJSN6dZ29EkB5R/ijsp
TZa3MJzvD0+mH5/ga+I5AOZx8OSkVshr7r6Q5pIISfl7AhshrSCTBeLC9OmUybhZ
XU4SUL40nT2B5GfvBzd6l8Fa6wvfmFvyc/YiQyDBrWVdIMfpoKkM8PJRdec+YxPh
YKd/Csnwh5FPBuB64/e7Qj9GoPgL4O3SjwJ+R8+vOoEQ6VZAJOwpTdyMrR+vyBpS
q3iw/hRQRKMCl/zQAE6emWsOXiEd3yedOZfjRFzqofJU3uVnVHuGXiPgo+Y14PXv
CcSgsWQ6DpqFyB1LDWj1zH2kSzLK8ocKJqQU3omsSrxf0mz5Skaevb5CJTJ3VRk1
NNYTf38XMe4yOp8d1a/Vba/O5NouxzkPkT+iqmGtjjLP3kLry79xB9pcSP8mZeQS
yXTK9cjiPSeG8vACEsYETX/RncF1dLFN6ebCnTQXTXfiicQwuF10FQ/OBsrhXC5C
D9ObYMsvFZx+Mt0lo6UBGD9gb9AOE3wnDk/LVA9aloKHoTGGufAYRHY96XzgplRY
xrwomGI4DUiVsXyjb4uTqDnLeucFxC88Ua8io6Srnk7LE9Y+ewkh6Ixn2kBKZXDV
TfQ6uDYTluubkgk5rNPcwC/HSMtBTFstK4/obTWKZAhJQdoNw9fmJiGtxMTUjSuh
LDOhRR1u2zIiIc09F6TYORPSQPh8CjHUhIgXLfA4WvLSv4zcm0mmOMvQ+4pA1GKk
aoZ416FPJAjbSkaNCaoDVoBeXruaSTRNrlUtFTIOGGBWFUDM8ynUmaEU2Ml5rxSs
wgKA6/UhySTmRnb0QCidv+7NrKSXdeOImyylHPpcP/JcU6zqtcUA827V5PPZpT5H
7X3XPjZUzeVH06oU8/YOaCMkdj72EOpko6qoxSvubua4zwMx5gr8oe2Qz9HNsY4d
Z/e/SoJkXMHVvri9IaWVT7+Dzq83pdu0PiVE6adby00HYrj59sekhOIGRYBik7Xe
KjBLn/Cmnqzqce2lnHLVBSMUzGR6jdLXffoaik6j95rfW7tI2XgnOciiWO0j/HgQ
9YzhtTNQmtpGIMgO6gAPeS44M16ic9kOZSQm+yd+AwX0tIQBaVDi9njGHa36o93H
6SQl3rvDZ/rwDuFarnLP1BquOU3CH4qY6X5Kk52/iYo4+ljxOZVIb//jQRaBN719
mWvMa1LOcluePGaX8e7rdmjFlE4pHVUuGputoruWCjYnIW4G8dAjNvwMue3VHKib
UhnqMg2Zn5C3IkUjO1F/lkCbCsxhxFVmj5j5oGZxhgKXcILDO9zCnFJhWJaSYA+d
e6HsnLSg64ccwrlLARckWh7G62XZsqQUII7t+kzHY0Jtuacxqpj23c9mQE7HdgkR
hJ5JnI4pip3ctV3wp6pAbNt55DRr1SCRQCdTN0GeacHE/ZvIobGySWz9feXG5tfT
CWtqNTyLmbRH9QwZbBcrb2ScXYaz9Pkl1lWKRrJdvkjMJExVwcCFEbzaJmGREuKz
sSEAnqM5E7hLI6IWq3ps8YIOODKbuIunFkNYOPNQHkVapyKAQh5pdnaZAybGe5p/
bpYvVgGqETA0kSY2uCUDprPuJua9pwHMaStvIzaqCFf9CPILhRkAQMblelVJtD6e
BtvfH3CJA4mebWRHDeGybyyAHQs96umQNHY8nyBXI4xUlR+hHK2SxnxO1EffcNts
kgApEiAUePtx0hBexw+jGYEIzykBKBV/rr0Bg+MoJ4fqgJ2JMiYY8qkzB1ojYhGB
wzbO5oz/2tBYTa7o6AH6wKBA1oA2Du46+LLjDa0W4q211NT1gNsi9NoHLcF7fjFh
o3mrSdMoTewhLZV6m01nBrcdW371EHm0JnEPBmKg8QioLdFu1tw0xuS8D1poMFIH
K9msnwz2jPmRqXmaf12u1uyvqPnqvRVDsECr3KayxHgaNvYLXKR75E9bXYaaqAj5
FCQLyQ7WNDyv/ApXLjQqPsHsQ0wvvbPCm3CbIu+p7JXzIrsQlpy6baHIgAv/CLXn
3QX1YyaK0BU7M4KWZM1v/hXoCS4P/LUrG/3Xdvxn4ImoG8y1s9V50rD0AP91uCmN
7wat20qtNGr6RweZnpou+lCiFKGiaGRDafZAipn71ZX+Hd1e4rX30bHO/ZSmB60R
rMNEi8d4uy3coGOKLhUO6ujCmgh9qQvrWD38+9U4pV6hQw1ZZcOwwtOX7nit8vtu
88yTRprU1DacmMiQ+5ZUoeDFnNU9vkBbHvp/9caIuZVL3R2u02/aPqQVknPz+MYS
ozEhnG6b6jsmvAUrM07qTtMardOZc41yWkuk1ybeTt21wSo3qqcPTlSlzo5Y1Ru6
QykkAczKJ6I2HZ4ELMykWRiOpqnS/czuImTP4YLUGzkoTSxZ+kahVPU3zTAeqnRi
6CU8X2gfphFyvGobjlII2E5EYHriGRfuq+isMs0wrYA0Vlma0ZBr4qV0HTa7MmKG
JLTyP5dBqzq66y9OJl8jhb2MfEtnWkojtNxbNRqcLYR0uM5nbxdXgHszgxHHtmhX
HAOnO7cNKF4jq6IEL3S1HXkzAMFsslkMfJcROwn4oPWl55dxPzcH5SV9buuU0Q13
mPGpm2SWcCXMZiOkQ68x5W+VaRLoGL4DcIdc9r3K43AKDA8nNCzlGSZ5it2WUbHe
+6+t4YxEzspXZUHdhKHr+By1Ua08U/2gpGsVRoWXWoFDdxi4VOKH8zSkfhU8NGG+
i96HeKAHvPLa7fFh4GQimXfPNDAZNsiZmSe1s2OfLh/0Snf6/cJK5fegK7Ubeoh6
4u7ddBYtV/LmQHK+C57hosmDv0hV2MqlT1N53jUbj8ocFUO/Clv8/VuHMh56dJUE
i4B4RnRsBSAg6QC8t4wzZcazaMJy3eK5/q4wnYxVCYJkIiR+b9AEC9nrdpaZylkW
rOb+npWk9YTz0ptuYj7Su3jz0wq8faNS9/IEWVxy8wBuVDGR3kSMmBr+Z3+ihHOI
cjb25NqKzMIGR6UVEkvziyqPpwZBSXCWLYpPASkZEmABRqBG5uJGchIz6ICIOAap
k+a4tGiVmEH4sGxzLYhQMVuqiTdmc9W/xATGwK7vsTJAOCjQmyjuMrzfi36g1crt
fwnxABlBVNbDbx7dstww3xFAk6chlw/jEgVOpmknlNOfY24HH2es6jEPT/u5pBPm
LsPy2xUP+s0286hRC/MswBbUfJ8yCtlWTzemUTnFQCh2ZFF2Tf1vJ5AKGMGVJVBG
TaXBMpMsLJNDDPprTK9HT3Bl/HM9DHRAHPy0rneahL89a7NmFWCwRexUUxyaCj6t
wtQNgihU0sSV0NLbpp5/4kLSY3edQEM07R3wIfRv8T9bfZ8oREHAQIh24ivdoHVN
+oqXd9t/9UIeeeezX95/BM2vDN1bpJYxesc4x0rOJZtal4ylsdCRnDfh8Vg26Nbe
zJGGqhnqqzBhHdHQJ7grlQsRN42nY1pIzn57YXBBh2/0m5CtfiMZVg6PJw6U82Tf
SIc2Gyj4JuNPM4r+bIgBtTL3ZVMpAXgBaeCOk/PgCrIgLi+WFlvHjK90b8EcDshH
bUyDKj7EDsfRb7uvX+M7T9iudKpzgesoPEFBC4HUNyFQU0yPEWtEdJIFLQ8I2bU3
O1MLfp8M6eyRundkgItONUteKOBQgH2pEgvx4JuVhODJqvwZIgiEE3Jz5JBHq59F
3GX9DYsR4kB1SZnK/gDoI1ggNl6O7Rz4jAfQjD/G9Ml/xJQ21Fpypmvgs3biyKQy
qSibnV32vumUtPRW6WpTHEwsFc/wQg/bhbZLF7O/E1yZDxLjnGdLuRH7xtLqMCmW
5mNenojmJoFnmKHzLEQvuG6JredJT1oVvEdWEH1iHgLzf9up/OBsMQ0qrf3wlY20
sVeTapZYAwrmm5I7/Y9BWAYSv5s7chWMFFhcc/53CjmNpfxPJ7LHQynQrktzB23m
3/HqOxylkjOFo5yWT3R+b/cG0MlFKsOsVMpg0eN3EBT75ekMiKOifSa0/HhullQh
zrQPy5N5qmpRqmAQVAuL7l01Ac26rkINB67XjmH6wWOwvlVGbSsSjiZKC5+8whIx
hrmB1ee2DQJwNStqnOZTciu/0LP9DHwQ/PxvKOJk1hC77IRgUvcuKXyvJVr0sEYG
nPD6FokMCsrviTkagIcIohRslqDDKpwx+s17rw49W/2dzYjDZVafHApQDZGgsMdb
fodypuF3NrjVU4neD9U6+H11cNyQGjXKO7qNBn5HVV/SOOMWTgHau7oGTC3laHti
Lu948mIXgVX+kPWtc5DB3Ie4ZpVs/gHPkJo3xWs3Jxx6sXdlxjOj6OtYa1D0G6Gw
a27RqNXsOGJGeY42p3xakmT9lCCIRJDpiKZVIh3uNr+P8sHf7jOyRmUnVLxMzT6m
a0ASsEOBBL+jMUd3vIYLGDKk0Z+wR+zh8PpOI5w7KpZGUqYaeTpzfMRt1Cm22Pi4
0o/7klHvpi5lTlOGmZ0zIkMmOf0fDhgt9Hes8vHx9FdYrmafuqo0WC/8fJ9hfoT1
v3aKqIVNgOjucuzmLtu8QzN5lXuD+eq7Kz2FDi4wsdc3OwEI1BbaMogbfGAFD/7o
+DSViVoSvwZz6h7USDqKuyzZa/iLXX9Yky7kj6D7zQ6sFHKH1wpkleuJbbgFaWw1
biAUTFiQHKEvvbSCvWgQbOH6tCiffkp2B3EGZyjIEpaFkLc3i0Y2NYv3MnXfpvLV
Fdr1QkSNsU7JtnAF3miADH6H2Pap6YV0fgmAfFkhhUnoWht9Ud/jtHTf5aGw8YcI
lpyNhiJfTxbyCJmJ779eLv7MehEY/a5OGpYkWudF6K2HY2amq2tI6n+Oz21WsWQB
a/oOsbYYRIt6JPjv0EJMGjTEC9EFMcPUsA3mTrsNdP9xfZdfK464B5K/iwtS+rfR
0B90vOsTWkkx5z/yeWjEO1sQo1bdhbZqGfQy370hchZVPAupnwvRrUHEkE3PGdot
aKiZl2D7Z98kQrC1yBRIjHnKylxoz+s8564ags4B3/RerQtSmbfVF/sRUl9/0pFq
XENCkIIj7fbLta21ZmRnTeViemdduAxXXddhkJKD1yEqd6ZoBsuMhZ8lOxC8ZOP8
tSMlnsZPurs7DZHpPhPqGdZv14vkF7wY72jErwhsZvG4nK/Avpzn8fFRCscaPtsg
Rk4Cd9COgAZa9tiOTYvFv2c+fifLDPAruGQblCpFjC7qiflmBI1ZCrdFjB9CbfNI
T4gl7CMr/Ou/2WkgoC/oZZLb6wd8fnj84satVhQyqPusezCb9oJuF2tFwWLkxtIT
zLQ+pedhW1KgUhcFlCx+4gbYLRVuZAu0Goq11P0De/Vr7k0pouHtqhgn1c5owS2A
OEQKdUz56NKGm5SRw3S24kaIHf9PFQAHlICtU7WYOD1IWLuJeT7cWoOKEhm/Ekh5
k2wRfTx+HtF1qnGxT3v/8D/qB24mrgPBxnRoNOsn9VKUqHoYG4DAuHF9z9vy3p8j
/le5kPO97owfASqSL1KroAZUX0Zb/YSY+6kNihIuUbyyMIz9lgIrTN7XBSOYMecH
+HXKG2C1Cw6KgVjm6Icos2cEOk4DXMi5KPsfTPcXaPeyy1DSAVbcnIk0DroUQhC2
GucBhy22waqdaFom2+Jhdnhea1EhDnskV4unbbwHS3WOB/yGQRHZt5L39SE5dXIc
Iqi/pBkAFfzTJrNP7pJDl/iz3P39NJ19ehl8YYCJlTrtMe3DSfCde6/hwkDV2HET
u7esWSNS/vh5EfVWoOgPaHEZLHBBQRWS2sj1dfy7SQdp5YZKmZhM6NpFmIiUqdEa
XgHwuTAxzlDSgyRfaXdgfoYTc/0UQaICj6whOwl8Uoa34NheabBVzJfP0nl/q6Um
Z1qJwOh2/lsoLgR1WX9cKks4NKoXuIDCWNmcDQiDcFKehuo0BT/IwO739kR/y56w
zV4OxfYWyLbwyAtE8M5keu8s6KL/hoFt9D9kHsKQ0sZmJr/2Ot02lvxKkYVR7dQh
xZ66v2avgEh8/WLd4wv2sa/Y9RtD5BWB4KMOhO7oOmvnj2lhMdPzIIc0oS6eUPd7
emnD2DdAhe7geA46saX3J7wgOUxZLbYAl+MVYsJW9btrSXMGszH++0Kb+yzG2/Cp
+ntIuzqclX60F/K1xQRxOp8XzC3WPg4xp5Hpom1+bs2PeSae2PpTWIJNSNABPznm
kLWx814gzc9MIAOp2PVYNiCNLuybjYlwh21GBMWSMJIJf/nqPMyo9SW+0MJKDz3S
gu4zXwdLiXit2GuCMM3f30+FdIlPYZWMz56/lrtcA9qnozm7ZLcKJ05DqXuWa4aK
FCQXedgByW/PRUm3mJhHpUDgegWxrd4zEl1y6xKlXNsZocVusF9UStUNDcaRiSbK
9rHSqOFJkDq2DVIkcOCAgCoxfaMfB55io6r91xIwG+liaVSPZy5qW5st8UJZG9Rn
8Ed7iPUZZgzKrtrIAHKeaxIqIzcQsLmGrWfO6frF5ejm7f/vkHE6WavPGnUi6Riy
JIqM7sdTsT8lhdSUciqiwQAL1pjboQMxqXrWnyyVJfvb/iDrvJSXtqrhVjxOfNLE
AjrP6xiWSzRnqvcyCjdcANtFqwRFgZd0OZzGj2bFmbUGi+E7Fxs5tl2eKI6C86kY
erDupWPiyL/PgJTD8+hPZ0yzErrvjclK1v3FcQo4K5PegeVgXsW8mW8VCsWBJImh
l3AHoBZGTk8M4VJoc/tc6F3Z1wVf870K2NIaMHmpml/J1L+CjHI7YUUhECItx2Ob
FmMXGCVTNq/A8lJRi4UIrdDP/CSi8hcMbxR+vA62w86RVgX8QCmiP2kxqqGAp373
vU81xXjgzHBKEH58GCTfwBYC+e4QqUD0eOfU+nCncUujdS0sjVG5Hrslvt8DxH4e
SWy4j0okKckNbOxw8GsR70vLnRoDv50C9JF3YeAeRR5K2l/GE/nhQ8GJiUORtGHd
ewPNIbYrlNrx8j1lOcw509Zpja44kU1Ij3vFS2/MJRv8It68UNEQC4iVHIbzsowf
KZ9v3V+uTFg1FskIYwSEOcrSMd0LYzVRHxkKk7u1EEmi408MjMgZdf6ogQ2zROxW
rMXna6PAw7o4KmFhqf4kjLJO0EUaKV6N8kdrOO9x/yGjWkx1vDgvOSaoIU61wmZw
f8i7dbhrdFTTWfaaqnTcREXC0PwUZ6FLERn1gVBQ8aldDGI/BYp0fxz1nzfCMa/r
e/xeWpgm/yr9haoYs5w5Vp3+kH+e3iL2e5IOrVdIKpVBl95rvSs9lV27kQ2//6ZN
qKG9Pw/U/xqQ/zbhrmvxjuELIRkmgCo1dCgWGsRlI7CY3w6MWJgnmCl9hZKvx4PU
rDeW+rPcCM/+F7YrcrgyPwD1QK4f4sojyInJfV1cQIoUe14CxG8NjZYmNEp/NBco
o3Ix4VdJJHqF4bohALhypLyt5dFLgtdIl1nKNb7bT9M0truwqM/ZELC0LGeA0rHn
55tddpjrODfDUHhfAJz0PurgUbNSOU4MRoy5Gl+Bis+9MzGyAIoT/DaW0E+IG4Ku
89lDvn0aa1CAJRy80AtLehpKCzOHERC8kaHkoFIVP2p6YmGaqjLebQFOrij1qD4C
nalNO4bKu8Jvgv24FBLuG9V9UUGH47KuO8IkHQ0xD4P92J7PSUw8ZG5WKAfaUzxO
+f62YXwJFluUeGxN3hMafaS/AIW+vN24UFWxpAy42c20UQZ+SQWEzVrxYhe28Jfl
NM5m0uoNz3qS845dDeoU+lnHqZCNkTFyFEqosSAF5PFvWSmZSUjqspux/cMrXuxX
/bqXBn9+FbUD3VEyvORk9PGpJcUr526uQqiDJ3Nk1zy5NA49t4Q24iroHIFAALaE
38VotYbLY4BmfDeg6X8xpx8M66k4cjqkMg8ZHTHo4bltDwiRTG6jB4fqpB27dQBf
VL1ctlDK+damBs1UfFFDemXlTdMiw25Ux3Lwwu8OMAJKOYemlJpFGaFGHaNQozp4
oXDO5ZzcX1Auf3Ts5eOyVGHJMpLBrJV9eZ1lWZt8EDlmGvdEjykpsH/0PedOTa7I
r5Cbo9hj0aoIiHmYoQhvvnjqJyhKixXEqjVD5pvfMkAjTAgBtrKrW+7t+TBeFhEV
ngq3a26Yb6Qsj3rlTUxMLkn6McC/fXYkR+7X6iFF0y4sL6qK3xvUZjuES9D/H5X0
iWgmchkXa9/1zaX/iVocvfNwSuFdQbrLfSfSolNgcV9eFydLuTU+wbCpN2NYn63s
JzdHZljc8vHuJnul2fGEpdLXKkuRHBzH9qkBIdfkfTOOMWCdOEdAMA15XCZlMtkc
xqe+p7w01SMcBsjRY23u4dJSQ0Xa2FHKEy/ASXGy8Ghc511K0fEFwauNnt/jij8t
KeQQhTEJ0cKqeMJn6trF4KhOE7k6hFtW8d78EzVIbamBfhkEZlSyQWZ2Gjq7gFcq
QwWo1fS+UlrAhDtu0ECmAAW9vb/Q7CRz4LnHAEbhvbzajspcILwB//QGMXyLa+yf
nhPTklezeUHHZ6B5XlprjJrW7b155+C9XI6q9PwE2uBAQgc0xlCIjFD5L57thZ+K
YgY8wmt9rPzFf4beVFMcV4bV30czPTkn9Owip2p4UWRbqfxJaDzcXjYXjkWOvxhM
ZT9ELuyp0oK2IOITZkAmSYryr3BOijph/rgZs2POxk612Aq7JcGEz2FzovKm6lB4
cTqcBzrGDl5Cj+Qe0fzD1vz+OBMY3Bp5Yv5+rp2/pxDB/ScB5rTQ4cqY4qw58uEe
tdNbwRygGKU74hte1RSKjvbcxAnGVzxO/7wDJxOArguJrEHO8o09Yxrfo6Junca5
lgRYhqtldnVVnEVQJTa6+YJzOvkykQAyAxFMZyIB0mx1aEIj7qMahEVJuq4RnfPo
ii3YFSNnoLTcr4i66zS+fngDU5cQJds4LQXct+dpdq2i0qLoZUvhPWUfa87lwc7J
NxmH7rzN6qofHirVM6AQqUsgF5foxOd6bJOi5BMkTbrKGBURFp4dtc0Mm0AOTK4+
QFH8sAJ00UfGAaiJlVuKza8F/3RSaq3006xOwVpy6cYdwFUoOFlDT+ZIEXp1DrsJ
tlMNe616xvXQnw9b7Xo5QpuoXyA7554qz4jsbW55ftfMb8Zy8nHWc8wfRj/oxZQW
oUsWFYQxKFOaCqDuij1Dycukcr5qVLXP+1kgW7USNv/klYupiYG8EBaGmzb7rU8t
tUN6qbV0n+FqXmLhjXFlxpBqtanvxFI/jyoNBscdnJy3biUrTzqaG7tki9WWi5Fu
FmoulLUYhr9fgXmfdr2BFI4aPhub89EyNiRcXKtJVPiS0JwrHRIaafzNw4l3v/XI
15Qvljp8UCVk8TPwXQbCn/7TFxNOv6JQ2scGUgonsXp+O0t3puqz5h8I9KiXGpgm
XzP4aeZZ5B/ELFmvgKs/GOaRY3f54Ehwl5KlqbiJkpqKKw+98YJWQHfg4lUYhUd4
hWEDlyACHDwEvftMqzfhIRSgLwbUpnm3C/wOEcesACn9Lk6x4xATTp2tYmy5MKno
4/nbV95Pfjpt6bU286bJM0b+imW+K0iWTeptXDKWkcxLSuqZ8fghaZv99/MQ+7e0
wF5n1+zdzQAqXm3xJce4hIXnmAsZrj2ogdtkXWTEm5FqhGj3uzxRuU4BYQpGXf9i
v/UJJHds2lt9ORKntNS8+GZpM2OBIOqzB+0KbGl9Zcyld4mjUYP2i7V0EMu6A63K
Rz6NuPawsR+yXn65ZXYzuj37KwK8TzgMGrUv2Le60vGlqMaN87ZlzfHNoe6FYhnV
mG9o7fbh8bvQLMxoFxD+IXJTgApJHnwA7c9vq8oesGnLETvaVM3igXmpoXUYeAb/
idBUwhqYX/9uTfS0HUVIxLw7wfxKrmax6xNOmO/2YQ+mszKjwsGz97s8TVk1UN5J
m5C+dMihcuTufdZ3RntSYCYOEfafhh53WddvDNj8BjD+Pa3n0qJuLRfnmezukYsX
5w94+EKuGtimujG0CkBZWcaToyHeioQ+S8hqtKQx5BkH8/Ikc2DokhFvZ9frDGva
BzWYdosGx6KbxFbxyxKI526Uda/GU9xx+SxlYiYpPTR3K7GIOTwBLqkaqb8MbQBA
Yu8M0K4YLVkuaioVxDacDOM37rgQjaztNv90M8KlRrEVZEg33nFrGQeduGPRPmSx
vKnJ5he4af6q5sF7rg223bLxfYWGuYYXwBEX1CT7tEke/vDnj7k82/cKcCGDUh7G
sQtNnxxN4DLZcm90knw8iqm3vOHUbZbksVXQdi8mXrlY9uopuyAuxTGUQ7wKuaYi
Drm1lOOGyvgqNzmBHmbmK892EY5faFmR0I7W5UrdUJxKUeXTXMBiwyyUC0CQYmjA
b7YYYg3PwsT6hnYM2vilZfHbXKJii8CSQc/NiF8Ld2KH0GDwjNSGOeol0m80Gwz5
8SIWupaZxmrr0q/GffElVyih3Hv6QmybfQqNUu/1Q04eBlnPIDx/uQbRtKU4rBZo
jR/x/CDgXgMzqV0M6VinKXXRwUop+bhKzUp/66JbuSZ1Sf9SgqxqXKfyxXGw9x7a
jlTapMlgVawvYEE6yBPFl7JMAD0iJ7aaqA4qFT2O5gzHzBAhrkxcqCsFlNGzof/y
Kkfy2V7LjkgQSI73SVRbzzy4nC1LLeSsfVy1QNrnLk1TxokqyFH6M/1Pd0aPZiSn
75E+3LDy0zngyRpjM+jPBj9G36/VyrOjQMfwIyCz3LnbmGVV4a0a5KUVWHhASaj+
+hdC+miVkuF+qfY38ICR+/JCHoomT1r3Jg9//L0YUFST0JDvSn/kTQ6ZbyT8wY9B
8x+y+wvB3vxtGd0HTXYWQkrB0GuRSXychaLR/I0LPOQADQxLAq1082vw01RLfz8O
nMRsjbsXli+eAT6sg9XfdgaatuTS5a6ripePI9lA3vL7hOJas6ieV5eBRx7Cf7hO
D6Ya/vv5kw2iXah3P1LXVx7cu4fJehFiK9j2UCyzMXpyHhIxK5wxygBic+g1T+Fg
zxLs/R+KGsRTNp7N5tpJLUR/OKZi7fcZR+6vWdH5Qdp5r5JKW9kf5qURNvVFmhTB
JjC53djFNZ+l6VXbsoa+9wMIegV2DPhVgyzgoz1/FLBGlkrDAug8VC++prxINOR4
cQizOWEj0qPpnpcVca/VFxc/47c50nm35di/YRbydv9e5+TFVnk0isKwuc1kCBFh
2ux3OaZm2AJDmC0TR+xYNRijaxzcDoqIYEu1bSLsxtG8lrlaNpjowyQr/ggvs2rg
DtUq76LKB6av+DlB91v5u299HAr1zJiRrkXb/OZ8H8CepGGjmUcRiDDgR2fsI3tO
j7QGkRNgLKrI4AhB96BsHIkx62lE1a4DFVhrlB/zo6QPsEZkG3miR1C2wSCoZjYp
n5dHwNv9VC2zD+orPsVLtXLVjezKCMPtAy/GUv5EnVTRJZ/i7G76w010c5TjIQsG
++A65mpjxqbRN4eB2f5WTXvizBRH4qWwTHpMYu5zmQ1QOlng3AI8NTYt241aaMip
VPELBw4B/kPTxpz4kk4l+U1k9vnM4eGIXT7eL/EScgHXuH9Tez16cVFk5BrPrmtM
+mB3X3YSzKfnubYdjVuNwWQLgTcED09NiZqPP7zEleigGABWI9/TttGNig+B+0nN
oZGuieA3Cr9ZiKqb4RxwoNrmRS22t8GvnAHh/u1xzR0uHthmGkAY40oSSzAP99G0
y2XNYnw6jzJUuNJp7e/CeCXiJHX6vNdjt2WRxBByebgwEjLkBCEobA/WPurVKWBD
IuhXHsFNPLuvJQd20h1YG/n/wRCxGm5FUEWBp6Oh6dFJHCEx0o5zDBVIYXuCD0JP
i4GwcPI/lymok1rpHG1hkhXhcll8g9IxEUwyMbbvTWyCgniGA21VaZHm8NItBKXC
BjlalgDLwRyeETxenLGwRblwoeMKbEVZq6FyGM5kx5cWe1tX4LhefhWJSq1HrDBI
3hVv1MCDYvzSnd6s7EsxmhyCAbQjw5BaDm1Cp4KLHuE+uJ6EuzWOnLsPHs2aXJ+k
WSTgWVZQkyuooC3Ft0ElxXNQ254124tPsCp0NLS1DGZc3ddlwszzQwUicKsqUdXF
5UrkKc58eoQgCAWBTzoq+Z5/wJiimFWmzcSpgBQphxNlP5pVqogevt+LOPNPjWBE
5/YjJCv32nGGqJyPIgdCDiyPfxUDE8XkLG9uln7yQietMkWtesq3gN3//ONFf1C7
LTbK+s8jO4+X9pVGtc4O/ildIsOQJdgd57cOiRdPso2ltqC2uamyMkJIsMqSszhs
CzLiDbK5YbNzbLVwkjHiK94WwmcIO4MmQQDHdgFJWZSSLPb8XaDjr7gpFeV+dGSq
lrCsmg84HZKUSSHCu7BSxYVYPxdZyafVxyUbOkTA0jMjuUAXcYZJ7Dlg+9xumJHF
iuJBI36rlREDRTRi+A2BD+JZNtvA0uDRRUtM3KFwdK/iJYmGGcVOUbQPI3zx/R3M
Xix0Ot35KC40ympn/xfGjmqCfp4l2GkUz9bKSrfLZF1Pjv7ELJWQBl0UBX362Gss
Yl8UME7Don6MIH1mFrKeLzDMaPhEp56lgOGcGazD9iuW3zOqnNotrSFVPWC1O6PV
cIY8X5Bc4+x8pXdfknkNpvTvR5oeJb3SOFbWqSIsYeWcP3m8WaKfbBl9Cuv/1fyP
eYEhX4BP+9zkOJZdNuZpXLne49v2pQkA+u8FAqmlfuzdP37V+b2CQTNOBLmuHD8K
c95fvyToZ7GVgPLO5Ji9yH7gp9XvjnrDaF+t6Aej/Eykz6bYAe2+zHA3RHaYTBsB
ClrA+/bQDf8Iw3vUrX5gXctSJBI3svjmfCAkyueCpBFjK+ZBdLmxnWdsCAYmWiCk
FR0Kb6ePODwV52Byo+aDUdqd2sd2frgqi3yrSSB50ZwiJPKhYE+j6D/mui3IPf1s
+Fi4xxuYOXB+SxpKUXrEcXupSP5C4gCs7zoNAzj2jgPknr30ZRmEKr0ovd4Uhp0E
EzuRcoYTCsAL6kNgQ7FCNGVI5vmMoqXD4ipPwaQDAfloIA8nsZHsCk8cXUkaySg+
az8kuiMy1jk65mRxqH/tdAaF0lvQyfOqEoUYOV9Ad7VMvj+BFcB3stt+UQ96KdhE
/7n819Gv6PxGGeqAt/eyjf3iDRauMnukm7ErNnICxTx4lg27a3sOJcowojR9j7wD
/artTx2tN4e2N5OxqySJ6ly537C6Vlk1COq5fB/skamI16LyCci6Ty8VUFUHe8x0
fDnT9UScxzqduM8xWelytzeSDsa3XLbnI9csox7s6P6T6uYiRkXMnB7VVMrdq71s
p7MT2zBgBZWWTT9FMtPeKah6A/6pl3+EBlMT+JHy7e/6jkvvPRO8Vrozk3oHUqyE
cOl98j2eFYpc4sbiUvq/iaESrOhTwRVc7bfGLV1h4pqcxgo0Ja0mDinT2o2t3h2G
yyIGppG9DhRDjRRHlORbqvU6kOXo6sEiUUeOl2fTG1VX9ohZ6cMsJIVUDB9mg+Th
L8wYOlRqyNu0+JG3O9TD4iHEtNJ2PVO8z+em9Tb7oQ3XNqsoTgZgNtwFWWdDH5ph
LrVNfwxch+9G6L7+mGSzVFcw/AYn0IbV+Nkyssj3BHCB8/jmcewfdaqfaiz5V6VN
lX7INasfioVSIUNTVaNTPF0yXaVdG17ap5gduQRB8Xe/E+hyvwi+6qfdSDoIRnEP
edNq7bSUrMawOMKR4CfWeuTcjS0Dty1vcPTV7C5VvPrmRKJ75bXuHGR44HW+2224
RBL/nQDGdszUV3YsyLuFxYkH9v/UIlnmqaskWarqu3J3hastuGtY3xrFLixAvP1t
sQo62RACuGUg0dA0aF0MKB1lamZ8B1Og3gOjN8UrRa2DTVvS1QwTWrDawz+jBkcb
l1C2ptWC8yh2tR287N9BBq5tlq5nQITDrVj7gw9eedug8WfI9r/uwj7RC0gNqwG/
ZejfcVSjOsGxAwq0kvPUwNKf6wu1Yr4qW1/cvo8diEHyBPtg31diG9hZFmeQuKM0
1TZLKLU8u1/mUuarhQmbk6HfLu+1q3uYbpCAAv4HiC8esxk08Ae3UahN9LBTiWmW
MWon0PmwpQQjJw0cbCgAOoBbsh2cScqm3PlEmkvZ/03TcIHyhKvhg1WLL9NWPNRo
PUuZ4lf09kN3yCpI1V9VeX3pgiDEI99/gWNlNE8MTNcLt3VwG7O+YROrVHhyI/bW
XDxFxkhTKbt7yZQEJ5fALg/YpFG/2amQoP6ptLodi8B0n+URysuGPtIr6kNNhNY3
VIXKN0lDPP1N54IPwQUvXmkljdlwbuGQ3fzFMwmsPnXEBiGrpHdpTqdS0LBGyOqO
rhmOPDu5KbZ/qGUlFh6X9BocrJhbVutmMPpiSFXyQjvRlY5Heq+ERziImDMbe3Tt
E7ssxUiwERAmmpBIBNPMLL+HpKnUidTuypZUpq0Xz5XI/dhghUrkRqFvHEsnf0hn
57jdRJB1cJZo+g3ZXPC15lmdM9Ej0QtojoJQUPljHqkGXxg2GvfhHC026AF3Nd3K
v3gmVb+eQBAFClmNra2EPqwHTYj8QQGh9NIyf48ZyXQfV3ueHbVhGb2kakaUVoqR
18IeUhEdNQrl1OQnLrev/UrXRGioBiwjr+jo/oInbrqoS59wPSPFAr4DuFL/LF9o
lklmgQKM+VM40VABXpddbenocRVVJHtbEg1AaajPrki+eGRGJ9xd4xgJwhA7/TM7
0DTvVeR+88iElHqKjWfw95r7o/m3PrqxyZrvfutLauGcuvTGF4TdbrQXkIN6J2KU
tdILoO5msKXsKMOJjV+UKsise7SaRwsf6TN3oWkQNWrdZxkW5K6K3gSL8ebY/PQt
TOSHDkHqyxql8c00cYiNLTWBi9TpnoNfgnabZbZQ7cX5ZwYn5AiJHQzZV4gZT3YM
xLGwwvvov9POryQEVVqDZ/v9WpdewQwhdHLv9fTupSLvfXw9CWP81Mx5DzLQs29l
tBQXAyVUDVSwQV/aA2UR0peZPLHD9sHqeo4VtVQKJsbcrmfJlb/bBNgfvSuww2Ds
f5dxf8F2sgUFkE5lyZdMrQ9NJhUvoIaIz0oP3Fm+YYd43dw+d5p9D2gvETgmAP7F
YeKMad24mXnh+Se4gdEs1QhntuW2VYYr6keMExeCDfSnJ4DdT/DGN7oPRBwrFHbJ
V/RhtcTbbBexE1L/vQXzd3yjM/ORAhDlX6LLxu25/ick+68HHQp28cq5VYGcLiTV
WToubKquB6A1I9g8nuvoCVcMHWrhhWfH5z6Ny3rFuun+m+D3vDJyhvRSVYnrM48Z
11U7tl0KVPAJzhS6bBIKvrHWH3DvseGS8P9+lf2H+HN0zOEwDbaloWtXv3Z+Hfnr
j9WJwzYtDB8ZTsotZX0XE2uAtIxVsf+bRRI4fXIQ0LgYKR/tigNl5bSGhouniUm4
dZAmgPVdi8D0ubZDCLalVsuaqPIWDtGBaWCnCV9ThZRljgEmWrBqUrwaHsdTvVjE
C06/pv3jCoiBZ/pSs2j4gct3nbsg4Ops04bhUZ4Rcqxhxq0FC+noN9/Jk7xnapG9
NJSjV8ZXjMpuqm47QYQLTaQ7OKGbhtrCbgA6dERGLI6NgnFhS8xMHDL0O/721BS7
pMigIANRZ+1+i6CN0qROpUVaJbUxd7u6Q4I4r0UvmZ2k7HhaqJzsT7LdXIfyRBH0
4OPqRKPw/+CcHB5MBHzBZCc0bNuYj5gS3CGVQ+TB5CSFYrC1Io5n03yWsJDgNuTu
9eAtp2eIdnDDEkULrMSsqgd78Hx76wQfuoKkNEXljegh1rosj3UAKLRMktsnEpr9
64rVppBO9r6robWHnGTc6InoZml/5dLFhbz8+7UIVmbBdoifGqjIZeMAs8H2MDDc
168T3AFKZMFZKGQHYx0DCCVyzVdpoNmShshBSujcG7F/bhpL7PgTZn9QeVY1otQy
Fr22eYM35Ere4vkui7DJn3o9mUO3K+2B/NGv3YNya3zK3EeUZ1rZdAZvBudI0WYe
dj0ZCEGKNJWYKMvW2NjZdnQMwFOrd20FETMjaG00bW5ybYQv3SdvAVSRa2g9XNfu
4EDN/tqV60khZnwkT5RqTpCbZQifcxeO5eqk+C76qh1FnmEWD7JTaaVi4KLMG2hN
8BZ9UmHGSUqzQj8ZwqiJZBPdMTyRBj16Hu4l+rS81KjhcxjTV4ZqdYAq7mqA0YDz
AZxIyFOVjyfnq3CiQRT1SleWmmJKFDj9pGjao2nQkome1XS91Jktjf2PlfmNnF7i
ZrdK3B1hrY0QYrt2Gv11Lg6VC12qRY+r3aLc5JcvgP1JmoH2xm6Q18uWSjwd4QK2
eaQRemf7k8CdN5VKZXhzhQavPHo1toQCgSUSqjj5nVvSDhWJPG/Etrxf6K14nM2K
x1BbCidwv9wwWYXmK6Dw6JZ2zGJaBsSrIedxsIof2BDT049Mk49P8mrh7IaLuGXX
ApqMAwCDyLluzjVzalFCgyGTnwxrJrJJLt0MxA5tzYZyKTC+oApA6guh6r8E+Ite
tyiw8YyolcQhjpPJxWJrdjkInrHuuted9HT5/tDgokDwtt29So1mB8KCI7tDQdfb
dHI4AyzinIu29xH0fIFtdxnZ+X4TxsKtuG5kZRIw3mWrPq+FWxglZM2HbT1pZoDp
CcgZj+drgvKoubzjVwpgKMABqus5VwuhgOutbPtCdrhn22xndMqb7HhDvPKKQ5H+
QPaLopz/2+gpCw8dcRynwq6UeFUcgKWa21lIjfriIw4ED5xULXIvgiKPiiUFyT4o
TYQaHFu2DGRDrqD5qD8kTfFxpeH1rmGcNh042Whs+LArCyHgIgh7R1Lg2fc8vtHR
rrINaJcHummaJDj6XT/RgrXGjaGicJ4eKimNJ+NOaYO5iIHTW0+mO9mMpUiexqkI
Wj2Jtc+txA5yid8S3fKk+SawfykY58/kMalHESpMyY/dKNM04UVDqc+N/ikCXUSt
0Qt2wbHZ/02twXP19KePElrv5oV9gW4w2hTmmvaUymtXKvxB/AdPPX/0QeMKOx/C
ibUvk+Cn6w/EGoysKk9C6aA6cQbux8LWmVavq78+o6EoB7aKy73irL2GzdUxcEqG
b/JSur7vW2ei1wXFOf3b/xA/ljM4L30Q0WNlUN5JEf4qkcdCDybgksJ38DzRcUmU
dne5bF3c/wtFKyFOGtugWF6c9HBwRth6A31xeYbjHnvNu2I2yFCbLjVtflCAmXGm
BnDMIl+U6k6AZLcq4OqQ05bnvMs5/h+QK1IboJssd/yG56XZJu+HIe2WHciVaMKH
+EEB85mjCE9rEQ39zUalAy97ReZp8hq01DKbbRqDThqaxPw3aO8fqr37MeI7WsFQ
QfULb6YIBKMXI0crAfPLHO8yppxLEv69mvyTRW3HNkcXH6p1nRLrwU1Rl0tlNQsH
NrW33nfiTNPP/lWDcTjRyFC+UAKm15fvkdSNqBnDpPbBRpnZQB8RXtCzAGAb+fzZ
grSdQExJJFgh55U72O3GBF8PNIAyRbF7FeyBbbVzMWuxJ5UwaXXR4WBZZXxez/Do
JEecY9FrDr4Ff+84X1kIplrBwae7HS4pzww0NOWfhaCBDFBbvHuxIAsY/uEZrr2G
C766E42ffVtdd2rPxzU27r3QlqBEKB8x9hrskxsFcFuwVLxjZIAeBrOgw8L/aRN+
n7KNfcwvlwmWEVwriFXo0o6YgQ4HMbuIOcj3OKLD55n7RHVvY9E5mzfIc9S5UBFY
XhamuE2WCqbfff3EpbKWdFISOGRLf1ZqnU9R2JasbdQlhPgjv1qaPBLnif+WK7Rc
atpJpnrye6+cI7SRkBIjcJ4/ZPtIWZNS4yW0y6rhOnd71EvIg1ualVyJBRna+7F7
gwXb3Nf+TZh+tbxOMR65l5ux0e1vA3Gk6BO5m9TSby9kxOikKMHDPK057HAn30oH
wCodFNzbEur0JNe9NW2mqEJQELMPhuXh+dYmTR1S4GWaQ8ivY5S10r9SYtQZzNCe
hCnfMW/fj6SNQGFaYH6Iy8sZui7eIqKMdCwaVRQ8C+NTQrrMaxDTDBw7wpnJeqt2
5Dg+7ThxhU9JR8OzlH5rWsIoLGlPfd3O0VFbVdqJgYqtrx0ibhyFGWe1YBY63S9C
yiVjmmHsNiheID1lCxAXLBSnpG1BbdA3RELNJazWfa+ThAtcpNgeBKWvI3JfxDYm
b3q/1FNj5RENqRNHCmOgpnfBhkGtoNiIam7V6SYQi2HdMwZMPW7h8oyphBxW3MqI
yNmeB+zhjq2MdJdWZeLaDlSkGLQOXrqIxhU4gA3+IlzPNJ4VGBIoTPmuQpfzqUZl
LKSbez6dHzkxCcSHO5H+72oP5b0Y3LN/rj/NPn6nzvhdjl8lftdkC7DD6ahIYOIP
eTHVMWSxkDwd449E/3yYaLhi6AmMn6tcm5cIXrtE5VVSJAFYiIVkHD36kwadUfTc
1dd1AOrxq0/2IqwQn3JIohyBxT3jm1Z0HYQt5nyw0+Gni9jDeUTyRZ0e46ENZGiv
nmOhifRf8I08bN9WtlKjWpKGdJgBmUEZ1E2KI09G1boL7ykE9FBnUF09l+qBKG90
TSl6RAeVYQhMIWtTzl+Ki2rWJoX3N/aCbHYqUmnuYUPx64r3Ceo9WJsAmkAu3gv2
YyIrKKlXCBz2g9bGgSNmnlCpxm7nYw0404fRuJrBYk1fq+CVOwn6rRUqlnXePFL7
fBGvZ7zYhpk4iOOYFBNy5kr3gOrWyFw8a8kr8gQSUviCprLWr0RyWrFn/2eHHUsH
IZ6p+PJunMHgHPvzXlJwPioQ7pS0lTQGIa7FQ72TNCfZoSVVdDw9hBm/MJ4tXynn
2m3Qg1RQh1BOpPZlwFFCQYhYDH3v5oZVjZFJ2nKxLkFhvlFjw+b25tP3B9FM8j0k
npnazyjXF+WFtAlZSbiQmpK4qzq6VZCTHprlFzyjr8i4cwcp/HNPl91z1tzU2d4v
BKIZR2CLdCz9RATU/7z0Fk50BNofMru2ygDehxrQ3bpxc6vUInMNBf5p9a2y30tY
qaurs0HpKqWh5mBHYqZQTu592yc7YXojQbu6c2oRiLtjJ5vsdVHniKQbN6l23Y5l
JJF3xEKk7w/UN/tOALZB/WEhLKONMS9M/ztcyLqcbGDOCwvGkfoFvkJpjdU/OM7T
Es4W71nXLJ3WveLJBxXzntOiipbqQ1NYO0r0C7l7GTlKIQrYudIZLGthnwYk7o0/
/7DqO6DxWxtwH/k/mWYYnmQ72exVkbX9K+3W4dVTQFpInsnXCqi7NvqF/zPHT8H4
+YOLOr1M6cmYNwAFI3+WASo3gWRywV2Fe7PhM+HkBQf+k3onvT7KpRWv59b01E6W
O/fAAhhbmDI6GV9fkmUqs8ckTe1vhHztIcDOE9AiYNTGpDsiAhRK5I1nhtjv3fV7
NHhcnLQokanYHXHnq3Cf9NVJalaBpeRLMkBVn8flHxK4Qht0DhpxFNcSAVhyGmYg
6WmpFw0aG1J040iJXtQZ1dEkPHenFlnMUl/DTXA8ZeOwnI6sJNn9t8LJFYS/UfRu
NE2izA1Dai+u9UVzQkwl+ysb/BB49TAYudrK34Bn1hmHh6eC8ZFkrhKpd0mPAzxI
4sHlsuEggBi9xZ8D4I4lhaiDWaNP+kkMkjDUUMQIT4OXYQ0hW8VZvwQ6nSvGDpla
xCsO2JHm61VQhIv0axB03Hbxp2oPybI4K1dKU8rXV8Xig0E0oc/cGttTbSB0/PEo
Nl1J1CZuBN6UtJLooNg4TkMNgV8VJzrl56FLn+ddlGcAKO+BF5Y6RSceUzlWwDdN
hH21TVlwBc5Zw+/uD9Br2pE112bLuyrBmQIuHgKNMGNDAegPrHv3aADa+u5ImAfA
Kd7LkiyY0m7IsonVr2f1wy8AmA82S4yS5ssB1mqyGRs9ltoXRS41ON2gugYXkzed
WbDIYdD9+/h4pJtG6Wy7lnsHAQxxmLYBk9uKYhwxPWSLJKV1q50zvchc1o26IjqV
JXSx1hCr5O6nPCSZCGb4fVCWxQclEHI4YBy5KQyEA9G+ob40fFtcO3Zr+RH23w3g
erB2BuvqrD76fzY3HNwhxu1RY22NzE+GTX9x3SmKwKpi1M5nZxQtEcEX9hs5iqqF
3VV/s8WFEz3esr4g+n63A9x1EZqC9cb7tVS60oMzy7oH+skDChhO3lT8WuIwOFrC
zE+zvUncyiur5XNvxFvCzvNz+JIeHwryqfC+pjsgILJFv2VEY4YUCjpVEL6JGGa5
nWc4CYcUXR/sOCaiKlc4tx9jqQGRSJy6iVezSmna6dnZyTBb6TwtbyZCWTYIvfdb
Wqtms5OIO6DxDdBOKWfEsbH7mFbbtgtSFtaVR3cyFBcJaAW1tfWBbSX54QtaU/Mf
gfmFQ30gLpHAQAAHWcjSZJ/oBK4QPySmkkbudIOCM53qc9cO8zdtrZVXbIPG7rQ7
h+4JIe8UGDxggnvNkvBNVCp35XiVN3B5dD/6V3C6QNCixsW4aNlPfKiTpEUOvKOE
0gu+AZky/D019zAcjFOYQHxtbK48DCJWJ05oPMPnOXakMvk40Swqi2STSaBfudG+
1b6UQqib9TVcpZURhHHUDMuJrTHUX36Si5leP4vkVfh72OcdJsj4An3DAL0/E9oE
jNWlR6q7tL5QRiz6aaMFnodZ1Xs/5Dc+vToti9IOqXkwcKURVjbW4Tg5mPobDu9x
432k7sBrRc+dtnpSuUdD0tAhDQBWesScTWwXLEJ6s3eL00oj20DKPpGQGaDQwYjw
JjTGonN5frd2a2GJZyyww8GyZGkY4ZI2nw2uje0kOQ5j/NO47XUvHh5rPb7yp1mq
zNQVxI+5lrRdsBlCT7f3leYWlxOQChs7ibcUr7/aINpw/GryOwJ7mTgOU+KA9IGh
YhyHIqSuaLB16KccmGmE4lD6wtFeLbX4DtvtNMSF4zWtr4gKdl9oZeihviFYgs2C
ShKE7kHMdOpfWKUBcoiTNOXNl8T/rQfk6xpc8XVtXi1FWHY1jxAItXTGkcYnd58x
uB/ZXUr/T2b8NjNrCC6eUBTqVc7eIQQqHSXLtCoddP/vPFkNXrt6CIddrhkHMSNF
EaqHB3CycqW4mVvB6uecdkrHnBFq/N1OkrqLl3LFHblJcbD7XmY2fagshlaH5ac3
1Lc5P5mydEePn2hZsIWQqaOxeO+MfMPNn78RnfWkvT50hJ9PRbU7/6EVUXQi5VUd
mb46noJ4Z1egvAm6sNGOSdXpq15AnSrhLAZBoR8NlKpZGBhQIWe94ZF25LGIBfHj
M0cONXma5q2p9Rrq9auaooi5ZLBtFyllOFtZueo6ljl1X603opbJZn8h6yUR7w4d
txMBk9c8K7sMD1bk6Jy4y6FNJk//aZoeJyFq3wlRZ9WnaXryajs1MKfLXQ2Yvq+6
YTZVfETUWv8sRIZbPo/PX4quplJosX1tfjAfFMiVy+JaCB7l7G8mHMcYLPCWoyst
wShY4MBsA9LH7nLRofZy/33U2SgW6phIUxJQeWhT/NFioCM7hDoVIbVzhaIWIaF4
ijSJ7GnPGYw9B4/8PY3B2VUWMsktj/qMB/MQuxsVFlGXy9SkYVuuK8t6IPdc75Ug
jFeJldV+q0GvvCBHyNe4Gqw41LCenUYZTHAbbEoFNjpWTNNAFh4ivJJbjhDoLyvG
hima90j7YGIC0MG5EDmMWPWoM3LxdnbbuBlFjQJUTvF1kHxLQiBwZiQY0U5HVsQP
75PEdyMv/HnIJsuVseGHbBr8jb6IoL4A4V4GX6mXjd0mfxc6Ws2bpxC1WwL0q3/J
4Va8nCTptztEK9Ykow7Vz/tvl0xcDYioxNuBjth2p3M2mVwzDSHat/DMwcIhTCVo
YRpHfpzkBoZobfmH/1sC3gEgzHVzq2npS7frAKewLAJRSniIVu87usoUn+TwuZOL
b5iu8M8r8u/yTjMBVel0cAJh+NLsnF1fmb6QT4GAdN0D02tySFlWF9MUTDjgHebN
F+Dez/5XRae/PTlqsdDkiiUUORmX8SIDZLXx8/d7hrTE3ddoOVMkXHrRMG/PAfde
nHb3G3/MJDT+noGnq//cQKZSaMhgCvRFDxtoXRVZz5XoPGbCol95JqzQ5BwXkrjz
dB/bQMGGbhkrAi2WrB4lkdaO8vnTTbBC2dL933+J76ElYf18vXM4ugKlWse0xdOZ
yBD8HFX6QKQovuiz0HJw+TQd5qTMAUYp9zuxliMLglACH8/f9BmH6Fpt1ezEXcX8
jXR4QDCxpU+8lvrfs3L5pKfhAykW2tYhHag585BpyCRmTYkE7YZNpwNIifxp+HXD
mVWvJnQZXf61nE/XJZX83RDzFBSFx4P9puhsCDiIsVzMVZIvd/RIJKrXvIqqhHOx
LwMS9ZmNeCywxr2fnBnaQfUgrU8TSasKwlRON94lx/Y8MN8E/X10QfZpXFa+yQgi
t+kyzAD7lHrIHpfEExfkeZyg1G6eAyLgFSP+4+Gy5E1zaXvoqTGNl+1XCee0Cgkq
yee7wg8OH5DfrZLS5lFQE0Qaj7VS3/HVXftHQ8xkSeJ+5yTcgMqGaWL1Vb3fJNeG
ZuhALpvGNxfeV/NsMzpgbN8DkAvfMekIm7SZBmseRCW3+DppJcp8weGHu4S19Y9c
4qF56mmRt/kRc5+2LMKeyIyD1rvK4nPMYsjG0FRdZ8iwC1R1ETACoiO1r9TMsPJ6
0DLKmEU/218lHJX16Wi9fu6uYrl1a7pLpi0UoLvU7wzHV4CdYrAvYr52RfP3Rrjv
LagErBlzA+f7nf9GwoUDmf7WII9W4FL0M+lUbhtLUG5nWF3VQ1BB1ZthYzNl07/P
ZUecuWlceBS24+yQhKOvdTyuTMZQl6+GZxjTSKl/NCre4h7c/KuRelcg27BjWU91
qf/tKnvEufYbbEc4kt7oirPyMQZdfQBS74vcls4YoJJtOsTNksUYxKqVRBg8LzMN
47186e9w9LRyCcFJHLOwb87iaX9ql18ZhZej+/zHK1+KZdq1MsGc6HyqowHvHnWE
CKu4+3c0gT2/u6/Ga+HaM1SOFkgn3gozdcNU9fEUYXyDFlvoC7EKoEz9m2Lksdet
hT4CDcPB3MGdT7FOdSJfvjF/nFvGMD/E+C/XrG1vkuOnF+IEw4t83Eiu1Z0eZFVO
qNytikiQnk/HzOpXlh44m+l0/1h9gKsMHuHya6rRxej+8F33lU9K14P9gexhvsIu
UhrXzS3FrVI/+yxq0Gss59w2nC3AXAbtXsccRdpg4GSyGFs2Zl6GgJbKpxFjS+2J
tZMaCZgmjgzrXuw9Y6bOWt1+uotTayT9luWinyEy0ezk7JgQNi44lydvy0i20MyU
fGgVcyth6Lredq4BmZ2ZeHiUihLYVLV2cd/KViNn8rVqeUbYEy6mX3ASSP/uX/AX
QSvXQR3McuTK+MNrVC2a0wzkblfzLz5i+5ly9AdMHlZty0/fGF+wlwWZcAF9FB6x
cp5iz+qDpZDnQgbDrYzvpEbXbwlqfSPH4irauevblc4xBuM2pk39bDa5fXkCK9TW
LbKnk0PLh9rjjeMteOHOKbRiDkyzNZTBWmu6ySXag0FfR3TdXh9H49zQct7iofY+
jX3ok42v1IscQQN1I02Biwe+J0EpHtGFs2MO/6jdqbc1SEFbILcUt+6kBT4UTjFb
MnHK2T4qAFzba0e46A4AZJG/Jl1AE4umnFumu9SCMIQg5LI1y00L4QVZTZZgRrMM
CdmPj6NeqpPuhs9gryoiatM3YiQiYymcST+LeUIQ0aPKq0WueFVe5O95rBcmT2Pz
6cy47C8ZLoMMxOZpixGaFVhG06//vH19dIz0qa+JhW0z6tI/a8oPMDCWdRZ2UQev
ePyAEaxGEZ20sbvUYAFP0T3cjaPNHdYFFeT33dZANsi/FbzldMTOYz+rEC7g/Hhh
kkBP6r4ZFAeH4qFkgKv1A82fHCOCMd17RCate/6h4DciCRXxJru5s4/GU9CwuYz0
YdlirI7CuIsaQh5GvXZxTFZYIjvmWDe90BAquZfw/ayM7mKpO3Izp1vo61nlRWIy
c9CIjNSPAa18Nq13aQGLjNgCaFVn/P53YE3AGAXsIjGuBVzbTlKAUw7m/aPLaNjZ
a+GbACd5/hR1q5BRjnql0wHqIXgzZLYaEcN/GsIpMO7eU1N6GDnbQX1+CnKNXXqd
r9RrFAwfgoSWmhxE/kitGHAqvO3x/c4mQBb9T0JErV4ewbzh5IKOyCGGlK4EGbRq
UpX8WJ6FbzB0mcp9fOyG+mnEtVwl+dB4yArQcH1Gf0zhkMH/Z8n58ej1wVxwDerB
QNqNDjDTYF3Ns1WASOdlsy/o7ZWYMqtXIsqmthbAsVGB0Z5Bw+C4i5fJJCLMKVuS
9I4+v5OoJzp03Gp03kC7FHZvufSvoY2yANmO3hZSdFi//S9DYzDJ2XXRQgPwkhKd
oeIMR10g5yn11tYX6Y1COdpZcXzjpYwZbTOd1v9juVXFBtyYbH3ncQBdOZnX3/i8
XssJZ/FXZBpKCTDrtjAXE6OSTKdltuiAvY9yfgyXzMUMfWCf17OCwGFzIibGm7fB
CE4zubuiX/Ck5ZIhCEua/kVii1fcl4+o/g36yjsoDlrC/vTqkvg4BFigADKI4QQG
nmXMuYZSseA+EZmeIGpIceOC1gVPHmJwW0j2uit+RduYth0o+8BE7P8Y/sciwBz7
5vauLrC97K+bbdObzcg5w//vc7Q86EkTbOT6TpKmKJAdimr5XRKEx6XEcYtmYDD7
Ke4V4IhlP3vAl4aMpTsYu1azOTHJDFO47ULBbg/jzO/Hq/qcpe4qX+Spegl3X+h7
OSKe3aYaxOHT2faxnA1BG1CVUOBDPPsvzbUYTOVX5qszZ20q9YQmWQHkZa9olrmb
Zn0MLKsBnZuR/uu1n5iq3fzmTTinnKvCJdFU36uvRcfKRETgRVBFMb5ouvBaDHDZ
Zy09q47PgDD2T4Kid6KXCoX61PoO1xCFVtkn14Z9/A12Zx01mKhuIfxp3SKHq2M0
Jyl4XoCrdCIUN/qD6yTc20+TrpeXtgXHJbK7genFdnr/4VkHQB5fuLqDFaz5+8R9
DO3gmJG8ip7qdI3bqop/940JhGrR+MtqH0atPHErkxklekTllk7k61n2rjCSfx+g
YfsNJFH2L1uh/tEBP5JkunSdYeAH5NFsso/gBMRqXp2sAyHqZ7NI8qMPT8jj4D5M
DcRQDMccR2qOwIqLwL4UDe+hI3OPIiLZgEiAp1kUgPGjOa8s+u71jw6fmdVS3OxD
5vD4vB1gUapLt6l9ejHf4pgSi7vmW2arVwz6woV9+1WlDhj7rTxI07hl3Y73I5nl
LRO6gukTMlaglxYeftkiVgZnWnh2oYQKnPVBh+xC5/XLN6V95BMhoPG/Mq8UkIi1
GEhgFbbloZz9whTYhAQIHELm4AdJAWcoMLClebXNRMkvQC0nTpsm0Pl+RutuVCTi
YzGK91nzjvH0gnO5xLNG1R6Z9zyzpXEPxfRfH3HHXO5i3z/8JW83QHc8rKxSb2Zq
fRDBjQM/IrR4vKOsSrTTqowzebaengMcCOAcVZCQqgqVx/4gKKSGzf4dQunfbScU
X1buiTdwgljEQhoT2ZKthOKvrw0FyS1egxzEl2tVEIk1YMtH5BnqiPC7bNBJWX7c
o/O+4wj4AFAi4q6ro0t9SjKbQ5xrscFAaLJ0Fs8l99gdXon32a90FjbAeYTj2olV
JYWS7mEqL+NJ+0F0hNPIv/Q/SPobTYg2M0F9ZY3DAcRLFqJGaADe/FoIPW0Y/nm1
kISTkbw3DoGJ57iJa2vsMaK0bMlqRXO63Wc405cPoDVOAJ3pVkZpHeP6Rnuk7h2Y
2jzo4vbx167cOqAD07xhYY61CiHKMaDSiaBG6UQdlKPGiySLv4HXxtva8ZEBq9Vo
3zq2qCL2t9JuTrALbiI/L6Btw14v8RCogGChIHFqTlwMqI4NnzqWKHu/pG1/zgt/
UKAFf5l3yxFTJbbMyaojR2SL5RzJW41xw8vQoL5HxAus9HbieR+1EPTzZwjXn275
xPZCvVSg3ZYqZuLQ+u3hbC/HIIZcYyUtnZ5MZNi33JGITzHN6tqg2VFl72TlrRcR
7s2mo//ZFIxdPp2b7O0/jTX6IzwtmCVFFemfLAJiMSIREiwYnbJhvL7lIJDtPktV
Qf/imoTiSpBMTW2VKM1cxBJLxgTl4ILSVz71V959koF66xYTSQdt+8gfQ+kPCuUH
jQXE4j9SyCiBc7Mnb1H5Hj+mgyls5p20dOu8DTa+CuHCHzYrsjus1L890q6ZYVmf
mcH67XSEIbqw14c+acTArcCnUqHUM1ZDtYgr6Qd1abWZfZRSzduwiMPbihYRs7+r
D6DFQcbBO7ofQWRaaNmvhebzksZHs/k1u857NNYK/mhgQOAuCqoaoNFEAv9DDcbT
lp94uGf8iO8lAXDElxdkFn3Tj7xrz8AKHBwFncxy1xoXuvE/JjtTWNYr96xzsRlq
O7QPagx2v6Zax6rvmq05SUjmdy3d6kCYrmVmoMR0+d114TDRwDtnP6VerzV/GsPJ
4wzX46jxStXPkGi9wHjw0jNVHiy0Z3j9QoNq2dWkP5R/0VdHldx0xoxg+wQT0UKF
/Z4heiOhfg0fjT2Sm7jioeKKcgR9Cudq/y6LUFwrLtWs6IVVJ4YVqJUyFdqwRb8Q
D+dLoFfFSVV8NklwgGcFdQfl7v0NZLFaWPRotPpKjvx4weLhnS16HghRDoV28VVQ
n1mdgZg46/zZSqlaBw1QODK1083v8Zzc8dTZIt/HDkz63ZOzytD439jUOVJ5cvoB
4BSS7vVFxzSs1N3uEUNa97xyHNx1segXsxPsyTJ+PwizkASTeiL1AgGggjeEBsFw
7DOlSx0I/6ptODEwxI3HQfAA4VPIxRarJy7L5Uie/WjCcRYyDJ8fdFJHqAgt9L2p
0Hu47NVwpfw32Q1CdpvNKrZiLIFCZR/dqK26HDZhd+tqGqmuS74Rajj7BomkXoY6
lPOS3zzP493eGa7VWQjO30kWEP229FQkre6Nn96akSiIuEKhUSHCfhHhhDfJdJdC
HN8wgai8mJW+Y98K2/QFLwC9E+nLuxKVX2lmeo36CqQW5Py4CXrYCNCU43NqPzhv
xKxlEL/8khltwutgVbihgbvUr/GA4dphiaF9/mhGxO/iCBCtFt7av4EGSS/mn08N
xQl8HR4ZmV8zSHOkG77B34f33R+Brr1BPsNNFlfB91H1Ifjm2vR4tKBGYv/gaCEr
h7Z7fDmIjT+u9EYpVM/Mzm8ldkjOhu9zoCL1fhTMlmkWgLe4PJTkBa8wvki0Rqv7
LUrZidEfwHUVTUUalpwYHDhgo6ZuQk2h1g+H+/wHQvllA0ZTNxm4flAtjYalPifH
m41gXUwpTR1jRmm9OENmq9Fz5U5xL1wWSF6/l2SijOCFo3dFim1ecYdGkGsX3zmR
8wJFjqMr92KAlJywZOEcu1TUhmOhrNJes256hzeg5UMlvszeVLG7U8wk9JIIFUUW
9RBvit2cgdsTwWj075t9YdLIsx5PH/XGhGDhhFFb6yVWknmhiKZ/+3wvG8YiAB4+
rWqI7uCWE6r9YcGPPYb2hrNPydniJFQ2vPBcsh18PmBf4Ah3QWdGYae777phnlm2
5zPsf4rk9edeBEAuUMew6wFditWGy41rlIDhRcTQoZjdS+7PUVfSv9Ep4Po71PLZ
oTUBspaLUCDP5uccTaJTR/teTHLBSqUFOcATqymrUMIyihpm8zceJqhfhMrtfxcy
ClSg+Wz3hTHuWt+JLcUjiDJjxJmma726PWmLzy9lmKjYHx5K6lCc9ZvZuZfVNOxU
F7BfcDVV3SiHiJ13LVeoZ4j5bfKJZZ26c4Dvn+RwfZ88r6wSviQ2sWw48m0QoSY8
MYMx/f1dg1znzSTcxLDEFPIloYyaBBCGg76I5XsY7kvfoud6CCczqKa2W87Ibiz9
QDttpUwGDB5PFuX87Mz8DB27KswaPo2i4NsBWEwa3kPtREtmoEHf4mOOhwaxFTm6
PGJpt6WNqHl1ZUNCd0hOCKCM98VEBX/EUNudiW+5lGeuvEa6/PDoUeXKxExYy1Yf
Tc1DzODdjcdpaTrEOC0X9fKowSh5ZWtRn4kDcPNKE1RNEAPzArZ/vF6N+L7V01wn
ti2Qa9dDhv0gKB2I5ubs6ORinpIFxw0m/7ToNaR9WEIypIYH2NQwmVwc7aaDo9sk
PQ6JG7utT0zw/ZA/KYps0507JwkRz8eSVu7k/0D8vTBPg3U5G5+0f0TG3NSPfQif
WSzWvIOuuT8YmyVu5I4BoGAW90HIGXHXMZSt3OoFBT8WVMnD5hW8Ywn8Kpp1Pg+0
5NGxQrXSbLEAKrtHOlvyENH9oYRliH4MXLj/ysqIWvX8JLiuIihXdKtXRnwzkSnc
ffS99zp6ILbCF/g19TBn7TN6hEUGZDjRenY76233h6uALjV7LI94G4E/CgL5hEoA
mpos3tPIkl0KqQgG+MkBcruYrQxTEDURdfbSjhq3KOmWp8kdS6feLgAh1f0cDo7S
eIVlvHyUmcTBvwNkFIR/srIPErcJJKyAHdz2+LAPDWDd4VnN+6mb2gYn0aU+6TUb
dbeQpHjAdIohZQaPU5HD7lcGUvPqmi9Eij0R/Ll3bxM70QbJymIPOGQVky6KbLGm
qDvrvbw1MVaCkZ4GCei5vPT9cZiT1nKameTKuN/7iTCrk6Ofysd8KsfgjeWtPQKw
hMmTZ74i+bKA+R4WRWu2dqvywxlEAS7lbMFAcHifZUdRFiwmQ2oThUshoFFA25tr
5EFa5jPo2m6//Ubo6GgpcDh6G/sJUuGyKguPZqh1yqAwjpIjJjJNtls4WcElj4jb
e62UoQ6831fkS7n0U2VNO2UHgcL6TKNKVAQ2njrQmM6yl59eFT8RSx7LBwSH67LC
Gn42IOES8nS1IjSTmB/t/11T4lKK3bbHSW7+s9jDYwYZKa/SEOUFkKa9wv+MppZS
3HzP6QcE2U3cWeWUeQuVgkRvgy2vlSAr4h12sAix9QptMG6UcsiUKojiqRYOdD4W
3oTAPEbMGqNZ88svkFdyQc4Z0rni9yegEOqpkgJpvA+uadCchSvxGf8cjKqrLQ7F
ibMzwNRbji/x3+3l6AFoK7yuf1lIS7ywpq152x1RNS6EC2QNm57jTGC4fg0DJWhb
dLN82R4pzifOonAn581YuGtZVH4D+38oQcZyTzdrtYPupI9OZtdC3F52WrWJoInQ
glhWhFauBijiRC55oqKlFss+8cccuuiVSpsE6ejsCbthuSVHLmeV9txE/dUcRzcG
IqT/YyYGvonbcVt2WZq3IWoDCV23f1n58/CemP8D7NguUz09doxKqclnAFjC9NIf
BFfKbHU+J+Zod7LD0oK4gsCIUJ1F1cUNkkQUdM7nD54WJhxrVisXpZ11t5kgyhqc
P/7ZXSE28Vm7G3QCBrrljk43LoIXPMKChfc30sr0XgnslgcTV6T70Iu/6y16aRSt
iHD+KpGxwlWoQ8m72SOxDrTwo0c+fS6KwUPEDxnwMxmu0arf6p+2odvrgeCXhhok
+81r08a+2AgYH9H7SdsRINl8wCwqo9jPjFM8WTNlV8iE2DYddtFVLqjXNizA/mEM
f+Bf2avLzjexWIL0cTNlB6qVtWH39WSGUblmSbw3emmTRClBK/Myv25c7kf4Km7D
U1wZIrnY0abWnY9GUejoY0Q/kxwlPnb2J663QlwH1lTeI4IysMANiUZqYXDHmUbh
hwJV5ty+D26Wkpm0eOZLkqzhygGCowbTb4PZDYe9dvLcT+9hhYok9FdT5d0gUpHl
e6ZavpQRp+9aopPNpYxQdtx4We58XjsQqRNVSqsfMZIOoc1V1Irc/ues0KgJzaG4
/mlJz5YJgqkiGmliTJFwLDSAZoqH5tgAiQO0GNQxnpnKP5V7DF1uNth9DdcTbG/4
OcpCSGQLKzQ1MELhZdrbjc5yJ6w07yX+Lcb75uXsB++GGAuQRnKKCT9GuywBgivA
+N7SumsuaXg7Dj6PuKpkLfWMGfCyGWYbPeUeDIVyqVodHN19gd6k3cFUPWAlVgm8
3DUOQQ4Se2AV3fSzvt3m/vKy4eSyJRB3C5+EoY4DKl+6Aqd8fsocwKK5CtMnuXJe
Z7dcRtonGyscUmGKZWg2hPN7gkQfvKtOWKANK1awK48SOvCJ/bLk8jfIusbh9Zgx
WOZM+vxXbtl85Uqg+EdSQpLP/JEJoB3QUViCTWSjQbv+h3FAx27zaDPSVTIbWA8O
WmwLptzRlkriEu8otX8wlTAzKIEVqfI2mYROnDDxX7KlxaeN7XSFn8KpVlj985kt
0dlZ3t3T4RcObTOYg01E/YWei2kwbUWPs02tYQelp2oKFZWQyQNYvGvTtR7YDkW0
TUGB3EWorzHh6Pwey9a6sNEKt0GwGvHG+uTW+7hZ4DOWjY4iuVn4ZNAT4FJ7SkOd
8hnLq9fJ/E1Th8MTrY0T3dQxgKU0Tq/oS/iuBYwaa1l1Zz6saKd/UTYoi2HpmhpO
eoQ/G0hSBhngf/hcUYIGhwNEaMWf26mO8k6WkNt2Z5neq/TfmDP2VnKbSMOfU8/B
p5VgCKViKFEFKW8GgmuaBAuw6m3udg5kk/rEZy/okyWKIAlbXcRIRH1UplORERsG
Ba0+pxSqJXVWoKSuZziCPwnJd/Hq8I8aLkNVaD2ay+YAGXGD8tkcrUW1wPXC7OUM
wehhyEAC+3vZZWz/5lL4JroBjZt0QvYeU5qAwV5Eq6j5lhFtsGndPI5kIIEqeiXh
W88X8FG72krvZmeQcwilNYojfl519DawfGLE7RfWEsCs2D/jlpyyWyv+AbDTli7f
JBejxh6LH0zZvByOg0rT5XGPxSodAU/vA8PsU/aA3+s4HRg2Oq8T8+tOh426+Jbd
LWZcsjFm7q7ZAZQMVMfPalVgq35TZYJT9oeupbxxQcqwB8XXyXPcGMoXSh9NEmL9
+bzT0H7q9nYiTEvcGuYvf5TC7P1iuxK4Dq5MmsACAUyrKAraGFQ7C8xscTnpTGHL
lN1VNhqiJ6qcLOgvdEfCYK01TlOR+UeciqGxjcbBKnoosYAn6JNnHWWuDtF3vqSV
Am4bNIOgk7itSC2m9pyoVAYjapmHHnhDXbn+kOBgrGehOeQbhd2uAqf03ZgYNkj7
A9Y2NC7Y6fKa77IO/oDtF/976l1nJvcivVueZ3yzbsjtwRZ2yCXwGiyYsA43RzPR
euqVbIPPWNWDo/oD9oE9RizTgxr1mJNJVmBP8N/Tz+kBxGlopS5J0q1kM3jdDN2H
kfGS7P/GdT3tABh+AjTVr3H17rrqDXdQwcBdrLwKXeEAnIqZqzubyjou6SELxsvN
4ugvzqawKUy5Ly5BQDzz19ITnzLufjYoRYQHErk867XfyzPJ8h6/3y88wuQeflxz
niYtX0Os4Y6Eo8Y7HoiNwAihqXappHgAo5zRniO8piEuDxRPjdXokSdi0g22YyhJ
YRhbPujFEPIS+ncsu5ySAXdVvlldLjKie/z1mm9plimS3hB1uRyAWYCm1oeD7UgB
vaLvsj3FZvmaleOB5QtQTHt8UQnMku5FFPke9cf9wV/+eA/qrWQ8ncFtsPTaH5S+
wUc/9dpaTG6YFf9DxTT80PDgi/1b4ikPyFoP3cJfoeLGZIqeqJnYpqwII4wjr9a5
Pe3SkUOaeoh2I5GahZjY3XmKtaXpuK+dtQn3CuL3lJemOxnYiXoDdCRz1lW+x3V2
Mx6O/2NkZ/7z/JK5T8PIiGcJ3XfYpn0eanc7ED8No0/6GMzVAGdd3KzWXkCKXyv4
ufEGn3bSC06a4RNE5cgf7DJvwx/Lu/CyGrPVw0owT1zgRVhz3L2Q0JsBSMGiqdzJ
GPz5f+80wjCKa6rbFkldBUNaMsISziWMHU1N4Ak1FCWJZMckSMg/7Wlh7yLgbf3y
jB2b7TVt3ffbEqqaD5iuHLGWPEmgaUhLNtlDMK27Do6N9BYBmqvRM9cU/V+jTabz
Kmqd4mQh3dCOt38Wv2BS/WfS2dcLTB4QVIXMWRhkKD7SWBOuYsimDa1opnD7sqib
zM9iwWbh/2nSxwWx6K07lk3Ev3In2R8lDb3ZYGhbKAW6j1tvFYylLhU8JWtxlXsW
/9wPRO14putvdH+kaCrJx2MVEFKK3XGVRwBSxkFpWZU6XwN6Lm15AYrAzyL65KEJ
wWUZWIGLdIW/hhMylZv9pSRBpCJIHZhw88rgLmzK7lQTLADtkEehNpvL4FmNoB6P
BzAQ995nSGIn9CzXGGDI/9pX7D3eVwWDLnNxh6oYENOFoI6BJjTI0WlsZgGk/qdM
4ssq0bk6+jabFH2VIseOABgC+FjoOTPLQRMWh0IlI/lVPfz/GSvnbc92wGUY/VMt
0fIb8NoXx7fJ6oJrOYm1BIjp2F5FGgtRYwa/UJCsOrgDjIl1cVerI6j2qwmeTo/e
dktBREIwjtPI0NTH7qJqIdfYQuqNs6tT5L8tIU83K7F9/TED1xqmZ1q78aqfPu9u
Wtk6XwmZZxY4bmARJBM74mU8Tiueq4j/f6x+z8Bg1CkFUJiTsjFe42lm73zAlCvN
cqej4GllJbV02ORmw29DQixJ3b+KHzY0y4XlN6DwdpHumk/r3EK6zFAnuKEpIsTE
ikNevnyGjooLZqhyUc4i2qvVAFq3slRAXfMfMA/YHjBAth5YWXsHpmo6KwaCAEsT
jWg2Jv5Ytlp0Bb/ssW04KJ0lUtEEiiFAdiUDRtWDwBFksvGIOZKOyawtiQVhNvVa
Io41q9ohy9le1O1Uhpy4DX4MKaKgRJEzpahdrk6NF7wcpBhNkTlZeNKX9GTITv9J
H1IGCf/Rmha6RcZaA5OX7wpwlwaewkD8CRyqlagb6a6H3CUORE4Nx/RajOVi52Qm
97okLqijaBjWbcsMvKppir8GEIMacea0hMvdPxu0f4glXdhcpjCoT4k4xMKiCcrN
H8qRC+zQmv8qDoyGeaa92SutgPs2ZDB+s8mRTiV1YNzX0O58I70gB0etJ9GGhreg
iH4brn01PjceyFgTMV/F6Vz+mn5oF9r7eO3BVR6cpasum645OqzzmP0VKYay3Q2i
dbHNG1GjL7DUw/jF9AtBg413+SGR+/7B/Ealyx/irmaH6n1eSy9rLflx5cg0cOoz
jv9e5yzRQ9SgVMVHaGFutOxV4f5itpgiLkAfrk6vTlvOszc2ftAQpCXVzc/29Fje
f91/9WR20U01yMpmmN0GvFM5oZyD5ZPlcAq5Iy6Dipl1V1zXxCs+1RKDwWrV7nPA
ABwOgeHkF5wdSYtWWllBsm7ruvf8AXDKHJXPOXSwXP9savnmbYoDb0C9T22Te95y
vm2zQyiIQSqlGpE8P4OADBFxwJSehpaijVovmZKo6qsHnZblizL95PSo/vrsbxR2
qrx9Ii0qiq/RvFN69JUguWgVT1u85yNg5dmWUjlLV3bpb288z7ZIt2BdS4jcthqH
yzcojOhd9XvNdi89WJkMc7WblzPfNWVVV1UXgKYnnjGXx+VcR4TvKixAltmf/zoT
E8pZhw9hZ8vDRBkLrfCuAbrPCr92qmV5CfgymfDYgRS4GEiLsfKMk4SxQAq0Agwn
cfZfczrMiiJvQM4Snrg9TsZc5zeQpBuBsDgT+BLvT8ozmb1UwyOmaJNyNTNiX0Wq
cmebbiROXi64KDS524Y0QJBH1bwvbXNDMQzZQRF86jtJ53kl1ECfHkVpY2z5HhOz
Uea38N5UGGPFyT3rkG6nJit00PorvA10yrZMuh/r+BLQhqQRc0uydUhbi5WAT7Fi
083mxWJdJhvzWWCDhWu0U2kjfUBG5WZm4h8oPc7O+NvaFyCPWqJMu1XsEjqE3+DY
jzkWDRnJ45IluM8BsKBeX4N3wMNbv+pUL+FdwhvyAlDeKLOOKLp1TCqR6W/FJLLj
eLSWTyOomfQjpoEPS0SrOK8JWkCroe2B/mdTI+FOpnNMs9Jsx0uZTnnBVxDSLlgY
2WqWTv7YccWZeBXFJwwOGu/MTvj+tY+L+XRStjXn40qXh/vsysrn4hH47/MgdhK9
MgOsSClQHCak3QKUknJWl85jYFafH3QOOkpJH/NrsPMnsUlA4OJ1id9HWKwW0iiE
mSeUdcTnngcIYPt3jjT0WUmk2YA2kpCXUvKuOPgM1Sbkp0HR+Sw9vyolT9i2gom9
Wfsx5dVZ07bG8oWxxkpDJCCIlcx8YVcdJK5TwdDPh4HZRYhbt6BHFsmBvyFXSUvd
/CG0fOrphKhpxKxVUw3hhtYl2FpqBOUkn3g6UHgu1XeokRc4MQjBIsO7wHuzSvEg
618+EwuCy4IqKlszbL+aru+1za2ZftXRr4n2p5ZT1PZwZOvHMcM2aOFifdWqlRFJ
ByTSIuXkmQQT3lKEwvAnvXfQRh9oVfpJiwDs8PF0c7d0J+Ey5vFax6Mmyf0cCqqs
UJXHsWMa92SwgqWvAhuG4ABgALxRlEfZOwzXk64zYW2ROwaLt8zRmsUrF3Bwu26B
EEQVju28eF7PbTofB4vxIjAnARc0MRKkqUuSLhkPzW9NegC2OBPVS2Ud1GyTy5kF
YPeJLSXZmdwPPN7mvygQhfkBGW0x0+O63HrpRTYf9geuvBGv9NkIPsfoihblVpXG
GrxfLiehjfyMwbcqlRaLJJWjH2UKXOYkyeTTKsPyevA8k2EAsu3eFyK0eLSpyHBA
XTXQ28s8gBkLXCFKDIkOvEPo25Trw3bLmR8PBaKgsaHYs4LIyi4JmJxkhoN6QRvs
We9PDGDTFmyk0otXGyIhPHMO+t7bM7I6AqUc/VGjDDRazddTMhEiJOrZ0cb+jLFG
CCMhKr3EoN8WS5hMs86jt3gPWUXdNLcg7JeSy+duBxZVfIWDmV7/MGrtuusn4/sx
bb4fA2+QzDeXBynOWKi+AuY/d797YZsh5u2uXeRGel1hPchUO3Q+K94yQrBKCTeg
fM5d8vEKF2abIIvauqxdnjnc8XBzaxP8NE/9HeIK8cyKI284zu8mMtSAfsB3/vjz
cABJ6srOGJQWal1g2BRBmWJJpTHHj2glyZdn0NySU/dCfqSRTMg0CkCXdXeX44Yq
9b0nf2VuXmIzbeYFtJyrgOoLTY9KnHuPJku9zBBZGA3awFrtx32OiPYOlje7BMnm
G5985GLvyhB6E1T2UMrtmBxtlMQq1UDJfIe43XteUmfrTfeYLQ3CiCZ8DO9xYoYG
8dnPGd/ARrzoS9ywr1LbBwygCtA5/Xzg7cfGMxtSw5BdvvX6GgW2AMvbKHhgOC5e
Z03Po0argCFNhf/F8axInHxv2QTzPj2/boPVHCuWvDBIjyBCaSrYmG3vNkRAoSWD
LHWNJKRQn4L6E9b2Mkk50//32RIK3TEVMHrF5W73Z1R553ceZqB+0qmLyg8jTw8M
s0HsONo7ZL0a+ujDIZ6O160FDZLYOqf9w6B35JwLUUop/xb+/but6md1xug5VBgf
gnIZKsH/fsf53C33y3js+4RDt0GYyzlD6f2iDxB1HsM2P/Szoe+M2bdP/6X714Ay
hiEIXfClCwGtuIH39yqmtwfgjpBLyJFEqpespFdApgmMtXmhBw1kBthLcPcBVKWq
pux/oIGhwObLXKJblqEefbICSZ0/KZAFu+MRPPMinfcXB3q2bB/Q9GpWM495Jcr8
9RzIKGzNSHWbm8QjGUdoaXBPAzw6I3MdysQENFAFd9EqCs9AlFkZgZEl/qjJy4KH
YOEbHuw+HEjdgPFyigqCcdhSwQ+I3mxKVsadpR7yz1makdPRH7SXS6wqog2vjgzi
QgviGldbzQE3vVFUBKNOBMkrwjzowGmpq+ElPlKFWGmZ9L4tWGq4L24FMD773x5/
+jncZdRX8n0iVfzTtGHFjSTvebsFHODhNMLfedm1KIcqcchYeuRYTtTt85IOPY0p
iyL/Gkpvyv5tdfqXu7CX/HZhcn7saELx4jtD2D4EfnKsluQCFkeJtfX5Polfqhr7
34n9F+IwLAH0ajUMIeZnHaInlLErqUruNJ4ye56+unjLFycRKNbuf2fPND6+bnLO
cAlmdQWIkLo2lOngG31TwZKWrwpYAEshfssG32+Duvnn5RNFkF9kTXFMgh+m7UzY
hH8jfp1kn+A4Uuly1hgqWfF9jDPBIrf7CmCG9xDF0u0VXB+LjgqR0ZY1tpSIBjNy
BDC6x4beT/qiiE+1Sz7NVrKMjxJs2GRNU/U30ajuatZlSbvCTYyFuRM76HFOqHkV
WZkXp8WJ1YaI0HXCaA796RdkslyCWsJ941a4RmiyQiQ+ifutOOCoPeXCMx9c5Dvc
n//pMRsWYuz9nHOyvZ6W6jTdvXRdN0Reuy+dUOxuaByJFa1a8l/KItPD7TducT4D
l0j93L9apmfPJJBqi7snBT2evrLWm7SF5yHCEB1nST/2LmEyF1QXKPP9EdMdtFD/
tz6HL67fk9LfPAmaSngzQLQi0byA97raFoTQug0Y9IcpSBSZzDmra5BHyWEDPDu2
aazbpVVuOdasTd25zKkO2e/dE+SLaeG/MjQAjuXevETYimh5VoG9U/fD0xezdciM
AblTWyWvINBHriV+2dmnAQ==
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:39 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
icmIjluVq/U1jSKP5/9IcddxrQEEjn4Md/aZPYLxJbNYIIaI+gw1fJtZ2bS1En4x
fj1lxczqjzT+8VgqQT+OxHFl+EncB8vhuuPXmSwIra8LQick/mDO8vW4SohyRPQ9
ZuSuMqhetZHjptNsZUESpA3ti/Kedx/fGcZHDujG9PI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24992)
h67IADxHB854zP2oe0sowZ24wDNWau7hHx14wgLrRmxFvJeyAWVNM8uXUCcN9TWS
pGh6cS22V2WzC8KMQBHNeCGJrWUbm38vxvJtMG6N2STYgdcvIrmLeInBUYUdZMwU
oDgsqrAeh+xcgzI0DTEX5anA5DK2TDBnRMSUKXXZzNNKl6hJXVq8voNkKcByyvSu
QilmJPh9vqcLeRPZCh1xAq9rhMMQ+cNu3NhncGzdcPI9p840WOZDGFh2BN/kHcPp
A5GkQeT6mbf24uwoC706MqI1emdoLUfRtE5bAQPv6s3OtG+3AdcKK9/yoHCGbQFn
yIb/5usBM1BgX4/wXj5cIAw+rVB12GcoSYnloK3I/LV9Mv65l0UU43BCZFQoiYO3
rC85KtdxdBdGjinkJ0yK3IDhYB2yKzNXFGUBDuPjX/emet29zoB00iX1cJq+K1vC
lcepvN+9P/3ViIt6s4x9qt7MJNpgYBsoQwaXGEM0iFx37/2BqjIAUCxNJSx6Fk42
/jo44cFZ4NCmREwOym+oaa3A4bgEfsJOGIpEcOnhNcvEmfvbWgwkYrcQN2CTXVcJ
xvsYBK7KsGIHbC7ZSAVh3lnyvCYNDV7yZ7v5C4S6gPm7vRe6RsMxn7pI/oqLfZ72
h561RdFzrLbTRrJXnotlxrOFHDHAx+CWNFKk6tniCHLbjd+oecCpaxh/rtDbovcI
wkjb5zPG+qdBSkwILDpOWzKUnwHggV6otxxTYJubi0oaVKhMlw80naJ9tglPeVVx
/4BByxm/slp9Si3H3f5wVoYfoT4J8OqimZS2h/UyN3wjJMF5KK5EcRB9z/kiWU9K
A5RqYIE/4HRaPR5Aui7762VhRdOZyRU1rHz87fuRx4GlwPufBn1Psz+OBEpZdXdu
M8td4sAroTjAGmY3eVSMUo/8TgLfkXkX8dlHVS4xA3oGSZn8wJEuMqoVwk71t5gB
b/vIdenzoDAjh8fZEhCzkxEL4I2J6TrmEwsCUqkubRJLnU8m8JwwIz1z3723pgGt
fX+riSDbuaRW0Sa8ZGueHCRf2N4RCLgtn4gy9UiW1TivT6E97n8l0hn36jQC0EgC
N7YFKZdPAe77JbFkYlv34GYTVb0cJjBn2SxrMJwO+2pwF+hTkBDJtpU5gVi0KG7b
/H6crqDZM77PRcbkCVO01SQkeCakuGG+R87mjqr13ZQrI42t928++wmFx7+/4D84
a3cAVOhgjnewYzS4Q8ZirOkCuzKftXNyCxXRuRRaVMmbB2qYiC8aNFWP07Tq1trB
IUQ7EfaCRBKXIw61L5Usugd2CE1kUKh8Gtg9Hs3z++nWQ3NHpZYKKseFAZuK2GVh
H5iDShhQxwWQpeqySLAFNLS3teqzfK8zbI/tvqUipljVbk5YoMK/mFdm7pkrFsUq
8kzE67vgeE3ZxXWsmKpj6LmIp+gW4Wag2heKAacjIRMKgHJm/A50D3dYiPaR4HFF
C9fCSeqEw3J4gOWNn7nTVTO+dBQehrKm63GlL+2S96v5wZSG+u0TVwTzaN9fc0Cj
ufGmyjRsyaYBzRZxauzrV3tBwmo4eXI9EwByKp3+ekQHsFrO3snuXoX4NTUG+PMw
vUWfmDO8TbhehyCZjUtzq9C5LTgiZUQ1wAta3ziPW8Gv9fIbdwJIhoTGqbmV0DXG
wgL3nT2xa8ZdV5Tlw/xaR4GIr3vH8+pMUNHyoAImeZBxIbcyLDoeqH1nHzSgq1Vj
xJnOU3OSuX/JtnFgfucZgc6XCnwMepkMQZ2+eBBxl9q94iPkiWamtNhXj55iVl/t
dY1DmiUn7BbEvxT8smfJtcRy2e7QJ7V0LFAdkQY4Qm//7JtU0OLFqwK0ptTD6g6u
DbNAu6FPoLSZ8VIJe2hT7MoCe5LsdmipbGb8/o4u16O/nfs11d3WkR63TQ+2K/oB
G3XnHstPjfAbKCCjKtgeLmlU9aX9fLF9qV6GLGB3n+4ubBsWhFIVahWRV3vFLLl0
LxF1gWv8VfG2EwOLsRlR+I/ouphoxYycLy+Od/2Gxw+5fI+9ryV0QyGl+weNwmCJ
82Wkc+mijEUx84d72LmDatPCtS4o/BMK2U8F8h3g6y8tQu+bJYCps/dBLufi+BHM
3vZaKmDh1MmrUhZPEdBiGZJZUxUTBMQUhlQM+VQUPtwuTKHrgJcPECDabIQvBXwy
dN9Iy+ib/PTsmsC8zjrW3ZR1ZWF0eGbdIq+bVK6jNTmPjzno3e8fMpLzMjFdTCM1
opnQHu/v80TLxaZxI/IkFV8UdL/td3ZFANiQ7uIjHg3AsppUsGo0T78BtlOPkgMH
ZCmH9Vq/PIZxeKf9l7KSyy2Vt3jJBZdlaqsUgK6hAZ+bZ7jzKkor3o7/AOW5GIlf
ezwMDthfTtCFIicE8mVjxOEjU+i/SPtOBMAN9AtsGyfH4vH7Mudoo18IY+oc618Z
fMlq656j7eIuLEk+lPquwSCNgoPV1EpUpX43PCsC5FUruvANCZ6yXGcGddiE2NeU
vBpkoCZGP16+vpj+74FGHnQdI4GgD7rESmrOQdTsjqxorr7QrqH7vgGXVWrmB1hq
EJAB4S3Y4jQoHXKf3YoR7bXOlA5hNfmmhrTI87H7ENZ2qEOvr8hcU0A/gpUZ8by5
+otGEhpRRXZkC95+PGf45iAT8DdWNz5pgZtM+iuHfV6tOrnJfZKq+QfzXjgt028f
VH6m66hzX0dbLsf56aH9V8mNM9XW8OM9+qqW1aFVftAue3wSeLMoD2z22BSz955T
mmFK2hlBmit2OJGGCBacenXJAzNZ46wU8JQ4PchoiERYo3ZFQcDszdNFCcQQeR6T
h2egb/9BOvCHCNPh4p8ozwi6tSXf4XKKLUzahjWvUU4WcXWYBFED5tnfm5adlCae
XLY4NqG3EDhk4teEe3HWTaVSiIocKGvLozCjQu+TU4CcVTtOf/VEGwqyG5z+SETC
AGZn4KrvyWkFzhbKKJx768PApLDkNc3RZ1nD1YXsypPmdnSsRNhGzfsOAGbzGq02
naGc/GI9cC4v7LGVZA49cTg+zw+UKXTjrPN7bu4XEgifiUlqjdVshdV7e1kWHHCg
piZlKtSGDeJCUTqCSbwco0sUaaqM55iECpObSOcr1zbyMoVsGBZN3ulm6+QA8p2C
RgqUl7kQ88KVjlhe5a/QmgPorob+OxiX1CyKIOlykAVIkU2ZssX4cNi5rnfmPDVE
MFBUJkM9KzoAH96xMM8QjeMvyeq5VOAadWd/yzZgDdHX9ve5OJStwtuj3xmjdCiB
ey6hVaQSuXcXxKNbbeHKR8k/ediOARB9JBVDOAGvH0MPL+GD4cuQ7e0Ojqkh+Kmm
HRccHGdFSvfY75M5M7adhFy0bTKZcD877jped+K9Wo9XtS5xoz0whNMt2V37MxI3
S29wIQvOpnBRn1gMUXvGjaw/PahFuzdtOh5WAPO5ibychfHmWSO8/i9Z3JqeyqMW
pknU2DqTPwzXOAMQufxxiFYj7eOqYIvCiSR8e8bFbV7x7C3dWDeaXpJQM7JgroXF
8annBW0UphQ5i6+C7PQJdeNQ+N4MaVEWHuF1Xfw+mC5JDtDumrpfjPk+gyJtlZ3N
vEbuZqBQhvpTyIMe4ESxmEos6nKGmTD3p9GlrrI/8bKFiTgxD13+wy58hxahz7RD
nWktK5YfK2F+fiBL0MiTMg9jQXnNk8gWHLYBLmLFAKl/k5IhXMQ2pYTa+Rrtiaay
PCUbSJUsZsNakhurP2AlNY6RtLe8YbJz4Zv2ycT3KpMGwEt2UAsCZL9nVwibZFs/
oBlCUlmcaop8vo4pS+6lV8cM+Uhdpo8zeQsLVGOlQe1siSyY5Xjs96IIfBZbH8Pp
ijyRookCsf14ulWT4Q7F149ONo5VGqleashVYqB6eRmWoJURczrPqgQShLogaeM+
Tj7RUCqudJ0tXMyAsrRL3D6TReLB6RffkKY0K3aTJyNDdRMGrAjz8A0W6RPEtfUa
QOt/sbeQC/Rj1+jBKcE5RDwXVzCFDQ5BgnOQw6AYL/VvRvUqLLgZ7HEEk6OAahD3
UopgE0PdhRLQbvTB8gc7P1NzQ7+8dmAXRoK4+BeyRgrBZvvE8nSF1Qmdq+lXcuKz
RROzx2YSzQAEEg9GVIu5Wzjyo7N0e8RuaoxhzSF+09CefsWmREtUqdGhXuAo8NPP
1aYF0xR7wWwXke0AJQMIUR7jMwOD9scekB6vRcxs9wNXxPy4sQreOh2nB84p6AKi
8mOrZA0GtT8nLP7PGve85zzZJXTK6UILVTizjIBFRFiZ6RI5cjNLORRUMG5IhQFG
clj+jrG+7EocDkxc2P6u6kCsipK89v3LQDft0/hYvka6hoD4x+ZpwHGjg3h4MtEJ
0aTsiHoMrfjFlkllAoYjyYfvy/0XagPUdUbV71T/D9IuF7yG9U/SQzytQbOepqLB
HID3bK7a3rvPMl794Fcfr0Sc+5zpwvKyX/FN/0xCrx0nt0vjZMxDoSLD8coOtyX4
A9kgfbZt7VbB9i8uArD0wjJR0a6sBt0YLtrFPNyb2ksxzf/OnhcWC/JepGQ7EywP
8eyjtRxzAsKe9PE/zunTm0LyfPH2LD00Qt8MVcE5kO0ubShgu/MrP/cmmclbnirz
ttwShCJue/FtgJgiJc8K6MS+cRXnB41mdyXeIrbDBZrIjziVDVLJKmT3u8Y8/JRk
YkCJ20d4T6gA+N7Mf8MXSHuAD2/WC/i2poalnNKABhSVZgQEYdjbH+oSnbx+zZHf
nAVqtqFyM4dlfC5+fvkK8vkFY88gu4H4Xqp1y7TkEnxUmuzIPWqHeNyL9+QPRDCz
EmkZ8dkqQjMtUDlvUNsslvDVgabRLGFLqvxdRTSlFmFeBws9d1cOX73fRqcH5z7X
YnZj74nlmGBd4Ze/2b6dhY01h7hPpLBce9dqR6+Y9nJi3de3SPl9QujAXbRxtvIh
JWRSVoELtWaQYe97CvP5Gfwc0rtB9xqxW8wwCkkXaStcFghkisSG3PxwiSWfsGqz
GoHlkOIDPXU3VX7UjGZvvcjeon92qgA2SLDInTjbXGZGOUp4sXc+DpD5lVQaqH4y
D++v25/L/KOfGRqqV7T5C/QNs12yHCjXiH2UhCzk8nQEyGlqFA1bKZk1jalUCHql
V7oprfCFspafJnzf4ELbF5tLiWA56kmLDRDIRzpr5H2pEZlUYl2gszA1sbx7QODt
t61II3i2sWFSbWikTh61Xc8rGIpuAtKHYstIyC6PVZw0gqZ8EFJ/VXB4FXE6Xc5s
MnSx6LPhPBrVz6giWzl4L2hd8F846ERS2YEj0URfF3pT6ncxTVLWMD8u1InNMV11
U4+Kw16QiH/yaUEgomY9X3l8eOQ0G2uW9mQelqTuTyojihT8TpXjCB9p1ox82h8P
2k6O/yWsZ24/sUX7NeoLsde9FE3FpqaWm/oZkZBjjR6QSgmjjh12n1pCtUjs5nep
920vdyJZyZ5ra9zXQNabQrqWkRPg2IDCQg2Q4/boriexD8H8Na4nsDYeKReljfZU
JBmo0+eFBX0gqB9fUnRmq4RFXprJ6a7HchG+aUWpNVBv1JFZkZ/ki9C6HIPD+Uh7
g6/YEUtf1d1ddD0vUAxQe0LbeZxHOFowWbZV8wGU/gHMT0N1I/8sZBdXxkejceJZ
GAcyVNN9ktBpSmPSrpCqkazucJoOEeluTsumB2V/2U9y044l0D1lvWrAjzpYx0Pw
uckZoC8iiF/wm01MECviT32lJOC40XgwPnuy0Ln0OosapVilfroVEO6YE6/bt3X2
OcG0NqL2ZMXSdPiXVFO1OWMJOTvUsD5+NucCmrWJpFPXRQGNjhg2UnB+cpbbC3nk
4998E0L2oM1mOkZqwJly9+nNLwGJ6u5ntxdmfYs2rJAgY9Wf2DepeBkrW+LXRAaw
BFUnfGK8D1rCj8qdiMkNV3nnTOsnhx4KEzydRhSS5LyA4fZuIai90Gab7ujvP3eD
3XuHDRnXfpQ4DWAtaLSpObNCmZVnE5SxqwLshu0fmgwiF5K9Yv5qlkwOSSiIRqnj
4KtUGhyAzCQbX+1QI3DBTllUjK71mjDhbHy+bWMGwrwB/ZIwpgI6xFyECKxJ+q/m
4Cn7/SrbHs1o9vVIWMVug0AJn4VWXD2Uj+5khsdECGkraeNKQlaRTL6zR975zifW
d5P6hy6AavXZ3nfyjixOKPGkWaNCZLByLZHA3RXzA6Xh6G/Ad/qRvaQosnOIBZhA
xFRf2kxOf5TX9q3GqupyMar7UhPn0YOjS/gEl0MkrxGlPMgoyxH+X590O4KK2RZA
MhpQp5qZe8d/vzSlvQ3ffpmiifrummB4hHcVr8aOCOiwZHg2fiewlHdKzfC95z7u
cojepinLW1x64GMuvknf7JP3r3G4UtpdZs6mGz0/+c9DoM4pVeOdR0ChUdtbz7v9
+ab+LiEx7ypORE1ccDUUrG4MyxJHJdOh63Up+XQMKZ1DxE9aUjHtq8IsuO5zOyfr
1uuhiZaXNCKlhdXlzyif5TvYaCqzpVGdH608KewdqGl2CD0En0ZanHMrKllNjdYA
v477QNKrSFuQ7ua6qRBm2z76GBqVTru7mL6IaDy3i4Hkd5yG/8dga4NBkLkGpMs9
GMoIppamy2O1CBO2RbIGSjwhX3p5XG+QX3mXqFmd8zj/WRW4g5/2NM8bMW16PMSd
OJy+YcZH2pmIrBfEYUxG4x2g+xRP24wvIyi0MgaWix69g6ZLi1zsZD9TR24XoHPj
YSw/fLMbUhkhJrDqcTjvnbdgAD39eSaraHAz+ZjoknlvjBHtaOpjU1SCwUHifRcO
0O9g8rNTthyXn+lfkBvW9PMfIDTzvs8loxM49zc+AF/YpIaHDPptWrU4cUB1HnXY
o6EQUE7JWrqdMsJH7GkNuLXP7Giw7a1e9YOrTFxbnfoiur/ZiU96flC4ygBcP1qg
Iph5faUjU1HDvTQlCKJPJhPRiRUNYi9nqHehxylxtbGFr8j0BFIkpZH1cc1EPxMB
fL0KPDsAkcG2BQwJU1ppWQ3H5FNGXf1OAX++6gb3M2VuFT0Pp74eEpYLFZWTN856
gbDQxkT6fySmXkrkjZrDxt11OgjtxTNldBmNgWQb6YGl1XsBCH7qSnOQyp4dJz9K
c90ualmKGgZSy6UiLPBi6fwBqC6Wa+bmwlrsEO/Fg8nBKNtNDxitSI9cvT5Ny9Kv
oVCx1ywRQGp5NJwovAMLHSlHodhoWzfeOxT+wh+ItLprqmOt+QhLyoSZlQGmwihz
7w5K2j8+jEaNDtC5LNmpzGpzI4nr86tbV2EXt756sBf8XwVx7HgTwIZmEJNeERE1
OE2lUHgHzI+v2/L/4mWxWRSfA1GmbfHpaySQUbfiPjpXI6tqZpSfToAfydW0DaVW
wS77HQUykMyYwE+1Uub992l2k3ryk0eHOoX9Sx1VtL1LMawV2xzG+7D5qgjEh5ay
voxBLk28thaw0snpNORzbYZIsLpnhnxFIGjHiD/zndyViotRtNajjN67XTHtHkWA
CwgC2Oo0KxO7QIgNELHClMOnhXDYcuBl/5orJMwK9RoW6ca9lAG/bJ563vD4DaYN
wIz82FgZpXdmboMUVXsNcXsmkdYScoafcuIES9LIIL+WQ1FgG5f4P7/fZpdwIlZV
E8CVODfDROTALugs4moHYI8T1dW9Py5/3TeNk7DVqHITGoeUCdZrZ3HuI18rtdDC
Q++SuBV5Th4/09zgM+HZQl0ZDqfMsnrmNDv6e+GvM2fKyhVP8TALZ1uBjlbPAmJC
gv1adjLXuU8PBBJ1v70E3/E6LLFYl7tf51AGe9z1QGiTQoyZuaGEfkgDcF8vtPjH
1SE4vX8TzcZOIJg6W+Vlg4qc3iJp/8ukMVihVFKFTET9WJ6P9CgGLrMWWLv5I5e5
hdLgMoVr2tyYFLUEkwo9tAAxTjwbofTFwfr03gfcwy4cNHqzIUHPgzZFOvtvmgTm
ug/8/6k9cekDLzFIgOElvL/xZVg5n1vidiQV7DloCEvbUMDDUJNAxUIR6tVqNvp+
oRFfShjkbwlr8wtT0CQTu6QivO4YXztLp9o3Fpw6LKC6YOOkctpwjn1IS3YA0iCq
DMKt2bKwtogcpG1Oh5qktKb4UJv+2QJg8kfr1QUKdNvDe9S0RdKvh7MXfCrUXhh9
SnXHRD+QxW9xS/yM8+ATi7QMPVWm0z9Eo74K37HrdXOTNUKOt7Wrmf3MeBwqZ/K6
a8yHXYjbmiRSSXFfRbTqgXR388T5skYmoe+4KmZHaD+BSfD3rUyq0wOpnkYQMSS1
tN5CHLN8dBHisa03rMozRMWQ0BGfLkEr8Y7wmpkDt+T+oHh8vdlAiqZd24rUY6Rd
x4Wpt+JWawWKZ2KwhLpVV0a58h1+rydT6bMm0v0H6RP+V7Fd0WvV7n8HVju55TSW
DnlxhUZI6qxoVpPyVZ24CE+JvQf+G3ai/nB88j3am6eKTxhpzp6MYGUh/sdhJ08Z
Jiw9y9zhbqSa14izvUijpSMJdR/uxFaWWK+nSIKnYZU1R0LnlZ3oR06FeFoVnHhl
oQp6IBuVe+bpmng2BWcxnnTiirZoBQXSaMt/RVGWyBbbKf8177XT6u235EDtqhnw
Upa3L96AkpTgRAHKlIgWf5n+DrM86B53GNe4vcr0tQh0z6pugRf44HwZtdqcpif1
tjiY6V8YUt/EPME7pQeGSbjtpd5zseGuCqYZwg8XxbKL5RK5cFGWxu2AsFpi3A6m
aI+OTB816VIvPBLAbzhwWnAx4TcknDfvWScOgbW0mvn6scpknZdyKcNbbUU2f5mn
4pqGqqwZ0g+j0pY1X2hoU136LSmqQBXptsVNTVYtcY79RQ+G8X275EI6xr089fKL
DZcu/NaQ/ZGmaVEp+dxywg5YEf3KlOwYMiIun7Ir+08OQvQNftih10QCj2BqOg+D
442wooBQHoUmletixp0SGbDb6sH2gcpxMvD3CBsC1qG9Lzpk2dSrgsIvFCQ5BQCe
kP3qF8k7QHxuT3D3Jlvq9LkA5yQY7xMLASOsyRJVqNYhNSpJf1ktmDUpSMhL1i/L
OIimLiv63oq2kz1U/FDgG8R1D0hiqYldjZd5e+B9SdBoALpk4tjCQH0zGUDcnyZ4
xXD3oEbxaJKkXNo8LZgMRReBz8fAzsNWnA52FN1pDeQ3EyTAQ5mAWaz3Kn8G3c10
VVahETf/CHBq2SM96faELYiqAh0oVIjPIAQ/jvRTlC47GK9aGwneAn5nvyHCOgxE
40NDRhhzn/VusVWwJLvZ4VhjbU8aucSv1iIfURdZ+5hq4GWXqTcc+WPkmWVcmVMo
E5LiOQc6hjbKdUSU2qAgSLd27a5wLjPpawNINBmILwSXLbavtp1A7mRbZtj2lZS4
PPE0BNg88ou0GBee+E1+SE9G3OOMmLqG9anpvsbcNGkvHGHPRa456hDIiFjFEZ0X
zt8TVV7kSz6/Leq48Bt3TXY5BAqKkRvQvFdN/AMEP0wcv/Fofp7YEONmQXmXjGtO
FnXk93qxAjUy2dUyhG/tfrWGxX4X/63F2wXIXF5aEhhmxjDSTprAwRtL9GpILxpN
d9z+CYOUmFCJddJgbcXKBNCEhr4aVlCpIAtUko6MR7MfcXCUMGRl1Bg6RRixeTEd
WtRvR9kJx8ay0jLyJzTLnjkXpTd3J07zaBCdiE7mlU1/KeMU+jFL3fuGMwy2xp+n
RQifoZd3Kd0426G6n9vOtnlLWjeaCM4SAZkOC5US0eMQlQm/3yayJJR+LX8pIt13
M8o9u7Fbdgn1qjWACDToonJJdFXtZX9OH+3O6/Lvkw86VuKgj8PvneSkzw4/Pavw
UQCHB8oCGhDhOl3+tqkoV9jRSRoZF5/RCBELli8zUXhvLKQlpK3h+pYXTB2sZSNY
guampchTDeuDN3+ObXFh3GS2tRmK9fASR1j9+Je/C7exUStw1gC52P3X9SlBTBpi
6hVqdg2mzwc8AWzitrtW0pkCzb2e17wHgdk3FXfXk6jYhTkAvqFRxAnIIeZnfpKy
YuL3kyw64vBoZgGwSJ/HxkCjpe7aSQQQ7IiCOSa+6F8lz6XyjSycJijjrg1fYrTL
B2uqrTnu6QYqxrIAtl+mgza1swDlcfO7ClwaE2VdlITZm0b0nq6coP6iUEVYoa7R
W6BDkybfvtjdWNhKdtNvRww78fbOEyW4CFDlFMVEeUxh8qx92jcWzdxtBtW2rAq+
xtMf7SBABZaBq569ATdOdHM7Za1UiqD3+FHrzx11ITbiv/67Al90AkA4unmVOWNR
+h9fl2xy6/d9fV/CwVNdcnl25SbTmRz8f872+9vVZL8nyYE+5Ho4oZ0ARdZ5Qghy
dIMOQNPGZsIBxAUIxRB0To9qNl4f1IHkYPp0tNHT+76WO23A/IDgRzNF7+k8C7Fs
1GS+DZgK23TYBhqbj6oZ2t/jyxJPKqIOdQKZ0SqFJ1B3IPkxRKl4ASUzcXeF++kT
Gg+xEZUPeWC/SqUzTuSABEVajmT1BuKaR0OtuuLhJ7YajVvIwaDH6j4y/jqQgdWW
2YDZx369H7RJkhS0/2YGRXtdXduLp7LU5Bkdy03JLXL7ISGUrNDNCpOJFyPROiAF
3dfjIbKxd+tl+eeG2bL+dB6Mu11vYk1249iQSdudgMPUIkxm3AFuB3lgo8Ws7rnp
s0VmYfe+UedCGSV8UEJd1ITeYZ1/lronOQJ7GWdhVItv4a3uEtD+4UcutNT37xeS
moh2dWcJ9GhAHKdmAaSBJ34jltH685lUhNOba2txP2BGA0z+AhVCskm8oNKPpCGq
wKODh8/IHF6lRc7pu/7Q1Ub6lIqJ4qIawei72+tvtdq2jsUGsWV0eJf1z5xoZ2+9
9aGzdnHKnVR2SECp4gs9J386yMk4Mr9Tx7V0DQLNr8JDOSv2q4Sq1Mbd1Bv9IxYO
TDOhJP7j7leUMwT38allXeu7BVLGZJmWl5LQeQbFuMjyB2z1uejFCEvHUttZmzbN
eWJEPxluoXJf19s1MKNBzaNeGDXMq3cABEfzmYuy+REC6w6+WRbRCJwbj6aWyuBi
p5tMs47KQSP+iFClbVk77PxYozE9nLy3dRrqkWpv/+ffep7T0NRU6J9jrF4eYfzO
DR1yu9ZFxLyhQqmBXG30A+5j498kQ6Qhcu1Xi+7dviuUb/8wOzGywkwck4ljQM63
L0uySmI2vlNOmqM/yzDXVmUE7Ej+29WYIgZpnoUht5x6MRVVDd+grWkZXeOl+phS
3eLaMqksVmw00w1CDGP9VgE3IjIPdIAARZlsnio8+R/GSJ4kmIs7gnDqfJzg4UWT
HzDFZFQwDDQ31pTCNuxvbVkrZaQE2TMXCbhodz/ByY+tfK6N+Hk1NjdH/u61wmsR
BKf3K2V6tw1tH/MrIAOKBEFrvJ5fJLTU2tIZb11ZPaG2IeaIYLwWCE3JmiRuPFbe
BFXAKApUVlyeRvGs3UW9+pUfuhq1Geq+x8NB8kujJfP3r7yFshhl4CR/IaEDHQ+M
69+PgPiyJdmEH18uCgs5xhBU2/YFekntnHkG7M/LCQ0u3SVP9gvka6Iif/5pj2K8
2dC39u6xHre5GuwMpZICHI/DQYn6RuMECK9PEXwbl+hCVZzFbHbzQMMwokaSgNm0
3uE+Kz7TXQC+2417BxrpMMKuH47r+jwEwqU8L0Bnp69ktDwtq4fml600J0XJxhoG
Dt8c0hJt/Degt4G6s41CL7DDXkDJDpwKNs+xjh9vdxmaawy8TocY+CYCw/ILQDqS
5EYNEgxiDWJah08kznZ5IrD1ZfkzAoV2RzAL93xwSrK27h8PUdxhy9EFZcfAKWi0
fnAHmkfEvZ0gHPjQrduIqcOtsn8N6WkOSkKDhXYxOiqlfNvdw2sJKbMjqtjw3g91
C5BjlB4oI2JZ9iwPJEpLNiC6Xh9Ss0j8w8iDym4vFdFSnzbe9297Jnv45YQydCqp
pJXs1FJFz34m+V6g7mjaoDe2f7cQwCMsikU292ClrXq/0kcV7yFyNlMbzvP3Cb7X
4CrMIm8oBRh3UpsbYz7ksi9D9/vUODGI+EG04T6pwrGg5Bd3Q9c7cyFkmKMjWM1/
Pqh3MzvgwtYJQolKDmPxdYbbn6uOeQGcBlhWbP8YWzkTFdiMzqY14bZrBJBF9OMm
JEqaaHSsBlCCqQVTcSpZxr6D8HNFaM4Lsol9RlwBJ47R6WdROZ0U7dY9ILDyJUKP
3dExZv4HlLAbYNnseAfRz+16Aw4VeInlvqqlDb0bFEx777iq2YHNWq4i4PI2cMn1
U4j4vs3AAoZirpWa4DMk5NfMAujyFckNBd5S3ms2SMOKrLKo509bILTaaio9mvHl
XOyldKg5gTDq0K3eUTDu74GzpLVDjZuXOI0fB2OWNY2f+3ExqPDM19GUMZPaSmmv
aLJQKp1DYM+D1xKSagYYi+rrrY7sFa8ZTmRQxO5LVUAFC5u0epkRhc8Z/ujC7nwZ
6k37+gQnTq/KD+nrnxqxNNahzswA4LG9N6hV+XR5VGBh6WfFUcImynww/baaZ0cU
9TMbz96LmvDkPEZl1oQwqazdwuKCuDXifoAz0F3m2pcx7rsE+RsmW6SVgz9SvCap
IQht0DSqpxbtI++LcRltkSvVh3jypdREr1JqKb/2W5r6dbdQYt1GMf9n3z5x2RAe
FBqgaa21LtCatTvjGqdAehP+8pPXxuW+6Wtv4rcdAxlFDbocQqKxXGsDEcauD1Mo
ygVHTwV1+P99PgOXNvjo/wOqdqnHxl+BYcqxE9LSs/UkX+9ygrtio0WvAg8VPPx9
rPQ1RX9pVEPxT8SV7iUyF9rdf9D43t3m22zFrjasLAvgiSoTHs9As3qGEEv3REUU
xIG88ofaHowlHHMDYH7dcIjbKlO+SjT0KI/RGMMKUXoUcUIi8D7FES+es6TO68L4
7nzLa9nFak3f2dX4+fRFBW91dse55j/4JWegX+KviPRkYHogLiTyWYgWv6Bqfg18
jJ2EoWkmfK1UF0K1tNR/Vn6OgnnhfuZD+PxGm5tBP6IikYs/ADbQurUBzHOBoW1M
kBjbWbo3YMUkXg2Aq5IfgbZ7C39XW+ZCcWaDZs8EsjpDiNY+EO+EC2BjCVmtc58g
IRJZRSg6kFEgT1+UOJ1d0JfmH0FFborpjq6e497eTQe/kD9Bp4SQcVYQtYyPvQDs
pe/oS/tWSOOccKv2Xw6mACYeN+0CoA/fN2do++lDFVEm308BV2GuDib4Q9Dw+PcF
HiNwhOzDAyMRnUnmu93oNjZYoC6BhtbSdIyht7vpcqAH8mzu8fT2lenmEXwX4yT5
dduMcfuW+tBGH7+ZrW7UMuoAxO0KJWHgl80GdU2kjgOUQ8mzVdzRdxr7Ia+EjID1
PfEW9n46GFN5UMmis6EtVpRezf//B23SwtGdqg0ghbmRKPhCv79U0pNQJmp7jckk
KjjxjC+YtSiW7nwURGhih267l2EmcjdS+wo+JRwmOO0oaHSxuHORnpWIAkRszC71
2W3QFZGTMJSb24E36wShzc3p7OCy4w0PUBrDJ9T9dcxvNGPjyMGIHHildjHeQJfC
27Om68+nhZfucTqiJdnDUG9RkyrrlKpOjqyy7NoXMOxxX3aW4ICyxYSDnI8Z6nAo
3WpLu7yxhW/jZLKDeQAQ4uk/TQLpMtWo5sMX14lLDlIefiyXgLP6+dRE4ZVp2oCL
srksAof0IFfdQR2i95495nMlszxgiNPR7sJcn+mBFGIEHX5V0aEeFEPcOl5WgFpQ
LSS59zM7mR8/u8r2kMLlk4ybpUzTP7ZzrYBPzk9F5p1dAygiVkIh8hpWny+Krxmw
vzTbrAqiWenkQ2DXZ4xlphO0pebuYuzO+0OCgLLXPut9ZrtRCJsdnFIANGU9akzJ
fA7UFKXKxiRxMmeDfoi+rBPgt979qJQfcIykOsdyPH1HfMVjnTJ2yucPElfjyC+Z
0LcezyNDJQlhDj68lKR00r16h8EIzN6jmkwKRIvAhBlHpCnNztck+Q19NQsmDxPJ
RhiAEfFHi7w4KdmTqt3jENPzbDtXjv5/iaAddZNFbuDb8mmvs78tVF6zqq4vgLGz
jyOgjzLiyyOs3MCP6offj8v9OX7CpOSt6smdAwAk0vPVW4a7DHfdW53bd6qjbCBq
uHPW7PthLYApEPkEBbsFwgZLp2SeNqI2QrYNq4WaPu6W+egAQZDPFXQxkaAWSG+y
x06VGG1a1JpbkabFZ8jnkL3maAgklOPM0FmAn3SkrJ0H1iDUjB9h82ed4G68iFfu
afx8OR1OdMhPgNe4qrewwUT6g+73lXLM7Gjhu3iRyN61zoa27iKVebivAQVSuo6e
h5WaTs3fuuVX/eLoK1aEG14rpy3heg1e3dg41pH28J4BhClGpdqhVYMZvsgLMM9V
yFBKqJ2L/nwBNA0YK8/dnMS3WB4agVF605GQ8YhE+VRX/LS3dCpTgjkdKaW4YI8A
qPEsBGSa8K3QPPeEevghM2Ui8K6yUH/tl9dcojssutMmhe0wL7WDhtaJZ7qAeM/a
R4ZQHgd9zMAGkfmhER3HoawXOpXx8UvBWLWhX5ljc3BAZL9p2dluDTl9pZ9O+sG4
oneaadvoHyiDigIEM5HqxtWw926ZKGsl6lnHoX2e/y80KXSZOtGalRKKHkDLxT5E
9K/C65VmXJCcXUNzGT4Rhw7ymg9M+F/DdpFpX1gTRs3ggOAN00J/JfjISmYam40O
8IDa7LlmGxH0j/i7dE02YEMCEh1VuYcm9Fx3CjwWiuIqtA8dvHu7Sgh6FZrn2ZNS
2vgohHbohrQTy5MBKxvo8QzKmV0aRCN2q9M3locygQz7qr4XIwlWnO2jzA1/+g8R
cpcPpFFBVcVJ+xF0x4v6ycCdlj0D2j3F23LJBkR/b6PI7JwDS8E1xik27S++n1Rg
pq89YhoaLwww8BSmB3F35gZP1dGRALLUk22bOyN7DRsiv98fb2jFCOVX540QENYX
bVuLZxZVVxz0z5Ji4vIkkRzds6f9fjhQyrZ1IjyBUO3YqZBILoAXIawhLGkrmPIj
VYHbcvK/jrJgakdInV1dGZ18NL7KcIA/z9LedvK6I/umC3YYJpc/7TsvyiP0g5p5
UD3YhOF/IB6W+qk0z0oQoXPdmCCrb24njjQXSosOZbb/zPDJlPO3WebkEFoGxTBa
TDAI9eMmIFWpfXecIaEtfqDjP59gscn+HJgBs8kiaCjg/2XhZr15r0+Neql9eeXC
QV+o7uDzwPLvnvWA/jWxJwLvsn8tTr3ysT8CWatVobUkQfsp+UUN6dLUJg0vGcJv
RYCNZoRhh1kbxVd9clM9YSKKo1fcA9p4ve8yC/+ID+R2zLZmPDaIPdDc9j3ynksY
Wr4SM6hMoldm0Nk4+HsS4g4uA2pfg2kLjW+dGr5Mdag73Vtr/p3expOCyTWp65uO
fgw49GycP7DiDe8AHEMfcsu6XeIcpklDi4iCnHBErxkPzxkduucKqjX3/hJHSzBA
obeNhHzSdRm/YNkCbNGyCckGno4vfTy8oM/weTenmJUK0xOpVwbl0NCivE19Oh68
sUgEHK5kG7KZr/e2khi2+/ZDJsGmhDlAPmGw50K1m39Lcyu6gx15KRrsOLsHFEz+
xeXE22v7UtYgkETq4hIeq9sJVgBVAsbiItJq2AUdQ9p+exwy5x5LhpQ6AOP9Kxzx
PO/3MTP1bwEM0XCXYcOpsDBg5K29C3vL9T6s7PbZCQNqOgFdAmhgOJmTqN1Ha0ur
6iiRwXjXQz+7vzqqZP9U8FgCHFLQTpA2W5WiEIzMDbMRnBLDqqHV29HSGKv/eN6J
D5UBL8334k5HUTHAtTwZ1XM9q+uU91EbA5cUk0+CRauL44YpxqF/YUKcV/e9iT/p
uK/Z9/zPMubYkBX+kB/OIrCC7A6meZJrPt3MQQU3a58YofX6RBu3cpuUsvdGa/iP
dYF4cL97hbJH+p0EG2o5FiNqj3Uy0SxPKp7tQjRUlS51zpouK4tJXRa8wv6aKyCa
taKaCKUEUqfB5VoL1wuAckvndvsXMl22AgdVLftfDlhd1xWtjgK7Zfngw+YFe1yI
FrmZANeRVa27Ml1Hcgy+Q7/ltJEDay2G6jEF9Bv3Ew0c/f8FXQ+vRAvqewI3hD9s
fskQK2oR5jCWrW3CQyd73E5ZbIKgmj9rF2DnBcxzZ/aROF74FzWNkuz41F/cbkU6
q7kZdcWgkEuO7M5VvfZ9CzUn85Hi1wSw0+Y4WJr8FGj4cGmDTdptxPcZjf//Iw0u
yIC5ZD45CQ3cbNNMxhPtcFbiMkTEfwlKwUgXXmFMIG3pWlTyedMki77HLLRyVciE
JkAOHl4iqSCgPspV7DhdM/uzJUFU4d5vlBefGS+mq88vw7QMP2w8C9IsJOC6zzLv
n0IokdRmLNJucgYqgJkmwAt5wD2c+Jn1DfOI5qpT+ibNHK4yYylPvY8LNKFtuG4p
mJ0cpc4eToOtbyb5NvKMoI1vT85LlBU/cq7U2OauuMXXwrXAxhZSBavBdRzBIaHw
f6VLRwhIY3pzw3wNjMt6Cc4BO6kNyQu3t7D+s4RMeZTsMnV1x8iIFlB8h4vDa38H
DMasJ4Cppny8oiemhrfQiM7baOPichyBruHcCyYLRA+bvrbNgW6dSlkexOpOYqk0
7q4v3tBXYy1p8qRpyNPQ+658kqoMqQvsSnjG2hrrT2AC0H5/+MCJXADPpNm9zQcJ
AswQoVGMBMPvQKyUpTwddjM0Ap+tmwWOYmPqVjdR5EhDLDk+K11jExuKStmD3Fr+
r+aJGCWgo23nPf7bSmI822qHapTHMcvOaUz1s14RhRjAr5bXWqQI3Di8oSGbcS8h
Apa7LDDG0mCrL+743wBzoW0VxqT8fF7Xh0JX18Ju4drQ0RI5NoWgQ6Z8M7ieMAZu
9j5tgHeUoBPlg9ji/kq1JMNbYLP/xwm3vLWgzgzGkXaKqnBDqTmZiOs44mjSVmK2
BhWcmv1yynXyO+wn8zhGI8krW04ZM4ODmHn2Ybi/9cqssyktI8KfB/k+cI0uMCQE
ZdWWk6imRpedtf55Yy2mZxcHhHBXdp7hFGa0lx/J6R0iN6Wh4ecB25QGBjTXRjsz
dIvuNtNa+/ZSRMo/nRAfkZRo+JEA0sxBTva4HfiTDDryKmC60Uf8jdWfC5W0KW6N
Q8KlmAJZNvn9KUEATGLvcU/TN74TqKqiaTwmjAvudP03GR2/rEtTPrzIsPuWsoU+
UysBdFqniVdCFeuPDGtwAIYqJcyQJNCHo5t5T5L5PiYlq40VJzkAY41z/s7Lrkk5
XP65lSFqvXVb78oT+v2dHZsw4+VXGO5ovhS1/KZCh2MgyhSw7hXDEmVt1JLZ9o20
Ks7tiiLeoUasENdgCcfDvlGAjU3cezH861BpDfRDo00HYL5o46vCpJ9L9emCL5QZ
w5UJAqb5pMhZv5lVZBMU35ym5sKDHE47QxcUryEpum5m1dx0iAzXT+b7o67KuYRq
AbZLpdVs5zaMZUfnoDhG/aMbva0iu53cMWFA0K+H0WiEmAUqniHGj46Jj7/Ys4R0
zVsGy2pX0C2Y48Y0ukkCNY0A3Kz+oj5bMBkJD+p2J4j0ueRLW/r69tTTi8P3yQok
EyGjjgzCoqMUD0UesEG8qFiZADSnZFaJ6m099/3Nqa99rV2gmjn/o6pccgZETmxx
L3EGjtIMwM+O5TKBZbzFYNis+uOft0mmJtQuXOZQmRJzuHVS26/sG7++7Bsfc3QC
xa555ZmWebNhM6ualxbalgSO0faCjbJuUE/nYHmnnHP7OOtO0JeiEDXnBRXaDUWl
qrl5FSOPZX/jL23R+vUm7TDblOaAw4QwchwHABSfQyvZ+XUKTSJMdQp/rUHb1k7T
v2ebyvOZTHaivqSzTRPmh2NfD14bnUndEvenXMQoBFOZAO7wEWtLARtO+4/J69w/
eKCw4syxef1cpAWyztq30+zYCfgv9ZZ+5uy0mNAb/1+K3PSwx2UBFbbTguBRND81
bVYCmjPRG+dyRoR3Fb51uZOzy+akQZjOFVjh0bz0rs8y0V66zX8kAf9E276nPYb2
dXo+GjqRnnR+sjT0eqfXEvEjjKxqmxWkE9+PWjlDHgG8dXQjKgeN+8lyxInZxCUB
tls4ggEiJp7fRvWIXxQfoSSxGAs9ojMevt6MEhxZEDuMoIZxjtC+aEmukVpp59t+
DxCirEbRXukqPQhbRZzxEj/1fGJPq58x1HnkDomJNDv0EtcBgxCYv3DLHw3wQ3WI
foDA/NReAWoN5oZbd6P2bne8Mff6v6tVPLK9S57TDLfZK+5rMfqSLcZf2pWiFw3y
KqkMLxxD9ax4YBdp+E8C2Qq4TYKzeTwXUgwmHDH9VfkTcj8J7FZMsfJzzBSslaXe
8oNa37cugQYbHG51KW+NxgiKLvWEcBwzIwp1nR1eMSF6SoVbmSqZD12Ed1uele1e
0m04sHfApwzXbS34UMu2MYgYyEphx0cBg8oq5HPIrm7pO5SW8VGs7DlDDaKw9gZ8
iNPICwJqH6Rt9ERNCC+t15/mU8q1tdN8Sh13QU1+Mn1iU4CO6jysDmNTxJnzT1dJ
igDMMSrplmQTysj+8GcuIRdVj/7+6Xzxv+0yfEKZYfl4OzeFcSsHRXFUscPL8f/7
8byQSiiJ24r3n4vXSPVgaqQfb/JOPZqVxLGH3WEOsadeNOvZqrqitz2qVFI9K+iO
Ox7t225vEvuxlHgC0TWxYsR4cfuvuBZ4JfoEdGNL8Onf2OL4ZjMfv9VfpVrLqtXR
XOoAfvTjzU8buTfj94UDV9bgOPuNC2XiNfE7DYkrQIU9GXi77ade7wvFZ7aixAs3
B+8H1DQTh6M3k1FJnwgB2iXzfKshVknuxOUUR96/9e6baVhs4VpZGhE2xoxV9pyg
DZJOyvfNKjFF9hWNIG5QHrt7LwOTzd7IwvjsNbKtDGi73/+VwLBXmDSkxlye7xnJ
SzIrLkI92QTAsvLgn99AfHJC7xMd5wL+6H6rVh4m1miUmytUZ/jon4IZ8F6+5m8W
qC6RGQzuUFObDNFLJXoGKcKHBIihGAirqZNhPjfWlYQ+huKgeCc9qwQV93RmBqUl
Bnv+zWWCpGsKSSfO6HkyNl6cCHCxXdqO3QExToz8wEyEIXLo0VV/iuWKFu/Pyg5R
9Ii+aikRSJ0qGR8vqfnfFHxRu1NKQC1hGUGiIYMFlGduzfiElYa1+KYtOl+M2yu2
R2A9mSFMq0lZPjxSUSca+se97p22MUzPlxnimX3H6yFkyvv9bzc+nrg0+SETj9ht
2cfBsoZpizqwamMt4uyj5s/QNZKZnlujfFBIWY1djVXqt8/UQ7QKATD4lt7te6Fk
tthnh7ooOvRk7b9NCFOy5lIAYqd33fUUrwMk7uyBrxsQ+uNu0scBkx2PjykL3Vpv
J7Fb0cdbP+X+1dWY3M5g0JLQuEWzXox6Uz9SPFvr+cJ2otXTNeFZz+OQakKOa4TS
U8IinkBgHpbHeaUyqt0GEV+qfhZKXoLGW6tcx6vRbILtKhG3VC583lHvBXUB3OjX
eRmtkbNMTvZ/f2KhZzPIzndIPpeI9MGh+9fsYEY0RKK1dePNzSX8Pn/e8Rns7x+S
Rhf8etWB5Fzk/b3MryW/d5cpJyJYMQDTGxt3J1vgZZMxxBpsd2+NPu0k11cs2qId
cGbGOiYAs0Hk+lpSzbgSgq/aNh0uTIC1ePhPq1QDZrPTTRlOaTCZPP8ykr6b/X9I
s6XoZlDXTSPZ2r86XH7fazBC28tuYCgMoPUAsuh5UzaKj2/gT/MXpTTl64UA7jc4
43CBU+GOv8RO8GgJmBHJvxH5jTEvmIG12hLnNeTXsVBGRY5Gmkg1YwC8xvXbsSPD
n8ahyIqV51SPGAi/UDSqe9dn8Er0WGCOKIWxGQHlBqZrbV2tpxuPVa1cvm5RTAAY
YceX5n4FUsnJNkFpuDZpBZ4cct8wbTCsy4gMkCwz2cUGyAP+a4VKXnL/SsuP+CDi
7Ig4ZJeASN/9CXDTqF/HRPgfVFhJ9HaS8Q11ZUAzBKa0TY/ER7rQM1TMesjHEY9e
bJr5sC2npf+b7sXAaPyebVFhh1dTkN8Y8uBLCHytAFau2RZdW9IFiAVcMXJW5P73
7WuTdIPY5JckYgpWceiiBGTRQ9nHJAPDu6ypAJzBQFM566YOTWT6wnhH+BRfyRqR
R0y2Lo0/YRGV1+Sm5zjacQwi0SOMPk473EQrMayMnxN3JV1vNPDVHdobScBjV5WJ
27Qsg801DP155WupzYIwOEK665xKEv7u2Lbl29cfLqUajqISZtY2DB9BsvnAVuoE
a2hPL3iwnd/yxuX72Do2cD9D3as0Oo9QMlfVhSCkgPHgVd6d7NAlwZEtXe14ALAQ
AqRD9rijon3XHR7e8Il/CytkNcteP7lmvOSP8AtBR6bW5Ctqu8cpmknoVdZckEXu
L0nGxsFcavhR634BPmLk9z+nUlSo8/PXtQCRGDGWjcXeXykseExJgV+pcDR5hBOx
/PsZMyBYMVF1eptuqQ/kyJTT46K0xL38R6BHL1aoAUVC4i/XFudeBuKHXq9AeGDC
kKmIwcSB7Olbfry87qGdpFGX61O4V2tR5IYaGDcxV7LVkBIuy8bwcdobXdki7gMM
5WoE1/KnTNPaI5rptgdG2WxVSRGARcn+cj5gPxLCriY9S73B9uI5PCTsZBBU1bcE
Ck49pamzHA1u+A+gJLji9r+rO/IX56mMBMt2MZ5U8P2be2SlVrFwx+YvjdUN7wAm
Qz1sila1o20O537DKufG8bjc8s83NN6IjyYCOqtEHgpInp82tQrOSNf31NbKm1H8
bc1qG1f45miehbz2Dlt5Qd+c7r1XJMi9/uckNHICRO00LuGhN0/OjJofVF9lw3H4
Ftep1g/ZkCKoRKTtmg3WTg+hRU9EXbZd+Ho8RJPhdigderyo84fBGmQ5e2rC1F4N
0o9cArE0GlLDv8GpkLjE1J+8f+53W+/RgVpHcTbYEhuD3RZGChRK6bHHjIMg4Xm+
QpB+7tI9/1H+Je5YiPmEiXHEi+K54oPGJ8h2ksiWx9i65V0BSRcZP4jPeuiTHTpj
hm2VMQUWLfa5GTFhWjN2A6zsH44x0kKPc0uBoAj+nM+UmYfS0fk76veaENrsg0ku
2LWOfm3JJa4Zu+3ButswoMAsZeyE/4NB0B960NLhpt0yqN21drHn35VEpd7goDaB
97ZBDhWZR/AZBw5Ve1rSWjrBOWKK57BupN/AQ+0Ns4+pIPDiTHIo0Z/ZGiuKrf9n
T7slOwt0U8T15t4H/3UFPpw8oK+RBNlOrpT5bN/MwGVAZ2/dTUGSjoNdtxkjsFrz
XKN/vhTfrjrMSyJ/5V8N41qCUJi0pjP0LtjOQzYYzxE0xT6xiv+SmQ4u0y9N5w6n
/ox0rj4Jc7D47+iPBsgaRdYxxbOU8PJAD99SBjVIt/v/XQGHMiXKXsp4WBorelYX
AEfP/3SC9Zs4aKswGwjIN48glgCZGsjUGYa5uSRiu1r9pNA+C7osiQR43E//F5Ss
Rd+v8LQPZICDmyR7EnuTbubjWobAMyS9guYw4/RBURUTIFUCF5+cD7x4JHtV1TRf
HV9HSX9xr7bZ0rWNDse1aQat8ikXiTO/RJ3/pc+udgXqjOtNTyChD0e2TafMHK5P
HTsG2MeaMw+xhIeyrZsG/dC/aouZUXq7NbT18XBFHoQvXwKuGVL81NXiLu6c6bYq
zoggszFE7G7etjPmkREFFev/gLgSbOw9My7jTPcRWiFLgnL4bcgVvLwj6pKXJy8L
AppinMMHg4MFDir/uo8kO4Fyosb3bIg54MtH7f5w6J+TNPI8qWi53BLhTgvbfTNC
sufasreFW91+QGhdW+CLgTjw8rTH+ViDY6feSSmUOu1xG9CcPMGezWKg394/UBSY
KGOOEFNKbS619B762UkjrTF14T3ptuj3sPoz4PptLRkxdFJuBxbQJyZ2pGDPiVQr
T/XV0EKRcTz/UGYcFRA2/sb6qP6Mc0Wr9Iec283ACGlRAfia4QxMUFHvkZewSGJf
QXrLiGAhFYkLa/iloRWCAbSoYihhRDIzpvRP8y1Hvel7BTnvrrUjvAyUstgoEfVg
byKUeXDY2tR5Uwg2NIMGiFHqU30hGTGeblc0suzM+mmkS6fxl3pcXcbwUR+hy2Ng
1Evm4VVUKPyKil2nMohvSS3QVswyJVUDDsd+0UE4OxIM5fRBoa0WQH1wnxjbSSsz
8J2PfiOzq4Jfvz2LRdj5ShQL2YYN3FcYl7WoBQfQ+5FMdhNj1ByTGoalUqHH/58p
WQBPS3TY7ZC057BXZdQl6WuPUK0hdnLARZhbaNQtVhz4vNZfT6w9AX1BrDSezkqz
+3YOu9i612V4tdRSRH4roqtz7gLOwUfBVwgP3Q/J1IoenEJeEQ8sZt66vbmysJ6G
fcXKWD53YiAyQXRUCGBKKpgmMGDr4iCqAAwgIU1v4hnmpB9ABicc0lUMYKTsjTAT
/pIAjmsbEDEkOjmTCF2xQBSr/t/klAFHI7kyxzrGX/EL7Ww8EYGSvT5wWSsenCjT
ChJCRcnAliXhWi0fVDAtOCd8oAS1nDefSdQndtPYUqgaH5Sfn53Z9MeuP0WY+Aue
C+H4lptNdrF6R+GCFLkmpQdArQy/VF9vwmcWSQ/oIkXfLeVnqK6y7ns0b0ieBGHT
QVO2uyRU6QFm1tNYcGKPrQnAhPHGou6eCEJDFSlAFdQ3rReLASK2EeaNVhmWif2P
nlfGQFo1MsDrcWkve+gEVQFgicFz60ifllruCnHAS7QA4/39rQJsxOY8pylpeto1
cOTR0Fb8PJFUX6pm+u6Fonm/6/rUfN2tEXAAVqJjnPeb7nAq1IFUXzXSN0woYaif
qin+IAXU73pzLcLd+H75q+AptLVL/k+IeVhWHbgsOow+M7CyPAo3nv6fDWK35apA
OWmpaUIJDB90gbIYuDoMGFsYM/aJmIqGBkEujf6pJivgLjzqjnMUEgKJx29cozmY
KS3YPh+4SsizW9OSZN3leUnlfS+9DyVVRAoonntLeGz2nzwLtxmUybGnS3AX9JdG
h/y62JONH/XtGZdssaZgfuz/YNjHZWu+RT2axx4wE9C5Yr067r24AnyFHTl/MOS+
MdOlkywkR/bwuXNbQvxUwvqf9KMnwrVkVhvpY5mCXx9Kh/33yk3/ITYJhqjYWohN
uMoFf4Yl7Piol60nbuqOJYzlgu9v/TUSVIThYOgcPJxRkOCTrvH9/bTKkUF5FFDM
QMAeX3mB2f6nlItK2fcHfWE6oZoV88XAS9QTUJJ+3Cxh5C7BdqJRHOHs0vhCXChe
j5t4oh1UuGWnW3uXispHeeyOM342myrTMIaLvmF8vXpKq7+hTIhJiTFfYq9WuZXS
seo4qB9Mt3+hm3UwBAQMzYFipf1Ibkm8C6JRSZCckh1vYhaQSCS8dGHIkL2kWje/
d6MqvICANgUCTNM86NxrlAntqg23d0X3JismkgH44oJe0Qm1mxg3vcIGbP04aTP/
CiR4cUC3+vzQCnNJaH+I0EUuEZ56nxRikZHb0yqYWH7ByuyMS2+fJxS2s0hQtBWk
P0G07h+kQfpdm7zWHnyFeB6YcsoF2ZyzZucI4UNzXfL+vHqPYGMloVGA8EF/OxPt
ikoim5zpZktCiOkh6icQKrFVrhoECbshL3F4XHlAhT4+M1IEarocyOMCWckSFWKA
FTqCJn+DVu2osN9o9NmynrxOKlPASBdGCq8SMsNXuMG1RGyEE1LBtDapP1epCF0b
7UNxBcnYRLTfH/XbsPx680UeR2vh/ZSlBEcThJIfbDPrRcajm+jMv+6vsZur76NN
C6I3O9QnIYWvr2dgQqfHwWCTknjyWo/lyBb+QYTR6xKYxNy4y7KdG5RwegsEGDLg
ghpgBc7WuuTDL8pxwnreQ+6rU5zsvBEzeF/0dYpbDnYOUJzXyrXO6Uzovney4Upw
V6//uj2B15xpuSZwe9QB2xdjb3BvjJgyivV1X57bCTMQ8xf6gUio073HP1hBEJ71
YR0jIWzVwTrAPdfaZ+iMLk/kHbzPqQAqjvi6vQcA1TE/W8a8xwuiI7hVgEG3IWLk
B38hJqa2/c+DIaflj5/ZAqjot0Or36kwgKotLOEozQfkSxdyNx7T6zQ1VPo7nDm7
xUvxaNwq/qS8eMMhvbWQgZB+6kBGVcx7qHAW/TSnrJJLsige1f0NuuZ2MwA9pojI
983A9jFWqL7Mp3holCGGxjZ5NU8ecwh4u3tXtGyEl0heNCq7dc7xc1/rwd7qzF30
8vf37LQnc12LtpBhQJxprRTPoNwliAA6ksMvvpEQX4YQTRPcaT0k4iMkwr+9+zKL
Y9fo+8nWsg7wG2gTlCyNFQiySw+nWdUirSeuRZ7PobMxbZkpYGrTkSs/NZJsjEOi
iO23oq4LB6oPHX3dcsODOtFOi4xNHzJ53JOVEHzVhtTyXE6J21OgM134wTQbyIkk
UDDQl3/fuM9cPBi6BMfKAvs60PEwP+THSw3DQwf18xSYL70P5PUV83HYJhmLT7Vu
cvQWFk3rvfNGUvs4smOFis2BqOcX+MkMmYCAccj8K0MiW/A2QK8hzGCOwfpV1bHj
yFHFvwQOpjO8vl5PFUudThrQYX4OuR+7HfHW00SmhS/J/bxp5JeSC9TKZERlmAar
deaBi9AUZL6436NzxlJs6V0LfIs1q1EjgIOTZLk6W2Xa4zP9JzB2BI02YSa+Hmsy
5XA9pHrNEWZp4p/ojDGrBVb4Gho2RWNI8wtRbhFDMlMv8tmJc1PPTg3OLG+cvNnC
Q2x9CqEbW6Dm3/7E/BR4V/e3vzezjA6O5D78eHsSnp6agKj15BqH9rDhpeNxkKDk
mH+ojiMKz5EuJGA7FvocyDRV6xqhBN+lVyOpc04FVmbY/71IDbIyE463HVTwMNWe
Bbf5c8YZ8Yi+tP7BsRsEgVrOc2jT7+Q/dWdZ1z+m5kqqJU1iup0MIqKLa63KPOMk
vBbVd/coNsQLXr0AX+ZuApZEoD+xNKjZ7Tfps4E1lsnzQH7ijdpH2DS1fLyUsYu9
FVT8AMf9F1zHZSzZfXCaJiaLpcq3Bj5Ch0gw3nVk5oqPoml+uZf4kUO+c1OXjrPY
HKrcCOYtv7JrACS3UODYyKbHD3a94tjcpcPhvH3E3Xcb/wqlfj9a1DZRm4UF1KHX
Bul8pXkALL5ac34V2+Ge+h/R2xEM/R89NFoFZCmtAgWKa9oP7XiD+3PjI4w6J2RU
+PFD4TDUPZ2wxKO6N79DbhqkToGj5H34m7fsOnDonx0nilb6kYRPmxbM+2aH69WP
pOa+Ew0krgUFnvQSNp4U1O/vG1lInGEDx1mInsmbto6oNe3g7PAoF3hFC7KKQDtD
B72ncXQOugz13gVIZISDUoI3357xTypzOLlAukqgIe5vjGPgSuMEzo9PVgMz43kL
a3PjBbgmfBxMMlATH3A/JutpIqHvzsoCh0elw6T01vcCx3xPAkIzKASJ9ZEmC5MK
lCCns1Qb65eMnLjx+U+FN7dN6zVQt2kGx+c1YxiJk5voAg698lsC60rUVqztnOUY
476A6BtFkhbD95iQJKNY6bZv0QPbHl2eJnck1L2Ey/QCet6Wg/2GPideui6mgkGw
rxSzdrgwl1Rb0wtoIiLSBK0Il8F8TNky1Lvez1CjX62c6WKd1aUeeQg/k1xhIMdQ
bTi3BXekMaGvjN/CRwah67fTSZOJoiYAFtXYBcROdNH7SoFlmJXqGLMgtgJ1+fM4
i8qh1HUasfQ6TwoyBF3LCPVjn7yyRpok2AZZhZdoOGL/H0kRngPkR6/A6j0h2ZGp
NNey8fXJh44yO23Vi3oX03glr/RLg8gf4z8S2IkM/PhthgPNZfRKcOE0jvW/bQJV
o0U79AW/KHV5SCjYUPATmB7ZwpKIDLXVQwP6yQ8OsjIRncPdyGP7gdupcWW9I7AL
McXds3GUc7+ZGnOdpbNB3w0BiH5GmdAAlcv84BiuDlTWe6Gtiz20mrxy2z0OLD/C
lHpy9Kray0J9JwlW3tFuKMdcl2eO0znFINgtYudel77j5MrKzO55R9zR/nfsCUsA
4K3f89OJ2aqvfZXnCPaPydwAeergi6GiwKq+9GAX9NUR2moFvtRyUBohClbGE+vP
SSvHG7s7cyIdLgo8JIYD+rShWrYaaWpSFFuTB9SnYfe7AigENgW+8n7YdTTdlFjx
MvBqwZhTloH0VWSVB0WfDcEx8gFKAsSntWv//lVWtbIpzbZePJ54kn7BQKsHUx8q
GgtPtIVLsAgrwHGtCQ19TkEOYJzkAFFR1lxvoSavAEk3XtOeDVTxGMLafS1L0f/o
6rWox6xUKPCgUeUZYtKHSEyMsrYtO/JOm5X5I9RDSPMnUqbqOklw4UfvViTsT8AR
tC1wfCo7Vd5eSUUSAZ5riCNzILSaktHTxiMessSnDq6c8FJeAFVxsqgfl8cIw9Lx
KMFBqSpKGqy75+y9SNMlfItUUKZVnFb6UdIFvxe0nF6HMt+0hhc35qFjDKbkB5Kp
mVe1Wj++FxEAu7Ni3mC2s6gzGe0H+EgYPEtSQtEFDrEjpAa3ECqxCnwGFXFIDQ/+
zguIS8odtYGSuSG6JFNcfbABcWOhhw7WAZ6nHc9N+k81F8THD+6B14JwAr9s8HZ/
x2NRpz2eIb6MaDOM7tcriXq/eBZ/oqdfuI8TyA513hclAXw0NnANg4kFl/ZMeff4
o1M7n4VSqYD3c9ujdw34iKSDK/J0YzQtFhOzy98s5ESGqkWxQjpe64Fiel/HRgq6
J+lS/9dptxg8mClaLd2ybbt6t+NFY1XF98roeGZPb0v/tQK2tnrtiV9G2XkVnqyl
4hs+LrlOVOtvCuWixHk4GVvXKmf5wdjZYaGRVpAq4iU4lsRg6X4VUYRyalwyDQSx
IMAOKMaM1OcpH9NYKnADHeCpR+eP0LsXL8/xeGpMX/j7zieE+fw802CMTqp1J7GA
PzZrQ3YWtWXT3PWdotsSrD2FK0nHpGvCIsas4G7z7zznTcEvyXLswihuQOo8T0EQ
d3YT8C6nhDmjtwNegdNC2R05TQKBGuD5SYUdjC0Fvjbuc5+j6cJGcMB3RqcKGt47
6oeQe7Sxgna7dlXzH8BC3r4lFt2zcBcF2/oVfbIZ13utRJPwug2tnyGQFNihJDdO
gS+mBovpp0usv13ubtzW6h9x7It/cIpFbefqdDuq30jOwGaTKpMrBQMha9BfEpO6
cNxsTUYF5or8BYqymRl/Hn2Bx5chanZPEUCrD9qJx4N+xmUZvMD2f9gT0xx6T49h
K0uI4Wc1GHkW6vaeDnTT/mu7NvIqM+vcpAWPhwFMYjYK9KRPJhD4J/eOQ5/8USi/
Pr+oK1C0W1TjRRG1Wz2gIqrxPkbT632tNkMTumOIs+RF6nZ8qexOdt4P9atVka3l
aDRX/KnFyUrQeKM9qFOOU+iuIHVYPIYDMinTBbp9QKbR6vIlwftHQWjTnqhJW1R4
/VCwVFY9HKg2SfyqrHMQR7UOmnGyyQztFfzId5MOYTTfmzusXe7m0CXmnFc25oHb
sP8sM6eaWzb1OGKvwnAXXKKk2/g/D3WRp7i3sYfi+NfCmnkkCPxBK3eehSHroqLG
RwpLho7g9wSs15Nsu8V3lokwLjdFXjsmhvlJdRWyBR3vCAEdRZWCMBMWjUNxXgCq
BJGJ5HgYqyKtpScYcTYNAftZmWgbokBaLUxdPyDCKzl5dDjjcucDyorVugBZpSHU
m9rY0xoZkHjWzlf5XSezAmr8Qn+FiNzxkXbC+BYUEh3bCeLEcjXdxctvgYvBlFzf
OyitkhFvSoyYaLjRvtsXM6H/c5NktJrxfJI2mRLOmL/64gkWMIbc1P9cBFjqPGqc
Efb3L3dc5BMV3LIEwL9qT98FYZq9IldPyzSmzJ2e29YICODU/x1KDJmKObupt7ur
U4AGKg0oKUN2yWUKxizYf6QaZ1WYvxEvtfhZXXBlO2SN7cZct9sR8HBpFKbigmqJ
IRqFtTMdIgWHjo7XAPwTetor3W2XYM366+ztu0fKU0hcTea3ED+sZ/olstZUFjHv
a89+SNJK8nYcMoKbZSVGhtOZNrJQCdYychwjAoG6/oBtdmV2AaX98bIb9TPSL+rt
xwkzEjiKbpTsFkANq0luMyJu3hlQmbvlqH/bo/S+c1yIpg9NYBOA9547P8mN5E3O
aO5PP93dAL+pDoGBH2KDDzC3vGyxATp0iMrYTDXLA2+SuTU9fSFAOlvqnQPxC6Lh
dts7B4rUVdr7J/kWcWxSZL/CnrFdmGGe3MxmibMgM7vqXv3Gwp147DRLKMwEj7lB
tRN0HQ8bYz8Yvlox0yeNnmP/YqMNU1+pOtdKW0ClTMUwlkCxdve5MOCJ7x3Zs9qg
IIa26lIgW6LNcVIsx+DbF27QV8S282EKdRcm2yFloi0O9eWeuVWSHmhxqHhnL11s
n2ipYsIJrPkHHp8IXO7RHpNrw2V8gH14WHT19mKaso5aOJif1iWAVaa497lJXAZx
zZPkXZq4UO1C0Z5u7AFRQjzSSScFsJ2TVSt1/DV5h1OFAOoc2HXL1tS2i2Gz1n8R
tV+V9tsG8MbGQdyT5DXQtIUElKtBO/PIKIQ4ms30Ct1OFq/uTpwbf1qi+lphCEWA
DQ++YLO91Hd0oKlXn0+Rf/m3tUjr9S2mocAD/ixySGYp7uUiuDFNL66wLhuUuThs
H1shNTOzpmHNltOWHkWcACzFuGiNLu4DBvpTQgbx8y7p01umYxODRmZTsto/g2Se
XvwFQhu8JKUkQEkIOCKxGsp7BJLTXrCu2lxFbBrRs5vYXB7OCuHRdsOyBKkv34C+
hoVEUhEq5C/AgN5Tyv+8ZW+4L0GsyhIrGWE7FQbB8Sup2V8jpPYyFqm2hukTU1ZE
INwdBBOtsmQjGjDBhGsXrX1n8iW1nxTiU2YUYoFdzTKZJLDnMt4Q5z/j9Wxl2BzR
CH/XPEDkBZsOjHRH7IsTptQL5uaC6oZ6f9/JG1lG2CxhQRTv1zyETME/u7NSz82U
fLF41u6Rh8Hpop11RiZjqmxk2c7Amf/oGh6qTixlbVG0i/iLmIXpNu58NlYgq+JK
61qK5aP/xY8oFTA6dTSmUUovqQEH8MZXyGLknxsM9nXImLebrQE4jgMeOLabBR7a
7ztre7MDO66xbTXDKsm23Tl7aJ6QRk33mt56G5S3q9UuRyAyVybHiw1Uft058Ztb
/lP+fBE0k17o7s3NegoOFYoghjWTcpLU/3eoajSPhGwoBzGY5VMr/1j5kWrE1DD2
hZk0qy62ArIh4hDCfhxZXXsMhPx5QC5nEqi2N72KfS8/cnxbrFX143U8PoqMukug
ezZofBF6moy7LBjm7AgUTcEnf7ZdwqZPnmNnQgsx3EGfYoLKZqsjUY8GtwDSKiMG
15auVQaFtKYT5Xabi19xhAR33Pg8Zznr45/ANty1/+Er7jm7ToXD3jZO79RAvEDb
6DipsJOxiFcPoD6eAoJOW6E8SIiSTvpo4rNmwkvUvsPrsffJCp37KUqHWn9YVEzu
raEza3qJgMnWil6U2N/1mJRZln4vNTvtxFMjHH3qhuYKXL54HHETDMyAOn1wm9lw
1kl8LJnwCJ1LFGlHJej1rP3EUoaDFo0estXOTDFDTP9xMmRgirZLYXnCpTLcQwOV
IHoLM0i5KvVVmKErdixtHwt4VhwUCbnEV0UJuuWAEJtc/MA0JYFNhW5V5d1FpXjZ
Sj8AzSconD52ADZ4pLO+Q4AOQ/QcspjwpxbxrnC9YmzJu83h57LpZifwFQEim9i+
+6UtGpkceYO3807fJSxJe+rA5SD2P8+HivYuAEXov6myWBT3iqytKEzcS/0SJjtD
LtMkAUi01T2G/OJjttkJkNJipoCGPzYMSmiqSZ9gv7GxD2Feh5jsN17B+Psp6qXK
V6eKqrGC5/uuq4FzR7otQVV+PBqWE4Mr2R5w6oKIZn9q6KOjAMAuZSil/ajPglxI
q67UPjL0+z7w+oFZxPwM3dYuA2g0YWbjAtgNjLZQLHDNdi6Sk+62oIqkBgsshwru
TYYy71MTetxMV+ogRy2ZSbFyq7UydGmdOKGMY4QxpZloQqYZeDgwjwn6Wz+rAg8a
rQ6uqdNRtd9xdEKR0rPCxedEnCsWWXGPNK7GL5y3kSTJ5vcd47EHWtwum0ui7wGW
1NhSdgRcdP4EqfpFu2N9MOQRn3t1Nijk/V+EeSgJWYEM+ejShWZdVEqR4U48EmL6
4PSvc+rdMuT1v3E3K/DZR3yT2JTDvnJ1SvmKqzg5Ya1upwzCa2SXC2CuYK0Qfm/j
er1tld0Jg03kYWaOh/UFL8E53yqi9+l5W/XJL69prEgi5x30uvcreZYYgBF4jWP+
RgIjuGLTMHu1uijeKV8VeRJ4X4MlgaZVklVCQ5QpQBYgaWQ/LSN0ecil51MMjNsg
c5xi5EInAg5rWqO0xID/Hm7Z76HzzuY4jlwvwY3tjFcvPp8daikRxnfp6cnQwxQj
y5Y3CaW8PH6a4ijjpsjFAgOTmdGuAkdFiGTYgMp5/mFfPOMPuTSHwCdH2JRy26GA
KZ4cE0huY2UF40GGrWFpfkdsC1EFMG/QBE/2xdj7pDMVb3WZWUOOxqc6jCrP9Zs8
JLaBmVz9/E9azZ/SN7taWtLYJr/hHa7ki+jLBUKbtfHVgShMym2kD5fFRKJverej
Mo9g1E5XhpwXeaAl94HyGbDaUck6KLEKqPyRlOTZnJmzd0pnzd7L3RIWKLXSFYSJ
6p+KVI6dv9mF3aItkfB3Y+1FN16B4k0uC3GLiDIKIJQQgE9agXeXZfaoMZKMIJi/
ua9q5bMKvWAo0bpLyRrTpohs1YgrMBzEOLwnkWKGKXOaovvsQeFgi2JgSkc9Jjo0
/UB5NTBgub6Cpt3o7F1BVP/WsyjFTRZgzmUQkjsquYSF8Gk218FCro+na26UdVW2
7wdMlFxsviYA5kpRFpn/y/Z3/YvbFou7ACoAFOYCYzGJkVMdiqf/6etsck6HaHoj
r5DuIMEchwi6iNHmC7oqu2WTbvCMGHV8EwIm1ntrD1fhrXVR198jyW1VWXUgFWiE
RDxtcjE7ehkJCG8nnpGAArlrWKM5hS0RCPD4N7hnbYeAxt+Rrf/4d2HMYgUdBpnE
PSjOgEZiLPKabWCylNKCma2YehARAihVlp8yUKlUWQ6ZtreD7yE1GSNBAKFuDzLP
fJxIkCguoQf5Ml5sDSnm4RwzMKAdhrdEXioDKTI4Nt9JxHiZr2Ev3demyDHoo0dP
CB1pv8Wt7TdIdTB87QuMFPrJLUZgz7rRPJH542P4K3KGCI4X4yCqvWyi02O2Z4sl
WnT/dMz53L2+Y1F0E/GPCYWpVR2WvgGGSrmTHjJf5hOSybFjlGImVtOCstlHfqrQ
dwwqX6QCaEBMuUxJb7StF+VrTAr7/ptDp878aBBNZbKLPk03GPt7MH3IkvZrX3UT
dIcHW4undJeXHAsXCmtDVbVMpVcYpRECsWBXhplmIA56qM6ZYrcJNe++BNuo7/nT
aMivds9eUCi8fP9mwR3/wEWBafn2ujmmZx/HEPnmc1m98UaIFZcd04rOaR77zyIl
7E2o/SWarlgJC3slrqYtOFL+jRGk3/hlBeMNyafMBwETeRohLrAqwKW3aRuJXEV+
3yEVyJW3WMqLn8xyXGDJ1l9D13XzD+BH5NsF9Q7pcKLHIRCpIRROQKPgMALz2rUq
cAtuAZ+hLU5AEFmm+vt7eevBnywJhogpMWWX1Xiiow/LNIpn3SNK1qwIH7t/LUfi
lEWkMTuyycfSLd4L3b7RdvWvCJOiVhRLLELxagn69dIdkd8XahEe/S2UJcWSfz78
/mqZIFos/m53/3AR+mBe8Hz+7Al5OPTUD9k4TnOIF5b+6/jv4w/zCSpquE3hWOiB
NzVvAemeJ9gDWYXZ8xgS7TDojqPlD5YbOVeZkVSQbGoCbg0SEVeohju2nJh7pKoV
nlkdyFiv52S3VA31SSg90ks/zfyQdJdJf/Jhz8hxx+lpd1bKa2kU/X/izn3jAnI3
r5HfJEU0AR2GjlWvAixvq7bCG/xnPhEbFsYP2kYpqKJJ+DSiTDtcf1qnFFG0I6au
xf0WGbNo1K+3K66AeyuRQHYi7u+U3yD1xBp2ANUPzHTRTaLKoPw0alUcrJrpsLEK
MbFW3vCPLSJny0HNjvblYezPZ4k3uk16X9w9xskF8DL0Li+xQaO2iVH43I8i/avM
hcaHwdHf6UcUqrTWKnvPpvyOCemEeEX/VCnPdwDQkVtPsldSo349fcwUwGUldLGz
6ITp/7L/qnBbAAtC3QB7TW/bgv2nMiOoGN3xyLNI8kp/4KlxvyS+qNki2teqAlXb
wvk8IUE4cdmcDoRPvnFg3NakwGCHjOw6bLFJJIFiSMMJlxRwVPB5Z/+GfnbcrNJu
Q6fhPM1TMNtYgFS2K2et039z3mxRktGA3+YfnVweoku1CszRgPzY+qy3yHLITosF
MYd0XgDJMy/5bh5vobh803pIT5l1iNfDEaY6RmPmp7fY91/yj6/oLkROIlbfY5vJ
l6N7O+MiFAzi7NoOl7eYhgd2FL2EXw4wtozRPLI8x2cQXa7b1zbEK2QI9NnzIBRu
0LtfLPDV4eGr2/SrBnJ4Tf/KJqfJsbmSWhNXXIlEzJ5iGgDRN4cKjktWrhF5pasz
WyTu3dzhg/NSS4apHxjGhGjWn2gOCUrvwKt0IkFvApy+z/DePVmItWaO9icr92r9
XKHD741saIVcfwzPmG9OBMRmpTPM/Hb9uYes9oHGg9eC26FjljABHZpHc9QbNgIt
07WGyMY2ZlRdy6dah18YGUPJB1cB8zkG3VGibvvuXyQSEUJcLGxVklmQYUtTKGZO
atrn/xcsArASqAPiFcSsThBMAsjiHWrXpVoatzi04iOsTS+k6i9j86xRtht5Yi4H
HrAFL4uhimDBLbh2dYGLn0EXXEelCKu8vaQInutIADzhHfogY4RGGNx9jt6xHv+W
9DOXtYTr2kCUw+UAsbjrr0UVsrii+BDG7BOD2ZMT/bMys0Nm4t0HJu1cG3rX6+Xj
RFRUM8WsrT6qmeUZ1ELa0rWlROWfKRDEQsaog96u0nhK2z+OLABS5IWZ+96izr47
XvGTvAIesS0m35tH4vMMwDft5TSjV04AzPIRJzjcfXfQX/9RbY4Sybqc91hBR24P
TRe3Cu15atc28z66OuFX7Lekgnwa/ucDBpd9kFUVW13FVBVPHmtfjgKOCPSEjlQC
U6gi376f2J1oDlJ3M5RXNqKKmnFiYsS4OwBK48sOqymPBHrwqcX+RheSMS4VCXut
BP3r3sJcFd3EzNISw+Qba2Vos7GJZIy5CcKgrnHxp6bsZ4OlKZ3RouxuOzFahSfF
kc1D8wecLQXkziVO/SlXw8dJZkboyhJMH4Ey4fEa9Fw=
`pragma protect end_protected

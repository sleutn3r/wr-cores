// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
AtfO5F9gz5rqKQ7iOinM79w3sDT2OQ+qzXX4g0WjPNFqOAx/cXMxfS2fKachwwe+
/N1GxLcIMLs4QMTIn44GmW4+jnMMcDlbKnqP2nLtdfHwOMt4HIdpAMdfhalPu/i8
uHy22czykxV86TXIZX/2YlYRXTwioKtS0PJCsW3A4Eg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7984)
LUqsmJGuD8ocCd0AvBtp3+nCe1IpnxGJRRtiHcsjftbizVpC3OdTfFXEeig3Sqo5
sNA9u603P03bh+waOhP/DcGn2RPRobUd5yznONFkuB9gy8QZ8YvkWxjNIeVo34vD
AYzOnm+QA22uYUSW45hQXUZuoORY2pVYBPSZ/9K8a7Jbi9qLJUlTeoDaCfgSThm5
1RbkT0OzLoMGa6jlrD18ERtW2TcZ3w2XZDFkv0BA507zfICbHgtMZra6FZIurB/N
Qp8ZObccbw+in0i9M4Nw1NMLTpCV4dZmiZZW4QHp/xA4haU5sNfwIqazZqT4sNzR
b367X/tqHjPjOHLmaPgQ8884uUL9bzlh9e/i0Xz+YqKFvcAOAApqGRP1OfNR54gZ
48Zs5qkQURRl7RoEv2vUxxZ8f24lK7rpiHopMPVn+x5oIlgVCDgQ1SbRL8ZyDgna
/MfInQPG4YYqErNXAQI6T+9QjOcAeyF6LhPQmm/VRZ3Ql4KTS0KQLcdG77HZ4fh5
BAETaXP0BFX9AUa3Is4s/suRwJnesIQtHW7g4w7Jy9fWrT6Bqafqx6FTFpFSolD5
zJAVv8EmT9XOI5czcWV4Bs1hFcIYvsxni7pH/N4XniZ3UV/+4OZd9E3aeJAQ7RaB
24dJVcAO2frOenKBmDBCtwy4Zg/SpqnPmoPxj3+C3Vt+jKQqxuLK6ShBl/ARI26S
4JL+RWKjR1PKJ/VG8ROgd7DAPT/KHsZWoLUYWqd8z711/skdnit7CgiCnLY+8QG7
B3MYN5zx2pScDVnFH9/8zmghMsIKB9sU/fxlPeKmRIh0dHv7vIwRcDORKdYJhY9E
lS8JlLZ4gCXBVrEcM6W9MzUA0LWk35hEqgskYqbBjxa+s9oAymB/sWFNLqN+4gQf
vYjL3Vq+Kkh3pz7FK0yUv0+8iTNJLDdEZbHyUzJKJMRvKGeA7JFD2KB+SlAwitJx
bTeRp4c+2IRiz36U+/5+m9v8mWuJ7bRAk5IW32jjJM4vDy2Kk8fEzQe2jiw/W7zE
ksWq+JJbtjr/CaMUnU5CsrAr4BkOwnVrVFIeOKXAXVoYhPWYkzozGhTxDdho3CZ5
EVHRDzzM3fLMMBPbMkr8iPUzSV6krVNduw8968leNGuY9TFx9ckfURJ8sM/R1Hny
/GWWJ4QE2TUbxBQu9uAofLLjQxoO4vZplXlBg98EMsgxMABUp0MKAhDhUwtxuSbP
IJbtBAgOcp5eoh5e1GV3ym55b2GPGYlOVb9iSqvJCdXdi7bxmkUNsyuRLaGxnqTe
rcUEQxEGxf2hnLuW7yDgXnaiBLlGeVRwD4Ww78xlMQmZywpXECRiKe0yV/PGwd/f
Gymwu0FuGQjh9ztKqnTw4rY0mL4eNX/AjlUy3K9x+N7Qoj+jpiEQSOyE3kz9dhRM
Wl/3WSVWVc1fCBzkxcPETufuFb8f6k5jvXcMOm2hn6jipC8PkjxPKYvwKYcOMWC3
5szzZ1Cj7s5gkMs33G6L12uYut9qI7TtZ1/wAIFa7uzbrJA/JKx5Ai5WSBjz/OcB
1ULS5ptRhjyo66Qf6kN+IyHPlWrSjFnQFXc4nulHfU2aAKTIXd5qXpronxuACJRd
au0n0pIdd1RW004ehVTW+Nx0y46l4J7TuWtEzGLP9HK2TcVfWt6rQk75htT4rXIP
urqOIc8tgMLJ2mV7A3/UUpRh+BMLQKftJHUgAPPbt5eOi71QARc444c+0IpKWvVK
ox3/oRmqnfwTSDREJ+NlnGCmkmwnkxYVvsmhT9kLbY/KSv+QBBYoqQJ0I6jlqjlA
2sVxwPPXXWpI+2IQKyprECAkfYesQ0mo5AsR+WqWafmnI5/pwreuQzAAgOSVUYGt
eZ+z/XcNpCr78q1e8o7ScNmJA/Al7oLrM6qvJxnukfVMIyA60CpbmwA438JKOHCA
F+uuCKLeD+j/8j45M6DgNpQZuGYYLW+f2kFthlR2dHeqohSFM4MdrbghHwYIQYeC
YTeHQg5HfL09SwFf8gANLz4uydD1Wt/wuRchMKZ0p0m/MTTzmn6iuNfrX8/MrEeH
7FPBWVTe2ICTQ2N0JEeQQSCvTl7YaB0i3KHeviHE7mJn3mZT8OlJME4z6gxQJjzH
hd8Cjtol1w6QK4B24eeeR/Comm5HhfsFMzD2jfG73eNh9kr0z3lH2O7Ufxmr3Tdq
9Yc2/hNF2/Xq1/WP/EVdDz3QpEGpaxKsPiVez26EYAXiTEjThzTr4cp0vJLDo8zL
OR2jy1NH0o/6pV17OjB8A6Wi3K6AazClQqsorjmVobYXh9as/OSalWLp2Z3OK5uJ
ECsODuAxaIZfVpTKmz9gPVRw/7ajFVGSAgvSdQN5Dt4jMOmVnUmyKTE/orXGtHQ1
RuZKERJseoVYCXD3WpTrUIWluRjwN+D49JSbwSZ4WxkF1p3RrfzGklMB7jDaMmDM
Tqm7AgAEyv8bwf+TT0S9EH6geoWyHAS38MKCbI6k7ooJmRBzmcAmYcCDdG2gW8hN
i2YIwodAbq+pXV0aY4HmonyPGhHzTgB0YlckCv7zFkw5JMaqux9h20e3vO8PDrPu
VwgG1zyueie4JRfXj+0mDcRSYfk9eaT5XToYAXRskYnx28pOkKXSANrPiD2dI8FT
sheAGYIZTXM8UA48VE7PFsmMiFsav7g1DE8AN1b6TLuP2TPRwmmAMqvYqviQUUlD
xZwOMKOFjjbY67C52dVFY05Vjo0JdT3vKcEpoRkE80QYwiVHV8mMlgWPe10X3Kns
dMIxLuzcJPlL/OrI4NMEtVTx6TgwyceA1+Zg/Ujzr6mScCiRxi7p2ZOolBF258J4
sTxuEkIrf2OGW/6ULRtjOe3BETgkySF/IeDJq/8YSyJrxRqmS9ihYSn3XxQJpMCW
tXMeuSjbTFt5FUGJX9wvZy+PEcv08jirbUPj0QTP7LzTtXqxmHeIP0UrjGqwWoDj
qu/MUonjP/E9dx+t260YkjoRBUufsILoqlFrkX2F68yQyFehmIaraZfJT6LGPcEb
povc9zFZSClixCnMa6shQEhQsWcFHn/U3/3GynwdAutrMBOMQXVqwIYaOAm8rnOX
T4+2yQZXr4DPvKFfYhQb65/XmdLZrXHKGKfKLJJyBsKee2H/rbb717RwjSrqfHSm
/u9HOEnWcwHF3TMNOQ94e+St9XBSCPQan5c6sDdvm7I4sVLb1YQ6Qfp+UTdxQrMQ
Dtj0WhVO42TevTuMAZ4znRqURWUAMm1DlVA4p9iffAwpML12o0V/gWX2DVBv24Hk
mgsi2JWh/mi+vsSXE7h7zfS1HYykMawOVcuImAg+DtAtnuawATFn+C7XNvsUnhus
Wg4aQdCyJydQNOvzpPmCCOgxsl8iC3rnOr/gXgDhViCgrVP5VG5/poxviJv4p298
XSdtmi1IseWMAqVobaa5TcItiFDL8aCevk77Aav9EHl+kGzruvVGcGTkf0jixBjk
tx5UmOr4VbM/TSh+Do+ztCNAtjREqE8ggAUCiTUmS7PSSlFv6u9CQZo8gKKFmbxy
FRsTq6A6KHPZxaNqcwoFWLWj+a7LwcNBTcul6BJWZV3S9rmRQf0Uj4E7Uqc2ha9Y
1v8O9Y9ITQBSYHC3eQJiPgaxE44Pe24NPEHb2W7+bb1dSA08wgpSh4UausHyEBFZ
OB0r3/uO3Vb8ql5ozXlXxgfLvt9+1I+tTB/zcComW++R5rl2JbQzB2qzY5fj1jQ2
muwzZvX6kiZO8rTfzhP+tf73zpCakEiI+Fyi4+GRt1dVuA0YYAvTm02t867WSalz
SNGCYFIhSy44RJ4erHJQYwJa0PiNeShwj+k5tDoPGrcyoSfwG1FSDqTbwfPqPfVz
Zb40FXtrrCZXyRM9EMpPvIImj6Uk2nT8gKxo13YIYuOiG1uwi1glwbAW/ZliwJYb
27GKOUuLM+6v6gXxMcA6g6RVP4GgPtUNG+dX8bwIq9i/C6MGiakgwpmzUvTw0g8l
pt9lZCRzupvDdnQvM5f9FdJTIkdabPZQov6t4B7M80zjK9QJCcTKEKl+ut5KLxTf
T7dzvjw6/f8IrZrorXOAH2V/0sE3Ja4U1HE2fCA0uLi/uGiuU4xxL6U9m2W3yJN7
90OztEoRFb5UOHLVEHlKYTf1Co46VAREWlaHcKh8ngO/VPdU9fqujUs7vGFpQkUp
a9iGO0IDgIBMRaErCLND/6jA9EGgDt7cEYR5A8KhxdSMkvjn/St4T5o/Q9QU+1tr
DfgyclKS9YPk0IiUGnUuXr+bWt9C+Z773DnhTzGqpGVVQoz5KDsgJ4J9SIlAl4dy
u1OcdIlb3FL+z/IeIsCN6igg8dBMNd6SXvjMiwsY10Ri3jN0z+GAqhcvX50UvXQp
tl0lD90HCGEdWg2dXSoptRS4QZDn1MmeKjoYsESEnimoINe3PSTnJNQZoC7k7Ifz
lBWKOllvVf4jYruZBH5zwZc85RukIVAOyUkgxRlf0b9z+3Ul0RGEyw8mNRP4G1bV
y9dGylIFDn/yGmA2DJqNTuInj37GoW9SzoGIYIuoDs2xDD2/gu4IsKaSWEoeS3/S
V1AuBTsg0NtJrXNfXjOVfAQZ0MJuxo9fecCpiOm7zqIoQsbO983rZGzIYGvFFkom
hVcV+vGcuPjf3m5s2bhwZ5OXW8qs0+1ggOqS1yGm+cZLTs7eSK9eDpw36JgRvvYv
TiDFJfaYUpqR20flBMwhxa6cwriRJX4igCbcBylECVamqYM8r83K2YfP6JzuDWg/
1kXeETh5Xdwf7Iim+yi/UImw/tnTg4zsfwwYQLGfR4FPqhCdMU2fG3XCqCjiVE3L
MH6g1swd/8RDG3qi9Ku2l/fcq8ABp7T6cRxiyHJ6jCF1C6YzmMLpEVb/1+BGLn50
3Imtoo8wexQLs0J0f844NIp9DRnDS6ZQgWEwv5uGitbAwqHsTqGSW66iLJb+smVI
xx+K+DLgtFJDVRiQ5D6zCxECQCxAEbzY7V8G+idOL+Z9CWclSoSIZZfVcA2pwd0d
d3l6mqvuciH2Lu6h+zopvPI94uWa3AQRg+cZceOalfrowOSLiPx3OYXfcV/QIuzl
8tfvCp2MxAQIkhuqAGCW04+CcCQBj+XrdvATjXsQeNs0TV9vqXaSuWYwPVhBiI7p
zUdpXz2mlpLCOMhPkbe1dU9yb0L67eEC0Eg5DcnGsEDy6Fgq4FackbA0AWDOuth2
D6tqfacED26W1QHxeGNhojPi+VL7AvPKefsKLpk//QP6zdcltSIduKKD518Ctkqo
KnwBc5ENL1wkfZlAo0pDXWF+nDFG2Rrwrv8TvDsc+GyqDp117axnovvHhTflShC3
x9UpehuiDevi/zNZq5RUA7rHsPTyTEkyrFVC/P+RKcXQOS3eUPhEv+Y0rdKSl579
EmIMV7buOxG9EtSS6ffbTQPki3JcdFgRqyJhoKFdVXWyat8rmur9/XsQq5u/WtJR
bhsKeJNZlsp4P3qJ1BcDyuQSIXLyWd71ab6s3EFp9VAIcNAqUkffHw9gz0rSpQdy
82ZiwB4wDVaszNiRvZ9jk9anJXHJhxmmUQ9NzsnqOVNzUKTZ87hNzsixsqjIPxSj
zRtri8QQ1ujFLaKxX9P5bg7A/aFle8ddsWfFNkqQnNaKqvxj+HoI58IoUr9mhknn
w2gN1DUioLwiiMo/LZzhUiCDCqdcXElB9V1W10Zrk9Em8E+F0Slhfo5S0nXgso/U
9D8DRDYljeX1rMVqBIEqLFQvtM0Wojrt7Ip25/IUAGwgrWy0A187WIYnCUGodOQj
gaa3LfzIeihCABzCoCJW4tTiHNtNfHE5jzdF0/HCrusR6ovjD70GcggWF8VMnOQz
T6GBX58kMUUyRHFVWWwFGLY/e9bZ8G56ndU6el4plUX7u7IneTZbaRWAiQpryqdo
P0gKijkJy8THiq4dpLSDo3Nd2g9iiMwWkhCmCW0oyGhUKH4gnDxNHv8ZXgcc9fvR
ZOyUG7DbKRpG+B5xINcJGgM/nTM7tDnFOlAuUAs3hjOWnAb/16LjJ1g0+f7eBvwJ
scWDNLeCY/lqAPpu+QZ65tUXc/geBVXRI++RLTTMiug5uJ9wPUWCDBqwF/w3BWv6
9zbDoIC5Vy8AxMlOtflqtkg5cJbx2VRRBZW+6CNkXT0kXzLQWYrSjEmQv1j3cQjU
0eErfkM69PtvEKiB7ssvU3z7Is7qgwjputhUFtDeHQK3dqii/qSo55HtA0XYAMXZ
rczMh8gpTk4Ox6RZk6zK0xggOSBs4m1SWdfins4vG6jpnj2IdOI6Ur5AzrcmJ0ne
MK3t8TyS9c7yGz0Y44Plekvfe4pdO17Ir/mkh8YRLfy3SDWXE5NpkyHaPpvSYoPb
iwqn+QbPXuR7Mb9GJmpum0qRjsmWOF49xuyX4cHXmVz/dmFFiUpuGlXFd3gAuAxp
v76pLPQALOIcjfaabofW4jLX6vw7H/h42gBbabyXSfToWPtVj+ogZJX9E9HbDxUi
TT1dy/HgBpnJnvibBT8Qa130nPinc3fk/4FRPFdxH8nCu7KEXA/UVuCAzsFzXgKI
L9ljF40nRBM+RRZbS8X4LqHADG+M9MxsMnTzFHBT4HsLJ2keuYX5HiPsvjEwi8a9
7zJtbVR40PdP/qaPOE8KkBnH2O9Ypv9raAK0PgxakUX/C1GpkG6PS7/iBkvSAlKP
/cu6APyDE6SaoKiYT/CHI6aPOkd0ICLvco965Wtf4xcxsk1gsWqzKvS2hVO43FtP
SXj+0tqdN1AShypY9E19F8pul8GJ+wCMGTc20lmwaN7IjDVhRrlPrk5GijgvXKOL
pXCe/bs/eyaSJog492hZ8NZ5u/yZDI0zIGxV5HuUInxL9wdmZ8kfaMfuIznz2EU7
KjpS1ZO7j/hQoyttCmLBZ9DooM+1kVHbe44aBQMdAoyZgKtvWQTStGELEP00ktO2
GA9BZLFtc2Wf0qdv2FLY64j7fLbo61v3W124JGYG4ZGSgbqwhejvcpCaRVsnmdyn
A1R+NpsnbcUFuU5SfFl/0HBUmoNA8oGQ72dFjMMOrSzuT6FOnh+66tJe1fXkINlO
/E4pLUq4b3kptXAxxL5sWB9SATD93Uyunz0slGL+oZv5cnqSrdsAAbj44dLCrZGy
kAJGOa4cy9x6l9y2UPJfs1jlfZ3FGFfEK7KpSKH4m50jKFQ+/iYkXFghPtSXMTKx
XXv6ds7tfKguvsLzgRJoNcRfoTSxxaEnbSxS1A1WOn30jhRZu/oN4kZh6HAfSjbu
m9FJiDQNmjvTEo17n3YWvYJs4z9VEwrx36dvzDEZG5e8v095FEjTsZ1hycLgbaBo
yg1yP0Yl4E+5aWKB6Qs5AD1CTZGR4VWhV4Uj7d9QW7M4MTFp71ISH8cJnqR8BrgN
pPnH1Z0yGy70q5lgQDUJE08BvI7M8NqSP+6Sx/OQqJKv5VwrTizSzYeMgyvl+y6f
28MBD9p/x53yJ7w0rmASmSXXVlftDPmsC9QLcwNVEkE0rIsiknZqoDaToFwU1rDN
OiZn7G75A+1Kr/HqAL2k2KUjG4zYFW1ip76+oUWaDJ7Zs4pjuWz/Wz0VevR1OnX3
bp3+ubUDeXt3FGj48EfJKdoZQkRSrz4ACOopy5YNn1DiiYHTyO0s7ZhFJwzMI5Di
SY3YoSoes+IO/emOqSlZJHRXWe1R4LIwdyK8H5UIrbV7edhmumzusbqwOtfO3EUz
Qbi3VzID1tiVzoPi9hTzW24iho/Mz1BfSxo9bINIMa3B+4t0lsp5jzuFU/UCtPh9
WLLCshS2vAE9txJmLsin3XfreKEr0jSjw5/4RslzvThFNEuqqlhLVvrg/tm58mzb
THFeCTVOjN/TUQJTu5YShH6PUIUwOUHX/C7ktDb+dmSDRCQsFwYVR28igCCqPIzb
JmGGHjeMQt1o6UAYHmSwrvQ+p0mR2lZK+0N7kgqN6+6RcY46hcTzKSZdbSPV6dDs
HsjzXPWt+bAc5YsLhcVfZaf7mHxRDhvLZtnq7JgUYR5kXYT0ef/Du55ipS1/X+AH
Uz1FqOKpEIokhwitYK7kxOGQNkR6z7RZdixm65qT2JG7GsrsmG5qaKuCuj4a2S9I
3KRVsCJ67PnHSLuKx8CxCuoxcqbZki8Cq337v5Oj/vTKLXBXjR6da9GehkCNOsEM
orFks+IqtoT/10M8oGIHh8cWfbxn5ypNcY23P/YIjXG7jwD5AdYoxTNTsqGRwRHj
8Q7DZh5i6ifrrtKWnmKbdAqFeRTKz6Sbse8zYMNhoU1LzWrYbCgpq5iFBpJKrk0m
tt2ChxniuiKpluOMSVp8VYmshMgDl+KlHiQw3B0Wr56ru0CvVAl0I0RH9wQOiX2i
CR3Zog86rZjuZta8XfvWBKheY1VmeX4czQzS59sxF2oJPNEKT0JDx+7v4JxX1N1h
//dkf/c0mXvTTER8PjTQXeVb0d4iQ/EtWKkDwzMTW62Hh6IHlfDBC3U7HupsXQGy
G3fBD82i+nlxqKOQWL8JqTebKnVHzMioAB+1p6+vWoYJrZ4GoQGB37m86h4bQbO5
ToCmsw6Q5ID5HSgfbi5oPb9ElgBRFnQPyVg11HuYb+s4RX6KZTsdYp+ElJuV+Hq2
ClUub9ZdwzW18OmLghNQ9zz2JPATqfQo15qnEY0Wf90b5KWz3zJcnbrH9Mgmfc12
gg9AoQReb67Jk+gqAp7dLqORIPoQ7KzGmzHeKXiHk3c0mJ1kugegl84xCiMKVBGh
BfgUOgmo4/GJmdxsuuvShqMIwaVZ+Mj9BU8e3BczZJ/7u6Hr0eSQhiTpeBYi6EPG
xR2IJJbP7fjCunax7x1iEFejh2va1ffGi33rF1/6VguifQQ8abbG24oNl2HPVh3e
kqB4gsI2mUlLnFRuXAESZtDEQyvU4k05KzNCDdItYGt3TcXubG/4bAsAE6GGSnu6
Qfy4KO3yN0MdjS0EmpDqvayFwuOnDjjjBC9U2s2TBGEjw6nHTohHYUEMmM0Yrm1C
mIGSEgbesBMq2wVYRYiUYmdE086Ppoa6P65RQ4nIukTzzrM/DBK4Bj2WOd0rFtan
58ytH/1SZ+c1xjlbGk5jvSm5Csdm/73/nwGPjimJh1GiLf8x5Sq4Pjpp9a2nPFVY
gP9ov2w9XYOVNNOlr5i2c/qd9977LrfpSBseiDd+u/xcHNNxjSD55fbCOm/bIY0/
n9dLtD6v/qwHuC8HjTE5KakLxikUYoKJwj9hxxw0aw2mYBGxGrMCZjv1mpCbPkJU
09LZAGtY8srjaeqhyV1jE21IUGvAZxyb2WiuVpZfGW7YJZxebZDAcD5J4rCEkwae
FfW76AzkJPE+2rx6cpIA//EAcGzvC5rRISB754Gvb+25mhcoFnpYKV9s3mHe1mRn
0q9PjHHT5u38Gb1s1m4sKlzXyrBhbux67hR0h+ZTGtWVMTnivSjy0fOKh2igULVE
Q70GlcqvasmcyDZGVb3u18epyh1M9nqLUyTfizBgYQ3Y4TwvJf4D/MrIyk4rbFDp
dKTVdBpk16ooO213DGzPL5xshCtL2LsuUNPcAmYjDnpihh0EHIg/7u+tfSJj1mga
W84N/MRvmaYr9FBZT5Fh0pj2maFJKHUk7aJxPqap9tNW+sZJ58+SUoqDwYpEub4V
gXJbmEMxpi8fD/eill/eIAOShfX6ueiJADpV/j6u3YxEsAERbQjO6r+30WipELE+
lANQ5qlVnpEI+Bii6oJsoX03Oe/Ijd3pFFZWCn7j31Ky0bAfx/Mom9Vv48Ts8cTG
0jZbHb1G1mYTd9sE2HQuAY09Vlu3rB+Fyo5m/Ip2UW6HFpFlI8FpbfYrTeU3Olcs
LnwKHhPfFwsoXXp5feXVKMZnNCxwhh+DVAVaQ0E98tyiXDMUQhJTM3e8xoxlXb/A
xRuVGE9zCgMiwE8kQ7D51NrsPhDiY+onB3XO5piJtE3NO4OT1NAwZVaf0uu5rXm6
fZs5HgilPlKECnPaDcyFSGuZ++VO2bw+OvYs3wKwG71VQRc+NGHPPnT2og1Cf/uj
4x2R0Xj4f8gXN4t4HrJk+JYX0P3Aqu7fsIc158GZgm2uLFynGDhl7iwQae7K1Nvi
iwwZTbinjayU1ykL/F7aSfU4fhI531mLKzb7Sonq4/Z6gsYDEsLFSfXPgPLM5NsI
6OFjNCoXdopiA8YlNnxXWHkO5jOhAJSv4FQuoYcbpRhGNHbCF302xXES8GN0ra0T
HpKNvgD/3w5TO31j3BQp1coUZ9SGfmuM+oWNiRfCBsVtnmwUJhr7Q1rSkFpDZDkl
jP2IhDFCaRl8UctPfVRM1mGz2vWoH4FZzE8nPpgPPGKzUn3+zCoSKZhn/1qGBOJz
4uIZem9hxmsWJCEJ3ao2vmXJ7B7IjFD6EqHGst4XEtvOExW4hS21ARhLWUWVDPwh
PtxOxH+0wGUlwYv4hcDh8p2ECkRhod+RY0X9Ca199dQHu6ouj53NQObTw3qiug8h
xSfPP4wMoBA12EVF81vWGj/pQ5jdlk18JM13KxP+ek7Cieg2jkKznVboGs2rwVKZ
wXaow6x+vyJV5vi9fcrT2qSV9i9Zy5ShfJZxKJMJ8cEluTpUOQpyZ62dkUWc5rR2
cGVcXqEOC0vTkdjzwMGh4xtA3cbYR4u60/7WFn7QZk862aL/ziipzGAOI4Gs4yD7
cEoQl8oL1Mu9ssOLOzvpRQ==
`pragma protect end_protected

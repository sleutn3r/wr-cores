// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Tsq3lROa96flnc0o9fbLjZuYN5GTI2jYPhfRWrtqlU8k1e6nqvuGRZZIrGyIfqpB
DsV970OR4b1JF+IZ0ha1ghYYjPQ4EbFNc1g6WWWqg4TTWiDZHthcC0RsYJ1epvz6
3152xyzaDJNSOnGH17UW/AIoG574Nn4pxPwCZl2nYyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6944)
UW7kgGsoV75p7Fw6okwKMVPkO704PpP8wrpMcNmmL9RZKNPN2io2OYlur35GQ2qz
/dKkrFGp36fkBxrFyGmCHH1dEAGTW2YAAqD9zep7IsyFL4VK17hruPPqpBepYTq3
5M0+RqVB49/1DP6GHInHslNth6IgQ+P+moG6woK2k27DW1nAvSmxF/jnkzNd7VgS
+59VpQfGkXuwNTRAUf+czUeCoJTM1aVujreO5doqFP+cmTYEsAnW7uYCmzuN5v+e
eXwUpf/zUCGJ1hnUIGWflqz3h41/AucIwVcSKRM+uCp2xX7wd1LW6mhBCZ45uRQx
oqvOAcn4mk/ZPdQCwi4DywnRjVNIT2oeybb9yyqr1R7tmk6ZLpVzo/IiZeN2yF0m
pws473dZm0iLnBIvVuqvKS1eOaDsNpzC+M2G2re0n1NgtYejO8Az/8aTm02XnXLQ
Do04nfja1sQtmuB1dgLyYo7u6co2wiOisDGBbwYtTEL4LBPS0SiKq/QtmRrMiBeG
nLgIov71Ky9gdcfti9RdoYhGiz7ZoF7ip0SJtAS3L1LhlIuXw+H/Nb51kl7Lb9uU
sMZ/215j9t1w7qx8X6Nk/jMNj5vSEm+hRMTL1wRQbyO+BFxFFvwqlulBocg6D9I1
MbpgShnZt52HCwXTbxjGCvWejj4oL6+BGT9zMyAPVOrxFKZepAOsLgA5Jj4p7asY
jLHBP8Dr3pvl26jGcXOafuFEcKugwVuearwIzuAaUvp1V7KyU3Mceq5xOMi1VQz/
CxijFO0nim+XNb0GrJtj0XG+jn1EGEwG74j0MhKOnUMTGq2zscmHFKUSa8NVjoYx
2a3csB+YfcgvgA3tVchJaLZoRfBDe258rDTVXVQJ+jyMt+GKI91ODJkKxNtMpPPy
w94Sb2Byh35I/HUmF/s1YmBpMCgvnQirC6Ggo6KMFITapbE9TCaFnknwpFH3HyoG
bt2igQbDy0gqY7BfBPsbcIAXF6NDczusdC3hrX+f9vcVOFeLLycWGFVBDPwDqH+o
BCk2EYFFa1oXiUqrIWBN54swjzXTZ9HRKHvEPxkjtDh7Em3W35PZbDBhupnUtjAL
Wg779uGWID8fdwz+PAQJ8ZW5gTut2daUUak/E9VNiXfgXAdEiD/09HhbP0Dg7tY0
0o46S1PxtKq8H4ZsPlX45ev1qMKXurml3MDmJM3MJ4Rmiw/z+95g5934uU9MXoS8
Y0y1MktPMh80uU6le6jkidRFrPl2OQsoIohHxXg7k2KGKakZOor+ggjCxeaqKgjc
GNMSkgkNP+IC5pjBZALsZTdsETuUXVyUTcAnvuxmfm8etMuN1pHkoRqtj0Cgwvik
NskBGa4Nk+WOnP9peRwuDMAorlzcg0v5iu6xTli/qfodr75zMatL+b3cHyPV0cIQ
WfrtIpEpREompHj4xdyW7+yzkAtJKYpD7y2Dp8gnEJSy0o/U0k/LwffxgZiNBUXb
gANpuHn4sdB08XU5L+KaYpt2mkA53XrcuBxTdK3tBovOur/1QD1MjXhXxsiebp8K
eJjPkiQeG0NoHzbeFpWSzUhgbm66JiEcLQied8gYS4vxc0ReTP9mvVGawPBwck9+
+1eZyQTREBO7c5GeuLbP5PNexzNzG4DoABnhHcD9c4mzSi664VAUB2Yw+WvISWLC
Cj2+9icQoDjfR93x5sCylOy8Y3UzG5wEWEuYYCum5itLcQV1RKL5In6oAWFokVXp
WE0Hsv7zU3ftqXjK/aYkF+Lfo0bNwF6bSELD1yWb+IejnZa24EEqCV9Z4MXj+stF
Px/0XHPPXE5sKVG4nHx/T/RX5hn4p7+Ec0/Yvnbw1t4I1HnG+P1jOnCI8MvauddE
0JbeDasjAngTicKsML0Mk+pFMEh3tVlB/BbgM+PrkNkniPg1BWdTcBu+FwXMajWb
jp1WDXw1s03pVXoqzBx6ndx/2ijw9pY30jSOi2ape5m0uB6PudSzuoDxptRKdrIb
OTXFs40DKqO08s/rd5XRsA4ECyjE2Xq2h8zvhEZfPlur+w9h7bVSijwoGLXAm/lk
unWGqgATIrGGAnbMh0Y1s+hDUlU/VCpI+t968cAOZabOstclXjqFYAuBSLcy6GTr
S3aPGMFE/GLqq9oWKcfo7eCiRhiprWvUWw+i7WZSHvwe5eUx7YVEczi0jycjAgiK
y1F+BqTyNPwfpPKoy0F/MwWqDrzG2buDNt1lLlSYNxHJdng2wTakyGd9HmkkHcz6
37qfbvbcX6fdy+GqLNsKDBwBZE/zaKM0Lz/vP491BSQTO581D1uXLYB2Ng/lSK23
zH+UR1fjpSurgugtV/b1YT+Qr/ZjEQUQsYydK2/bZS02pQzf9G+gSyELPBQk8ECW
xUVm/qRRIav+VCa+CGZoQDVyTTMzOXavBX8wPBqIPeJW2n4c32G8zdhxOP59F/G0
fNRZufaH3moJoaE6sVSIlSfeq1N3YNytvfOTGvdKRD9YsEMS5NHd6eYhQY2FuuPh
oRsaMu9ghfGayT9y2fId4lSrK00FdfdbOYrY1AScK4o6YGdlCFJ3JlZXqsEBnEVx
Eg/KB1cNZ/lc7GIVmvUoFsUOdlfu/MLpbrdShdFebC5xJlNXWHdZ8nmm12Kx1gRM
DuMOrLWUSHZqbFivbeSqjTuQ/yZ2AdYe4/JQkVzi8FBeRawIJWVXdTHlBxraBPoT
MM3ekKAgMH9ZEnSXDwZ1Alr1R+UId2aVS+uidV4Ni7ooe+uY+ehEek9Xdctg6Ldk
hPLXArfw8JLdPJ1vHM5UpM+89hSr/O8cpnLKdXf9lBaibvuWF2XzJrTtjy48w1yZ
4yCqbtBi5YkjH8KG/ggQInDVoenADVAHRUUlYwqOXlPGjEgiNdKp80oIgtK/X5/u
YjMDxSUlZwpCiJ+MXK3PMKj/1+PjIK0V83++/liLqT33luj9Fz1eg1IWc36fbdiY
JCObZqRNYKp6F2NR22n30QIY70N9mXECog+7d20SOA6cLI8aKJ2W+wL/iPBRtiNY
ViPDmdOkDZMB8gvcMg8YIEeyeXezzxfGFwlVDvYU4dw7j2BDzgSx20f2tDe+448e
HSnFGbxQY5ok4ABzqui0xdL2AuHqfG29Y4SmzFnRWenCK2NavDxXCxc0S6guXMjt
oNFSAAkCs0C9Iq98PCcFkQziM7nkwUjVxQpCBOk3V0VMbqjqmAZLHZc69KB3h4CX
zHpXd2oZ51tjHxxAETaElRa3hFN2o5HcjguXOIzDXpj68Y23ncW3+12nvUMfSL3B
JTjP3EFBYpIgdFpU2ZwLeZvvLRItgv65+V60S55qho8r17zzOQehsQ+duhFrjc+u
0haCHAcFzLHHRAlJWaV+HPlJoFxFwtQrYROB/f9pNPIlk5j3tugI/hXIYUo3fEPx
tcIckEq40QhSnxLMV/wwOAFumKivzmO1xHCWulsZMcjiaOasfLVMcF1MR4ypbZCo
Pm24iT1t5VqW/WgM+xgkVXa+Zy55r+kWwtiXFzz5jsB2l2sPEfyWHyfHyl3qCtaH
pfQojr73ittpGhljHZ2vExVfVCPT4nflPWgXgvT4sJt/wUhbg+IPI4CSSr2tjzKL
E5pS5SmaU/k1awOBdUEDY98Hd0GdGrStacKTninJOvzJl6MiRqoy5aqk5W97pZ7R
TnE3lEWD8KTQ35kVnWZ6BiGW8aX1+CclxfAy/S3M0xBcWBKptxtPDOpApOUMsT8I
CaeprOG6EGZIHkZeI+Ugnr3i6tTS/xRSV8/ulic7lxHcyeQ8uGhS6DdDqDy+Fz12
wDW5wzdPMXIV4JYb33aBKc3rA7PNW2j+6eiv2eL78H7nI4FvKwfLFao3cQCzX0iU
AL0NlE0c0zPDXKQ8gXyMKoRRxEdfYjI9yMWqETsQSZx46zn7szHYjBaaUYckMqEO
s9MN6KfrMnSotuf/gd+ESiDZkI+Gs103tdNpgLhewDRgutu51bW1CK8NlGjcOBUh
YxdZ5f/xp8AA4EGxBmU1sO2gBiyWYUe85QWY6TiqJkOZ3QMTcLLvM8BP+PETF8Nu
/VhPbUQvk42h2m5HoIOCokK7OjIeeej8jiPqq5XzXjd2unTBZIl3Is+LD1uBPayC
EKzU9Ncp6m7F9tKglyrFVb/56OtYjH+GGrPK6iM+u7mqpkVee1plq3477kca9xfe
aSpNH/3+KMd96QrEGR8jd2AZ0tlvQnzTng1zZXTi+fhf+7hF9N/AXJWOe1oLasB4
9tlpBDsXJQS6fnUrnzg1ohKGqqVxf0dt3hYM3Gu4ExUIQoOQGMrogO2CIgkcLadL
2aeBAKiv4gfISPM3zQJN72aG6juAWMZqNpn+I6NfiN3qP6J2mHQG9C+/0N12rmgj
jXnIH3VvU56lP0bLWlnm02jB79KkmIWQUCiFaE5U2FcTEgxnbhGc+3d8hcI5ITrQ
Ite1t7jigEd38vHP+CNVjTv5hpvYmi7v9i3P3JQDxf1vxdfrs4UpHi6/MmPy9jpJ
u0mIXxqHB2dQhptxe6LFGfFXJrvaOOvQNbzVpvSWXV3DjbtUlzaA5msfDNagbX1W
DpA9WHMoAF4wZk6wm68qscPGKXrk79w1vUc4G9rwNDfkhW8vxG1yNzVc3umUsxF6
tDOLcsvFty/XGpAj4TnywxiT3Uf4nWVl0iTRna90cM8EP/a/FjqjLdwWA7Yqjz1z
yW9QTdjcTXJZKG1CnUviz04vy3OHP/u9HyGOjJe0PVJNlLSUbDpR7T7agw45Tec0
apVVcZc+qGeRB3y1PpVLuEWOmY9K6+IRcmmJ93yHHL9mUEEvX6BJbBP5i+X2r7jo
C/WSTZR1lOKnmuigdpRajZtuckRUKbxXIRrsLbJehrbgvPWGQMeKz98x7MMa/z+l
YxCzrZmIlk/dXgMIuKQSH+lcbOLWV2ZXyJsLgBuEGCzoCR6hN/f9gt+P75SxTlG0
4WolHdOFD2T8wbkM9pJ/TU3qnOMdtLZjr3j4iUaiFTWKNwfaKhEo5EDb7pZxt9NH
dd/SPfiJjamPnR/bm3kI92y+gKSgCo3ICWelOwf72Cf4dMT5FIFToOD1pK3kLE+x
sJ1F+yvTlQcZ7RdlehSYyRrWEMQDcyxICFE/ydXET0KdQgLyX5wkBIrADFoLRVb1
CO9+D0ZE8fXTqUjt8L9dtmyKA5b/5eBohAOlznJdU4fjPES9AN8q7DGuNU+ACvbM
LVNnWVPq7TXHOQpaWLgon2VPVrVaq0Mt+lJv6z87w3g/hP11F3eeNA0Kc/ebN4UO
x6/6QDnLe7syuvT5Y73vhZRjip9Lof32X3QIAsSNbHIVxUMO10eKc1IrYvF0NwuG
vy7C03cz1or3+uDSI8zMyPLLiM4PwE1PIGiZTmtws1PjxRCU1PRF7jY82ZQlbahC
AZZ2DsNBEYq8B30En9uaJP0DewTqUhccARz0g2888a5t+zqNRfRT29bYBoRv9376
ch9vbDAoR1wom4w2Qynl27tdCz5MbTKrMeJDo3ij+0x+EBvPUZPosMZc4pWYMscz
/oTuSe+AZWTWx12zF8koHlNswBoQ2lfBvaMUU1XFtkoLVdOGYA7b3eqeE8ocD8h4
u6ZcvoY2YynxZ1Q/TJazQVaS3nLfOKg6CrHI760EwDF9jYsDe4H8t5kXTZwrr7NZ
QHwnQKdp+NP0KO/Inuk7oDRLXvaJ1L5d+QCPrnIK20mNRIV9WFABxzBfpaY1lHJy
m+r2YQLey61QEw9BWhxux7xgUFmUi1hm5VmOTUPYTJjb+8LuUs7Wi7eexEXLQ61p
uuN4pwUGuJorzVHAzCjVLqxItTD/FKDkUTgFRjfmPO1gVSVs65b2fKbtN1MJmWBx
f5j5VJadmAlmdJwTTMAnZCWWIglW7lxCmivVcZLl3Jtv+nAJqzV961RxNhxgvy3q
hGBx9l4d/mKPC1/jvjY7GYZbrNzRkqCrw76ZhL4IIlszzJ0mJWU6iwIn/gsEzuQ3
thcfPHM4qHPcPewxT8jdBNVhsPWp2pNZGaapiFQdEOLiMI9ZXmGpwLyX5Fum378X
Pa/pSgGhrD7vxWJaA/XnqnO0IcXsf5xfCqP5d4oHLDiTY6daHUDrjbCvTRcy8mB8
vriYbqIrY6peeRkjBNC8PBseZsiwRrW6qA0dHWa6KMGBsvd+4/x2B6me0hOa23OA
STt9YgTtoKf8BEcVGZLTPJSaIoHzitalNvvUKzBudh1UcUkliUJ48FWhxjEQ9dvr
VB70H3cHckEeHm0s0N/dUE5+tBYjD7JLklR0OxQPx1npHaL8HD20+lqplviwAANZ
GHlmoAUeDQBq22XfaKdWfl7C1i0Zov/F8/TkrtOneUWmvoroJZ+BAzm0Rs8/vawy
tiohDt7GjigP9A43e6gypH+rp5MggbLKY9IcMTuuJZOp5cuO53sijjAf5qmeph7d
EsV8daqn5XF8TMMce9EBriK92H5p/Ui6rEIpwewM+90mRdA71vzv2tnUm41pvYFe
SgA3YyRFhxS56j4ngyOBNuLoJvLJQnBYyAumnCq/CtF1nTWqw/etnTJg9kRfJMAN
cpOehVCSDNrkEPsSt178JRy0SGfPZ03t/TBzxb7D8W6Pzfw7udjbIwShmeDZhYtm
f1kXX6OSKFYu9tEehh/W9xw757sa5Etu35TMVdCJUbuJCQ6kMpFkpt2SNLvyuMup
Uo9n8q4uHWI0K/5YWiDi9mX+ZeVMrQRt5+FFdlzMuIY3Zg9tsGQRmk/+9TLm4F5a
WNjgcajgvyBCaFsynuUOXmm9n/sEqG3PUinqZHNm9FLCeftRYOHznETB7TvGTi0W
AdFYAPLNjUL/BOK7ufdJC5S+1pAVzLZLlZd6jDcvhqBs8o4GQmhJVYa/6G6OcJpU
rLZpyqv8/frsbN+PAew2y0J3THvKB+yZopNEb8Srcv+RxqK7VknJ5B674tanwqwa
SU8SjWIRRu/D+M6+bDtgoPkMvUmcvHl5+/AQw2iZeBwM8jVBNIXdN04AlwJSIqRq
9Ea6tiA7WmBJhng7NZJVCEE0GNYCfO+i8g8emayT7wCY2VlKxLk+3kRgDmO8GD2B
uN+GGD26nrL119jNjBaUmBFDeDBjeuX8nzGGWMYs0CD9aOs0zKEBE2TQmAmn/w7Y
joKsYqfrtJ2lywnMqT92KXJFECiv3c554WgY2VF8/Em0KrsVh89ubIltZhedvJA2
YCNQpJ7U0p80eUITlCQSk43+lw3tY8GlHa2t3GjPGidIMJosKK6w+cZY9QHWncw6
JMnBagh5Ywq5vH53acT79oidwKRoUUijygb1WAZIUeDwTggQMjA5Hmt4AAR9A42W
06324tAzO1GkfCGrZHiX+ASNvtH829n/U0rilSNZu1rPxhIIS3mL9wBa9h7GIB90
LycF/8LHRKU9ByIUCV64uBb0mOqwE+zyIyI/XmSoOObOzmoxI+5VNsKDEstE40a3
rLsl4kZBFcNusQVEEEYJMcX1kHPsK3cbjnKGAuEReFLwg1ilQ3GCAM4ElDIXUfJC
6fSODX94KaF85Puc0UJH/S25XcdZWiWcIRHhCvhoEiVZWl7eZez7Y/5ELb/kVd/Y
pMwmIivxrWk7O0pG5JpOmVl73NSBMW8aqv9wJYdCYFwziCTXngxVOBR9R/Plnt8M
X7wXq3zzrxkV3xkHRTcYJL9wzuy+1tEEu5dHTy5EcvbUG/ZV06C4GeMrbAG//Jgw
2mOeoRQqaEeYhS7rsjEKryYckTTTb0jLpHZvXrVHH7myGPO/NdivHsqBi70Pruvh
Wu5AGaq/KvmMuyBTTBl5KPuW3yA+UlyvZ89jJsZ5R+uHMD4cujnwII9X1v1scny9
KX1FJmBn4H9oTD19pqtCulz1/3aEm1bQoAChw8DYHGwLZPJqRfjh6F10owODGyY/
1nZ4WnZW55gn5Z8vZCtFKRY0kOguchPy9h1k80YTex/CeefAGesh3QTMrAR7uC+b
tNZ3V5XD1HuXa0FoXs2AXt52kxww3qK0CllvMA2ddANlqqXTgKC0IfE/Uzo11nt/
AL+nsBQOX4I0ve5dJckf/UcckrJtPtbx49Lf4TecENfhdDvO7BotodDz2BFjQU8t
OFG31fSBneHa8pxUwIYiWLUIAlFeGs271xxkazxkNBQS2yeiOh/jikxuwJThEhKp
XIB4ou2jVaUYBFN3FcQAERRZwCVml9r8aiGv9H4MGhOOp0kLfzV69VWfKgvnwz43
GjfLjcx7ubjIXwsugvwlNEDvIjUYCECwWCshiESdp61qMYU2B1K6kNWMUq44nkKA
aW7msnRQYW1yqCQW/XEygJ4YOxf4J2Goz/LyZLqnzTrbJ+vR4sou03480CcXft6Y
Spe1Ywp5A/S12Zw+PZm9dlGVYO5UZTPgvJYdHh90g0LBz8UHzwaC90ykqGaETvxv
xyE/cYNxIcWovHihlt8x9QlubvDaz9ppoewIJhjxTg68fkOyO5dShPndvdHOihlr
2XlJvQ1vDSu0j6Gn/PGdOUepXC6C5ToCmBQDHKqKFtidCrrtxjKu1u2sZ5/6BmAH
ULHzOiD8wMFYQ/lfFa4JnQTL1KVyGUERP+DcOrTAZQtEplAbjw4DNHypjciSdT+W
5v6pZFvgK6zUYa3m44/Kn5AaMB6JN8IT3Llx2BMGRPozczdk9Vh79FKD/8SaNOc7
7CfOoGqprcsToJ+rHVeMsmx+PxBDf1f81rWbZuZdi8NBObGPBY+R5gzsMevoSMWw
gdnqyQvtLWEYO4LbaYHVxbwHHSEpugf/Zb/XlDhGiPMrbCorNvkgPllF7HDFVu39
AeQKi2n2EvnikjCjIcUZMuRN68Ukh50TS9CD2GWsZ9B3Il6j+OaKIfKPd68gjvyo
7IWYVfjIcMNpFCD9JDjp0CGD9vMgpV8opJKheiQUQbcfsyNpX3iU4d3dUsBONa/R
fN57/kG83vtrJ/aseqQG33fkR3/mDilZpsmR6OKRRVtAtdjhq59tSi63b55O2mEt
ZOlSNZEZ9z+eTReGCv+7vynJZx618H0gY/y3ptl2n0bRkVEmP1hHAY+Ic9nCU85X
hd8HEd5Uw+WBHL53QJzhUiJfwosw6A59vPkX6qtBTdbPoNUPTe3PrLL6GzyPzMoF
NASxhVT1/CPmTDhlVeooRp6s0LdZP9ylw0m0udERtoPtDKnJyUBfBZTqi0zj9JOR
P9Z/YfG8imjeGwpqv+MFHdKACd8d0wrJKxeehziLM+IZ/XXE6TwQ4A47EetFA5C5
Vjjtt994SKko47lL+re4dO/TUBBlvPScf07zfbHXX0k=
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:38 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DL5aCKF/3wYHD9ZuBeZSnuGcbb1WulfT2R0jtsFuxiubwa2EJyMqJrtMJe/7deUf
3IF36sOTP70UOw/CMmO2xRi0WjETkHt7QriHxgIifESyIiSl9zV1OYMJtf/SRHTh
tBbyDvEgS2mEF96jVE2pSd+o/5sjb3m6zX6PT/xSq8s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3216)
QdoPWNu5QvcRxhnciAOivBilcq+8xtn9uTc48fTIoX5MYDDuhwkEkhSRpvmOb3O+
+RSOCBREZE4QOTCQ8ClovDB7XDEJb/QlmgLLT6omlWYLwDCXCnFCLMi/TYDwXZIY
Mx2ksvLbzoTl+JuMPBWXVYLASHJGnMLugvmORSk2P7dOk/9t68ZQkhl8R+3QUnjr
MHGcrE009z8MQD3ad7ZzgfWKW8xjzYBKn/Y/UUDLtNed33wh+1KwMv4s7GpYL42O
oaoAC/GU4huRlJUpfpI/MdZMH4Hd4cbB/yVEm3M+Qa9tT75gpsmOIK7wn279aEB6
ACMU9rgZ4JtzXiIwTmzDNLx/WivquBRzo0+hM/97xL8lzVoKFQc0NZ1KmmxmiJ5C
Xt1PmdFu+rpImcwXyWZ/0+lKdqnAGuLfGGVghEuqOQIbP/E6Kkhsy8H/RKbZBkRY
3KKsA1G/sHltZdcYm5ifTkNjsJyXkN8DejsQGj4E55ipGVYw89jvMTTnTJwZujwj
HBL/MSgQffE+sx1hpNWyGHb5PRWAlZ7WbexiFmKoXDjeEewWZ6XEuDGX3LanpB0F
9R+zwnh/q1fTmw5/t+90Es6hueBYlvUJNqGCb6Agz+bCS/2JqZkxdrZhqzDi9s0l
+TWujnhiKZQIkVaCRFur5X0s0COJscnxkJbc6KKm5xv4LB1fqafqgtwp/9SJ5BhA
bSXHia2b14WzbmbMMv+jIYx9FtkG41QEHNtxgti3FElhXc/JPR/Cj6xlzlQX6gfr
j0lDYzy8cLxGoQe7+hFk1x6JPPBG15CUNgG2fHqIhRvDz16+gumz31CQfTM3xI0J
wWu0kuGUs69ZvJLedhOMdvzDw1vPgVc+Vwu0/eqHmFmff8CnV9KFKFIv/BfRBBzj
FRAHfIfvpBxdUUifMHf11liXCVpM1R5D37N7q70QY1lU4H3JRnlgwlI94FddWDTF
89sc3jHREA+9rpf4vWaKeXhfaFEzMNwUqQQKnWIdG1NXScr2mijYr5qoIsNpfY7g
oZsSTEccC+sFVKAIjGuDHgVC6hGLR5WWEpmQgtHocgrgHMI/DcsYDw+j/BdzQa3M
1zyDiYDtYkOpP3Mh2qUrh4SFSVWLD+fn7wFzTEtJQs2jsG+RF4Ifca1Wc/QZhwjl
qBk6NPFp+tqs0FpiDKY4jMtfaHuVnsd/2Mi8qSK7ISqsBLZC6p1CbHNlUOyYzty7
QmTDLbaGjZOsyYR6FRl3nLVPQwkmAUoTarG41QipYEJopUWb0a6wmZPMPwkXaNGl
BWKNWtC30UKgTn4vsxbju5/n7jybLkp9644mB2QRNl4IWsSTOqugLHbC04NK/8fh
jNzKmG+4zcG0QQvfkQi8vQJt2tCRIVanj4RNW12hw/WrvSYBzjbLhQxGIaxiKdyC
ZcrcGUnxpYdorIZVewjEMwSiqWXc1ygJ81Mu8oHytCVGQUJvfcn5hkSgl2sbvYiK
kH3Ft9lQanRaBMekJkalkow4vF3a2he4am8jy0RxbfRtkZttlqeqNxH4eE/LMlvJ
KTvWO+5FbAmaAKqcPUnqiasDax1bvC6DDCfMjsFmnRTGQqWjhVX06DxVMddqtwL+
4//Pl2ATKALd7owjazCHFl3SdbEoaQd5TNB7zbv1MsOWdvh+tj1QXveZbeZTS7Ul
i+k/9tzyyNoDPYbzxUcO8YLutaGF5Q+WzNH2/8A6plBLnj8X/d+85icUDYmgM/Y8
lL57MBtHqpEhoPM16Xg2Zjvd9XYpUQrY3um9fxM5pCD+0Y+hVYbmPb6kQYektz5c
SvYbEdt6m56N225Nc+kyDErEq+hlel9oVyLTixypX4sJmEuv/d6cXywYS59PoTHM
P5woGi62H1FwVIAUtbmxPU0ve/oLVlbJW7iqNUDJUOZMbe7hJaRQyNTzlXydcwxy
UaBunkg013mkIRsLcQtVsSyr//pdSdPf96YlZcb7xtxJYKvXXqDKMJLucdQIsHfL
W8CfzTaBNSwFHzyILXTZ891HetvNmDT46pH1QLXiuReoGN/kYoVLfAN/1MrrmGay
ElmA6uLGcl55Dl2e5PHmLU99xFKLYgnJhJjeomyaSztVgC9R1EQcX7/0Wk0voJHK
SJbqraLS/O0DHfIYBn+Jw4JRtjvmc3GQSp+D32bYv875SU7CwYs+sZd/bCcQjr3Z
5nA20tTtoX/qqvBxXBTXlUad0/TQ3Oopeu2aR+xMFpXVs2axZk4qkZ0n+27T2e72
ojC6syTYZtlDrBwf/xUksYmPWlW8YaOa55viKduhGLgqwbxF1YsfpbS/+C1kxLft
87lHFIvhptpqk4A7Fany9UEaHIp+pKj1v7VRPhD1feDBDc42AIxOOVj3jDzMWned
iW6xjt9pa77J2p4DYg0hrCrojqDRpuGQv46qySC5DppRV+Ce++Cq49AoBVpmpV8t
QTIV1hpWgka5R6vX1WeZJRQn1THkLHxHztH1DJDZDIf8e6S0lAFd2BvSPI39ERZ8
y+fZO4x9p19QQFGhisqvXUvfs+bas3VpGXoReJoLgHxBZBAe9xStqeXy2Um6Gy3d
63sclNTGGQL8cCS2y332Xeb3rEuOKIefXi3ES1WjQ9mBAQoFqBV1v8ynE+O0Supt
s0LES1nJiU4IhCQlVhVLgs8jmLws5vQvbWFOUp/joblVXzoombM5UUSZ+tfWOxFh
Vr0GHCd9whhBGSRGCA/BhPcu0UxEy3/5THztHYf4gvimVPiIjFo/pCV0e4WeDa1z
FKDzP6qTK7Em/sWSZOcF9Pl5TQ4kn1p7qyLLwOZ1ufqQ0pml3BXIOuHsBSNxHGzM
JHjiML+SqwtZl1pf9rPedVWT8cFAuuEt8xcf2Ko5hS3LuQh2UUbkbBzS/WWt1GMj
oT6jWdQ4iOJxBK9DJClHK1bl8ql37EtHvzMYCXx1atH5UpPrBMFDgRaZzhWKz5bG
c8+B1y6EWXguCgXqFB+H27Z25wSSJelHpuQ1jN2NnokEL+uefG0MWt9vWCnX1N3G
IAMYSDCqopjilv8fd3hDPT0JyjEFHXnz9O7dUfMeYx+Km5hJgH9lobrwUjnungXu
Yxx2WJbxQt0CPQcn6bevEkUWW18JNA3xbnvMnzYXI96e3i7AtlmPZJtm1AjvDTr6
w0UCfHJ4Hy3pc1nG8SVEUORGDnAuvosUfHnPKizhC5FR7JqxAit/16iiO3b63yIM
X6P+9YAvPjb3eYckJ/J/bkA0ZoNssexJ+C5nph/adxEBIgElx5kJ0uy1w+hFcbv7
UsKyGdJbqtJrpGqsI3b4xaQMDNKWFB3BdjOz4iAENGaZ7hutP4xAViqHV807o6Wi
kerMbzQ9WWoXj95zQPY+BVzXG0e3rFt1h7x+Ql/d+BMrpo3jilmyAgxTcwi1uNqM
P6IbsWPfxzSQNmU3E31JTSK1h5Uy9eVy7PyskVcCicT7XHJ4d5HXfkMtci2sLYxe
8HJUowP81Uza63L2cycq78T5J2BopMaf3YhxO7oDXniuao7SsQa7CwCujiMnAtdp
z/gio5J03xFmSd5TGRTlcXqFdGS8qxZnfm2uIK/MMxKfS1tYoCxFi1icOhQN90pZ
TzseL+4qmUTjeuRxZqBS71441kn2Yn2eVnFB/nfToQ97/73Ov7OCZGX5bmW8m6pA
Ln5kqTkyN0IRJFrnajPjBGPFOJE3S5UvpEbsKKyzmqxQaDx9+wUnOLI+QVc9iqR/
AKQaVPowUMV/7I21qrJxXmJuYVQ+ESb1G4nSizDib+sBBuXDKjhHZa1QX2dTZhsQ
C1CLE9Z+N45xZkbnOgby8HwHe5XUWmIVUcCD4WL4hPE/GqfByOyVnwnWpuSkanK8
9jNV5b2N3zhsqw1YvVcSXtxKrwRre2SS68+ydNbS3SX8L0uBABYUaCSjyigCfxbi
XDM0yfZwc1XaX6Euxe8nRCtZi0o+ljtvNL4Hts28E7IyZKMm+YuN7K/FWvQopnWv
wcaks6tE6Tc2NRrcvbzyFoWjVeHc2/HG95Pesm4d/JgIzmnswcQBUgLEyuNAVFmK
m/a+xaWoGRWH7WCQMxtS9AnnYjfNTNRx3AnXPyZ3svav2uUKBQizDOPm++AP785x
Gpdz8EIbWLe4bV/PbSx7SIzlZgkhqE96ExyEVh3lHsCI1QKFZXTdGTBzug9P4xqH
wsD4uZiRAE8qizTfDIUyrV/8M5nzim1PhJBAFSodyi6KklpO+JXNsT7lnfqWbzvj
72iILocTewW5M38O+3Y9/8Y5Q6dr/4KLPMgjQtXbwIvNCMd+lgDzcMlFKYuOBi5g
`pragma protect end_protected

// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0.1
// ALTERA_TIMESTAMP:Thu Jun  2 05:35:37 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
oL2gUULlvoreXAj98/1BulcIT9gfWMriC7f2DDmVWkyb/CUMwGBcn5Mn7kEYOvC7
0sWxMA1CyqNVAMO97ITNcbTRmq19Ml7XkH3BleZNWrJqmZsiDcRCl1ZfGtWmjTud
ZgAO9eArgp8i5oHXk8a/qfNWq1vHtPffl/ysn164mBE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 1728)
CBbIFTl+HDxXfF7nAinQCdbiGQ2xwKIOa6XJNcrN//Lu52nrRdilft/zgmj0AYhn
2NziZ8IBHOWiGUSBPbF0BapMcJJmIyApErfM7hNDkR0QlpMsWJpVGOuf1XHPElZZ
L97drqFGqHjCqLIifyjSva9+3OnzJoFYlDtVzTWj/x+27xrihNC5+u+Ri8ai7RGb
MyTBzSJ+lGGdJ/rJ1TBgpSWXVjxy6/DpqmMLUnbEFA9iSQYHuHbv847Vw1w6f4fC
U9vX4QwQ0D/JHT9vZzcMedWJCoCpIADAetBe7sMhnthRYng7rj1SX3JYAGVRk/Gz
G8q20TCPgaVRcWIk8U7TKsJShwy3bN6f6bcsN3oeSzX4PbuBC0c4Vm09OEV7/BYI
w/GGw1SncamP+UlhwdcNUZa7kix9rKHyOinENg+HE4pESz6e0mbfeKXg0GDQmZo2
3S/LckLGWzoHHpTfIZvG9B0HnTMl4bjpVFwA4V8TMsvhnMBoXMuBgLH0qDIUBO3B
aeu4ERWkTPI9kdHesS9piWymUzFJBz5ZADmVBhU3e05Obcux+5m0/6PlsiZ7S/t2
l9ZON0ArqgKnFUTTbEY2JYFbtYrWdsCkfafNAr28dA972iqvbepeXqqZwmZgYsDV
8pQJOq/MIg3Cv1zb2GizCX9POMMq2nM4EKXRhFo+HZ15DmiPaYAkXQyZBoMBF8id
DNq7/0YReX7oPrNGvPSlI7C7+ylMbfWVSal5DkxQaO6wsJa5dg38wA7PpVpH1rAH
QEUVWTG9JvGVEDXjyGsdegkQhetJcVS7D2efsdo2CJG41fFDSGD9EWuX4HfGMsrR
3l2HCJ0Aot6AArTHalBSYpNlngCnzJCg3RUlZUE9ll2LUHYDcZb2aYYuC2B+vuvH
0kD/T51IabQZkq8Q9cVxyWxgk5PTnTYROIam1NWsmfmAb+fZn1nLg7JI2A6yOfhI
M928V+HpuUbasmSTedogGYCRMGKHWAhSrOvV1DzEsDv9JRRJGg6IC+WwDu3n9+t3
d4ITsTjwM0rnb/IkDbLboHJvAZuCauK3FqlaUNSs/1wDpi5C8MbiF/8w6MLOCKW5
OneTm6JLv5GKcpuutHWp83w49bDBbj0/HLVT60N1FLHmB0TuZteN29koRyT/a42o
jVWVnnnvSPtcZGWhhF6hYaI+MVa95UEuUftvTRk2UnhM+AZ0LUJON5KG1GjUPY3+
iQvWtVRgssofw4WGfkk3tKOs0gGWRQ/e/Kpo3iidEuXrjX2h17UyBwbHg8JW+gK0
rMdJNQlCTjahSSsQcBebf96CfDGj62eWEdqGhDImf2DMp7SkNdS8Ppzbv531Rysb
EAnkEI7vmHYw8XtcULou43N8B1vGQWkKhNPhkyaieOg7z8j+cHvaU5Mu7/Wun93O
muK0wyvDAC0wUWP8+RdHHGEEKtT3yo9lr9mUZn2Ky9fqRMXPjQIwC1IWR1FQPtxY
gt9K0q+7EsBG9qFbya85JoOsj105U3TC+rWWqykbeQAzLWIYEhivLlpr2wrPf7XM
bK1/dhyKFXpB90/Mkuf3KAgdR13p5NYCH4gkT1j2w/BEo+HwbaiPie+yVlKd5nr3
HIWmyJVV2qcBUfSeX6L7g5m70YTit5zhu7mvm71kMzNMdifchCWte0aw0aSBPl/x
ztSrEu22Z+07Xe+kW2jFUOTScR+rnB9XHACgaHVdzbJYc+M6q7ZHuts4Gd50iOKL
3LwR3WeXfIXpwhwaMBlK7p+7x9inezQbFe/l4jtDh7KJefHvpOUlQikjVn4f1J2l
kBpogiSY4hz5iwYbZZJBaGWkEPZRuVy8YrqRk9hnM0kuTyssvLggUqw1OwP5nAe0
IACAibyuXPIoseLzQZh2J/0odG7H8aDSeyJ8wMqVxtkovYSJo3Vncb8BjGxR3n1g
5yMtLn5efMqWVq74iaSGzWf94oOsEkwdFmGF2z9Tl+UQJbTiY6kO9uCuX2wRpuof
icMMYt+yGMEI5Ur1QS06TWOx0VeU9lbuat9BNVallonDsHVrzW5jdGsv4L2YlN4I
bUysjU/8Qy9aH4bGYayh34cOnqzqUNAibB/rg2CzIOCi1wTPd2VKdvOzwgUC7gnn
Pz0TVphKSCzeTMGV8bjJooWPAc/rKxHgiO/EYul2pqljYDzYcUmmWIOg9m/iKoe/
AmJZhYXsm2qt3ROMomCQxWiD6fRZxHzWHvRQJkIlbeaKsYHigPRoYztFvI/v818B
pfiNxefnNfs0fYArFZFOuucr5YGH2IhJPXPnn0wA7YyGuVuVrDFqBg7YRkrXOdFX
`pragma protect end_protected
